module basic_3000_30000_3500_60_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_1155,In_1720);
and U1 (N_1,In_300,In_2082);
or U2 (N_2,In_450,In_84);
xnor U3 (N_3,In_143,In_142);
nor U4 (N_4,In_348,In_2274);
nand U5 (N_5,In_1016,In_464);
xnor U6 (N_6,In_2836,In_1413);
nor U7 (N_7,In_2832,In_1925);
xnor U8 (N_8,In_885,In_1697);
or U9 (N_9,In_423,In_1133);
or U10 (N_10,In_1173,In_2233);
nor U11 (N_11,In_419,In_1663);
xnor U12 (N_12,In_1354,In_1539);
xor U13 (N_13,In_2901,In_1807);
and U14 (N_14,In_1646,In_2934);
xor U15 (N_15,In_2382,In_769);
or U16 (N_16,In_1740,In_2606);
nor U17 (N_17,In_1027,In_2527);
xnor U18 (N_18,In_890,In_2138);
nand U19 (N_19,In_174,In_2314);
nor U20 (N_20,In_356,In_1296);
or U21 (N_21,In_2491,In_1287);
xnor U22 (N_22,In_2605,In_960);
or U23 (N_23,In_1000,In_1426);
and U24 (N_24,In_479,In_1398);
nand U25 (N_25,In_2219,In_2120);
or U26 (N_26,In_2347,In_2738);
xnor U27 (N_27,In_355,In_2391);
and U28 (N_28,In_800,In_21);
nor U29 (N_29,In_2542,In_1323);
and U30 (N_30,In_1896,In_2511);
or U31 (N_31,In_2764,In_1943);
or U32 (N_32,In_1914,In_1862);
xor U33 (N_33,In_1144,In_280);
xnor U34 (N_34,In_825,In_2018);
or U35 (N_35,In_1057,In_546);
nand U36 (N_36,In_1954,In_2506);
or U37 (N_37,In_525,In_2717);
and U38 (N_38,In_1606,In_2869);
and U39 (N_39,In_1192,In_520);
and U40 (N_40,In_30,In_2766);
nand U41 (N_41,In_2486,In_1972);
xor U42 (N_42,In_335,In_1736);
nor U43 (N_43,In_942,In_919);
or U44 (N_44,In_2829,In_2621);
or U45 (N_45,In_2865,In_133);
nor U46 (N_46,In_1803,In_2243);
nand U47 (N_47,In_217,In_2355);
and U48 (N_48,In_2648,In_2841);
nor U49 (N_49,In_236,In_812);
and U50 (N_50,In_1864,In_544);
or U51 (N_51,In_917,In_2248);
nand U52 (N_52,In_2808,In_1630);
nand U53 (N_53,In_1279,In_2263);
xor U54 (N_54,In_2239,In_1153);
nor U55 (N_55,In_121,In_1224);
nor U56 (N_56,In_106,In_2064);
xor U57 (N_57,In_1719,In_2696);
or U58 (N_58,In_724,In_1592);
or U59 (N_59,In_668,In_2266);
xnor U60 (N_60,In_2848,In_879);
xnor U61 (N_61,In_908,In_526);
xor U62 (N_62,In_1686,In_1995);
or U63 (N_63,In_781,In_549);
and U64 (N_64,In_2455,In_690);
xor U65 (N_65,In_2323,In_933);
xnor U66 (N_66,In_1613,In_1198);
or U67 (N_67,In_2207,In_2653);
nand U68 (N_68,In_126,In_1231);
and U69 (N_69,In_2745,In_480);
xnor U70 (N_70,In_1145,In_934);
nor U71 (N_71,In_1077,In_1432);
nand U72 (N_72,In_707,In_2468);
and U73 (N_73,In_224,In_2060);
and U74 (N_74,In_1301,In_61);
nand U75 (N_75,In_2163,In_2927);
nor U76 (N_76,In_2538,In_1861);
or U77 (N_77,In_113,In_1724);
nand U78 (N_78,In_1434,In_1572);
and U79 (N_79,In_874,In_2693);
or U80 (N_80,In_1271,In_250);
or U81 (N_81,In_1588,In_1444);
or U82 (N_82,In_43,In_438);
nor U83 (N_83,In_2695,In_1766);
nand U84 (N_84,In_1113,In_1851);
or U85 (N_85,In_157,In_789);
nor U86 (N_86,In_1614,In_1635);
nand U87 (N_87,In_35,In_261);
or U88 (N_88,In_1787,In_660);
and U89 (N_89,In_1919,In_93);
xor U90 (N_90,In_468,In_1784);
nor U91 (N_91,In_1013,In_2994);
or U92 (N_92,In_1523,In_2032);
and U93 (N_93,In_147,In_1496);
nand U94 (N_94,In_2657,In_207);
nor U95 (N_95,In_2877,In_44);
xnor U96 (N_96,In_2666,In_979);
nor U97 (N_97,In_2533,In_1062);
xnor U98 (N_98,In_392,In_1639);
nor U99 (N_99,In_1875,In_1424);
nor U100 (N_100,In_2598,In_2311);
xor U101 (N_101,In_1343,In_1473);
nor U102 (N_102,In_2188,In_2881);
or U103 (N_103,In_639,In_2985);
and U104 (N_104,In_1440,In_2281);
nor U105 (N_105,In_2579,In_2958);
nor U106 (N_106,In_502,In_823);
nor U107 (N_107,In_1723,In_347);
nor U108 (N_108,In_2780,In_1239);
nor U109 (N_109,In_1928,In_567);
nor U110 (N_110,In_2149,In_2061);
or U111 (N_111,In_2814,In_912);
nand U112 (N_112,In_1429,In_1642);
xor U113 (N_113,In_1662,In_2264);
nand U114 (N_114,In_397,In_656);
and U115 (N_115,In_402,In_1753);
or U116 (N_116,In_2931,In_2249);
xnor U117 (N_117,In_2576,In_1876);
nand U118 (N_118,In_1560,In_2801);
and U119 (N_119,In_2171,In_2582);
and U120 (N_120,In_2735,In_2842);
nor U121 (N_121,In_1268,In_2936);
xor U122 (N_122,In_1286,In_1699);
xnor U123 (N_123,In_1061,In_1566);
and U124 (N_124,In_2275,In_1237);
nor U125 (N_125,In_506,In_437);
or U126 (N_126,In_86,In_808);
xnor U127 (N_127,In_1500,In_340);
xor U128 (N_128,In_867,In_1311);
and U129 (N_129,In_1958,In_1508);
or U130 (N_130,In_852,In_1615);
xnor U131 (N_131,In_2057,In_1240);
nor U132 (N_132,In_530,In_2493);
nand U133 (N_133,In_2262,In_291);
nor U134 (N_134,In_2119,In_2078);
nor U135 (N_135,In_1438,In_2000);
nand U136 (N_136,In_1172,In_860);
or U137 (N_137,In_279,In_1879);
and U138 (N_138,In_1392,In_197);
and U139 (N_139,In_131,In_1107);
nor U140 (N_140,In_1273,In_2840);
or U141 (N_141,In_1859,In_2652);
or U142 (N_142,In_1945,In_982);
nand U143 (N_143,In_2822,In_2310);
nor U144 (N_144,In_2379,In_1880);
nand U145 (N_145,In_1507,In_2101);
nand U146 (N_146,In_1718,In_2234);
and U147 (N_147,In_2287,In_1364);
and U148 (N_148,In_1481,In_206);
nand U149 (N_149,In_2041,In_881);
nand U150 (N_150,In_1357,In_921);
xnor U151 (N_151,In_970,In_949);
nor U152 (N_152,In_1217,In_1589);
and U153 (N_153,In_1658,In_951);
and U154 (N_154,In_2410,In_2727);
xor U155 (N_155,In_2369,In_1380);
and U156 (N_156,In_134,In_1041);
xor U157 (N_157,In_2482,In_2459);
nand U158 (N_158,In_2962,In_292);
or U159 (N_159,In_2919,In_2940);
or U160 (N_160,In_2467,In_278);
nand U161 (N_161,In_2589,In_765);
nand U162 (N_162,In_2245,In_2307);
and U163 (N_163,In_1253,In_826);
or U164 (N_164,In_740,In_2267);
or U165 (N_165,In_1490,In_2296);
xnor U166 (N_166,In_2202,In_1556);
nor U167 (N_167,In_2004,In_1583);
nand U168 (N_168,In_219,In_2981);
nor U169 (N_169,In_2403,In_1281);
nor U170 (N_170,In_2327,In_2671);
nand U171 (N_171,In_1199,In_977);
or U172 (N_172,In_706,In_2448);
xnor U173 (N_173,In_1325,In_1913);
nor U174 (N_174,In_993,In_1968);
and U175 (N_175,In_945,In_2599);
nor U176 (N_176,In_550,In_2117);
xnor U177 (N_177,In_1608,In_1540);
nor U178 (N_178,In_2803,In_25);
nor U179 (N_179,In_67,In_2546);
nand U180 (N_180,In_2535,In_824);
nor U181 (N_181,In_1255,In_9);
or U182 (N_182,In_1361,In_2744);
and U183 (N_183,In_1670,In_2989);
nor U184 (N_184,In_725,In_1801);
or U185 (N_185,In_1294,In_1877);
nand U186 (N_186,In_571,In_2445);
xor U187 (N_187,In_117,In_178);
nor U188 (N_188,In_2331,In_1136);
xor U189 (N_189,In_2887,In_938);
xnor U190 (N_190,In_501,In_723);
xnor U191 (N_191,In_428,In_2402);
or U192 (N_192,In_1466,In_2507);
nand U193 (N_193,In_418,In_2385);
nand U194 (N_194,In_1030,In_2209);
or U195 (N_195,In_1550,In_902);
or U196 (N_196,In_2799,In_2604);
and U197 (N_197,In_372,In_1739);
and U198 (N_198,In_1180,In_1681);
nand U199 (N_199,In_2480,In_474);
and U200 (N_200,In_1819,In_2356);
nand U201 (N_201,In_2601,In_523);
or U202 (N_202,In_955,In_1883);
nand U203 (N_203,In_2408,In_665);
xnor U204 (N_204,In_2297,In_1601);
nand U205 (N_205,In_1482,In_1822);
nand U206 (N_206,In_183,In_359);
and U207 (N_207,In_2324,In_1549);
nand U208 (N_208,In_2087,In_1993);
nor U209 (N_209,In_2626,In_2012);
xor U210 (N_210,In_611,In_1285);
and U211 (N_211,In_1134,In_1414);
xor U212 (N_212,In_1712,In_1967);
xor U213 (N_213,In_314,In_2269);
or U214 (N_214,In_184,In_1421);
nor U215 (N_215,In_2492,In_1352);
nor U216 (N_216,In_1634,In_2173);
or U217 (N_217,In_590,In_500);
and U218 (N_218,In_2484,In_1114);
xor U219 (N_219,In_1236,In_80);
or U220 (N_220,In_1014,In_587);
nor U221 (N_221,In_60,In_1329);
or U222 (N_222,In_2271,In_950);
nand U223 (N_223,In_682,In_1229);
and U224 (N_224,In_2757,In_1905);
nor U225 (N_225,In_1502,In_2022);
and U226 (N_226,In_1138,In_754);
nor U227 (N_227,In_624,In_75);
nand U228 (N_228,In_1729,In_2030);
or U229 (N_229,In_285,In_1810);
nor U230 (N_230,In_39,In_1375);
and U231 (N_231,In_2990,In_1671);
nand U232 (N_232,In_2583,In_2650);
nand U233 (N_233,In_1382,In_1289);
nor U234 (N_234,In_1351,In_2871);
nor U235 (N_235,In_2893,In_1394);
and U236 (N_236,In_569,In_210);
nor U237 (N_237,In_2319,In_1940);
nor U238 (N_238,In_2145,In_1341);
nand U239 (N_239,In_2608,In_385);
and U240 (N_240,In_686,In_645);
nand U241 (N_241,In_1707,In_1528);
xnor U242 (N_242,In_1988,In_1979);
or U243 (N_243,In_715,In_1125);
or U244 (N_244,In_1820,In_2575);
nand U245 (N_245,In_1445,In_1800);
and U246 (N_246,In_1403,In_442);
or U247 (N_247,In_913,In_2134);
nor U248 (N_248,In_1321,In_2270);
or U249 (N_249,In_1183,In_2165);
and U250 (N_250,In_274,In_2072);
xnor U251 (N_251,In_1152,In_2007);
or U252 (N_252,In_2798,In_536);
nand U253 (N_253,In_1001,In_1812);
xnor U254 (N_254,In_702,In_2733);
and U255 (N_255,In_2894,In_2140);
nand U256 (N_256,In_154,In_213);
or U257 (N_257,In_2065,In_239);
xor U258 (N_258,In_2363,In_1338);
or U259 (N_259,In_2009,In_1959);
nor U260 (N_260,In_2059,In_354);
nand U261 (N_261,In_33,In_717);
nor U262 (N_262,In_2587,In_2109);
nor U263 (N_263,In_2616,In_1513);
or U264 (N_264,In_806,In_2882);
and U265 (N_265,In_1885,In_167);
xor U266 (N_266,In_1577,In_540);
xnor U267 (N_267,In_2995,In_252);
and U268 (N_268,In_2923,In_319);
nand U269 (N_269,In_2602,In_2531);
nor U270 (N_270,In_1872,In_2150);
nor U271 (N_271,In_2945,In_95);
or U272 (N_272,In_2752,In_244);
xor U273 (N_273,In_2008,In_2913);
and U274 (N_274,In_37,In_349);
nand U275 (N_275,In_746,In_1866);
nor U276 (N_276,In_1625,In_371);
xnor U277 (N_277,In_978,In_1911);
xnor U278 (N_278,In_1672,In_2183);
and U279 (N_279,In_647,In_1711);
nand U280 (N_280,In_79,In_127);
nand U281 (N_281,In_2104,In_2558);
and U282 (N_282,In_2867,In_0);
nand U283 (N_283,In_1735,In_986);
and U284 (N_284,In_2859,In_240);
or U285 (N_285,In_1948,In_559);
xor U286 (N_286,In_393,In_731);
xnor U287 (N_287,In_1304,In_898);
nand U288 (N_288,In_1019,In_1007);
or U289 (N_289,In_2663,In_972);
nor U290 (N_290,In_2665,In_884);
and U291 (N_291,In_1998,In_2838);
nor U292 (N_292,In_363,In_815);
nor U293 (N_293,In_2147,In_538);
nand U294 (N_294,In_164,In_515);
or U295 (N_295,In_2485,In_2332);
nor U296 (N_296,In_2815,In_2335);
xor U297 (N_297,In_1282,In_1368);
or U298 (N_298,In_2774,In_1721);
or U299 (N_299,In_577,In_2386);
nor U300 (N_300,In_2896,In_1936);
xnor U301 (N_301,In_2083,In_282);
xor U302 (N_302,In_1814,In_2103);
nor U303 (N_303,In_1011,In_2702);
nand U304 (N_304,In_235,In_1999);
xnor U305 (N_305,In_2337,In_1499);
nand U306 (N_306,In_565,In_755);
or U307 (N_307,In_2776,In_357);
or U308 (N_308,In_1761,In_2729);
nand U309 (N_309,In_2443,In_772);
nor U310 (N_310,In_1118,In_203);
and U311 (N_311,In_2196,In_1599);
or U312 (N_312,In_1617,In_2211);
nand U313 (N_313,In_1763,In_8);
nor U314 (N_314,In_2224,In_966);
nor U315 (N_315,In_518,In_201);
nor U316 (N_316,In_1568,In_1318);
or U317 (N_317,In_2187,In_1660);
nand U318 (N_318,In_1966,In_420);
and U319 (N_319,In_1272,In_1710);
or U320 (N_320,In_1750,In_2873);
xor U321 (N_321,In_662,In_26);
nand U322 (N_322,In_1344,In_1230);
nand U323 (N_323,In_2892,In_1946);
or U324 (N_324,In_2942,In_336);
nor U325 (N_325,In_51,In_2953);
and U326 (N_326,In_1664,In_1110);
nor U327 (N_327,In_2603,In_557);
nand U328 (N_328,In_18,In_2094);
xor U329 (N_329,In_2552,In_251);
nand U330 (N_330,In_1785,In_2641);
nand U331 (N_331,In_900,In_2170);
and U332 (N_332,In_277,In_2600);
nand U333 (N_333,In_2179,In_925);
nand U334 (N_334,In_1074,In_1543);
or U335 (N_335,In_875,In_1363);
nand U336 (N_336,In_671,In_654);
nor U337 (N_337,In_2557,In_2959);
nor U338 (N_338,In_1816,In_171);
nand U339 (N_339,In_1702,In_1504);
or U340 (N_340,In_1553,In_2823);
nand U341 (N_341,In_606,In_2878);
xnor U342 (N_342,In_78,In_103);
nand U343 (N_343,In_2161,In_894);
nor U344 (N_344,In_408,In_110);
nand U345 (N_345,In_975,In_1990);
nor U346 (N_346,In_603,In_1379);
or U347 (N_347,In_2691,In_1745);
nand U348 (N_348,In_2433,In_935);
and U349 (N_349,In_837,In_2759);
nor U350 (N_350,In_2352,In_2855);
and U351 (N_351,In_1532,In_1692);
and U352 (N_352,In_2724,In_2849);
or U353 (N_353,In_287,In_185);
and U354 (N_354,In_1124,In_1257);
nor U355 (N_355,In_275,In_328);
xor U356 (N_356,In_1298,In_2374);
or U357 (N_357,In_862,In_2763);
nand U358 (N_358,In_2441,In_1211);
and U359 (N_359,In_2019,In_1598);
xnor U360 (N_360,In_1025,In_2155);
or U361 (N_361,In_1258,In_853);
nand U362 (N_362,In_1371,In_984);
nor U363 (N_363,In_631,In_2407);
nor U364 (N_364,In_1068,In_927);
or U365 (N_365,In_2864,In_773);
and U366 (N_366,In_1593,In_1232);
xnor U367 (N_367,In_2571,In_1857);
nor U368 (N_368,In_1595,In_2537);
xnor U369 (N_369,In_1336,In_2929);
xor U370 (N_370,In_1526,In_600);
or U371 (N_371,In_946,In_2731);
or U372 (N_372,In_1396,In_1600);
xnor U373 (N_373,In_1427,In_1266);
or U374 (N_374,In_2023,In_2843);
and U375 (N_375,In_2761,In_1640);
xor U376 (N_376,In_784,In_629);
nor U377 (N_377,In_1644,In_1569);
xnor U378 (N_378,In_1410,In_294);
and U379 (N_379,In_2711,In_2223);
nor U380 (N_380,In_181,In_1373);
and U381 (N_381,In_2883,In_1808);
or U382 (N_382,In_2642,In_1402);
or U383 (N_383,In_1887,In_1985);
xnor U384 (N_384,In_1039,In_1687);
xor U385 (N_385,In_1505,In_827);
nor U386 (N_386,In_1043,In_1297);
nor U387 (N_387,In_2740,In_161);
xnor U388 (N_388,In_1997,In_316);
xnor U389 (N_389,In_721,In_2193);
nor U390 (N_390,In_194,In_1397);
or U391 (N_391,In_1903,In_2437);
xor U392 (N_392,In_455,In_1034);
nand U393 (N_393,In_338,In_2939);
xor U394 (N_394,In_253,In_1604);
or U395 (N_395,In_2156,In_2976);
nor U396 (N_396,In_1415,In_1462);
or U397 (N_397,In_696,In_104);
nor U398 (N_398,In_695,In_1722);
and U399 (N_399,In_2862,In_2452);
or U400 (N_400,In_2471,In_416);
or U401 (N_401,In_2753,In_2438);
nor U402 (N_402,In_1349,In_1035);
or U403 (N_403,In_1189,In_1576);
and U404 (N_404,In_2305,In_537);
nand U405 (N_405,In_1770,In_150);
and U406 (N_406,In_512,In_2474);
nor U407 (N_407,In_2858,In_1078);
and U408 (N_408,In_2384,In_2950);
and U409 (N_409,In_528,In_2213);
and U410 (N_410,In_2144,In_2830);
and U411 (N_411,In_594,In_1131);
xnor U412 (N_412,In_722,In_1970);
nand U413 (N_413,In_2148,In_337);
nand U414 (N_414,In_998,In_1833);
or U415 (N_415,In_2473,In_2525);
nor U416 (N_416,In_2501,In_1483);
nor U417 (N_417,In_1117,In_2536);
nor U418 (N_418,In_2077,In_1377);
and U419 (N_419,In_2522,In_92);
and U420 (N_420,In_2886,In_792);
and U421 (N_421,In_965,In_566);
or U422 (N_422,In_1216,In_196);
xnor U423 (N_423,In_31,In_1983);
nand U424 (N_424,In_1381,In_38);
or U425 (N_425,In_1973,In_2820);
nor U426 (N_426,In_1616,In_2365);
and U427 (N_427,In_1992,In_257);
and U428 (N_428,In_2258,In_1835);
or U429 (N_429,In_96,In_1503);
xor U430 (N_430,In_1652,In_570);
or U431 (N_431,In_760,In_2760);
or U432 (N_432,In_2162,In_358);
nor U433 (N_433,In_1147,In_1020);
nor U434 (N_434,In_1701,In_1900);
nand U435 (N_435,In_368,In_2645);
xnor U436 (N_436,In_1837,In_2351);
and U437 (N_437,In_2965,In_1732);
nor U438 (N_438,In_737,In_1939);
nand U439 (N_439,In_623,In_2315);
nor U440 (N_440,In_241,In_2056);
and U441 (N_441,In_2649,In_1071);
nand U442 (N_442,In_36,In_2227);
xor U443 (N_443,In_1706,In_1174);
xor U444 (N_444,In_811,In_698);
nor U445 (N_445,In_2817,In_1425);
and U446 (N_446,In_2212,In_2590);
nor U447 (N_447,In_2902,In_238);
and U448 (N_448,In_339,In_593);
or U449 (N_449,In_2787,In_295);
or U450 (N_450,In_2679,In_1442);
and U451 (N_451,In_487,In_2450);
or U452 (N_452,In_2635,In_595);
xor U453 (N_453,In_633,In_937);
nor U454 (N_454,In_813,In_2837);
nand U455 (N_455,In_1292,In_816);
or U456 (N_456,In_1079,In_787);
and U457 (N_457,In_2282,In_1531);
nor U458 (N_458,In_1752,In_2964);
nand U459 (N_459,In_2826,In_2508);
nor U460 (N_460,In_669,In_302);
or U461 (N_461,In_2014,In_2758);
and U462 (N_462,In_1251,In_1220);
and U463 (N_463,In_1933,In_1570);
and U464 (N_464,In_1838,In_602);
and U465 (N_465,In_673,In_2159);
xor U466 (N_466,In_1264,In_2002);
or U467 (N_467,In_844,In_1278);
nand U468 (N_468,In_77,In_1535);
nor U469 (N_469,In_1175,In_872);
and U470 (N_470,In_2669,In_848);
and U471 (N_471,In_2749,In_1865);
and U472 (N_472,In_1263,In_640);
and U473 (N_473,In_574,In_198);
and U474 (N_474,In_2510,In_2771);
nand U475 (N_475,In_2701,In_2722);
and U476 (N_476,In_40,In_882);
nand U477 (N_477,In_2035,In_254);
nand U478 (N_478,In_1085,In_1097);
and U479 (N_479,In_1121,In_470);
and U480 (N_480,In_2251,In_1917);
or U481 (N_481,In_903,In_367);
or U482 (N_482,In_2982,In_2475);
or U483 (N_483,In_322,In_2736);
nand U484 (N_484,In_422,In_1406);
and U485 (N_485,In_182,In_2366);
nand U486 (N_486,In_1476,In_1555);
xor U487 (N_487,In_2339,In_763);
and U488 (N_488,In_1827,In_222);
nand U489 (N_489,In_1157,In_2080);
or U490 (N_490,In_907,In_1771);
nand U491 (N_491,In_2052,In_1858);
or U492 (N_492,In_2581,In_2998);
or U493 (N_493,In_2076,In_1485);
nor U494 (N_494,In_1194,In_1498);
nand U495 (N_495,In_2095,In_2130);
nor U496 (N_496,In_304,In_2232);
nor U497 (N_497,In_1728,In_627);
and U498 (N_498,In_1886,In_1957);
or U499 (N_499,In_2206,In_1162);
and U500 (N_500,In_2739,In_2908);
and U501 (N_501,In_909,N_146);
nand U502 (N_502,In_953,In_1026);
xnor U503 (N_503,In_2131,In_55);
and U504 (N_504,In_2545,In_1395);
and U505 (N_505,In_2127,In_1405);
xor U506 (N_506,In_2413,In_105);
xnor U507 (N_507,N_92,In_148);
xnor U508 (N_508,In_1095,In_854);
nor U509 (N_509,N_449,In_28);
xor U510 (N_510,In_1053,N_485);
or U511 (N_511,In_2241,In_1488);
and U512 (N_512,N_217,In_2951);
nand U513 (N_513,In_176,In_2856);
xnor U514 (N_514,In_2152,In_2948);
nand U515 (N_515,In_928,N_367);
or U516 (N_516,In_799,In_1717);
nor U517 (N_517,N_371,In_1447);
and U518 (N_518,N_38,In_2721);
or U519 (N_519,In_195,N_200);
or U520 (N_520,In_2276,N_442);
xor U521 (N_521,In_637,In_1391);
nor U522 (N_522,In_1449,In_2543);
and U523 (N_523,In_2426,N_175);
and U524 (N_524,In_1383,In_1537);
nand U525 (N_525,In_863,In_2672);
nand U526 (N_526,In_2325,In_1953);
or U527 (N_527,In_2198,N_170);
and U528 (N_528,In_243,N_345);
xor U529 (N_529,In_2349,In_2852);
nand U530 (N_530,In_838,In_146);
nand U531 (N_531,In_228,In_2143);
and U532 (N_532,In_2833,N_431);
nand U533 (N_533,In_1359,N_77);
or U534 (N_534,In_876,N_45);
or U535 (N_535,In_140,In_388);
xnor U536 (N_536,In_2265,N_347);
xnor U537 (N_537,In_2520,In_2559);
and U538 (N_538,In_697,N_34);
nor U539 (N_539,In_2102,N_372);
or U540 (N_540,In_2361,In_1780);
nor U541 (N_541,In_2024,N_324);
nor U542 (N_542,N_103,N_86);
or U543 (N_543,N_102,In_425);
xnor U544 (N_544,N_247,In_1310);
xor U545 (N_545,In_2454,In_1791);
nor U546 (N_546,In_2903,N_340);
or U547 (N_547,In_1805,In_471);
nor U548 (N_548,In_904,In_2516);
or U549 (N_549,In_144,In_424);
or U550 (N_550,N_409,In_153);
nor U551 (N_551,In_989,In_1051);
nand U552 (N_552,In_296,In_2811);
nand U553 (N_553,In_680,In_1303);
nand U554 (N_554,In_1386,In_138);
and U555 (N_555,In_2534,N_254);
or U556 (N_556,In_719,In_793);
nand U557 (N_557,In_2659,In_1208);
and U558 (N_558,In_2720,In_1314);
and U559 (N_559,In_1629,In_1842);
and U560 (N_560,N_139,In_2949);
xor U561 (N_561,In_2818,In_469);
xnor U562 (N_562,N_98,In_1126);
and U563 (N_563,In_1922,In_801);
and U564 (N_564,In_864,In_2394);
xnor U565 (N_565,N_389,In_775);
and U566 (N_566,In_263,N_135);
or U567 (N_567,In_1704,In_123);
nand U568 (N_568,In_50,In_2425);
nor U569 (N_569,N_197,In_1109);
nand U570 (N_570,In_2136,N_313);
and U571 (N_571,In_1002,In_1165);
nand U572 (N_572,N_395,In_1849);
or U573 (N_573,N_157,In_2747);
xor U574 (N_574,In_2750,In_642);
or U575 (N_575,In_1319,N_422);
nor U576 (N_576,N_180,In_407);
or U577 (N_577,In_2792,In_797);
and U578 (N_578,In_366,In_352);
nand U579 (N_579,N_8,In_169);
and U580 (N_580,In_1099,In_2926);
xnor U581 (N_581,N_329,In_1952);
nor U582 (N_582,In_1668,In_2299);
nand U583 (N_583,N_427,In_962);
and U584 (N_584,In_2544,In_932);
or U585 (N_585,N_472,In_2113);
and U586 (N_586,In_2214,In_227);
or U587 (N_587,In_1374,In_794);
nor U588 (N_588,In_1904,N_32);
nand U589 (N_589,In_897,N_430);
or U590 (N_590,In_2132,In_2066);
and U591 (N_591,In_2909,In_2383);
xnor U592 (N_592,In_2638,In_2810);
and U593 (N_593,In_956,In_1221);
nand U594 (N_594,In_747,In_1901);
nand U595 (N_595,In_1094,In_2597);
and U596 (N_596,N_408,In_1517);
and U597 (N_597,In_1202,N_296);
or U598 (N_598,In_289,In_2001);
and U599 (N_599,In_1070,In_361);
and U600 (N_600,N_292,In_976);
nor U601 (N_601,In_1225,In_290);
nand U602 (N_602,In_850,N_250);
and U603 (N_603,In_2081,In_2775);
or U604 (N_604,In_891,N_252);
or U605 (N_605,In_703,In_1591);
nand U606 (N_606,In_1137,In_2096);
nor U607 (N_607,In_2490,In_2164);
and U608 (N_608,In_618,In_1902);
nor U609 (N_609,N_365,In_1365);
xor U610 (N_610,In_1176,N_234);
or U611 (N_611,In_1867,In_2250);
or U612 (N_612,In_922,N_482);
nor U613 (N_613,N_11,In_72);
nor U614 (N_614,N_223,In_589);
and U615 (N_615,In_1302,In_1561);
or U616 (N_616,In_1510,In_20);
or U617 (N_617,In_778,In_1267);
nor U618 (N_618,In_2655,In_68);
nor U619 (N_619,In_2218,N_244);
nor U620 (N_620,In_233,In_2944);
xnor U621 (N_621,In_920,In_1860);
nand U622 (N_622,N_407,In_2489);
xnor U623 (N_623,In_802,N_18);
or U624 (N_624,In_2458,N_233);
xor U625 (N_625,In_1200,N_95);
and U626 (N_626,In_2819,In_1977);
and U627 (N_627,In_324,In_579);
xnor U628 (N_628,In_2988,In_1305);
and U629 (N_629,In_1521,N_266);
or U630 (N_630,N_46,N_67);
and U631 (N_631,N_448,In_1684);
or U632 (N_632,In_1056,In_2743);
nor U633 (N_633,N_460,In_1870);
nand U634 (N_634,In_899,In_2178);
nand U635 (N_635,In_1935,In_2368);
xor U636 (N_636,In_514,In_2230);
nand U637 (N_637,N_83,In_1385);
nand U638 (N_638,In_496,In_683);
or U639 (N_639,In_2399,In_299);
or U640 (N_640,In_187,In_406);
nor U641 (N_641,In_2322,In_2421);
and U642 (N_642,In_2075,In_1163);
nand U643 (N_643,N_391,N_113);
nor U644 (N_644,In_2067,In_2046);
or U645 (N_645,In_6,N_274);
nand U646 (N_646,In_258,In_2681);
xor U647 (N_647,In_1203,In_1045);
nor U648 (N_648,In_1367,N_414);
and U649 (N_649,In_2345,In_1506);
or U650 (N_650,In_1863,In_597);
xnor U651 (N_651,In_2139,In_1065);
nor U652 (N_652,In_1758,N_253);
xnor U653 (N_653,In_591,In_1965);
and U654 (N_654,In_2118,In_710);
xnor U655 (N_655,N_309,In_2362);
nand U656 (N_656,In_1777,In_2713);
nand U657 (N_657,In_1423,In_2956);
or U658 (N_658,N_457,In_2416);
or U659 (N_659,In_2754,In_1743);
nor U660 (N_660,In_2115,In_1300);
and U661 (N_661,In_1622,In_2698);
and U662 (N_662,In_636,In_1912);
xor U663 (N_663,In_868,In_1441);
nor U664 (N_664,In_87,In_1811);
nor U665 (N_665,In_2040,N_71);
xnor U666 (N_666,In_1450,In_493);
nand U667 (N_667,In_1734,In_1187);
and U668 (N_668,In_729,In_2016);
and U669 (N_669,In_2053,In_162);
or U670 (N_670,In_1128,In_1690);
nor U671 (N_671,In_1299,In_849);
or U672 (N_672,In_507,In_829);
nor U673 (N_673,In_1420,In_1725);
nand U674 (N_674,N_14,In_1665);
and U675 (N_675,In_916,In_386);
and U676 (N_676,In_122,In_2827);
nor U677 (N_677,In_2415,In_1547);
nand U678 (N_678,In_658,In_246);
xnor U679 (N_679,In_2045,N_271);
nor U680 (N_680,N_301,In_1915);
nor U681 (N_681,In_1641,In_1850);
nand U682 (N_682,In_1283,In_1448);
and U683 (N_683,N_127,In_11);
or U684 (N_684,N_129,In_580);
and U685 (N_685,In_48,In_2567);
nand U686 (N_686,In_326,N_215);
nor U687 (N_687,In_1086,In_1340);
xnor U688 (N_688,In_1038,In_1270);
nand U689 (N_689,In_969,In_681);
nand U690 (N_690,In_170,In_315);
nand U691 (N_691,N_28,In_646);
xnor U692 (N_692,In_866,In_73);
and U693 (N_693,N_47,In_399);
and U694 (N_694,In_1491,N_191);
nor U695 (N_695,In_2451,In_1135);
nand U696 (N_696,In_1309,In_529);
nor U697 (N_697,In_1518,In_1115);
and U698 (N_698,In_2172,In_115);
and U699 (N_699,In_1328,In_2495);
or U700 (N_700,In_2106,In_2011);
nor U701 (N_701,In_2680,In_2851);
or U702 (N_702,In_1342,In_739);
and U703 (N_703,In_193,In_1726);
nand U704 (N_704,In_2521,N_193);
nor U705 (N_705,N_177,N_419);
and U706 (N_706,In_2796,N_231);
or U707 (N_707,In_2654,In_841);
nand U708 (N_708,In_563,In_2308);
and U709 (N_709,In_2013,In_2277);
and U710 (N_710,In_151,In_2797);
and U711 (N_711,In_2676,In_199);
nor U712 (N_712,In_1262,In_2303);
xnor U713 (N_713,In_2595,N_286);
xnor U714 (N_714,In_1227,In_2631);
nor U715 (N_715,In_220,In_1797);
nor U716 (N_716,In_1960,In_1755);
nand U717 (N_717,In_94,In_1345);
nor U718 (N_718,In_2993,In_132);
xnor U719 (N_719,N_394,In_2273);
nor U720 (N_720,In_98,In_762);
xor U721 (N_721,N_9,N_474);
or U722 (N_722,In_1047,N_190);
nand U723 (N_723,In_1996,N_285);
and U724 (N_724,In_27,In_2300);
or U725 (N_725,N_318,In_2528);
xor U726 (N_726,N_425,In_1235);
xnor U727 (N_727,N_93,In_1909);
xnor U728 (N_728,N_3,In_2824);
nor U729 (N_729,N_241,In_809);
nand U730 (N_730,N_126,In_2392);
or U731 (N_731,N_91,In_1238);
nor U732 (N_732,In_2329,In_2667);
nor U733 (N_733,N_325,In_1890);
or U734 (N_734,In_329,In_2404);
or U735 (N_735,In_10,In_1493);
nand U736 (N_736,In_1714,In_605);
or U737 (N_737,N_349,In_46);
or U738 (N_738,In_2555,In_2084);
nand U739 (N_739,In_1247,In_439);
nor U740 (N_740,In_2318,In_2429);
nand U741 (N_741,In_741,N_5);
xnor U742 (N_742,In_2825,In_632);
and U743 (N_743,In_108,In_1619);
nor U744 (N_744,In_666,In_2431);
nand U745 (N_745,In_2295,In_774);
xnor U746 (N_746,In_889,In_1751);
xnor U747 (N_747,In_276,In_318);
or U748 (N_748,In_2607,N_147);
or U749 (N_749,In_2194,In_1320);
and U750 (N_750,In_2333,N_240);
nand U751 (N_751,In_2259,In_1624);
nor U752 (N_752,In_14,N_263);
nand U753 (N_753,N_436,N_258);
and U754 (N_754,N_218,In_309);
or U755 (N_755,In_2462,In_785);
nor U756 (N_756,In_1571,In_288);
nor U757 (N_757,In_1607,In_1463);
or U758 (N_758,In_477,In_2313);
or U759 (N_759,In_1759,In_1525);
and U760 (N_760,In_2068,In_634);
and U761 (N_761,N_196,In_1150);
or U762 (N_762,In_2704,In_1829);
nor U763 (N_763,N_12,In_822);
nand U764 (N_764,In_798,In_2237);
nor U765 (N_765,In_2306,In_2866);
and U766 (N_766,In_1050,In_2904);
or U767 (N_767,In_12,In_1778);
and U768 (N_768,In_1818,In_1458);
nor U769 (N_769,In_1694,N_403);
nand U770 (N_770,In_2261,In_1206);
xnor U771 (N_771,In_2794,In_779);
nand U772 (N_772,N_384,In_483);
nand U773 (N_773,In_2707,In_1470);
nor U774 (N_774,In_1245,N_276);
nor U775 (N_775,In_1122,N_165);
nor U776 (N_776,In_1390,N_475);
nor U777 (N_777,In_2062,N_61);
nand U778 (N_778,In_307,In_699);
nand U779 (N_779,In_1197,In_957);
xor U780 (N_780,In_1930,N_51);
xnor U781 (N_781,In_2205,In_1609);
and U782 (N_782,In_2005,In_431);
and U783 (N_783,In_748,In_2376);
xnor U784 (N_784,In_1454,In_1501);
or U785 (N_785,In_1132,In_1633);
xnor U786 (N_786,In_1171,N_115);
or U787 (N_787,In_2509,N_80);
xnor U788 (N_788,In_2301,In_175);
nor U789 (N_789,In_1316,N_17);
and U790 (N_790,In_2656,In_1558);
xnor U791 (N_791,In_2456,N_13);
nor U792 (N_792,In_1713,N_65);
or U793 (N_793,In_156,N_357);
nor U794 (N_794,In_2640,N_388);
xnor U795 (N_795,In_2184,In_1104);
nand U796 (N_796,In_2560,N_62);
and U797 (N_797,N_306,N_462);
or U798 (N_798,In_360,In_1339);
and U799 (N_799,In_1416,In_2946);
xnor U800 (N_800,In_1004,In_2200);
nand U801 (N_801,In_22,In_2279);
nand U802 (N_802,In_2380,In_1796);
nand U803 (N_803,In_2453,In_1884);
and U804 (N_804,In_2682,In_2488);
or U805 (N_805,In_734,In_2574);
nand U806 (N_806,In_586,In_2684);
nand U807 (N_807,In_2414,In_1944);
nor U808 (N_808,In_209,In_588);
and U809 (N_809,In_533,In_2872);
or U810 (N_810,In_803,In_2524);
nand U811 (N_811,In_467,In_383);
nand U812 (N_812,In_858,In_2809);
xor U813 (N_813,In_56,In_947);
nand U814 (N_814,In_179,In_1874);
xnor U815 (N_815,In_941,N_387);
nand U816 (N_816,N_468,In_1347);
xnor U817 (N_817,N_24,In_1009);
or U818 (N_818,In_556,In_5);
nand U819 (N_819,N_312,In_226);
or U820 (N_820,In_1685,In_564);
nor U821 (N_821,In_948,In_1961);
nand U822 (N_822,In_818,In_273);
and U823 (N_823,In_1974,In_362);
xnor U824 (N_824,In_582,In_674);
nand U825 (N_825,In_85,In_1775);
and U826 (N_826,In_1467,N_162);
nand U827 (N_827,In_2290,N_308);
and U828 (N_828,N_239,In_1478);
nand U829 (N_829,In_1067,In_598);
nand U830 (N_830,In_652,N_235);
and U831 (N_831,In_2690,In_2292);
nand U832 (N_832,In_2513,In_230);
and U833 (N_833,In_1366,In_817);
nand U834 (N_834,In_2585,In_1156);
xor U835 (N_835,In_2889,N_150);
xnor U836 (N_836,In_1795,In_2189);
and U837 (N_837,In_2031,In_190);
or U838 (N_838,N_21,N_156);
and U839 (N_839,In_1637,In_2033);
and U840 (N_840,In_1480,In_1715);
nand U841 (N_841,N_189,In_1716);
xnor U842 (N_842,In_687,In_212);
nor U843 (N_843,In_2221,In_1130);
nor U844 (N_844,In_1399,In_2633);
or U845 (N_845,N_154,In_1891);
xor U846 (N_846,In_2915,In_1871);
and U847 (N_847,N_376,In_1815);
nor U848 (N_848,N_176,N_257);
nand U849 (N_849,In_2079,In_2943);
nor U850 (N_850,In_2021,In_2364);
and U851 (N_851,In_441,In_57);
or U852 (N_852,N_495,In_395);
and U853 (N_853,In_2785,N_278);
and U854 (N_854,In_2541,In_49);
or U855 (N_855,In_869,N_142);
and U856 (N_856,In_615,N_264);
xor U857 (N_857,N_443,In_415);
nor U858 (N_858,In_2952,In_343);
or U859 (N_859,In_685,In_465);
or U860 (N_860,In_320,In_1789);
and U861 (N_861,N_237,In_71);
nor U862 (N_862,In_2564,In_255);
or U863 (N_863,In_482,In_2039);
xor U864 (N_864,N_305,In_1971);
and U865 (N_865,In_2069,In_1618);
and U866 (N_866,N_121,N_49);
or U867 (N_867,In_2216,N_72);
xnor U868 (N_868,N_320,In_1731);
nand U869 (N_869,In_610,In_1586);
and U870 (N_870,In_1494,In_1170);
and U871 (N_871,In_906,In_1451);
or U872 (N_872,In_1358,In_2353);
or U873 (N_873,In_2784,In_1093);
nor U874 (N_874,In_1369,In_2715);
xor U875 (N_875,In_851,In_2176);
and U876 (N_876,N_109,In_1411);
and U877 (N_877,In_541,In_2125);
and U878 (N_878,In_2907,In_1627);
nand U879 (N_879,N_496,In_807);
xor U880 (N_880,N_52,In_1994);
xor U881 (N_881,In_2098,In_758);
or U882 (N_882,In_1741,In_2238);
xnor U883 (N_883,In_1195,In_832);
and U884 (N_884,In_2093,In_2419);
nand U885 (N_885,In_651,In_1956);
xor U886 (N_886,N_298,In_214);
or U887 (N_887,In_2286,In_1783);
xor U888 (N_888,In_2427,In_1559);
nor U889 (N_889,In_2912,In_2038);
or U890 (N_890,In_373,In_2449);
nor U891 (N_891,In_527,In_321);
nand U892 (N_892,N_280,In_2502);
xor U893 (N_893,In_2624,In_2795);
nand U894 (N_894,In_2048,In_271);
nor U895 (N_895,In_2377,In_1688);
nand U896 (N_896,In_1223,N_352);
nand U897 (N_897,N_284,In_2596);
nand U898 (N_898,In_936,In_1024);
nand U899 (N_899,N_437,In_1899);
nand U900 (N_900,In_2628,In_1412);
xor U901 (N_901,In_2358,N_369);
xor U902 (N_902,N_440,In_2569);
nor U903 (N_903,In_286,In_657);
and U904 (N_904,N_364,In_2341);
and U905 (N_905,In_2342,In_2291);
or U906 (N_906,In_592,In_981);
nor U907 (N_907,In_301,N_2);
nor U908 (N_908,In_1519,N_134);
or U909 (N_909,In_2839,In_1679);
nand U910 (N_910,In_1191,In_2124);
and U911 (N_911,In_2991,In_2816);
nand U912 (N_912,N_128,In_914);
xnor U913 (N_913,N_361,N_397);
nand U914 (N_914,In_303,N_455);
xnor U915 (N_915,In_100,In_810);
xnor U916 (N_916,N_141,In_828);
or U917 (N_917,In_2664,In_333);
and U918 (N_918,In_1044,In_1921);
nand U919 (N_919,N_315,N_294);
xnor U920 (N_920,In_2137,In_2523);
nand U921 (N_921,In_551,In_505);
nand U922 (N_922,In_1955,In_2070);
nor U923 (N_923,In_508,In_2469);
nor U924 (N_924,In_1106,In_2190);
nand U925 (N_925,In_1653,In_1249);
nor U926 (N_926,In_873,In_1037);
nor U927 (N_927,In_782,In_466);
nor U928 (N_928,In_1594,In_1991);
or U929 (N_929,In_888,In_1834);
or U930 (N_930,In_23,In_1651);
and U931 (N_931,In_2611,In_2683);
or U932 (N_932,In_3,In_2111);
nor U933 (N_933,In_584,In_1705);
nand U934 (N_934,In_128,In_1219);
nor U935 (N_935,N_433,In_2228);
or U936 (N_936,In_630,N_188);
nor U937 (N_937,N_63,In_2692);
nand U938 (N_938,In_2788,N_158);
and U939 (N_939,In_453,N_316);
xnor U940 (N_940,In_1512,In_387);
and U941 (N_941,In_2845,N_159);
xnor U942 (N_942,In_1330,In_628);
nor U943 (N_943,In_1964,In_1185);
and U944 (N_944,N_317,In_1782);
and U945 (N_945,In_1256,In_2688);
nor U946 (N_946,In_1333,In_2773);
nand U947 (N_947,In_1167,In_1573);
nand U948 (N_948,In_924,N_351);
nor U949 (N_949,In_2737,N_383);
and U950 (N_950,In_2247,In_200);
nor U951 (N_951,N_89,In_1821);
or U952 (N_952,In_693,In_910);
nor U953 (N_953,N_94,N_69);
and U954 (N_954,In_1682,N_195);
and U955 (N_955,In_1605,N_155);
xor U956 (N_956,In_2781,In_19);
xnor U957 (N_957,In_1578,N_463);
nor U958 (N_958,In_1516,In_1923);
nand U959 (N_959,In_1188,In_2802);
nand U960 (N_960,In_929,In_2968);
or U961 (N_961,In_1052,N_444);
nand U962 (N_962,In_2910,In_1932);
xnor U963 (N_963,In_2226,In_1643);
or U964 (N_964,In_1087,N_255);
nand U965 (N_965,N_205,In_2321);
xor U966 (N_966,In_562,In_2071);
or U967 (N_967,N_392,In_1475);
and U968 (N_968,In_1693,In_619);
nand U969 (N_969,In_2639,In_2614);
xnor U970 (N_970,In_2278,In_1906);
nand U971 (N_971,In_1648,N_123);
and U972 (N_972,N_262,In_1813);
or U973 (N_973,In_447,In_2609);
nand U974 (N_974,In_2085,In_2847);
or U975 (N_975,In_1580,In_2129);
nor U976 (N_976,In_771,In_2411);
nand U977 (N_977,In_776,N_227);
or U978 (N_978,In_2027,In_1083);
xor U979 (N_979,In_1049,In_1841);
or U980 (N_980,N_230,In_32);
xnor U981 (N_981,In_552,In_34);
xnor U982 (N_982,In_2505,N_379);
or U983 (N_983,In_444,In_2086);
xor U984 (N_984,In_555,In_1276);
and U985 (N_985,In_2705,In_1215);
nand U986 (N_986,N_118,In_2778);
xor U987 (N_987,In_141,In_2180);
nor U988 (N_988,In_599,In_795);
and U989 (N_989,In_177,In_1102);
nand U990 (N_990,In_2418,In_757);
xnor U991 (N_991,In_2126,In_2922);
nor U992 (N_992,In_2182,In_1676);
xnor U993 (N_993,N_54,In_1306);
nor U994 (N_994,In_887,In_2463);
nand U995 (N_995,In_2343,N_178);
xnor U996 (N_996,In_202,In_2010);
xnor U997 (N_997,In_495,N_402);
nand U998 (N_998,N_76,In_575);
xor U999 (N_999,In_218,In_2963);
or U1000 (N_1000,N_533,In_2186);
nor U1001 (N_1001,N_642,In_1924);
and U1002 (N_1002,In_714,In_461);
or U1003 (N_1003,In_430,In_959);
nand U1004 (N_1004,N_684,In_1878);
nor U1005 (N_1005,N_366,In_2899);
nor U1006 (N_1006,In_988,N_466);
xnor U1007 (N_1007,N_728,N_657);
and U1008 (N_1008,In_1497,N_591);
nor U1009 (N_1009,N_339,N_385);
nand U1010 (N_1010,In_2442,In_2632);
and U1011 (N_1011,In_2231,In_1088);
or U1012 (N_1012,In_1772,In_394);
nor U1013 (N_1013,In_2357,N_497);
xor U1014 (N_1014,N_268,N_766);
nand U1015 (N_1015,In_62,In_1190);
nand U1016 (N_1016,In_2791,N_473);
or U1017 (N_1017,In_186,N_57);
xor U1018 (N_1018,N_668,In_617);
and U1019 (N_1019,N_779,In_2428);
nand U1020 (N_1020,In_1546,In_2550);
nand U1021 (N_1021,N_58,In_375);
and U1022 (N_1022,In_967,N_936);
nor U1023 (N_1023,N_882,N_256);
nand U1024 (N_1024,In_1733,In_820);
nand U1025 (N_1025,In_1552,In_2789);
nor U1026 (N_1026,In_2973,N_981);
or U1027 (N_1027,In_915,N_512);
xor U1028 (N_1028,In_1059,N_680);
nand U1029 (N_1029,N_943,In_2446);
xor U1030 (N_1030,In_2123,In_1666);
nor U1031 (N_1031,In_2255,N_878);
xnor U1032 (N_1032,In_893,N_222);
xor U1033 (N_1033,In_1703,N_906);
nor U1034 (N_1034,N_894,N_15);
and U1035 (N_1035,In_1112,N_692);
xnor U1036 (N_1036,In_1802,In_1226);
nand U1037 (N_1037,N_22,In_1947);
nand U1038 (N_1038,In_2777,N_140);
xnor U1039 (N_1039,N_601,In_1742);
or U1040 (N_1040,N_166,In_2378);
nor U1041 (N_1041,In_1484,In_1937);
nor U1042 (N_1042,N_715,In_643);
xnor U1043 (N_1043,N_921,N_64);
nand U1044 (N_1044,N_413,In_306);
xor U1045 (N_1045,In_2984,In_2476);
nor U1046 (N_1046,N_506,N_808);
xnor U1047 (N_1047,N_933,N_173);
nor U1048 (N_1048,N_82,In_2756);
and U1049 (N_1049,In_732,In_1040);
and U1050 (N_1050,In_1620,N_543);
nand U1051 (N_1051,N_360,In_2916);
and U1052 (N_1052,N_830,N_70);
nand U1053 (N_1053,In_2397,In_944);
nand U1054 (N_1054,N_265,N_210);
and U1055 (N_1055,N_641,In_102);
nor U1056 (N_1056,In_211,N_838);
or U1057 (N_1057,N_108,N_880);
nor U1058 (N_1058,In_2769,In_2105);
or U1059 (N_1059,In_1265,In_1907);
and U1060 (N_1060,N_125,In_434);
nor U1061 (N_1061,N_521,N_941);
xnor U1062 (N_1062,In_1127,In_2006);
nor U1063 (N_1063,N_956,In_2051);
or U1064 (N_1064,In_2622,In_1845);
and U1065 (N_1065,In_1111,In_1422);
and U1066 (N_1066,In_2153,In_2548);
nand U1067 (N_1067,In_1781,In_2389);
nor U1068 (N_1068,In_488,In_1680);
or U1069 (N_1069,N_800,In_2577);
nor U1070 (N_1070,In_659,In_1455);
or U1071 (N_1071,In_353,N_967);
xor U1072 (N_1072,N_675,In_111);
and U1073 (N_1073,In_2401,In_847);
xor U1074 (N_1074,N_337,In_1536);
nor U1075 (N_1075,N_221,N_901);
xnor U1076 (N_1076,In_1116,In_2677);
or U1077 (N_1077,In_675,In_478);
and U1078 (N_1078,N_525,In_1362);
nor U1079 (N_1079,In_2879,In_2512);
nand U1080 (N_1080,In_1927,N_214);
or U1081 (N_1081,N_970,N_622);
nor U1082 (N_1082,In_2479,In_485);
nand U1083 (N_1083,In_2549,In_2741);
and U1084 (N_1084,In_1667,In_1417);
nand U1085 (N_1085,In_310,In_2897);
or U1086 (N_1086,In_2225,In_443);
nor U1087 (N_1087,N_832,In_612);
nor U1088 (N_1088,In_2992,N_480);
or U1089 (N_1089,N_23,In_409);
and U1090 (N_1090,In_1548,N_760);
xor U1091 (N_1091,N_580,In_522);
nor U1092 (N_1092,N_922,N_975);
or U1093 (N_1093,N_534,N_929);
or U1094 (N_1094,N_398,In_401);
nand U1095 (N_1095,In_2050,N_321);
nor U1096 (N_1096,N_354,In_2444);
nor U1097 (N_1097,N_640,In_2160);
and U1098 (N_1098,In_2911,In_2185);
and U1099 (N_1099,N_749,In_2304);
nand U1100 (N_1100,N_209,In_688);
nand U1101 (N_1101,In_691,N_711);
or U1102 (N_1102,N_559,N_412);
and U1103 (N_1103,In_1557,In_1312);
nand U1104 (N_1104,N_513,In_346);
nand U1105 (N_1105,N_723,In_445);
and U1106 (N_1106,N_979,N_652);
or U1107 (N_1107,In_1479,N_647);
or U1108 (N_1108,In_796,In_463);
or U1109 (N_1109,In_2996,In_1597);
xnor U1110 (N_1110,N_910,In_1567);
xor U1111 (N_1111,In_2805,In_2770);
xnor U1112 (N_1112,N_202,N_691);
or U1113 (N_1113,N_116,In_788);
or U1114 (N_1114,N_476,N_461);
and U1115 (N_1115,In_1436,N_467);
xor U1116 (N_1116,In_1847,In_1790);
xnor U1117 (N_1117,N_839,In_1169);
and U1118 (N_1118,In_1184,In_221);
xor U1119 (N_1119,N_927,In_491);
nor U1120 (N_1120,In_2393,In_1139);
or U1121 (N_1121,N_713,In_1443);
or U1122 (N_1122,In_2539,In_2340);
and U1123 (N_1123,N_721,N_955);
xnor U1124 (N_1124,N_996,N_374);
nand U1125 (N_1125,In_705,In_2861);
nand U1126 (N_1126,In_429,In_2334);
and U1127 (N_1127,N_619,N_386);
xor U1128 (N_1128,In_2107,In_1241);
xor U1129 (N_1129,N_768,In_17);
or U1130 (N_1130,N_544,N_549);
nor U1131 (N_1131,In_964,In_1831);
nand U1132 (N_1132,In_2966,In_1581);
or U1133 (N_1133,In_435,N_947);
and U1134 (N_1134,In_1433,In_2617);
or U1135 (N_1135,N_722,N_560);
and U1136 (N_1136,N_406,N_500);
nand U1137 (N_1137,N_751,N_332);
nand U1138 (N_1138,In_2762,N_584);
nand U1139 (N_1139,N_434,N_624);
or U1140 (N_1140,In_1196,In_412);
or U1141 (N_1141,N_514,N_605);
nor U1142 (N_1142,N_323,In_312);
or U1143 (N_1143,In_1098,In_535);
and U1144 (N_1144,N_269,N_208);
or U1145 (N_1145,N_849,N_702);
nand U1146 (N_1146,N_1,N_892);
nand U1147 (N_1147,In_767,In_2687);
nor U1148 (N_1148,N_629,N_259);
xnor U1149 (N_1149,In_2236,In_1261);
or U1150 (N_1150,N_952,N_338);
nand U1151 (N_1151,N_863,In_2935);
and U1152 (N_1152,In_578,N_579);
or U1153 (N_1153,In_1582,In_2844);
or U1154 (N_1154,In_2396,In_1307);
nand U1155 (N_1155,N_267,N_644);
xnor U1156 (N_1156,N_548,In_204);
and U1157 (N_1157,In_330,In_1356);
or U1158 (N_1158,In_2689,In_1767);
nand U1159 (N_1159,In_1856,In_1534);
nand U1160 (N_1160,In_245,In_708);
nand U1161 (N_1161,In_1756,N_735);
or U1162 (N_1162,In_2504,N_976);
or U1163 (N_1163,In_2779,In_2961);
or U1164 (N_1164,In_1234,In_391);
nand U1165 (N_1165,N_536,In_770);
nor U1166 (N_1166,N_477,In_1290);
or U1167 (N_1167,In_2169,In_1779);
nor U1168 (N_1168,N_144,In_2914);
nor U1169 (N_1169,In_489,N_451);
or U1170 (N_1170,N_33,In_622);
nand U1171 (N_1171,In_2658,In_2367);
nor U1172 (N_1172,N_870,N_851);
nand U1173 (N_1173,In_2863,N_248);
nor U1174 (N_1174,In_265,N_60);
xnor U1175 (N_1175,In_1023,N_530);
or U1176 (N_1176,In_2918,In_1565);
or U1177 (N_1177,In_1737,In_2317);
nor U1178 (N_1178,N_825,In_1487);
nor U1179 (N_1179,N_606,In_99);
xor U1180 (N_1180,N_6,N_132);
nand U1181 (N_1181,N_564,In_325);
nand U1182 (N_1182,In_1931,N_869);
xnor U1183 (N_1183,In_267,N_593);
or U1184 (N_1184,N_300,In_1623);
nor U1185 (N_1185,N_279,N_494);
xnor U1186 (N_1186,In_861,In_1975);
or U1187 (N_1187,N_302,In_1522);
or U1188 (N_1188,N_731,In_534);
and U1189 (N_1189,In_1984,N_968);
nand U1190 (N_1190,N_182,In_901);
nand U1191 (N_1191,In_1951,N_938);
nor U1192 (N_1192,In_1962,In_2373);
nand U1193 (N_1193,In_2285,N_876);
or U1194 (N_1194,In_448,In_2986);
xnor U1195 (N_1195,N_958,In_323);
xor U1196 (N_1196,N_596,In_2578);
xnor U1197 (N_1197,In_1786,In_1277);
nor U1198 (N_1198,In_1063,In_2730);
or U1199 (N_1199,In_585,In_2586);
or U1200 (N_1200,In_626,In_2768);
nand U1201 (N_1201,In_655,N_551);
xnor U1202 (N_1202,In_1826,N_761);
xnor U1203 (N_1203,In_1551,In_2983);
xnor U1204 (N_1204,In_24,N_917);
or U1205 (N_1205,N_216,N_19);
xnor U1206 (N_1206,N_786,N_643);
or U1207 (N_1207,N_163,In_994);
nor U1208 (N_1208,In_2257,N_499);
or U1209 (N_1209,In_1647,N_523);
nand U1210 (N_1210,N_322,In_311);
nand U1211 (N_1211,In_119,In_2636);
xor U1212 (N_1212,N_172,N_452);
xnor U1213 (N_1213,In_2933,In_269);
xnor U1214 (N_1214,N_421,In_1817);
or U1215 (N_1215,In_736,In_545);
nor U1216 (N_1216,In_13,In_2466);
nand U1217 (N_1217,N_27,N_411);
and U1218 (N_1218,N_220,In_1656);
xor U1219 (N_1219,In_2417,N_980);
nand U1220 (N_1220,In_1201,In_553);
and U1221 (N_1221,N_575,In_2500);
and U1222 (N_1222,In_709,N_962);
xor U1223 (N_1223,In_1538,N_904);
or U1224 (N_1224,N_891,N_243);
nor U1225 (N_1225,In_45,N_677);
nand U1226 (N_1226,In_1092,N_623);
xnor U1227 (N_1227,N_848,In_2381);
or U1228 (N_1228,In_1326,N_664);
nand U1229 (N_1229,N_359,In_2938);
xnor U1230 (N_1230,In_1248,In_2400);
and U1231 (N_1231,N_84,In_1514);
or U1232 (N_1232,In_2835,In_1892);
nand U1233 (N_1233,In_1149,N_859);
nor U1234 (N_1234,N_903,In_2613);
xor U1235 (N_1235,In_2175,N_812);
or U1236 (N_1236,In_344,N_595);
nor U1237 (N_1237,In_1949,N_511);
xor U1238 (N_1238,In_2424,N_630);
nand U1239 (N_1239,In_2496,N_864);
nand U1240 (N_1240,In_1254,N_861);
or U1241 (N_1241,N_966,In_1636);
and U1242 (N_1242,N_923,N_775);
nand U1243 (N_1243,In_1769,N_873);
xor U1244 (N_1244,In_308,In_2283);
and U1245 (N_1245,In_1794,N_290);
or U1246 (N_1246,In_247,N_994);
or U1247 (N_1247,In_2941,In_114);
or U1248 (N_1248,In_1100,N_827);
xnor U1249 (N_1249,N_520,N_37);
xor U1250 (N_1250,N_940,N_445);
xor U1251 (N_1251,In_1575,In_996);
nand U1252 (N_1252,N_602,In_1696);
nor U1253 (N_1253,In_1468,N_884);
and U1254 (N_1254,N_149,N_990);
or U1255 (N_1255,In_440,N_319);
xor U1256 (N_1256,N_353,N_862);
nand U1257 (N_1257,N_73,In_1331);
or U1258 (N_1258,N_7,In_2043);
nand U1259 (N_1259,N_381,In_1669);
and U1260 (N_1260,N_920,In_2972);
nor U1261 (N_1261,In_896,N_396);
nand U1262 (N_1262,N_246,N_571);
nor U1263 (N_1263,N_446,N_765);
nand U1264 (N_1264,N_853,In_158);
or U1265 (N_1265,In_242,N_198);
nand U1266 (N_1266,In_2678,N_554);
nor U1267 (N_1267,N_915,In_1524);
xnor U1268 (N_1268,N_708,In_1179);
and U1269 (N_1269,N_576,In_97);
xnor U1270 (N_1270,N_527,In_2700);
and U1271 (N_1271,N_841,N_562);
xor U1272 (N_1272,N_333,In_2898);
nor U1273 (N_1273,In_2167,In_840);
nand U1274 (N_1274,In_857,In_974);
xnor U1275 (N_1275,In_743,In_1213);
nor U1276 (N_1276,N_745,In_648);
or U1277 (N_1277,In_389,N_510);
nand U1278 (N_1278,In_29,In_498);
nor U1279 (N_1279,N_456,N_637);
xor U1280 (N_1280,N_729,In_334);
and U1281 (N_1281,In_2782,In_1650);
nor U1282 (N_1282,In_83,In_991);
or U1283 (N_1283,N_342,In_2978);
and U1284 (N_1284,In_2430,In_1509);
or U1285 (N_1285,N_106,N_4);
xor U1286 (N_1286,N_330,N_971);
xnor U1287 (N_1287,In_1853,In_281);
nand U1288 (N_1288,N_718,In_376);
and U1289 (N_1289,N_772,In_411);
and U1290 (N_1290,N_207,In_1244);
xor U1291 (N_1291,N_989,In_66);
xor U1292 (N_1292,N_899,N_303);
nor U1293 (N_1293,In_403,N_358);
nor U1294 (N_1294,N_124,N_304);
or U1295 (N_1295,In_971,In_2293);
or U1296 (N_1296,In_1210,In_2530);
xnor U1297 (N_1297,In_2620,In_1006);
nor U1298 (N_1298,In_2565,In_1376);
nand U1299 (N_1299,In_2728,N_504);
nor U1300 (N_1300,In_2420,In_1075);
or U1301 (N_1301,N_378,In_1228);
nand U1302 (N_1302,N_423,In_749);
or U1303 (N_1303,In_596,N_991);
and U1304 (N_1304,In_672,In_511);
nand U1305 (N_1305,In_1854,In_159);
nor U1306 (N_1306,In_2042,In_830);
or U1307 (N_1307,In_2563,In_2054);
and U1308 (N_1308,N_416,In_1120);
nand U1309 (N_1309,In_1372,N_483);
and U1310 (N_1310,N_908,In_952);
and U1311 (N_1311,N_809,N_930);
and U1312 (N_1312,N_186,In_1612);
xnor U1313 (N_1313,N_542,In_805);
xnor U1314 (N_1314,N_507,N_681);
nor U1315 (N_1315,In_313,N_249);
and U1316 (N_1316,In_248,In_1987);
xnor U1317 (N_1317,In_2793,In_554);
nor U1318 (N_1318,N_238,In_2260);
and U1319 (N_1319,In_2554,In_1246);
nor U1320 (N_1320,In_1355,In_601);
nor U1321 (N_1321,In_954,N_545);
nor U1322 (N_1322,N_639,In_2435);
and U1323 (N_1323,In_504,N_796);
or U1324 (N_1324,N_187,N_522);
and U1325 (N_1325,In_939,In_1407);
and U1326 (N_1326,N_598,N_707);
and U1327 (N_1327,N_117,In_2203);
or U1328 (N_1328,N_26,N_911);
nor U1329 (N_1329,In_609,N_926);
or U1330 (N_1330,In_2375,N_738);
and U1331 (N_1331,In_2360,N_450);
or U1332 (N_1332,In_2174,N_826);
and U1333 (N_1333,N_877,In_2619);
nand U1334 (N_1334,N_957,N_573);
or U1335 (N_1335,In_130,In_1823);
xor U1336 (N_1336,In_2716,In_2592);
nand U1337 (N_1337,In_2718,In_700);
nor U1338 (N_1338,In_404,In_1700);
nor U1339 (N_1339,In_995,In_664);
nor U1340 (N_1340,In_2294,In_2309);
nand U1341 (N_1341,In_2097,In_1089);
nor U1342 (N_1342,In_1243,N_90);
nor U1343 (N_1343,N_501,N_35);
nor U1344 (N_1344,N_183,N_410);
nor U1345 (N_1345,In_2974,In_2168);
or U1346 (N_1346,In_2553,In_1036);
or U1347 (N_1347,In_679,In_846);
or U1348 (N_1348,In_1910,N_334);
and U1349 (N_1349,In_1621,In_1456);
nand U1350 (N_1350,N_592,In_583);
xnor U1351 (N_1351,N_368,N_791);
and U1352 (N_1352,In_1148,In_1469);
or U1353 (N_1353,In_1746,In_786);
nor U1354 (N_1354,N_524,In_1461);
or U1355 (N_1355,In_53,N_224);
xor U1356 (N_1356,N_919,In_883);
nor U1357 (N_1357,In_1387,In_735);
and U1358 (N_1358,In_2629,N_961);
xnor U1359 (N_1359,In_750,In_2215);
or U1360 (N_1360,In_2570,N_283);
nand U1361 (N_1361,N_799,N_382);
nor U1362 (N_1362,In_382,In_649);
nor U1363 (N_1363,In_492,N_784);
and U1364 (N_1364,N_245,In_405);
and U1365 (N_1365,N_362,N_697);
xnor U1366 (N_1366,N_100,In_112);
and U1367 (N_1367,N_714,In_613);
xnor U1368 (N_1368,In_225,N_348);
and U1369 (N_1369,In_548,In_2637);
or U1370 (N_1370,In_2662,N_792);
nor U1371 (N_1371,In_2612,N_951);
nor U1372 (N_1372,In_297,In_1457);
and U1373 (N_1373,N_667,In_2440);
nand U1374 (N_1374,N_432,In_2957);
nand U1375 (N_1375,N_620,In_1938);
and U1376 (N_1376,In_1350,In_2288);
and U1377 (N_1377,In_59,N_343);
or U1378 (N_1378,N_404,In_1809);
and U1379 (N_1379,In_476,In_2999);
and U1380 (N_1380,N_101,N_829);
or U1381 (N_1381,N_582,In_931);
and U1382 (N_1382,N_143,N_856);
xor U1383 (N_1383,In_870,N_390);
nor U1384 (N_1384,In_859,N_965);
and U1385 (N_1385,In_172,In_558);
and U1386 (N_1386,In_2930,N_913);
and U1387 (N_1387,In_1730,In_1981);
or U1388 (N_1388,In_2967,In_2900);
and U1389 (N_1389,In_1168,N_529);
nor U1390 (N_1390,In_2725,In_1031);
nand U1391 (N_1391,In_2312,In_1428);
nand U1392 (N_1392,In_1186,In_2436);
nand U1393 (N_1393,In_2151,N_974);
nand U1394 (N_1394,N_946,In_1844);
or U1395 (N_1395,N_505,In_1008);
nand U1396 (N_1396,In_1346,In_231);
xnor U1397 (N_1397,In_107,In_1010);
and U1398 (N_1398,N_764,N_815);
xor U1399 (N_1399,In_880,N_689);
or U1400 (N_1400,In_2246,In_2372);
or U1401 (N_1401,N_621,In_1275);
or U1402 (N_1402,In_509,In_573);
nor U1403 (N_1403,In_2703,In_992);
and U1404 (N_1404,In_1708,In_2932);
xnor U1405 (N_1405,In_2338,In_1918);
xnor U1406 (N_1406,In_1046,In_513);
or U1407 (N_1407,In_82,In_2387);
nor U1408 (N_1408,In_90,N_834);
nand U1409 (N_1409,In_1054,N_819);
xor U1410 (N_1410,In_886,In_417);
xnor U1411 (N_1411,N_328,In_635);
and U1412 (N_1412,N_755,In_2568);
and U1413 (N_1413,In_2091,N_900);
nand U1414 (N_1414,N_823,In_2439);
nand U1415 (N_1415,In_1164,In_1744);
nand U1416 (N_1416,In_1096,In_1178);
and U1417 (N_1417,In_1727,In_1584);
or U1418 (N_1418,In_1205,In_460);
or U1419 (N_1419,In_2917,In_1980);
xnor U1420 (N_1420,N_801,In_923);
xor U1421 (N_1421,In_234,N_700);
xnor U1422 (N_1422,N_875,In_494);
xor U1423 (N_1423,N_399,In_1159);
nor U1424 (N_1424,In_2116,In_1101);
xor U1425 (N_1425,N_821,In_136);
or U1426 (N_1426,In_576,N_895);
and U1427 (N_1427,In_2133,N_375);
nor U1428 (N_1428,In_1762,N_212);
and U1429 (N_1429,N_874,In_2610);
nor U1430 (N_1430,N_767,In_819);
and U1431 (N_1431,In_712,N_698);
xor U1432 (N_1432,N_663,N_87);
nor U1433 (N_1433,In_821,N_464);
xor U1434 (N_1434,N_577,In_727);
nor U1435 (N_1435,In_1757,N_48);
xnor U1436 (N_1436,In_2906,In_457);
xor U1437 (N_1437,N_272,N_883);
and U1438 (N_1438,N_701,N_470);
xnor U1439 (N_1439,N_370,In_1489);
nor U1440 (N_1440,N_153,In_1564);
or U1441 (N_1441,N_807,N_673);
or U1442 (N_1442,In_1709,N_555);
and U1443 (N_1443,N_793,In_2686);
and U1444 (N_1444,In_720,N_400);
or U1445 (N_1445,N_493,In_2128);
and U1446 (N_1446,N_712,In_1542);
nand U1447 (N_1447,In_1579,In_2634);
xor U1448 (N_1448,N_179,N_942);
nand U1449 (N_1449,In_1799,N_586);
xnor U1450 (N_1450,In_410,N_634);
nand U1451 (N_1451,In_2821,N_881);
xnor U1452 (N_1452,In_370,In_895);
xor U1453 (N_1453,N_932,In_192);
xnor U1454 (N_1454,In_1563,N_588);
and U1455 (N_1455,In_2980,N_710);
and U1456 (N_1456,N_487,N_610);
nor U1457 (N_1457,N_68,In_1252);
nor U1458 (N_1458,N_0,In_1181);
and U1459 (N_1459,N_174,In_1611);
nand U1460 (N_1460,In_1069,N_756);
xor U1461 (N_1461,In_1437,In_1689);
nand U1462 (N_1462,In_1941,In_2204);
or U1463 (N_1463,In_2854,N_822);
and U1464 (N_1464,In_1628,In_2969);
xnor U1465 (N_1465,In_761,In_1839);
or U1466 (N_1466,In_1042,In_561);
nor U1467 (N_1467,In_293,In_1212);
xor U1468 (N_1468,In_1142,N_785);
or U1469 (N_1469,In_454,In_1439);
nand U1470 (N_1470,N_699,N_50);
and U1471 (N_1471,In_1654,N_837);
nor U1472 (N_1472,In_1293,In_1585);
and U1473 (N_1473,In_2618,N_581);
xnor U1474 (N_1474,In_1460,N_811);
or U1475 (N_1475,In_2551,N_607);
xnor U1476 (N_1476,In_1182,In_2807);
or U1477 (N_1477,N_781,In_2920);
and U1478 (N_1478,N_750,In_678);
and U1479 (N_1479,In_456,In_490);
nor U1480 (N_1480,In_2697,N_736);
nand U1481 (N_1481,In_653,N_184);
nand U1482 (N_1482,In_332,In_790);
nand U1483 (N_1483,In_1545,In_272);
nand U1484 (N_1484,In_446,In_317);
xnor U1485 (N_1485,In_215,N_168);
nand U1486 (N_1486,In_398,In_1003);
or U1487 (N_1487,In_2694,N_99);
nor U1488 (N_1488,In_1655,In_1889);
xor U1489 (N_1489,In_987,N_670);
nor U1490 (N_1490,In_1515,N_912);
nand U1491 (N_1491,N_649,N_242);
nand U1492 (N_1492,In_1452,In_2100);
or U1493 (N_1493,In_2088,N_43);
xor U1494 (N_1494,N_160,N_889);
xnor U1495 (N_1495,N_752,In_1882);
and U1496 (N_1496,In_2114,N_753);
xnor U1497 (N_1497,In_1477,N_635);
and U1498 (N_1498,In_2191,In_1291);
or U1499 (N_1499,In_350,In_661);
nor U1500 (N_1500,In_2047,N_1346);
or U1501 (N_1501,N_1385,In_481);
or U1502 (N_1502,N_995,In_2017);
and U1503 (N_1503,N_1212,In_497);
nor U1504 (N_1504,In_753,N_1387);
nor U1505 (N_1505,In_2708,In_1544);
and U1506 (N_1506,In_4,In_878);
xnor U1507 (N_1507,N_860,N_1178);
and U1508 (N_1508,N_1225,In_2344);
or U1509 (N_1509,In_2813,In_2876);
nand U1510 (N_1510,N_725,In_521);
and U1511 (N_1511,N_1137,In_1888);
xnor U1512 (N_1512,N_1382,N_1446);
and U1513 (N_1513,N_1214,N_1072);
nand U1514 (N_1514,In_1177,N_1152);
xor U1515 (N_1515,In_2350,N_1439);
and U1516 (N_1516,In_16,In_1154);
nand U1517 (N_1517,N_886,In_1836);
nor U1518 (N_1518,In_1218,In_1327);
or U1519 (N_1519,In_1082,In_2481);
nand U1520 (N_1520,In_2154,In_2370);
nand U1521 (N_1521,N_704,N_1185);
nand U1522 (N_1522,N_969,In_1562);
nand U1523 (N_1523,In_2547,N_948);
or U1524 (N_1524,N_1005,In_2975);
and U1525 (N_1525,N_1200,N_1409);
and U1526 (N_1526,N_417,In_2498);
and U1527 (N_1527,In_1384,N_1163);
or U1528 (N_1528,In_1748,N_56);
nor U1529 (N_1529,N_762,N_1291);
nand U1530 (N_1530,In_1393,N_1041);
or U1531 (N_1531,N_693,N_1443);
nor U1532 (N_1532,N_194,N_1058);
and U1533 (N_1533,N_344,In_2765);
xnor U1534 (N_1534,In_2302,N_1028);
nand U1535 (N_1535,N_55,N_75);
or U1536 (N_1536,N_1146,N_1026);
xor U1537 (N_1537,In_2748,N_744);
or U1538 (N_1538,N_1162,In_1435);
or U1539 (N_1539,N_655,In_2348);
nor U1540 (N_1540,N_1268,N_1353);
nand U1541 (N_1541,In_2880,N_1195);
xnor U1542 (N_1542,In_2280,N_810);
xnor U1543 (N_1543,N_616,N_53);
and U1544 (N_1544,In_1530,N_1413);
and U1545 (N_1545,In_1969,In_2503);
nor U1546 (N_1546,N_251,N_1490);
nand U1547 (N_1547,N_426,In_52);
nand U1548 (N_1548,In_510,In_1222);
xnor U1549 (N_1549,N_1318,N_1400);
nor U1550 (N_1550,N_488,N_1242);
and U1551 (N_1551,In_433,N_982);
or U1552 (N_1552,N_1244,In_738);
nor U1553 (N_1553,In_843,N_1033);
nand U1554 (N_1554,N_1467,N_928);
nor U1555 (N_1555,N_1455,In_2643);
nand U1556 (N_1556,N_1176,In_2644);
xor U1557 (N_1557,In_2037,In_484);
xnor U1558 (N_1558,N_741,In_839);
or U1559 (N_1559,N_727,N_1001);
and U1560 (N_1560,In_351,N_626);
nor U1561 (N_1561,In_364,N_1479);
nor U1562 (N_1562,In_1638,N_887);
xor U1563 (N_1563,In_2406,N_1150);
nor U1564 (N_1564,N_1397,In_1603);
and U1565 (N_1565,In_189,N_1025);
nor U1566 (N_1566,N_1106,In_2073);
nand U1567 (N_1567,In_380,N_1078);
xor U1568 (N_1568,In_2398,N_1272);
xnor U1569 (N_1569,N_600,N_201);
nor U1570 (N_1570,N_1464,In_877);
nor U1571 (N_1571,In_1408,N_1265);
and U1572 (N_1572,N_1222,N_1149);
nand U1573 (N_1573,N_898,N_614);
and U1574 (N_1574,N_503,In_2483);
nand U1575 (N_1575,In_2465,N_618);
and U1576 (N_1576,N_261,N_740);
or U1577 (N_1577,N_515,In_1691);
nor U1578 (N_1578,In_1308,N_1006);
nand U1579 (N_1579,In_374,N_1282);
or U1580 (N_1580,In_1765,In_704);
nand U1581 (N_1581,N_918,N_1300);
or U1582 (N_1582,N_1349,N_1412);
nand U1583 (N_1583,In_560,N_1125);
nand U1584 (N_1584,N_1248,N_732);
nand U1585 (N_1585,N_1419,N_418);
xnor U1586 (N_1586,N_1238,N_858);
and U1587 (N_1587,N_1303,N_1416);
nor U1588 (N_1588,N_275,N_907);
nor U1589 (N_1589,N_852,N_1076);
nor U1590 (N_1590,N_1016,In_1123);
and U1591 (N_1591,In_1017,In_139);
or U1592 (N_1592,In_1683,N_964);
and U1593 (N_1593,In_2519,N_1166);
nand U1594 (N_1594,N_1275,N_469);
and U1595 (N_1595,N_597,In_2298);
nand U1596 (N_1596,N_1086,N_1255);
nand U1597 (N_1597,In_1982,N_1018);
nand U1598 (N_1598,In_607,In_614);
xor U1599 (N_1599,In_616,In_2268);
and U1600 (N_1600,In_472,N_498);
and U1601 (N_1601,N_1083,In_1072);
or U1602 (N_1602,N_1371,In_2229);
nor U1603 (N_1603,N_653,N_949);
or U1604 (N_1604,In_692,N_479);
nor U1605 (N_1605,In_1401,In_1760);
xnor U1606 (N_1606,N_1428,In_2395);
and U1607 (N_1607,N_1186,N_373);
xor U1608 (N_1608,N_1350,In_905);
and U1609 (N_1609,In_1986,N_1022);
and U1610 (N_1610,In_744,N_119);
or U1611 (N_1611,N_1220,N_1068);
nor U1612 (N_1612,N_963,N_1009);
and U1613 (N_1613,N_780,N_1174);
nand U1614 (N_1614,In_1978,N_1157);
xnor U1615 (N_1615,In_2253,N_1285);
or U1616 (N_1616,In_2977,N_1327);
and U1617 (N_1617,N_705,N_1289);
nand U1618 (N_1618,In_1511,N_783);
xor U1619 (N_1619,N_1363,In_2593);
nand U1620 (N_1620,N_986,N_1417);
or U1621 (N_1621,N_341,N_730);
xnor U1622 (N_1622,N_1048,N_924);
nand U1623 (N_1623,In_1143,N_1029);
and U1624 (N_1624,In_650,N_1460);
and U1625 (N_1625,N_490,In_1554);
or U1626 (N_1626,N_1399,In_1280);
or U1627 (N_1627,In_2423,In_2532);
or U1628 (N_1628,In_1587,N_1240);
nand U1629 (N_1629,N_1309,In_378);
xnor U1630 (N_1630,N_1378,N_984);
or U1631 (N_1631,In_369,In_742);
nor U1632 (N_1632,N_1065,N_1205);
nor U1633 (N_1633,In_1465,N_1404);
nand U1634 (N_1634,N_1474,N_526);
nor U1635 (N_1635,N_627,In_1824);
or U1636 (N_1636,In_1848,In_2432);
and U1637 (N_1637,In_2786,N_885);
xor U1638 (N_1638,In_2971,N_896);
xnor U1639 (N_1639,N_1056,N_1253);
xnor U1640 (N_1640,In_475,N_327);
or U1641 (N_1641,N_1140,N_299);
xnor U1642 (N_1642,In_2885,In_620);
nand U1643 (N_1643,N_817,N_1160);
nand U1644 (N_1644,N_203,N_1144);
and U1645 (N_1645,In_1806,N_1478);
nand U1646 (N_1646,N_632,N_1414);
nor U1647 (N_1647,N_1306,N_1354);
nand U1648 (N_1648,In_2089,In_701);
nor U1649 (N_1649,In_2201,N_694);
nand U1650 (N_1650,In_871,N_1322);
nor U1651 (N_1651,N_1420,N_1143);
and U1652 (N_1652,N_1204,N_1062);
and U1653 (N_1653,N_1122,In_689);
xnor U1654 (N_1654,N_447,In_2028);
nor U1655 (N_1655,In_1,N_820);
nand U1656 (N_1656,N_393,N_1325);
nor U1657 (N_1657,N_934,N_1047);
and U1658 (N_1658,In_2354,In_2651);
nand U1659 (N_1659,N_1117,In_1898);
or U1660 (N_1660,In_116,N_1377);
and U1661 (N_1661,In_2800,In_2734);
nor U1662 (N_1662,N_866,N_854);
and U1663 (N_1663,N_1148,N_847);
and U1664 (N_1664,N_1120,N_10);
nand U1665 (N_1665,N_380,N_758);
and U1666 (N_1666,N_1039,N_1499);
or U1667 (N_1667,N_1110,N_1415);
xor U1668 (N_1668,In_2723,N_1184);
and U1669 (N_1669,In_1060,In_1788);
xor U1670 (N_1670,N_1074,In_834);
and U1671 (N_1671,N_1426,N_625);
nand U1672 (N_1672,In_2674,N_1099);
xnor U1673 (N_1673,N_1142,N_1492);
nand U1674 (N_1674,N_902,In_503);
or U1675 (N_1675,In_1288,N_648);
and U1676 (N_1676,N_835,In_638);
nor U1677 (N_1677,N_845,N_1448);
nor U1678 (N_1678,In_1855,N_1276);
nor U1679 (N_1679,In_2141,N_661);
or U1680 (N_1680,N_1132,N_1280);
or U1681 (N_1681,N_1264,In_2673);
xor U1682 (N_1682,N_1061,In_1260);
xor U1683 (N_1683,In_2289,In_2572);
nand U1684 (N_1684,N_872,In_89);
xnor U1685 (N_1685,In_958,N_1401);
nand U1686 (N_1686,N_1328,N_733);
nand U1687 (N_1687,N_219,N_1246);
or U1688 (N_1688,In_2874,In_298);
and U1689 (N_1689,In_414,N_1284);
nand U1690 (N_1690,N_1396,N_1043);
xor U1691 (N_1691,In_1250,N_1046);
or U1692 (N_1692,N_1069,N_1271);
and U1693 (N_1693,N_888,In_2699);
nand U1694 (N_1694,N_1456,N_199);
xor U1695 (N_1695,N_538,In_173);
and U1696 (N_1696,N_1436,N_508);
nor U1697 (N_1697,N_1097,N_1105);
or U1698 (N_1698,In_2464,In_1370);
nand U1699 (N_1699,N_914,N_111);
nand U1700 (N_1700,N_1095,N_1229);
or U1701 (N_1701,In_1678,In_284);
and U1702 (N_1702,N_1057,N_782);
xor U1703 (N_1703,N_1389,N_1342);
nand U1704 (N_1704,N_1273,N_1410);
or U1705 (N_1705,N_41,In_1207);
xor U1706 (N_1706,N_1197,N_553);
xnor U1707 (N_1707,N_1266,In_2890);
nor U1708 (N_1708,In_2955,In_427);
nor U1709 (N_1709,In_2477,N_950);
nor U1710 (N_1710,N_831,N_561);
or U1711 (N_1711,N_492,In_2584);
or U1712 (N_1712,N_1362,In_2562);
or U1713 (N_1713,In_64,In_1160);
or U1714 (N_1714,N_429,N_295);
nor U1715 (N_1715,N_1441,N_1129);
nand U1716 (N_1716,In_2905,N_748);
xnor U1717 (N_1717,In_2199,In_1768);
xor U1718 (N_1718,N_484,N_879);
or U1719 (N_1719,N_1201,N_107);
xor U1720 (N_1720,N_535,N_1224);
nand U1721 (N_1721,N_137,N_1488);
and U1722 (N_1722,In_532,In_1080);
nand U1723 (N_1723,In_1048,In_421);
nand U1724 (N_1724,In_2924,N_742);
and U1725 (N_1725,N_1254,N_509);
nor U1726 (N_1726,N_646,N_1181);
nor U1727 (N_1727,N_1338,In_2561);
xor U1728 (N_1728,In_968,N_40);
nor U1729 (N_1729,In_69,In_1430);
nand U1730 (N_1730,In_1963,N_1216);
xor U1731 (N_1731,In_1431,N_1236);
xor U1732 (N_1732,N_1015,In_2591);
and U1733 (N_1733,In_2025,N_850);
or U1734 (N_1734,In_2710,N_1249);
or U1735 (N_1735,In_2242,N_1481);
and U1736 (N_1736,N_678,N_377);
and U1737 (N_1737,N_1180,In_2709);
and U1738 (N_1738,N_916,N_568);
nor U1739 (N_1739,N_1116,N_1131);
xor U1740 (N_1740,In_2240,In_718);
and U1741 (N_1741,N_1054,N_192);
nor U1742 (N_1742,N_204,In_2630);
nand U1743 (N_1743,In_2804,N_615);
and U1744 (N_1744,In_676,N_1356);
nor U1745 (N_1745,In_2235,In_836);
and U1746 (N_1746,N_435,N_1310);
or U1747 (N_1747,N_1147,In_2891);
nor U1748 (N_1748,In_1055,N_25);
nor U1749 (N_1749,N_1383,N_1360);
nor U1750 (N_1750,In_2514,N_336);
nor U1751 (N_1751,N_1241,N_130);
nand U1752 (N_1752,In_1315,In_1881);
or U1753 (N_1753,N_1316,In_2003);
nor U1754 (N_1754,N_1473,N_1053);
xnor U1755 (N_1755,N_1036,N_1067);
nand U1756 (N_1756,In_2055,N_746);
nand U1757 (N_1757,N_1252,N_66);
nand U1758 (N_1758,N_114,In_670);
and U1759 (N_1759,N_633,In_342);
and U1760 (N_1760,In_2660,In_1404);
and U1761 (N_1761,N_1476,In_264);
nand U1762 (N_1762,N_686,In_1474);
xor U1763 (N_1763,N_1207,N_1398);
and U1764 (N_1764,In_1158,In_2647);
nand U1765 (N_1765,N_1115,N_1021);
nand U1766 (N_1766,N_1175,N_331);
or U1767 (N_1767,N_282,N_739);
or U1768 (N_1768,N_939,N_589);
or U1769 (N_1769,In_726,N_1256);
nor U1770 (N_1770,N_757,N_1189);
or U1771 (N_1771,N_1394,N_645);
and U1772 (N_1772,In_155,N_1088);
and U1773 (N_1773,In_260,N_594);
nor U1774 (N_1774,N_1153,In_983);
nand U1775 (N_1775,In_270,N_836);
and U1776 (N_1776,In_804,N_1257);
nand U1777 (N_1777,N_1483,N_1374);
xor U1778 (N_1778,N_1141,N_1457);
or U1779 (N_1779,In_2566,N_547);
nor U1780 (N_1780,In_47,N_604);
xor U1781 (N_1781,N_1296,N_1100);
xor U1782 (N_1782,N_1344,N_1260);
nand U1783 (N_1783,N_1372,N_540);
nor U1784 (N_1784,N_502,N_1170);
nor U1785 (N_1785,N_310,N_1188);
or U1786 (N_1786,N_36,N_1259);
or U1787 (N_1787,N_778,In_2860);
nor U1788 (N_1788,N_1431,In_1064);
xnor U1789 (N_1789,In_1649,N_59);
xnor U1790 (N_1790,N_1365,In_1337);
and U1791 (N_1791,In_1661,N_1190);
xor U1792 (N_1792,N_145,In_2122);
nand U1793 (N_1793,In_1774,N_1337);
or U1794 (N_1794,In_2272,N_1320);
nand U1795 (N_1795,In_1066,N_441);
nand U1796 (N_1796,In_1418,In_1929);
xor U1797 (N_1797,N_1209,N_773);
nor U1798 (N_1798,In_684,N_1239);
and U1799 (N_1799,N_1032,N_557);
or U1800 (N_1800,In_2928,N_1434);
xor U1801 (N_1801,N_999,N_151);
nand U1802 (N_1802,In_2195,N_609);
and U1803 (N_1803,N_1055,N_1345);
or U1804 (N_1804,In_74,N_1392);
and U1805 (N_1805,In_581,N_688);
xnor U1806 (N_1806,N_228,In_845);
xor U1807 (N_1807,N_363,N_1407);
nor U1808 (N_1808,In_91,N_1124);
and U1809 (N_1809,In_1631,In_1378);
xnor U1810 (N_1810,N_1237,N_131);
and U1811 (N_1811,N_1305,In_1284);
xnor U1812 (N_1812,N_541,N_1321);
and U1813 (N_1813,N_1471,In_1695);
nor U1814 (N_1814,N_893,In_1659);
nor U1815 (N_1815,N_1281,N_415);
nor U1816 (N_1816,N_1199,N_1044);
and U1817 (N_1817,In_63,N_1059);
nand U1818 (N_1818,In_926,N_171);
nand U1819 (N_1819,In_1934,In_2831);
nor U1820 (N_1820,In_814,N_1442);
or U1821 (N_1821,In_2390,N_1183);
xnor U1822 (N_1822,N_565,N_1050);
and U1823 (N_1823,N_685,In_1018);
nand U1824 (N_1824,N_867,N_1339);
nand U1825 (N_1825,N_1438,N_816);
nor U1826 (N_1826,N_1380,N_1269);
nand U1827 (N_1827,N_1085,In_2979);
xnor U1828 (N_1828,N_1336,In_766);
nand U1829 (N_1829,N_1484,In_733);
xnor U1830 (N_1830,In_1081,N_1279);
nor U1831 (N_1831,N_1314,N_471);
nand U1832 (N_1832,In_1021,N_1489);
xor U1833 (N_1833,N_1331,N_356);
nand U1834 (N_1834,In_2625,N_1495);
xor U1835 (N_1835,N_790,N_709);
xnor U1836 (N_1836,N_30,N_743);
and U1837 (N_1837,N_671,N_1112);
and U1838 (N_1838,In_1193,N_1094);
nand U1839 (N_1839,N_1134,In_780);
and U1840 (N_1840,N_662,In_1166);
xnor U1841 (N_1841,N_638,N_1294);
xnor U1842 (N_1842,In_1893,N_297);
xor U1843 (N_1843,In_644,N_1487);
nand U1844 (N_1844,N_1087,N_401);
nand U1845 (N_1845,N_720,N_1127);
or U1846 (N_1846,In_2166,N_833);
nor U1847 (N_1847,N_802,In_2371);
and U1848 (N_1848,In_341,N_20);
and U1849 (N_1849,N_1156,N_1198);
nand U1850 (N_1850,N_1155,N_226);
or U1851 (N_1851,N_1194,In_2494);
nor U1852 (N_1852,In_452,N_528);
nand U1853 (N_1853,N_612,N_1304);
or U1854 (N_1854,In_2063,In_2044);
nand U1855 (N_1855,N_719,N_1493);
nand U1856 (N_1856,In_1204,In_835);
xor U1857 (N_1857,N_1121,N_1418);
nor U1858 (N_1858,N_608,N_1172);
or U1859 (N_1859,In_41,N_983);
nand U1860 (N_1860,In_2330,N_1452);
nand U1861 (N_1861,In_426,In_165);
xnor U1862 (N_1862,In_1738,In_1084);
nand U1863 (N_1863,N_1341,N_1326);
xor U1864 (N_1864,In_1090,N_1472);
and U1865 (N_1865,N_651,N_993);
and U1866 (N_1866,N_1206,N_1485);
and U1867 (N_1867,N_1070,N_960);
and U1868 (N_1868,N_133,N_1277);
and U1869 (N_1869,In_1108,In_2112);
xnor U1870 (N_1870,In_2090,N_776);
and U1871 (N_1871,N_516,N_1213);
xor U1872 (N_1872,N_1270,N_350);
and U1873 (N_1873,In_1673,N_16);
nor U1874 (N_1874,In_1596,In_1151);
xor U1875 (N_1875,In_188,In_2177);
and U1876 (N_1876,N_213,In_751);
nor U1877 (N_1877,N_105,In_377);
and U1878 (N_1878,N_1466,N_590);
nand U1879 (N_1879,In_2615,N_1203);
or U1880 (N_1880,N_1388,N_1126);
xor U1881 (N_1881,N_454,In_2110);
and U1882 (N_1882,In_2540,In_1091);
and U1883 (N_1883,N_225,N_1351);
xor U1884 (N_1884,In_543,In_2192);
or U1885 (N_1885,In_384,In_1793);
nor U1886 (N_1886,N_1430,N_795);
nand U1887 (N_1887,N_1064,In_2020);
nor U1888 (N_1888,In_940,In_120);
nor U1889 (N_1889,In_2,N_326);
nor U1890 (N_1890,In_2646,N_550);
nor U1891 (N_1891,N_754,In_1313);
or U1892 (N_1892,In_168,N_1019);
or U1893 (N_1893,N_1196,N_517);
or U1894 (N_1894,N_1403,N_1084);
nor U1895 (N_1895,In_15,N_759);
nand U1896 (N_1896,N_1167,In_1360);
xnor U1897 (N_1897,In_980,N_1136);
xnor U1898 (N_1898,N_953,In_191);
and U1899 (N_1899,In_2254,N_281);
xnor U1900 (N_1900,N_1011,In_2884);
xor U1901 (N_1901,N_532,N_1411);
or U1902 (N_1902,N_871,N_1491);
xnor U1903 (N_1903,N_1066,N_112);
and U1904 (N_1904,N_1267,N_1480);
xnor U1905 (N_1905,In_58,In_2732);
and U1906 (N_1906,N_1334,N_587);
nand U1907 (N_1907,N_1454,In_2937);
or U1908 (N_1908,N_1348,In_1976);
and U1909 (N_1909,In_2158,In_973);
xnor U1910 (N_1910,N_1329,In_432);
nor U1911 (N_1911,N_567,N_1243);
nor U1912 (N_1912,N_1262,N_546);
nor U1913 (N_1913,In_1324,In_663);
and U1914 (N_1914,N_1221,N_1187);
and U1915 (N_1915,N_1211,N_803);
or U1916 (N_1916,N_531,In_791);
or U1917 (N_1917,N_988,N_843);
and U1918 (N_1918,N_206,In_1269);
and U1919 (N_1919,N_1311,In_2594);
nand U1920 (N_1920,In_135,N_1361);
and U1921 (N_1921,N_1319,N_1231);
and U1922 (N_1922,In_205,In_2434);
xnor U1923 (N_1923,N_1444,N_1052);
nand U1924 (N_1924,N_1118,N_611);
nand U1925 (N_1925,N_1003,N_459);
or U1926 (N_1926,N_631,In_1012);
nor U1927 (N_1927,In_2623,In_855);
xor U1928 (N_1928,In_2316,N_925);
xor U1929 (N_1929,N_1263,In_2812);
xnor U1930 (N_1930,N_1215,N_439);
nor U1931 (N_1931,N_478,N_1287);
and U1932 (N_1932,N_1343,N_1171);
xor U1933 (N_1933,N_81,N_1423);
xor U1934 (N_1934,N_79,In_961);
xnor U1935 (N_1935,N_1114,N_937);
or U1936 (N_1936,N_1440,In_2121);
nor U1937 (N_1937,In_1409,N_1007);
nor U1938 (N_1938,N_1347,N_74);
xnor U1939 (N_1939,In_1146,N_1017);
nand U1940 (N_1940,N_110,N_945);
or U1941 (N_1941,In_223,N_428);
xnor U1942 (N_1942,N_978,N_1379);
xnor U1943 (N_1943,In_2987,N_1077);
nor U1944 (N_1944,In_1869,In_1764);
and U1945 (N_1945,N_1405,N_674);
nand U1946 (N_1946,In_1602,In_768);
nand U1947 (N_1947,N_355,N_1369);
nor U1948 (N_1948,N_1108,In_2755);
nand U1949 (N_1949,N_944,In_2529);
or U1950 (N_1950,N_566,N_277);
nor U1951 (N_1951,In_2742,In_2850);
and U1952 (N_1952,N_1000,N_1366);
nand U1953 (N_1953,N_1182,N_805);
nor U1954 (N_1954,N_1402,N_1449);
and U1955 (N_1955,N_909,In_76);
nor U1956 (N_1956,In_2099,N_717);
xnor U1957 (N_1957,In_2921,N_1293);
and U1958 (N_1958,In_1209,In_2712);
xor U1959 (N_1959,In_1022,In_1073);
nand U1960 (N_1960,N_556,In_149);
nand U1961 (N_1961,In_1868,In_516);
nor U1962 (N_1962,In_1472,N_138);
nand U1963 (N_1963,N_1482,N_211);
and U1964 (N_1964,In_396,N_88);
xor U1965 (N_1965,N_1228,N_1459);
xor U1966 (N_1966,N_659,In_499);
or U1967 (N_1967,N_1340,N_1424);
nand U1968 (N_1968,N_1020,In_54);
or U1969 (N_1969,In_2726,In_1533);
xor U1970 (N_1970,In_2461,In_777);
xor U1971 (N_1971,In_2870,In_1032);
and U1972 (N_1972,In_1486,N_537);
nor U1973 (N_1973,N_660,In_1058);
xnor U1974 (N_1974,In_1645,N_706);
nand U1975 (N_1975,N_654,N_85);
or U1976 (N_1976,N_465,In_1453);
nand U1977 (N_1977,In_1541,In_458);
xor U1978 (N_1978,N_307,N_1208);
and U1979 (N_1979,N_813,In_1989);
nor U1980 (N_1980,N_1498,N_1014);
or U1981 (N_1981,In_677,In_1459);
nor U1982 (N_1982,N_1475,In_2846);
nand U1983 (N_1983,N_1002,N_291);
or U1984 (N_1984,N_1298,In_892);
and U1985 (N_1985,In_237,N_1427);
nand U1986 (N_1986,N_1060,N_1218);
nand U1987 (N_1987,N_1227,N_1395);
nand U1988 (N_1988,N_1324,In_1747);
and U1989 (N_1989,N_1494,N_1082);
xor U1990 (N_1990,In_2328,N_1390);
nand U1991 (N_1991,In_1029,N_840);
xnor U1992 (N_1992,N_1089,In_608);
and U1993 (N_1993,N_1145,N_1433);
xor U1994 (N_1994,N_842,N_1233);
xor U1995 (N_1995,N_574,N_31);
and U1996 (N_1996,N_696,In_1798);
or U1997 (N_1997,In_759,N_1251);
xnor U1998 (N_1998,N_1013,N_1447);
and U1999 (N_1999,N_585,N_747);
nand U2000 (N_2000,In_1657,N_270);
and U2001 (N_2001,N_1375,In_2036);
xor U2002 (N_2002,N_1648,N_1040);
xor U2003 (N_2003,N_1799,N_1639);
or U2004 (N_2004,N_1766,N_1543);
and U2005 (N_2005,N_1864,N_1465);
nand U2006 (N_2006,N_458,N_1506);
nand U2007 (N_2007,In_1140,N_1951);
nand U2008 (N_2008,N_679,N_1235);
and U2009 (N_2009,N_1740,N_1592);
nand U2010 (N_2010,N_1570,In_711);
xnor U2011 (N_2011,N_1705,N_716);
nand U2012 (N_2012,N_1594,N_1098);
xor U2013 (N_2013,N_1030,N_1852);
nor U2014 (N_2014,N_1690,N_1557);
nand U2015 (N_2015,N_1955,N_1010);
or U2016 (N_2016,N_1610,In_305);
nor U2017 (N_2017,N_136,N_570);
nand U2018 (N_2018,In_1527,N_1315);
and U2019 (N_2019,In_1897,N_1866);
and U2020 (N_2020,N_311,N_1832);
nand U2021 (N_2021,N_1863,N_977);
or U2022 (N_2022,In_1792,N_1432);
nor U2023 (N_2023,N_1911,In_547);
and U2024 (N_2024,N_1728,N_690);
nor U2025 (N_2025,N_1685,N_1823);
nand U2026 (N_2026,In_1353,N_1004);
or U2027 (N_2027,N_1512,N_1367);
and U2028 (N_2028,N_1981,N_1518);
xnor U2029 (N_2029,In_2412,N_1635);
nand U2030 (N_2030,N_1542,In_400);
and U2031 (N_2031,N_438,In_1828);
or U2032 (N_2032,N_1038,In_1677);
or U2033 (N_2033,N_78,N_1590);
and U2034 (N_2034,N_1605,N_1894);
nor U2035 (N_2035,N_814,N_1667);
nor U2036 (N_2036,N_1470,N_1528);
nor U2037 (N_2037,N_1746,N_1716);
nor U2038 (N_2038,In_2573,N_420);
and U2039 (N_2039,In_2670,N_1161);
xnor U2040 (N_2040,N_1192,N_1049);
nor U2041 (N_2041,N_1641,N_1368);
and U2042 (N_2042,N_1709,In_997);
or U2043 (N_2043,In_2336,N_1834);
and U2044 (N_2044,In_2142,N_1514);
xnor U2045 (N_2045,N_734,In_1015);
nand U2046 (N_2046,N_1537,N_1128);
and U2047 (N_2047,In_2875,N_1738);
nor U2048 (N_2048,N_1895,N_1735);
or U2049 (N_2049,In_1259,In_963);
and U2050 (N_2050,In_129,N_1891);
xor U2051 (N_2051,In_990,N_1725);
and U2052 (N_2052,In_2210,N_1900);
or U2053 (N_2053,In_842,N_1406);
nand U2054 (N_2054,N_824,N_1034);
or U2055 (N_2055,In_2970,In_2997);
or U2056 (N_2056,In_473,N_1733);
nor U2057 (N_2057,N_1774,N_1536);
nand U2058 (N_2058,N_1853,N_346);
nor U2059 (N_2059,N_1974,N_1425);
xor U2060 (N_2060,N_1217,In_65);
nor U2061 (N_2061,N_1938,In_2157);
xnor U2062 (N_2062,N_774,N_1640);
or U2063 (N_2063,N_1797,N_1562);
or U2064 (N_2064,In_2790,N_29);
and U2065 (N_2065,N_1283,In_943);
nor U2066 (N_2066,N_1987,N_1323);
xor U2067 (N_2067,N_1734,N_1780);
nand U2068 (N_2068,In_2222,N_152);
nor U2069 (N_2069,N_1677,N_1611);
or U2070 (N_2070,N_855,N_1995);
nor U2071 (N_2071,N_1652,N_1051);
nand U2072 (N_2072,N_1584,N_120);
nor U2073 (N_2073,In_1895,N_167);
nand U2074 (N_2074,N_1751,N_1972);
and U2075 (N_2075,In_163,N_1598);
xnor U2076 (N_2076,N_1559,N_1593);
nor U2077 (N_2077,N_1671,N_1111);
nand U2078 (N_2078,N_1688,N_1539);
and U2079 (N_2079,N_818,In_1103);
nor U2080 (N_2080,N_1833,N_1880);
and U2081 (N_2081,In_2751,In_2034);
nand U2082 (N_2082,In_539,N_1451);
nor U2083 (N_2083,N_1193,In_249);
xor U2084 (N_2084,N_1232,N_1935);
and U2085 (N_2085,N_1930,N_1816);
and U2086 (N_2086,N_1445,N_1633);
nor U2087 (N_2087,N_1645,In_2772);
xnor U2088 (N_2088,In_1076,N_1786);
nand U2089 (N_2089,N_1907,N_1008);
nor U2090 (N_2090,N_1566,N_1813);
and U2091 (N_2091,N_1664,N_1616);
and U2092 (N_2092,N_1133,N_1522);
nand U2093 (N_2093,N_1739,N_1123);
and U2094 (N_2094,N_1830,N_1027);
nand U2095 (N_2095,N_1519,N_1576);
and U2096 (N_2096,N_1666,N_1796);
nand U2097 (N_2097,N_1828,N_1577);
and U2098 (N_2098,In_2460,N_672);
xnor U2099 (N_2099,In_2220,N_1589);
nand U2100 (N_2100,In_2895,N_1802);
xor U2101 (N_2101,In_1830,In_1852);
xnor U2102 (N_2102,N_236,N_1849);
and U2103 (N_2103,In_259,N_1534);
nor U2104 (N_2104,N_1352,N_1247);
nand U2105 (N_2105,N_1717,N_1989);
nor U2106 (N_2106,N_1151,N_1985);
or U2107 (N_2107,In_125,N_1887);
or U2108 (N_2108,N_1851,In_1129);
nor U2109 (N_2109,N_1837,N_314);
and U2110 (N_2110,N_1698,N_1742);
and U2111 (N_2111,N_1815,N_1722);
xnor U2112 (N_2112,N_1727,N_1948);
nand U2113 (N_2113,N_572,N_1726);
and U2114 (N_2114,N_1771,N_1558);
xor U2115 (N_2115,In_667,N_1682);
nand U2116 (N_2116,In_641,In_2108);
nor U2117 (N_2117,In_379,N_1463);
nor U2118 (N_2118,N_1023,N_1700);
nor U2119 (N_2119,N_1631,N_1591);
and U2120 (N_2120,N_1836,N_1560);
or U2121 (N_2121,N_1934,N_656);
nand U2122 (N_2122,N_1757,In_2422);
and U2123 (N_2123,N_1435,In_268);
xnor U2124 (N_2124,N_1578,N_1075);
nand U2125 (N_2125,N_1745,N_1811);
and U2126 (N_2126,N_1838,N_1601);
nor U2127 (N_2127,In_930,N_771);
nand U2128 (N_2128,N_1037,In_604);
and U2129 (N_2129,N_552,In_728);
nand U2130 (N_2130,N_1791,N_1914);
and U2131 (N_2131,In_1400,N_1737);
or U2132 (N_2132,N_1812,In_1274);
and U2133 (N_2133,In_716,N_1714);
nor U2134 (N_2134,N_1515,N_1081);
xor U2135 (N_2135,N_1809,N_1223);
or U2136 (N_2136,N_1101,N_1969);
xnor U2137 (N_2137,N_1609,N_777);
and U2138 (N_2138,N_1993,N_658);
and U2139 (N_2139,N_1629,N_1661);
nand U2140 (N_2140,N_1850,N_489);
and U2141 (N_2141,N_1627,N_1613);
nor U2142 (N_2142,N_491,In_1920);
nor U2143 (N_2143,N_1632,N_1063);
nand U2144 (N_2144,In_2719,N_1608);
or U2145 (N_2145,N_1856,N_1788);
and U2146 (N_2146,N_1820,N_1546);
and U2147 (N_2147,N_1810,N_44);
nor U2148 (N_2148,In_1675,N_1994);
or U2149 (N_2149,N_1384,N_1792);
xor U2150 (N_2150,N_1628,N_1978);
and U2151 (N_2151,N_1545,N_1841);
nor U2152 (N_2152,N_1940,In_542);
nor U2153 (N_2153,In_2783,N_1620);
xnor U2154 (N_2154,N_519,In_1698);
nand U2155 (N_2155,In_152,N_1520);
or U2156 (N_2156,N_1599,N_1918);
and U2157 (N_2157,In_1873,N_603);
or U2158 (N_2158,N_1210,In_2284);
nand U2159 (N_2159,N_1113,N_1764);
nor U2160 (N_2160,N_828,N_1840);
or U2161 (N_2161,N_1332,N_1922);
and U2162 (N_2162,N_1691,N_97);
nor U2163 (N_2163,N_1381,In_365);
nor U2164 (N_2164,N_1932,In_2346);
xor U2165 (N_2165,N_1871,N_1959);
and U2166 (N_2166,In_572,N_1944);
nand U2167 (N_2167,N_1391,N_1865);
xnor U2168 (N_2168,N_1614,N_1634);
nor U2169 (N_2169,N_1953,N_1926);
xor U2170 (N_2170,N_1681,N_1607);
and U2171 (N_2171,N_1665,N_1073);
or U2172 (N_2172,N_1521,N_1713);
nand U2173 (N_2173,N_1636,N_1135);
nand U2174 (N_2174,In_1942,N_1177);
and U2175 (N_2175,In_2888,In_2960);
nand U2176 (N_2176,N_1673,N_1588);
nor U2177 (N_2177,N_1706,N_1684);
and U2178 (N_2178,N_1956,N_453);
nand U2179 (N_2179,N_1461,N_1299);
and U2180 (N_2180,N_1708,N_229);
and U2181 (N_2181,N_997,N_1540);
and U2182 (N_2182,N_1683,In_232);
nand U2183 (N_2183,In_694,N_1819);
nor U2184 (N_2184,N_1191,N_1997);
nand U2185 (N_2185,N_1421,N_1903);
and U2186 (N_2186,N_1619,In_783);
and U2187 (N_2187,In_985,N_1672);
xor U2188 (N_2188,N_1169,In_459);
nand U2189 (N_2189,N_1219,In_2767);
nand U2190 (N_2190,In_2049,In_1033);
nand U2191 (N_2191,N_1109,N_1687);
nand U2192 (N_2192,In_2746,N_1753);
or U2193 (N_2193,N_1045,N_1468);
nand U2194 (N_2194,N_1762,N_1355);
and U2195 (N_2195,N_1790,N_1596);
and U2196 (N_2196,N_868,N_1966);
and U2197 (N_2197,N_1965,N_1292);
nand U2198 (N_2198,N_1941,N_1756);
xor U2199 (N_2199,In_2058,N_1680);
nand U2200 (N_2200,N_1615,N_1807);
or U2201 (N_2201,N_1585,N_1531);
nand U2202 (N_2202,N_1748,N_973);
xnor U2203 (N_2203,In_2556,N_1138);
nor U2204 (N_2204,N_1523,N_1831);
or U2205 (N_2205,In_2834,N_1862);
or U2206 (N_2206,In_145,N_1984);
nand U2207 (N_2207,N_695,N_1991);
nor U2208 (N_2208,N_1689,N_1486);
nor U2209 (N_2209,In_531,N_737);
nor U2210 (N_2210,N_1744,N_1657);
nor U2211 (N_2211,N_1893,N_1554);
xor U2212 (N_2212,N_1544,N_1676);
or U2213 (N_2213,N_1901,N_1921);
or U2214 (N_2214,N_1505,N_703);
nand U2215 (N_2215,N_1638,N_1517);
xor U2216 (N_2216,N_1525,N_1814);
nand U2217 (N_2217,N_1529,In_1446);
or U2218 (N_2218,In_1335,N_787);
nand U2219 (N_2219,N_1501,N_613);
and U2220 (N_2220,N_1750,N_1317);
xnor U2221 (N_2221,N_1704,N_1335);
and U2222 (N_2222,N_1012,In_1005);
or U2223 (N_2223,N_1765,N_1080);
and U2224 (N_2224,N_1787,In_2515);
or U2225 (N_2225,In_436,N_1042);
nand U2226 (N_2226,In_2181,N_1888);
or U2227 (N_2227,N_666,In_1632);
xnor U2228 (N_2228,N_558,N_1179);
nand U2229 (N_2229,N_669,N_42);
xnor U2230 (N_2230,In_519,N_1761);
or U2231 (N_2231,N_1130,N_1848);
xor U2232 (N_2232,In_621,N_1968);
nor U2233 (N_2233,N_1245,In_2457);
and U2234 (N_2234,N_1749,N_1945);
nor U2235 (N_2235,N_1711,N_1872);
and U2236 (N_2236,N_1526,In_2925);
or U2237 (N_2237,N_1549,N_1879);
and U2238 (N_2238,N_1720,In_2478);
nor U2239 (N_2239,In_517,N_486);
and U2240 (N_2240,In_1520,N_1883);
xor U2241 (N_2241,In_1317,N_1516);
nor U2242 (N_2242,N_1861,N_1597);
xnor U2243 (N_2243,N_1884,N_1970);
nand U2244 (N_2244,N_1707,In_730);
and U2245 (N_2245,In_1214,In_381);
nor U2246 (N_2246,N_1783,N_1119);
or U2247 (N_2247,N_1686,N_1957);
xnor U2248 (N_2248,N_1548,N_1843);
nor U2249 (N_2249,N_1357,In_208);
and U2250 (N_2250,In_2388,N_1079);
nor U2251 (N_2251,In_2947,N_1274);
xnor U2252 (N_2252,N_1469,N_1858);
nand U2253 (N_2253,N_954,In_266);
nand U2254 (N_2254,N_1637,N_1139);
nand U2255 (N_2255,In_2217,N_1919);
and U2256 (N_2256,N_1768,In_2828);
or U2257 (N_2257,N_935,N_1386);
nor U2258 (N_2258,N_122,In_160);
nand U2259 (N_2259,N_1679,In_124);
nand U2260 (N_2260,N_1530,N_1286);
or U2261 (N_2261,N_1936,N_1656);
xnor U2262 (N_2262,N_1905,N_1669);
xor U2263 (N_2263,N_1759,N_1587);
or U2264 (N_2264,In_1908,N_1571);
or U2265 (N_2265,N_1822,N_1776);
xnor U2266 (N_2266,In_1840,N_1775);
nor U2267 (N_2267,N_628,N_1954);
xor U2268 (N_2268,N_1600,N_1927);
xnor U2269 (N_2269,N_1860,N_1847);
or U2270 (N_2270,N_1869,N_1649);
or U2271 (N_2271,N_1804,N_1575);
or U2272 (N_2272,N_518,In_2447);
xnor U2273 (N_2273,N_1102,N_665);
nand U2274 (N_2274,N_1031,N_1892);
xnor U2275 (N_2275,N_1651,N_1692);
nor U2276 (N_2276,N_1583,N_1939);
nor U2277 (N_2277,N_1962,In_331);
xnor U2278 (N_2278,N_1393,N_1373);
or U2279 (N_2279,In_2252,N_1569);
nor U2280 (N_2280,N_539,N_1947);
xnor U2281 (N_2281,In_2405,N_1370);
and U2282 (N_2282,In_1846,N_1532);
or U2283 (N_2283,N_405,N_1612);
or U2284 (N_2284,N_1998,N_1781);
or U2285 (N_2285,In_345,In_918);
or U2286 (N_2286,N_1902,N_1886);
nor U2287 (N_2287,N_1715,In_1832);
nor U2288 (N_2288,N_1602,N_1743);
xnor U2289 (N_2289,N_289,N_1875);
and U2290 (N_2290,N_1496,N_583);
nand U2291 (N_2291,N_897,In_2706);
and U2292 (N_2292,N_1980,In_831);
xnor U2293 (N_2293,N_1773,In_2015);
xnor U2294 (N_2294,N_1946,N_1794);
nand U2295 (N_2295,N_1789,N_650);
nand U2296 (N_2296,N_1625,N_1437);
nand U2297 (N_2297,N_1963,N_1710);
nor U2298 (N_2298,In_2668,N_846);
and U2299 (N_2299,In_1916,N_1732);
and U2300 (N_2300,N_1477,In_256);
or U2301 (N_2301,In_2497,In_180);
xnor U2302 (N_2302,N_987,N_1173);
or U2303 (N_2303,N_1333,N_1982);
nand U2304 (N_2304,N_293,N_1988);
nor U2305 (N_2305,N_1857,N_1670);
nand U2306 (N_2306,N_1910,N_1923);
nand U2307 (N_2307,In_1119,N_1882);
nand U2308 (N_2308,In_2806,In_2627);
nor U2309 (N_2309,N_1695,N_1785);
nor U2310 (N_2310,N_1912,N_1618);
xnor U2311 (N_2311,N_1699,N_788);
xnor U2312 (N_2312,N_726,N_1313);
nand U2313 (N_2313,N_1897,N_1091);
nand U2314 (N_2314,N_481,N_770);
nor U2315 (N_2315,N_1071,N_789);
nor U2316 (N_2316,N_1979,N_1890);
nand U2317 (N_2317,N_998,In_1348);
and U2318 (N_2318,N_288,In_2470);
xnor U2319 (N_2319,In_1295,In_1825);
xnor U2320 (N_2320,In_1322,In_2135);
nand U2321 (N_2321,N_1842,N_1604);
or U2322 (N_2322,N_1586,N_1741);
nand U2323 (N_2323,N_1770,N_1535);
nand U2324 (N_2324,In_42,N_1158);
nand U2325 (N_2325,In_1749,N_1458);
or U2326 (N_2326,N_148,N_1777);
nand U2327 (N_2327,N_1873,In_462);
or U2328 (N_2328,N_1093,In_524);
nor U2329 (N_2329,In_1332,N_985);
xnor U2330 (N_2330,In_109,N_1769);
and U2331 (N_2331,N_1555,In_2857);
xnor U2332 (N_2332,N_1996,In_137);
xnor U2333 (N_2333,N_232,N_1503);
nor U2334 (N_2334,In_1471,In_1388);
xnor U2335 (N_2335,N_1758,N_1552);
nand U2336 (N_2336,N_1967,N_1876);
and U2337 (N_2337,N_1024,N_1288);
nor U2338 (N_2338,N_1878,In_2526);
nor U2339 (N_2339,N_1663,In_1242);
xor U2340 (N_2340,N_1226,N_1307);
nor U2341 (N_2341,In_1161,N_1977);
nand U2342 (N_2342,In_713,N_39);
and U2343 (N_2343,N_1230,N_1702);
nor U2344 (N_2344,In_999,N_1301);
nand U2345 (N_2345,N_1234,In_283);
nor U2346 (N_2346,N_1798,N_1846);
nor U2347 (N_2347,N_599,N_1990);
and U2348 (N_2348,N_1958,N_1844);
or U2349 (N_2349,N_617,In_1141);
and U2350 (N_2350,N_1662,N_1278);
xor U2351 (N_2351,N_1674,N_1975);
and U2352 (N_2352,N_1971,N_844);
nor U2353 (N_2353,In_2472,N_1622);
nand U2354 (N_2354,N_1808,N_1358);
xor U2355 (N_2355,In_70,In_2320);
xnor U2356 (N_2356,In_7,N_797);
nor U2357 (N_2357,N_1675,N_1510);
nor U2358 (N_2358,N_1800,N_798);
nor U2359 (N_2359,N_1538,N_1915);
or U2360 (N_2360,N_1942,N_865);
and U2361 (N_2361,N_1164,In_2685);
and U2362 (N_2362,N_1513,N_1795);
or U2363 (N_2363,N_1855,In_2029);
and U2364 (N_2364,N_1547,In_568);
nand U2365 (N_2365,N_1986,N_1668);
nand U2366 (N_2366,In_2517,In_390);
nand U2367 (N_2367,N_1712,N_1647);
nand U2368 (N_2368,N_1655,N_1899);
and U2369 (N_2369,N_763,N_1806);
or U2370 (N_2370,In_1894,N_636);
nor U2371 (N_2371,In_451,In_2074);
xor U2372 (N_2372,N_169,In_1389);
and U2373 (N_2373,N_1693,In_2588);
nor U2374 (N_2374,In_486,N_1983);
nand U2375 (N_2375,N_1731,N_578);
nor U2376 (N_2376,N_1580,In_911);
or U2377 (N_2377,N_1999,N_1736);
and U2378 (N_2378,N_1572,N_1541);
nor U2379 (N_2379,In_865,N_1730);
nand U2380 (N_2380,N_1964,N_1874);
nand U2381 (N_2381,N_1754,N_1658);
and U2382 (N_2382,N_335,N_1747);
xnor U2383 (N_2383,N_1507,N_1778);
or U2384 (N_2384,N_992,N_1509);
nand U2385 (N_2385,N_1500,In_118);
nor U2386 (N_2386,In_2197,N_1561);
nand U2387 (N_2387,N_1524,N_1924);
nor U2388 (N_2388,N_1818,N_1565);
nor U2389 (N_2389,N_1643,N_1502);
nor U2390 (N_2390,N_1937,N_683);
and U2391 (N_2391,N_1803,In_856);
xor U2392 (N_2392,N_1976,N_1563);
xor U2393 (N_2393,N_1925,N_1035);
and U2394 (N_2394,N_1824,N_1533);
and U2395 (N_2395,N_1376,N_1261);
or U2396 (N_2396,N_1913,N_1906);
nor U2397 (N_2397,N_1568,N_1107);
nand U2398 (N_2398,N_1949,In_1590);
nand U2399 (N_2399,In_1754,In_1804);
xnor U2400 (N_2400,In_2714,N_181);
nand U2401 (N_2401,N_1624,In_2146);
nor U2402 (N_2402,N_1904,N_1779);
or U2403 (N_2403,N_1573,N_185);
xor U2404 (N_2404,N_1551,N_260);
nor U2405 (N_2405,N_1650,In_262);
and U2406 (N_2406,N_1885,N_563);
nand U2407 (N_2407,N_1694,In_2518);
and U2408 (N_2408,In_2359,N_1973);
nand U2409 (N_2409,In_2661,N_1553);
or U2410 (N_2410,N_1308,N_890);
or U2411 (N_2411,N_569,N_1623);
nand U2412 (N_2412,N_424,N_1961);
nor U2413 (N_2413,In_1776,N_1678);
and U2414 (N_2414,N_1617,N_1867);
nor U2415 (N_2415,N_1642,In_1574);
and U2416 (N_2416,N_1845,In_101);
xor U2417 (N_2417,N_1827,N_1450);
nor U2418 (N_2418,N_1782,In_216);
nand U2419 (N_2419,N_1767,N_1854);
or U2420 (N_2420,N_1909,In_2256);
xnor U2421 (N_2421,In_1495,N_1504);
xor U2422 (N_2422,In_2499,N_1784);
nand U2423 (N_2423,N_1359,N_1896);
and U2424 (N_2424,In_327,N_96);
nand U2425 (N_2425,N_1154,N_1723);
nor U2426 (N_2426,N_1165,N_1582);
xor U2427 (N_2427,N_1606,N_1168);
nand U2428 (N_2428,In_745,N_1258);
nor U2429 (N_2429,N_1839,N_1567);
nand U2430 (N_2430,N_1929,N_1870);
and U2431 (N_2431,In_2954,In_1674);
xnor U2432 (N_2432,N_1928,N_1859);
and U2433 (N_2433,N_905,In_1843);
xnor U2434 (N_2434,N_1550,N_1868);
and U2435 (N_2435,N_1917,N_1889);
or U2436 (N_2436,N_1933,In_2487);
or U2437 (N_2437,N_1092,N_1330);
and U2438 (N_2438,N_1297,N_1508);
nand U2439 (N_2439,N_676,N_104);
xnor U2440 (N_2440,N_1408,N_682);
nand U2441 (N_2441,N_1527,In_1926);
or U2442 (N_2442,N_1302,N_1752);
or U2443 (N_2443,N_1719,In_1492);
or U2444 (N_2444,N_1952,N_1835);
and U2445 (N_2445,N_161,In_764);
nor U2446 (N_2446,N_1574,In_2326);
nor U2447 (N_2447,N_1579,N_1644);
or U2448 (N_2448,N_1920,N_794);
nor U2449 (N_2449,N_1697,N_1821);
nor U2450 (N_2450,N_1312,N_1916);
nor U2451 (N_2451,In_2244,N_1801);
and U2452 (N_2452,N_1898,N_857);
xor U2453 (N_2453,In_1773,N_1877);
and U2454 (N_2454,N_1581,N_1724);
xnor U2455 (N_2455,In_166,N_1696);
xor U2456 (N_2456,N_1511,In_2580);
and U2457 (N_2457,N_1943,N_1826);
or U2458 (N_2458,In_1464,N_804);
xnor U2459 (N_2459,N_1090,In_413);
nor U2460 (N_2460,In_756,In_81);
nand U2461 (N_2461,N_1817,In_1334);
and U2462 (N_2462,In_2208,In_2026);
nand U2463 (N_2463,N_1621,N_1703);
xnor U2464 (N_2464,In_1529,In_88);
nor U2465 (N_2465,In_2409,N_1104);
or U2466 (N_2466,N_959,In_2675);
nor U2467 (N_2467,N_806,N_1660);
and U2468 (N_2468,N_1992,In_2868);
nand U2469 (N_2469,N_1718,N_1556);
nor U2470 (N_2470,In_1950,In_229);
nor U2471 (N_2471,N_1497,N_1564);
or U2472 (N_2472,N_1931,N_1429);
and U2473 (N_2473,N_1630,In_1626);
or U2474 (N_2474,In_1028,N_1881);
xnor U2475 (N_2475,N_1295,N_1960);
and U2476 (N_2476,N_1096,N_1290);
or U2477 (N_2477,N_1250,N_1760);
nor U2478 (N_2478,N_1103,In_2853);
nor U2479 (N_2479,N_1829,N_164);
and U2480 (N_2480,N_1825,N_273);
nor U2481 (N_2481,In_833,In_1610);
or U2482 (N_2482,N_1793,N_1763);
nor U2483 (N_2483,N_1202,In_1105);
nand U2484 (N_2484,N_972,N_1653);
nor U2485 (N_2485,N_1453,N_1595);
and U2486 (N_2486,In_1419,N_1950);
nor U2487 (N_2487,N_687,N_287);
nor U2488 (N_2488,In_1233,N_1908);
xnor U2489 (N_2489,N_1654,N_1755);
or U2490 (N_2490,In_449,N_724);
xor U2491 (N_2491,In_625,N_1603);
xnor U2492 (N_2492,N_1159,In_2092);
nand U2493 (N_2493,N_931,N_1659);
xor U2494 (N_2494,In_752,N_1364);
and U2495 (N_2495,N_1701,N_1462);
or U2496 (N_2496,N_1805,N_1646);
nand U2497 (N_2497,N_1626,N_1729);
or U2498 (N_2498,N_1721,N_1422);
xor U2499 (N_2499,N_769,N_1772);
and U2500 (N_2500,N_2153,N_2365);
or U2501 (N_2501,N_2151,N_2064);
or U2502 (N_2502,N_2412,N_2070);
nand U2503 (N_2503,N_2321,N_2095);
xnor U2504 (N_2504,N_2167,N_2319);
and U2505 (N_2505,N_2189,N_2004);
and U2506 (N_2506,N_2139,N_2376);
or U2507 (N_2507,N_2446,N_2245);
nand U2508 (N_2508,N_2377,N_2201);
and U2509 (N_2509,N_2127,N_2261);
and U2510 (N_2510,N_2003,N_2390);
nor U2511 (N_2511,N_2340,N_2356);
xor U2512 (N_2512,N_2330,N_2031);
nor U2513 (N_2513,N_2076,N_2318);
nor U2514 (N_2514,N_2388,N_2483);
nor U2515 (N_2515,N_2293,N_2072);
xor U2516 (N_2516,N_2056,N_2424);
xnor U2517 (N_2517,N_2244,N_2240);
and U2518 (N_2518,N_2401,N_2339);
xor U2519 (N_2519,N_2152,N_2270);
or U2520 (N_2520,N_2267,N_2202);
or U2521 (N_2521,N_2198,N_2173);
nor U2522 (N_2522,N_2287,N_2096);
xnor U2523 (N_2523,N_2374,N_2456);
or U2524 (N_2524,N_2392,N_2482);
xnor U2525 (N_2525,N_2180,N_2233);
xnor U2526 (N_2526,N_2241,N_2498);
nand U2527 (N_2527,N_2486,N_2414);
nor U2528 (N_2528,N_2302,N_2348);
nor U2529 (N_2529,N_2308,N_2309);
or U2530 (N_2530,N_2024,N_2025);
nor U2531 (N_2531,N_2272,N_2419);
nor U2532 (N_2532,N_2493,N_2022);
nand U2533 (N_2533,N_2214,N_2236);
and U2534 (N_2534,N_2389,N_2200);
or U2535 (N_2535,N_2289,N_2310);
nor U2536 (N_2536,N_2185,N_2145);
and U2537 (N_2537,N_2147,N_2366);
nor U2538 (N_2538,N_2435,N_2011);
and U2539 (N_2539,N_2226,N_2393);
nor U2540 (N_2540,N_2301,N_2122);
or U2541 (N_2541,N_2438,N_2476);
xnor U2542 (N_2542,N_2051,N_2161);
nor U2543 (N_2543,N_2457,N_2114);
or U2544 (N_2544,N_2285,N_2124);
xor U2545 (N_2545,N_2146,N_2186);
and U2546 (N_2546,N_2409,N_2229);
nand U2547 (N_2547,N_2094,N_2162);
or U2548 (N_2548,N_2361,N_2450);
nor U2549 (N_2549,N_2039,N_2008);
or U2550 (N_2550,N_2467,N_2074);
nand U2551 (N_2551,N_2192,N_2363);
nor U2552 (N_2552,N_2194,N_2280);
nand U2553 (N_2553,N_2172,N_2313);
and U2554 (N_2554,N_2397,N_2341);
and U2555 (N_2555,N_2026,N_2141);
xnor U2556 (N_2556,N_2281,N_2158);
xnor U2557 (N_2557,N_2480,N_2005);
xnor U2558 (N_2558,N_2081,N_2043);
or U2559 (N_2559,N_2085,N_2378);
xor U2560 (N_2560,N_2357,N_2045);
and U2561 (N_2561,N_2443,N_2234);
xor U2562 (N_2562,N_2451,N_2336);
nand U2563 (N_2563,N_2243,N_2209);
and U2564 (N_2564,N_2355,N_2322);
or U2565 (N_2565,N_2274,N_2461);
or U2566 (N_2566,N_2103,N_2454);
or U2567 (N_2567,N_2265,N_2118);
nor U2568 (N_2568,N_2406,N_2468);
nor U2569 (N_2569,N_2324,N_2297);
and U2570 (N_2570,N_2104,N_2106);
xnor U2571 (N_2571,N_2110,N_2163);
nor U2572 (N_2572,N_2354,N_2065);
nand U2573 (N_2573,N_2246,N_2231);
xor U2574 (N_2574,N_2271,N_2235);
or U2575 (N_2575,N_2009,N_2062);
xnor U2576 (N_2576,N_2120,N_2463);
or U2577 (N_2577,N_2266,N_2166);
and U2578 (N_2578,N_2320,N_2040);
and U2579 (N_2579,N_2396,N_2416);
nand U2580 (N_2580,N_2448,N_2442);
nand U2581 (N_2581,N_2349,N_2394);
nor U2582 (N_2582,N_2328,N_2023);
or U2583 (N_2583,N_2470,N_2108);
nand U2584 (N_2584,N_2429,N_2237);
xnor U2585 (N_2585,N_2155,N_2410);
nor U2586 (N_2586,N_2333,N_2387);
and U2587 (N_2587,N_2427,N_2052);
nor U2588 (N_2588,N_2405,N_2013);
and U2589 (N_2589,N_2351,N_2206);
nand U2590 (N_2590,N_2136,N_2216);
or U2591 (N_2591,N_2224,N_2259);
and U2592 (N_2592,N_2487,N_2380);
nor U2593 (N_2593,N_2441,N_2307);
or U2594 (N_2594,N_2137,N_2431);
xor U2595 (N_2595,N_2303,N_2421);
nand U2596 (N_2596,N_2217,N_2256);
nand U2597 (N_2597,N_2129,N_2090);
nor U2598 (N_2598,N_2275,N_2042);
nor U2599 (N_2599,N_2312,N_2165);
nor U2600 (N_2600,N_2458,N_2157);
or U2601 (N_2601,N_2375,N_2176);
and U2602 (N_2602,N_2174,N_2057);
nand U2603 (N_2603,N_2208,N_2107);
or U2604 (N_2604,N_2082,N_2006);
and U2605 (N_2605,N_2097,N_2218);
xor U2606 (N_2606,N_2197,N_2038);
nand U2607 (N_2607,N_2087,N_2046);
nand U2608 (N_2608,N_2168,N_2179);
xnor U2609 (N_2609,N_2315,N_2247);
xor U2610 (N_2610,N_2425,N_2213);
nand U2611 (N_2611,N_2418,N_2131);
or U2612 (N_2612,N_2286,N_2019);
nand U2613 (N_2613,N_2092,N_2283);
nor U2614 (N_2614,N_2292,N_2210);
xnor U2615 (N_2615,N_2299,N_2066);
or U2616 (N_2616,N_2230,N_2050);
nor U2617 (N_2617,N_2171,N_2358);
and U2618 (N_2618,N_2036,N_2135);
nand U2619 (N_2619,N_2379,N_2386);
xnor U2620 (N_2620,N_2196,N_2170);
nor U2621 (N_2621,N_2191,N_2282);
and U2622 (N_2622,N_2495,N_2086);
and U2623 (N_2623,N_2071,N_2221);
or U2624 (N_2624,N_2277,N_2284);
and U2625 (N_2625,N_2462,N_2227);
and U2626 (N_2626,N_2187,N_2496);
or U2627 (N_2627,N_2228,N_2437);
nor U2628 (N_2628,N_2212,N_2353);
xnor U2629 (N_2629,N_2053,N_2400);
xor U2630 (N_2630,N_2116,N_2183);
or U2631 (N_2631,N_2475,N_2089);
and U2632 (N_2632,N_2474,N_2058);
nor U2633 (N_2633,N_2128,N_2238);
xnor U2634 (N_2634,N_2012,N_2102);
nor U2635 (N_2635,N_2035,N_2422);
xor U2636 (N_2636,N_2403,N_2203);
and U2637 (N_2637,N_2121,N_2294);
nor U2638 (N_2638,N_2338,N_2133);
nor U2639 (N_2639,N_2250,N_2258);
and U2640 (N_2640,N_2232,N_2331);
nor U2641 (N_2641,N_2477,N_2337);
nor U2642 (N_2642,N_2059,N_2073);
nand U2643 (N_2643,N_2304,N_2132);
nor U2644 (N_2644,N_2002,N_2264);
or U2645 (N_2645,N_2060,N_2014);
nand U2646 (N_2646,N_2269,N_2178);
nand U2647 (N_2647,N_2175,N_2067);
nand U2648 (N_2648,N_2248,N_2188);
xor U2649 (N_2649,N_2150,N_2385);
or U2650 (N_2650,N_2117,N_2344);
nand U2651 (N_2651,N_2242,N_2222);
nor U2652 (N_2652,N_2316,N_2466);
nor U2653 (N_2653,N_2260,N_2027);
xor U2654 (N_2654,N_2098,N_2279);
nor U2655 (N_2655,N_2001,N_2408);
nand U2656 (N_2656,N_2220,N_2453);
nand U2657 (N_2657,N_2300,N_2000);
or U2658 (N_2658,N_2395,N_2345);
xor U2659 (N_2659,N_2054,N_2428);
nor U2660 (N_2660,N_2449,N_2148);
nand U2661 (N_2661,N_2413,N_2257);
nand U2662 (N_2662,N_2335,N_2478);
and U2663 (N_2663,N_2119,N_2373);
and U2664 (N_2664,N_2254,N_2473);
nor U2665 (N_2665,N_2219,N_2112);
and U2666 (N_2666,N_2350,N_2306);
and U2667 (N_2667,N_2015,N_2360);
xnor U2668 (N_2668,N_2491,N_2055);
nor U2669 (N_2669,N_2382,N_2077);
nand U2670 (N_2670,N_2204,N_2033);
and U2671 (N_2671,N_2069,N_2342);
nand U2672 (N_2672,N_2314,N_2367);
xnor U2673 (N_2673,N_2100,N_2016);
or U2674 (N_2674,N_2079,N_2126);
and U2675 (N_2675,N_2317,N_2044);
nand U2676 (N_2676,N_2346,N_2370);
and U2677 (N_2677,N_2488,N_2445);
xnor U2678 (N_2678,N_2099,N_2489);
nand U2679 (N_2679,N_2490,N_2193);
nand U2680 (N_2680,N_2426,N_2369);
or U2681 (N_2681,N_2195,N_2075);
nand U2682 (N_2682,N_2472,N_2326);
nand U2683 (N_2683,N_2215,N_2091);
nor U2684 (N_2684,N_2452,N_2464);
xor U2685 (N_2685,N_2372,N_2383);
xor U2686 (N_2686,N_2364,N_2391);
and U2687 (N_2687,N_2113,N_2199);
nand U2688 (N_2688,N_2068,N_2130);
xor U2689 (N_2689,N_2381,N_2497);
and U2690 (N_2690,N_2177,N_2253);
nand U2691 (N_2691,N_2434,N_2362);
nor U2692 (N_2692,N_2049,N_2290);
or U2693 (N_2693,N_2423,N_2327);
xor U2694 (N_2694,N_2115,N_2455);
nand U2695 (N_2695,N_2417,N_2430);
and U2696 (N_2696,N_2138,N_2469);
nand U2697 (N_2697,N_2268,N_2494);
or U2698 (N_2698,N_2063,N_2021);
and U2699 (N_2699,N_2190,N_2154);
nand U2700 (N_2700,N_2276,N_2211);
nor U2701 (N_2701,N_2255,N_2399);
xnor U2702 (N_2702,N_2048,N_2447);
nor U2703 (N_2703,N_2111,N_2205);
xnor U2704 (N_2704,N_2288,N_2420);
or U2705 (N_2705,N_2278,N_2239);
xnor U2706 (N_2706,N_2439,N_2143);
xnor U2707 (N_2707,N_2088,N_2444);
nor U2708 (N_2708,N_2018,N_2252);
nor U2709 (N_2709,N_2037,N_2325);
or U2710 (N_2710,N_2465,N_2010);
or U2711 (N_2711,N_2140,N_2007);
xnor U2712 (N_2712,N_2144,N_2471);
xor U2713 (N_2713,N_2169,N_2332);
or U2714 (N_2714,N_2134,N_2142);
or U2715 (N_2715,N_2029,N_2123);
or U2716 (N_2716,N_2017,N_2415);
nand U2717 (N_2717,N_2305,N_2273);
or U2718 (N_2718,N_2343,N_2160);
and U2719 (N_2719,N_2291,N_2028);
and U2720 (N_2720,N_2436,N_2311);
and U2721 (N_2721,N_2459,N_2384);
nand U2722 (N_2722,N_2298,N_2371);
and U2723 (N_2723,N_2078,N_2156);
and U2724 (N_2724,N_2433,N_2251);
xnor U2725 (N_2725,N_2398,N_2105);
nand U2726 (N_2726,N_2223,N_2484);
nand U2727 (N_2727,N_2432,N_2149);
or U2728 (N_2728,N_2485,N_2184);
xnor U2729 (N_2729,N_2347,N_2359);
or U2730 (N_2730,N_2499,N_2352);
xor U2731 (N_2731,N_2479,N_2323);
nand U2732 (N_2732,N_2101,N_2034);
and U2733 (N_2733,N_2492,N_2407);
nand U2734 (N_2734,N_2411,N_2020);
and U2735 (N_2735,N_2249,N_2030);
nor U2736 (N_2736,N_2368,N_2262);
nor U2737 (N_2737,N_2181,N_2225);
or U2738 (N_2738,N_2125,N_2080);
and U2739 (N_2739,N_2159,N_2296);
or U2740 (N_2740,N_2207,N_2093);
or U2741 (N_2741,N_2041,N_2164);
and U2742 (N_2742,N_2334,N_2295);
or U2743 (N_2743,N_2263,N_2402);
xor U2744 (N_2744,N_2404,N_2084);
nor U2745 (N_2745,N_2061,N_2109);
nor U2746 (N_2746,N_2047,N_2083);
nor U2747 (N_2747,N_2460,N_2032);
or U2748 (N_2748,N_2182,N_2440);
nand U2749 (N_2749,N_2329,N_2481);
nor U2750 (N_2750,N_2273,N_2264);
nor U2751 (N_2751,N_2435,N_2275);
and U2752 (N_2752,N_2156,N_2030);
xnor U2753 (N_2753,N_2015,N_2070);
and U2754 (N_2754,N_2167,N_2499);
xnor U2755 (N_2755,N_2360,N_2120);
and U2756 (N_2756,N_2168,N_2264);
xnor U2757 (N_2757,N_2269,N_2306);
and U2758 (N_2758,N_2452,N_2340);
xor U2759 (N_2759,N_2312,N_2399);
nand U2760 (N_2760,N_2313,N_2049);
nand U2761 (N_2761,N_2027,N_2449);
nand U2762 (N_2762,N_2464,N_2148);
or U2763 (N_2763,N_2061,N_2253);
xnor U2764 (N_2764,N_2010,N_2222);
and U2765 (N_2765,N_2187,N_2333);
nor U2766 (N_2766,N_2486,N_2094);
or U2767 (N_2767,N_2165,N_2168);
xnor U2768 (N_2768,N_2309,N_2206);
xor U2769 (N_2769,N_2395,N_2411);
xnor U2770 (N_2770,N_2424,N_2183);
nand U2771 (N_2771,N_2125,N_2017);
xor U2772 (N_2772,N_2097,N_2447);
and U2773 (N_2773,N_2199,N_2055);
xor U2774 (N_2774,N_2201,N_2338);
nor U2775 (N_2775,N_2427,N_2273);
xor U2776 (N_2776,N_2097,N_2125);
and U2777 (N_2777,N_2130,N_2054);
or U2778 (N_2778,N_2246,N_2152);
nand U2779 (N_2779,N_2332,N_2096);
nor U2780 (N_2780,N_2345,N_2408);
and U2781 (N_2781,N_2223,N_2340);
nor U2782 (N_2782,N_2039,N_2478);
and U2783 (N_2783,N_2073,N_2365);
xnor U2784 (N_2784,N_2377,N_2417);
or U2785 (N_2785,N_2205,N_2441);
nor U2786 (N_2786,N_2021,N_2142);
xor U2787 (N_2787,N_2413,N_2061);
and U2788 (N_2788,N_2464,N_2322);
xnor U2789 (N_2789,N_2268,N_2478);
xnor U2790 (N_2790,N_2375,N_2429);
or U2791 (N_2791,N_2143,N_2205);
xnor U2792 (N_2792,N_2399,N_2343);
and U2793 (N_2793,N_2041,N_2371);
nor U2794 (N_2794,N_2175,N_2472);
and U2795 (N_2795,N_2391,N_2491);
and U2796 (N_2796,N_2413,N_2094);
or U2797 (N_2797,N_2259,N_2324);
nand U2798 (N_2798,N_2118,N_2315);
nand U2799 (N_2799,N_2068,N_2102);
nor U2800 (N_2800,N_2115,N_2236);
and U2801 (N_2801,N_2476,N_2122);
xnor U2802 (N_2802,N_2496,N_2164);
and U2803 (N_2803,N_2192,N_2449);
nor U2804 (N_2804,N_2450,N_2449);
nor U2805 (N_2805,N_2474,N_2243);
nor U2806 (N_2806,N_2246,N_2177);
nor U2807 (N_2807,N_2145,N_2242);
nor U2808 (N_2808,N_2254,N_2093);
and U2809 (N_2809,N_2443,N_2207);
nand U2810 (N_2810,N_2222,N_2040);
or U2811 (N_2811,N_2189,N_2110);
and U2812 (N_2812,N_2122,N_2436);
or U2813 (N_2813,N_2369,N_2477);
and U2814 (N_2814,N_2252,N_2262);
nand U2815 (N_2815,N_2102,N_2420);
nand U2816 (N_2816,N_2438,N_2152);
nor U2817 (N_2817,N_2446,N_2207);
nor U2818 (N_2818,N_2093,N_2436);
and U2819 (N_2819,N_2061,N_2224);
and U2820 (N_2820,N_2006,N_2245);
nand U2821 (N_2821,N_2359,N_2313);
nand U2822 (N_2822,N_2469,N_2012);
and U2823 (N_2823,N_2123,N_2214);
nor U2824 (N_2824,N_2125,N_2106);
or U2825 (N_2825,N_2128,N_2039);
nand U2826 (N_2826,N_2337,N_2466);
nand U2827 (N_2827,N_2205,N_2157);
or U2828 (N_2828,N_2382,N_2179);
nand U2829 (N_2829,N_2396,N_2310);
and U2830 (N_2830,N_2422,N_2009);
nand U2831 (N_2831,N_2388,N_2460);
or U2832 (N_2832,N_2203,N_2264);
nor U2833 (N_2833,N_2154,N_2278);
or U2834 (N_2834,N_2377,N_2172);
xor U2835 (N_2835,N_2065,N_2463);
nor U2836 (N_2836,N_2288,N_2043);
xor U2837 (N_2837,N_2434,N_2150);
nand U2838 (N_2838,N_2192,N_2372);
and U2839 (N_2839,N_2056,N_2085);
xnor U2840 (N_2840,N_2465,N_2014);
or U2841 (N_2841,N_2311,N_2094);
and U2842 (N_2842,N_2200,N_2260);
nand U2843 (N_2843,N_2155,N_2178);
and U2844 (N_2844,N_2121,N_2434);
and U2845 (N_2845,N_2080,N_2324);
xor U2846 (N_2846,N_2344,N_2494);
xnor U2847 (N_2847,N_2209,N_2382);
or U2848 (N_2848,N_2163,N_2087);
nor U2849 (N_2849,N_2398,N_2385);
or U2850 (N_2850,N_2113,N_2394);
nand U2851 (N_2851,N_2395,N_2313);
or U2852 (N_2852,N_2379,N_2415);
nor U2853 (N_2853,N_2434,N_2016);
or U2854 (N_2854,N_2205,N_2319);
xnor U2855 (N_2855,N_2011,N_2297);
or U2856 (N_2856,N_2149,N_2164);
nand U2857 (N_2857,N_2223,N_2088);
or U2858 (N_2858,N_2420,N_2116);
xor U2859 (N_2859,N_2057,N_2405);
and U2860 (N_2860,N_2029,N_2226);
xnor U2861 (N_2861,N_2176,N_2050);
nor U2862 (N_2862,N_2324,N_2206);
or U2863 (N_2863,N_2296,N_2185);
nand U2864 (N_2864,N_2147,N_2050);
nand U2865 (N_2865,N_2121,N_2298);
nand U2866 (N_2866,N_2008,N_2037);
or U2867 (N_2867,N_2406,N_2499);
xor U2868 (N_2868,N_2446,N_2084);
nand U2869 (N_2869,N_2269,N_2272);
xnor U2870 (N_2870,N_2400,N_2471);
nand U2871 (N_2871,N_2452,N_2300);
xnor U2872 (N_2872,N_2163,N_2093);
and U2873 (N_2873,N_2212,N_2032);
nand U2874 (N_2874,N_2256,N_2163);
nor U2875 (N_2875,N_2058,N_2366);
nor U2876 (N_2876,N_2116,N_2144);
xnor U2877 (N_2877,N_2273,N_2477);
and U2878 (N_2878,N_2366,N_2360);
nor U2879 (N_2879,N_2419,N_2453);
nor U2880 (N_2880,N_2382,N_2161);
or U2881 (N_2881,N_2463,N_2492);
or U2882 (N_2882,N_2463,N_2330);
nand U2883 (N_2883,N_2344,N_2499);
nor U2884 (N_2884,N_2193,N_2277);
nor U2885 (N_2885,N_2029,N_2052);
nand U2886 (N_2886,N_2373,N_2084);
or U2887 (N_2887,N_2424,N_2067);
xnor U2888 (N_2888,N_2029,N_2165);
nor U2889 (N_2889,N_2232,N_2293);
nand U2890 (N_2890,N_2097,N_2343);
nor U2891 (N_2891,N_2097,N_2242);
nand U2892 (N_2892,N_2065,N_2243);
xnor U2893 (N_2893,N_2057,N_2256);
or U2894 (N_2894,N_2450,N_2247);
or U2895 (N_2895,N_2352,N_2011);
or U2896 (N_2896,N_2210,N_2455);
nor U2897 (N_2897,N_2111,N_2092);
nand U2898 (N_2898,N_2178,N_2307);
xnor U2899 (N_2899,N_2208,N_2287);
and U2900 (N_2900,N_2267,N_2163);
xor U2901 (N_2901,N_2431,N_2129);
xnor U2902 (N_2902,N_2472,N_2487);
nor U2903 (N_2903,N_2025,N_2135);
nor U2904 (N_2904,N_2235,N_2448);
or U2905 (N_2905,N_2015,N_2364);
xor U2906 (N_2906,N_2444,N_2208);
nand U2907 (N_2907,N_2121,N_2023);
nand U2908 (N_2908,N_2330,N_2234);
xnor U2909 (N_2909,N_2090,N_2377);
and U2910 (N_2910,N_2337,N_2327);
xnor U2911 (N_2911,N_2249,N_2495);
and U2912 (N_2912,N_2426,N_2189);
xor U2913 (N_2913,N_2175,N_2215);
or U2914 (N_2914,N_2488,N_2299);
and U2915 (N_2915,N_2046,N_2316);
xor U2916 (N_2916,N_2456,N_2218);
and U2917 (N_2917,N_2204,N_2471);
nand U2918 (N_2918,N_2450,N_2195);
or U2919 (N_2919,N_2490,N_2083);
nor U2920 (N_2920,N_2257,N_2429);
xor U2921 (N_2921,N_2270,N_2188);
nand U2922 (N_2922,N_2051,N_2154);
xnor U2923 (N_2923,N_2366,N_2182);
or U2924 (N_2924,N_2268,N_2486);
xnor U2925 (N_2925,N_2421,N_2096);
or U2926 (N_2926,N_2480,N_2414);
nor U2927 (N_2927,N_2216,N_2497);
xor U2928 (N_2928,N_2192,N_2180);
or U2929 (N_2929,N_2150,N_2214);
and U2930 (N_2930,N_2470,N_2308);
or U2931 (N_2931,N_2295,N_2310);
nand U2932 (N_2932,N_2423,N_2138);
nand U2933 (N_2933,N_2018,N_2297);
nand U2934 (N_2934,N_2247,N_2106);
nor U2935 (N_2935,N_2209,N_2128);
xor U2936 (N_2936,N_2289,N_2161);
and U2937 (N_2937,N_2366,N_2416);
nand U2938 (N_2938,N_2003,N_2122);
or U2939 (N_2939,N_2071,N_2385);
nand U2940 (N_2940,N_2195,N_2287);
nor U2941 (N_2941,N_2402,N_2400);
xor U2942 (N_2942,N_2300,N_2066);
or U2943 (N_2943,N_2197,N_2292);
or U2944 (N_2944,N_2011,N_2245);
xnor U2945 (N_2945,N_2355,N_2459);
xnor U2946 (N_2946,N_2463,N_2036);
and U2947 (N_2947,N_2164,N_2195);
and U2948 (N_2948,N_2067,N_2440);
xor U2949 (N_2949,N_2452,N_2207);
xor U2950 (N_2950,N_2203,N_2386);
and U2951 (N_2951,N_2007,N_2164);
nor U2952 (N_2952,N_2012,N_2406);
nand U2953 (N_2953,N_2025,N_2323);
nand U2954 (N_2954,N_2093,N_2310);
xor U2955 (N_2955,N_2254,N_2019);
and U2956 (N_2956,N_2279,N_2330);
nor U2957 (N_2957,N_2068,N_2488);
or U2958 (N_2958,N_2183,N_2115);
or U2959 (N_2959,N_2117,N_2339);
nor U2960 (N_2960,N_2099,N_2295);
or U2961 (N_2961,N_2424,N_2305);
xnor U2962 (N_2962,N_2125,N_2388);
and U2963 (N_2963,N_2410,N_2307);
or U2964 (N_2964,N_2322,N_2469);
or U2965 (N_2965,N_2256,N_2035);
nor U2966 (N_2966,N_2000,N_2019);
and U2967 (N_2967,N_2086,N_2387);
nor U2968 (N_2968,N_2134,N_2264);
nor U2969 (N_2969,N_2251,N_2249);
nor U2970 (N_2970,N_2130,N_2201);
xor U2971 (N_2971,N_2351,N_2036);
xor U2972 (N_2972,N_2353,N_2097);
nor U2973 (N_2973,N_2251,N_2125);
or U2974 (N_2974,N_2333,N_2321);
nand U2975 (N_2975,N_2400,N_2002);
and U2976 (N_2976,N_2121,N_2135);
nor U2977 (N_2977,N_2458,N_2460);
nor U2978 (N_2978,N_2337,N_2360);
nor U2979 (N_2979,N_2188,N_2291);
nor U2980 (N_2980,N_2427,N_2282);
or U2981 (N_2981,N_2022,N_2100);
nor U2982 (N_2982,N_2143,N_2346);
nor U2983 (N_2983,N_2142,N_2072);
nand U2984 (N_2984,N_2230,N_2188);
nor U2985 (N_2985,N_2033,N_2463);
nor U2986 (N_2986,N_2267,N_2456);
and U2987 (N_2987,N_2272,N_2159);
or U2988 (N_2988,N_2168,N_2244);
xor U2989 (N_2989,N_2246,N_2272);
xor U2990 (N_2990,N_2492,N_2009);
and U2991 (N_2991,N_2143,N_2244);
xnor U2992 (N_2992,N_2268,N_2114);
xor U2993 (N_2993,N_2467,N_2247);
nand U2994 (N_2994,N_2256,N_2069);
nor U2995 (N_2995,N_2488,N_2497);
nand U2996 (N_2996,N_2033,N_2389);
nor U2997 (N_2997,N_2381,N_2125);
nand U2998 (N_2998,N_2058,N_2450);
xor U2999 (N_2999,N_2262,N_2324);
xnor U3000 (N_3000,N_2621,N_2816);
nand U3001 (N_3001,N_2878,N_2869);
and U3002 (N_3002,N_2752,N_2550);
nand U3003 (N_3003,N_2520,N_2740);
xnor U3004 (N_3004,N_2845,N_2798);
and U3005 (N_3005,N_2747,N_2909);
xnor U3006 (N_3006,N_2742,N_2912);
or U3007 (N_3007,N_2870,N_2688);
or U3008 (N_3008,N_2767,N_2988);
and U3009 (N_3009,N_2650,N_2834);
or U3010 (N_3010,N_2769,N_2733);
nand U3011 (N_3011,N_2655,N_2794);
or U3012 (N_3012,N_2914,N_2922);
nor U3013 (N_3013,N_2738,N_2517);
nand U3014 (N_3014,N_2866,N_2672);
nand U3015 (N_3015,N_2613,N_2932);
and U3016 (N_3016,N_2586,N_2971);
nor U3017 (N_3017,N_2986,N_2824);
nor U3018 (N_3018,N_2627,N_2998);
nor U3019 (N_3019,N_2590,N_2596);
or U3020 (N_3020,N_2846,N_2879);
and U3021 (N_3021,N_2940,N_2821);
nand U3022 (N_3022,N_2979,N_2716);
nand U3023 (N_3023,N_2696,N_2796);
and U3024 (N_3024,N_2825,N_2727);
nand U3025 (N_3025,N_2648,N_2992);
nand U3026 (N_3026,N_2566,N_2967);
nor U3027 (N_3027,N_2640,N_2760);
nor U3028 (N_3028,N_2754,N_2687);
and U3029 (N_3029,N_2676,N_2860);
or U3030 (N_3030,N_2708,N_2809);
nor U3031 (N_3031,N_2921,N_2548);
and U3032 (N_3032,N_2522,N_2739);
nor U3033 (N_3033,N_2617,N_2951);
nor U3034 (N_3034,N_2568,N_2856);
nand U3035 (N_3035,N_2811,N_2525);
nor U3036 (N_3036,N_2715,N_2877);
and U3037 (N_3037,N_2563,N_2573);
nor U3038 (N_3038,N_2820,N_2958);
or U3039 (N_3039,N_2502,N_2562);
or U3040 (N_3040,N_2658,N_2614);
nand U3041 (N_3041,N_2974,N_2972);
xnor U3042 (N_3042,N_2961,N_2585);
nand U3043 (N_3043,N_2694,N_2799);
and U3044 (N_3044,N_2891,N_2612);
nand U3045 (N_3045,N_2887,N_2864);
xnor U3046 (N_3046,N_2786,N_2746);
or U3047 (N_3047,N_2959,N_2936);
xnor U3048 (N_3048,N_2605,N_2862);
or U3049 (N_3049,N_2842,N_2636);
or U3050 (N_3050,N_2718,N_2962);
and U3051 (N_3051,N_2537,N_2603);
nand U3052 (N_3052,N_2651,N_2508);
nor U3053 (N_3053,N_2591,N_2557);
xor U3054 (N_3054,N_2538,N_2584);
nor U3055 (N_3055,N_2978,N_2950);
nor U3056 (N_3056,N_2726,N_2602);
nand U3057 (N_3057,N_2871,N_2513);
and U3058 (N_3058,N_2835,N_2556);
nand U3059 (N_3059,N_2843,N_2509);
xnor U3060 (N_3060,N_2505,N_2616);
xor U3061 (N_3061,N_2955,N_2714);
nor U3062 (N_3062,N_2999,N_2876);
or U3063 (N_3063,N_2713,N_2750);
nand U3064 (N_3064,N_2904,N_2963);
xnor U3065 (N_3065,N_2626,N_2898);
xnor U3066 (N_3066,N_2944,N_2934);
nand U3067 (N_3067,N_2966,N_2721);
nand U3068 (N_3068,N_2561,N_2949);
or U3069 (N_3069,N_2826,N_2512);
xnor U3070 (N_3070,N_2947,N_2841);
and U3071 (N_3071,N_2545,N_2819);
or U3072 (N_3072,N_2983,N_2987);
or U3073 (N_3073,N_2543,N_2839);
and U3074 (N_3074,N_2812,N_2581);
nand U3075 (N_3075,N_2832,N_2792);
xor U3076 (N_3076,N_2901,N_2736);
nor U3077 (N_3077,N_2753,N_2615);
xnor U3078 (N_3078,N_2772,N_2915);
xnor U3079 (N_3079,N_2822,N_2938);
or U3080 (N_3080,N_2528,N_2572);
nor U3081 (N_3081,N_2703,N_2674);
xor U3082 (N_3082,N_2647,N_2743);
nor U3083 (N_3083,N_2526,N_2777);
xnor U3084 (N_3084,N_2629,N_2649);
nand U3085 (N_3085,N_2669,N_2504);
and U3086 (N_3086,N_2954,N_2599);
xor U3087 (N_3087,N_2593,N_2861);
nand U3088 (N_3088,N_2779,N_2833);
or U3089 (N_3089,N_2744,N_2830);
or U3090 (N_3090,N_2882,N_2637);
xor U3091 (N_3091,N_2539,N_2797);
and U3092 (N_3092,N_2663,N_2722);
nor U3093 (N_3093,N_2677,N_2985);
or U3094 (N_3094,N_2960,N_2854);
xor U3095 (N_3095,N_2883,N_2991);
or U3096 (N_3096,N_2601,N_2570);
and U3097 (N_3097,N_2929,N_2735);
and U3098 (N_3098,N_2817,N_2785);
or U3099 (N_3099,N_2695,N_2923);
or U3100 (N_3100,N_2730,N_2633);
nor U3101 (N_3101,N_2728,N_2532);
nor U3102 (N_3102,N_2501,N_2868);
or U3103 (N_3103,N_2661,N_2855);
xnor U3104 (N_3104,N_2623,N_2907);
xnor U3105 (N_3105,N_2888,N_2927);
nand U3106 (N_3106,N_2996,N_2604);
xnor U3107 (N_3107,N_2928,N_2709);
or U3108 (N_3108,N_2618,N_2576);
nor U3109 (N_3109,N_2890,N_2507);
and U3110 (N_3110,N_2659,N_2521);
or U3111 (N_3111,N_2837,N_2880);
and U3112 (N_3112,N_2540,N_2549);
or U3113 (N_3113,N_2711,N_2884);
or U3114 (N_3114,N_2751,N_2597);
nand U3115 (N_3115,N_2827,N_2635);
or U3116 (N_3116,N_2808,N_2511);
or U3117 (N_3117,N_2719,N_2995);
xor U3118 (N_3118,N_2692,N_2948);
nand U3119 (N_3119,N_2981,N_2844);
nand U3120 (N_3120,N_2766,N_2790);
nand U3121 (N_3121,N_2840,N_2533);
and U3122 (N_3122,N_2579,N_2515);
nand U3123 (N_3123,N_2737,N_2852);
or U3124 (N_3124,N_2920,N_2857);
and U3125 (N_3125,N_2609,N_2682);
xor U3126 (N_3126,N_2859,N_2780);
and U3127 (N_3127,N_2705,N_2976);
xnor U3128 (N_3128,N_2514,N_2527);
or U3129 (N_3129,N_2691,N_2681);
and U3130 (N_3130,N_2925,N_2666);
nor U3131 (N_3131,N_2555,N_2541);
nor U3132 (N_3132,N_2784,N_2710);
or U3133 (N_3133,N_2670,N_2935);
nor U3134 (N_3134,N_2865,N_2804);
or U3135 (N_3135,N_2630,N_2910);
nor U3136 (N_3136,N_2606,N_2598);
nand U3137 (N_3137,N_2815,N_2917);
or U3138 (N_3138,N_2506,N_2523);
and U3139 (N_3139,N_2503,N_2667);
or U3140 (N_3140,N_2937,N_2970);
and U3141 (N_3141,N_2930,N_2968);
nand U3142 (N_3142,N_2632,N_2571);
nand U3143 (N_3143,N_2685,N_2699);
xnor U3144 (N_3144,N_2700,N_2639);
xor U3145 (N_3145,N_2933,N_2919);
nor U3146 (N_3146,N_2975,N_2564);
nor U3147 (N_3147,N_2763,N_2892);
nor U3148 (N_3148,N_2608,N_2587);
or U3149 (N_3149,N_2622,N_2749);
nand U3150 (N_3150,N_2899,N_2806);
nand U3151 (N_3151,N_2989,N_2600);
xnor U3152 (N_3152,N_2803,N_2662);
or U3153 (N_3153,N_2993,N_2724);
xor U3154 (N_3154,N_2690,N_2712);
or U3155 (N_3155,N_2574,N_2969);
and U3156 (N_3156,N_2720,N_2893);
and U3157 (N_3157,N_2787,N_2764);
xnor U3158 (N_3158,N_2642,N_2518);
xnor U3159 (N_3159,N_2757,N_2759);
xnor U3160 (N_3160,N_2838,N_2529);
and U3161 (N_3161,N_2628,N_2801);
or U3162 (N_3162,N_2588,N_2918);
nand U3163 (N_3163,N_2701,N_2768);
xnor U3164 (N_3164,N_2943,N_2693);
nor U3165 (N_3165,N_2946,N_2953);
xnor U3166 (N_3166,N_2765,N_2592);
or U3167 (N_3167,N_2810,N_2644);
and U3168 (N_3168,N_2973,N_2789);
nor U3169 (N_3169,N_2773,N_2660);
xnor U3170 (N_3170,N_2872,N_2542);
nor U3171 (N_3171,N_2558,N_2734);
xnor U3172 (N_3172,N_2926,N_2782);
or U3173 (N_3173,N_2624,N_2791);
and U3174 (N_3174,N_2965,N_2984);
xor U3175 (N_3175,N_2977,N_2668);
nor U3176 (N_3176,N_2646,N_2828);
xnor U3177 (N_3177,N_2924,N_2678);
xnor U3178 (N_3178,N_2664,N_2707);
xor U3179 (N_3179,N_2756,N_2889);
or U3180 (N_3180,N_2913,N_2858);
and U3181 (N_3181,N_2665,N_2535);
or U3182 (N_3182,N_2990,N_2895);
nor U3183 (N_3183,N_2567,N_2885);
or U3184 (N_3184,N_2831,N_2510);
xor U3185 (N_3185,N_2813,N_2656);
xor U3186 (N_3186,N_2836,N_2595);
nand U3187 (N_3187,N_2683,N_2684);
and U3188 (N_3188,N_2755,N_2762);
nor U3189 (N_3189,N_2531,N_2671);
and U3190 (N_3190,N_2800,N_2863);
and U3191 (N_3191,N_2945,N_2807);
and U3192 (N_3192,N_2939,N_2771);
nor U3193 (N_3193,N_2553,N_2997);
and U3194 (N_3194,N_2897,N_2781);
nor U3195 (N_3195,N_2582,N_2903);
or U3196 (N_3196,N_2788,N_2620);
or U3197 (N_3197,N_2697,N_2775);
and U3198 (N_3198,N_2689,N_2875);
nor U3199 (N_3199,N_2534,N_2849);
and U3200 (N_3200,N_2631,N_2725);
nor U3201 (N_3201,N_2680,N_2653);
nand U3202 (N_3202,N_2530,N_2704);
nor U3203 (N_3203,N_2873,N_2569);
xor U3204 (N_3204,N_2778,N_2611);
nand U3205 (N_3205,N_2931,N_2894);
xnor U3206 (N_3206,N_2610,N_2594);
and U3207 (N_3207,N_2881,N_2916);
or U3208 (N_3208,N_2758,N_2942);
and U3209 (N_3209,N_2544,N_2795);
and U3210 (N_3210,N_2547,N_2761);
nor U3211 (N_3211,N_2575,N_2905);
or U3212 (N_3212,N_2565,N_2551);
nor U3213 (N_3213,N_2560,N_2732);
nand U3214 (N_3214,N_2580,N_2783);
xor U3215 (N_3215,N_2774,N_2577);
nor U3216 (N_3216,N_2643,N_2698);
nand U3217 (N_3217,N_2906,N_2900);
xor U3218 (N_3218,N_2952,N_2805);
and U3219 (N_3219,N_2911,N_2776);
and U3220 (N_3220,N_2908,N_2741);
and U3221 (N_3221,N_2645,N_2729);
or U3222 (N_3222,N_2723,N_2964);
and U3223 (N_3223,N_2519,N_2731);
nand U3224 (N_3224,N_2874,N_2625);
nand U3225 (N_3225,N_2524,N_2896);
and U3226 (N_3226,N_2848,N_2886);
and U3227 (N_3227,N_2982,N_2956);
nor U3228 (N_3228,N_2589,N_2867);
nor U3229 (N_3229,N_2554,N_2851);
or U3230 (N_3230,N_2500,N_2546);
or U3231 (N_3231,N_2607,N_2850);
xnor U3232 (N_3232,N_2673,N_2638);
nand U3233 (N_3233,N_2657,N_2847);
xor U3234 (N_3234,N_2536,N_2829);
xnor U3235 (N_3235,N_2957,N_2994);
nand U3236 (N_3236,N_2619,N_2802);
nand U3237 (N_3237,N_2652,N_2980);
nand U3238 (N_3238,N_2706,N_2559);
nand U3239 (N_3239,N_2770,N_2814);
and U3240 (N_3240,N_2853,N_2902);
and U3241 (N_3241,N_2516,N_2583);
nand U3242 (N_3242,N_2679,N_2641);
nand U3243 (N_3243,N_2748,N_2818);
nand U3244 (N_3244,N_2702,N_2823);
nor U3245 (N_3245,N_2634,N_2941);
nand U3246 (N_3246,N_2717,N_2654);
and U3247 (N_3247,N_2552,N_2578);
nand U3248 (N_3248,N_2686,N_2745);
nor U3249 (N_3249,N_2675,N_2793);
and U3250 (N_3250,N_2808,N_2525);
and U3251 (N_3251,N_2963,N_2847);
and U3252 (N_3252,N_2691,N_2769);
nand U3253 (N_3253,N_2959,N_2774);
and U3254 (N_3254,N_2780,N_2836);
and U3255 (N_3255,N_2877,N_2725);
nand U3256 (N_3256,N_2674,N_2522);
xor U3257 (N_3257,N_2761,N_2655);
and U3258 (N_3258,N_2746,N_2505);
nand U3259 (N_3259,N_2580,N_2724);
and U3260 (N_3260,N_2888,N_2972);
xnor U3261 (N_3261,N_2609,N_2922);
and U3262 (N_3262,N_2712,N_2616);
nor U3263 (N_3263,N_2585,N_2858);
or U3264 (N_3264,N_2623,N_2946);
xor U3265 (N_3265,N_2592,N_2707);
and U3266 (N_3266,N_2513,N_2596);
xnor U3267 (N_3267,N_2890,N_2956);
nand U3268 (N_3268,N_2554,N_2988);
nor U3269 (N_3269,N_2589,N_2665);
and U3270 (N_3270,N_2683,N_2546);
and U3271 (N_3271,N_2843,N_2970);
and U3272 (N_3272,N_2921,N_2599);
and U3273 (N_3273,N_2748,N_2649);
or U3274 (N_3274,N_2853,N_2977);
or U3275 (N_3275,N_2918,N_2542);
and U3276 (N_3276,N_2994,N_2518);
xnor U3277 (N_3277,N_2911,N_2997);
nand U3278 (N_3278,N_2540,N_2789);
or U3279 (N_3279,N_2998,N_2875);
nor U3280 (N_3280,N_2792,N_2736);
xor U3281 (N_3281,N_2887,N_2588);
nand U3282 (N_3282,N_2580,N_2922);
xor U3283 (N_3283,N_2966,N_2996);
xor U3284 (N_3284,N_2973,N_2574);
nand U3285 (N_3285,N_2771,N_2754);
or U3286 (N_3286,N_2974,N_2647);
xnor U3287 (N_3287,N_2872,N_2957);
and U3288 (N_3288,N_2976,N_2819);
xor U3289 (N_3289,N_2894,N_2866);
or U3290 (N_3290,N_2531,N_2667);
nor U3291 (N_3291,N_2533,N_2774);
xnor U3292 (N_3292,N_2680,N_2581);
and U3293 (N_3293,N_2506,N_2574);
nor U3294 (N_3294,N_2582,N_2511);
or U3295 (N_3295,N_2607,N_2992);
and U3296 (N_3296,N_2771,N_2717);
nand U3297 (N_3297,N_2675,N_2576);
or U3298 (N_3298,N_2657,N_2789);
xor U3299 (N_3299,N_2853,N_2597);
or U3300 (N_3300,N_2603,N_2653);
and U3301 (N_3301,N_2645,N_2623);
and U3302 (N_3302,N_2670,N_2539);
or U3303 (N_3303,N_2502,N_2870);
nor U3304 (N_3304,N_2921,N_2631);
nor U3305 (N_3305,N_2609,N_2569);
nor U3306 (N_3306,N_2606,N_2882);
xor U3307 (N_3307,N_2624,N_2880);
nor U3308 (N_3308,N_2948,N_2719);
nand U3309 (N_3309,N_2926,N_2684);
xor U3310 (N_3310,N_2684,N_2943);
nand U3311 (N_3311,N_2654,N_2704);
nand U3312 (N_3312,N_2932,N_2693);
nand U3313 (N_3313,N_2861,N_2517);
and U3314 (N_3314,N_2869,N_2919);
and U3315 (N_3315,N_2516,N_2830);
or U3316 (N_3316,N_2605,N_2614);
and U3317 (N_3317,N_2833,N_2936);
and U3318 (N_3318,N_2635,N_2916);
nand U3319 (N_3319,N_2559,N_2903);
nor U3320 (N_3320,N_2634,N_2913);
xor U3321 (N_3321,N_2949,N_2845);
xor U3322 (N_3322,N_2585,N_2625);
xnor U3323 (N_3323,N_2890,N_2604);
and U3324 (N_3324,N_2624,N_2769);
and U3325 (N_3325,N_2565,N_2534);
xnor U3326 (N_3326,N_2537,N_2874);
nor U3327 (N_3327,N_2591,N_2637);
and U3328 (N_3328,N_2923,N_2971);
nand U3329 (N_3329,N_2889,N_2923);
xnor U3330 (N_3330,N_2767,N_2726);
nand U3331 (N_3331,N_2814,N_2822);
or U3332 (N_3332,N_2746,N_2707);
nor U3333 (N_3333,N_2626,N_2946);
and U3334 (N_3334,N_2602,N_2721);
nor U3335 (N_3335,N_2880,N_2905);
and U3336 (N_3336,N_2711,N_2691);
or U3337 (N_3337,N_2540,N_2818);
and U3338 (N_3338,N_2952,N_2580);
xnor U3339 (N_3339,N_2858,N_2996);
xor U3340 (N_3340,N_2580,N_2699);
nand U3341 (N_3341,N_2569,N_2637);
and U3342 (N_3342,N_2933,N_2817);
or U3343 (N_3343,N_2637,N_2943);
xor U3344 (N_3344,N_2713,N_2854);
and U3345 (N_3345,N_2529,N_2796);
nand U3346 (N_3346,N_2925,N_2537);
and U3347 (N_3347,N_2790,N_2851);
nand U3348 (N_3348,N_2960,N_2602);
or U3349 (N_3349,N_2849,N_2803);
nor U3350 (N_3350,N_2775,N_2530);
and U3351 (N_3351,N_2663,N_2699);
nor U3352 (N_3352,N_2762,N_2523);
and U3353 (N_3353,N_2927,N_2926);
nor U3354 (N_3354,N_2660,N_2855);
and U3355 (N_3355,N_2997,N_2517);
nor U3356 (N_3356,N_2668,N_2598);
xnor U3357 (N_3357,N_2986,N_2588);
and U3358 (N_3358,N_2930,N_2637);
xor U3359 (N_3359,N_2662,N_2583);
nor U3360 (N_3360,N_2959,N_2697);
nand U3361 (N_3361,N_2796,N_2509);
xnor U3362 (N_3362,N_2658,N_2815);
nor U3363 (N_3363,N_2902,N_2904);
and U3364 (N_3364,N_2836,N_2996);
nor U3365 (N_3365,N_2887,N_2784);
xnor U3366 (N_3366,N_2740,N_2774);
or U3367 (N_3367,N_2915,N_2569);
and U3368 (N_3368,N_2736,N_2641);
nand U3369 (N_3369,N_2823,N_2830);
and U3370 (N_3370,N_2901,N_2829);
and U3371 (N_3371,N_2849,N_2529);
nor U3372 (N_3372,N_2886,N_2762);
and U3373 (N_3373,N_2753,N_2650);
or U3374 (N_3374,N_2768,N_2839);
and U3375 (N_3375,N_2872,N_2632);
or U3376 (N_3376,N_2609,N_2818);
xnor U3377 (N_3377,N_2796,N_2979);
or U3378 (N_3378,N_2536,N_2922);
or U3379 (N_3379,N_2615,N_2651);
xor U3380 (N_3380,N_2703,N_2959);
and U3381 (N_3381,N_2870,N_2729);
nor U3382 (N_3382,N_2749,N_2664);
xor U3383 (N_3383,N_2967,N_2811);
nand U3384 (N_3384,N_2600,N_2607);
nand U3385 (N_3385,N_2748,N_2576);
nand U3386 (N_3386,N_2940,N_2681);
nand U3387 (N_3387,N_2809,N_2821);
nand U3388 (N_3388,N_2969,N_2984);
nor U3389 (N_3389,N_2671,N_2949);
and U3390 (N_3390,N_2958,N_2830);
and U3391 (N_3391,N_2725,N_2867);
or U3392 (N_3392,N_2799,N_2682);
and U3393 (N_3393,N_2640,N_2591);
xnor U3394 (N_3394,N_2933,N_2920);
nor U3395 (N_3395,N_2563,N_2604);
and U3396 (N_3396,N_2881,N_2733);
and U3397 (N_3397,N_2510,N_2910);
nand U3398 (N_3398,N_2580,N_2975);
and U3399 (N_3399,N_2699,N_2739);
xor U3400 (N_3400,N_2616,N_2938);
xor U3401 (N_3401,N_2598,N_2792);
nor U3402 (N_3402,N_2502,N_2933);
and U3403 (N_3403,N_2969,N_2520);
nand U3404 (N_3404,N_2758,N_2616);
xor U3405 (N_3405,N_2660,N_2650);
xnor U3406 (N_3406,N_2551,N_2800);
and U3407 (N_3407,N_2758,N_2826);
xor U3408 (N_3408,N_2802,N_2593);
xnor U3409 (N_3409,N_2866,N_2670);
and U3410 (N_3410,N_2829,N_2640);
or U3411 (N_3411,N_2954,N_2826);
nand U3412 (N_3412,N_2720,N_2654);
or U3413 (N_3413,N_2877,N_2902);
nor U3414 (N_3414,N_2942,N_2829);
and U3415 (N_3415,N_2976,N_2788);
nor U3416 (N_3416,N_2900,N_2644);
xor U3417 (N_3417,N_2656,N_2852);
and U3418 (N_3418,N_2728,N_2756);
xnor U3419 (N_3419,N_2761,N_2823);
nand U3420 (N_3420,N_2653,N_2871);
nor U3421 (N_3421,N_2925,N_2518);
nand U3422 (N_3422,N_2822,N_2825);
and U3423 (N_3423,N_2543,N_2651);
or U3424 (N_3424,N_2985,N_2926);
nand U3425 (N_3425,N_2723,N_2846);
xor U3426 (N_3426,N_2535,N_2584);
and U3427 (N_3427,N_2873,N_2814);
and U3428 (N_3428,N_2657,N_2958);
nand U3429 (N_3429,N_2797,N_2617);
nand U3430 (N_3430,N_2715,N_2583);
nand U3431 (N_3431,N_2765,N_2659);
nand U3432 (N_3432,N_2927,N_2870);
and U3433 (N_3433,N_2919,N_2836);
nor U3434 (N_3434,N_2856,N_2953);
and U3435 (N_3435,N_2839,N_2808);
or U3436 (N_3436,N_2926,N_2957);
or U3437 (N_3437,N_2587,N_2676);
or U3438 (N_3438,N_2509,N_2928);
and U3439 (N_3439,N_2921,N_2815);
nor U3440 (N_3440,N_2726,N_2958);
or U3441 (N_3441,N_2564,N_2910);
and U3442 (N_3442,N_2509,N_2533);
nand U3443 (N_3443,N_2653,N_2786);
or U3444 (N_3444,N_2875,N_2721);
and U3445 (N_3445,N_2701,N_2661);
or U3446 (N_3446,N_2724,N_2819);
and U3447 (N_3447,N_2836,N_2734);
and U3448 (N_3448,N_2698,N_2782);
or U3449 (N_3449,N_2540,N_2913);
and U3450 (N_3450,N_2769,N_2922);
nand U3451 (N_3451,N_2853,N_2967);
and U3452 (N_3452,N_2821,N_2508);
xnor U3453 (N_3453,N_2965,N_2781);
xnor U3454 (N_3454,N_2777,N_2557);
nand U3455 (N_3455,N_2732,N_2550);
and U3456 (N_3456,N_2948,N_2801);
nand U3457 (N_3457,N_2507,N_2847);
and U3458 (N_3458,N_2955,N_2541);
xor U3459 (N_3459,N_2828,N_2813);
nor U3460 (N_3460,N_2675,N_2784);
or U3461 (N_3461,N_2968,N_2565);
xnor U3462 (N_3462,N_2945,N_2982);
nor U3463 (N_3463,N_2512,N_2920);
xor U3464 (N_3464,N_2792,N_2858);
xnor U3465 (N_3465,N_2630,N_2666);
or U3466 (N_3466,N_2748,N_2671);
or U3467 (N_3467,N_2901,N_2926);
nor U3468 (N_3468,N_2877,N_2680);
or U3469 (N_3469,N_2742,N_2966);
xnor U3470 (N_3470,N_2815,N_2696);
or U3471 (N_3471,N_2720,N_2750);
and U3472 (N_3472,N_2816,N_2841);
or U3473 (N_3473,N_2884,N_2826);
xnor U3474 (N_3474,N_2970,N_2825);
xor U3475 (N_3475,N_2643,N_2847);
or U3476 (N_3476,N_2681,N_2577);
and U3477 (N_3477,N_2567,N_2831);
and U3478 (N_3478,N_2969,N_2597);
or U3479 (N_3479,N_2709,N_2504);
and U3480 (N_3480,N_2985,N_2928);
xnor U3481 (N_3481,N_2946,N_2822);
nand U3482 (N_3482,N_2561,N_2501);
nor U3483 (N_3483,N_2604,N_2557);
and U3484 (N_3484,N_2655,N_2739);
nor U3485 (N_3485,N_2969,N_2607);
or U3486 (N_3486,N_2740,N_2533);
and U3487 (N_3487,N_2581,N_2994);
nand U3488 (N_3488,N_2760,N_2959);
nand U3489 (N_3489,N_2990,N_2758);
and U3490 (N_3490,N_2551,N_2576);
nand U3491 (N_3491,N_2692,N_2659);
or U3492 (N_3492,N_2812,N_2592);
nor U3493 (N_3493,N_2600,N_2679);
nand U3494 (N_3494,N_2630,N_2618);
nand U3495 (N_3495,N_2748,N_2531);
xor U3496 (N_3496,N_2711,N_2939);
and U3497 (N_3497,N_2767,N_2626);
and U3498 (N_3498,N_2585,N_2811);
nor U3499 (N_3499,N_2522,N_2643);
xor U3500 (N_3500,N_3400,N_3406);
or U3501 (N_3501,N_3007,N_3333);
or U3502 (N_3502,N_3307,N_3204);
nor U3503 (N_3503,N_3015,N_3350);
nand U3504 (N_3504,N_3153,N_3098);
and U3505 (N_3505,N_3026,N_3415);
and U3506 (N_3506,N_3006,N_3221);
or U3507 (N_3507,N_3249,N_3326);
nand U3508 (N_3508,N_3446,N_3422);
and U3509 (N_3509,N_3359,N_3013);
and U3510 (N_3510,N_3417,N_3148);
or U3511 (N_3511,N_3374,N_3165);
nand U3512 (N_3512,N_3478,N_3185);
nor U3513 (N_3513,N_3490,N_3274);
or U3514 (N_3514,N_3432,N_3420);
nor U3515 (N_3515,N_3058,N_3358);
nor U3516 (N_3516,N_3300,N_3338);
xnor U3517 (N_3517,N_3216,N_3209);
and U3518 (N_3518,N_3441,N_3459);
or U3519 (N_3519,N_3010,N_3469);
and U3520 (N_3520,N_3450,N_3468);
or U3521 (N_3521,N_3346,N_3329);
and U3522 (N_3522,N_3484,N_3143);
xor U3523 (N_3523,N_3122,N_3294);
nor U3524 (N_3524,N_3240,N_3285);
nor U3525 (N_3525,N_3078,N_3011);
nor U3526 (N_3526,N_3072,N_3452);
and U3527 (N_3527,N_3448,N_3107);
nor U3528 (N_3528,N_3138,N_3395);
nand U3529 (N_3529,N_3392,N_3213);
xor U3530 (N_3530,N_3187,N_3247);
xnor U3531 (N_3531,N_3318,N_3466);
nor U3532 (N_3532,N_3370,N_3298);
nor U3533 (N_3533,N_3184,N_3489);
or U3534 (N_3534,N_3252,N_3278);
nor U3535 (N_3535,N_3291,N_3281);
xor U3536 (N_3536,N_3226,N_3339);
or U3537 (N_3537,N_3086,N_3167);
nand U3538 (N_3538,N_3473,N_3280);
xor U3539 (N_3539,N_3104,N_3408);
xnor U3540 (N_3540,N_3151,N_3488);
or U3541 (N_3541,N_3344,N_3389);
nand U3542 (N_3542,N_3233,N_3364);
nand U3543 (N_3543,N_3225,N_3066);
nor U3544 (N_3544,N_3047,N_3382);
nand U3545 (N_3545,N_3012,N_3287);
and U3546 (N_3546,N_3124,N_3057);
and U3547 (N_3547,N_3223,N_3376);
xnor U3548 (N_3548,N_3105,N_3203);
nor U3549 (N_3549,N_3091,N_3134);
xor U3550 (N_3550,N_3366,N_3152);
xor U3551 (N_3551,N_3429,N_3399);
or U3552 (N_3552,N_3470,N_3335);
and U3553 (N_3553,N_3268,N_3398);
and U3554 (N_3554,N_3243,N_3262);
xor U3555 (N_3555,N_3177,N_3372);
and U3556 (N_3556,N_3384,N_3352);
nor U3557 (N_3557,N_3355,N_3171);
nand U3558 (N_3558,N_3313,N_3297);
nor U3559 (N_3559,N_3175,N_3277);
and U3560 (N_3560,N_3436,N_3212);
nand U3561 (N_3561,N_3418,N_3402);
nor U3562 (N_3562,N_3327,N_3407);
nor U3563 (N_3563,N_3302,N_3462);
nand U3564 (N_3564,N_3232,N_3433);
nor U3565 (N_3565,N_3437,N_3311);
and U3566 (N_3566,N_3022,N_3260);
nand U3567 (N_3567,N_3306,N_3371);
xor U3568 (N_3568,N_3027,N_3331);
nor U3569 (N_3569,N_3269,N_3101);
or U3570 (N_3570,N_3017,N_3270);
or U3571 (N_3571,N_3196,N_3497);
nand U3572 (N_3572,N_3170,N_3354);
nor U3573 (N_3573,N_3121,N_3486);
nor U3574 (N_3574,N_3075,N_3033);
or U3575 (N_3575,N_3062,N_3083);
and U3576 (N_3576,N_3275,N_3120);
or U3577 (N_3577,N_3035,N_3123);
xor U3578 (N_3578,N_3087,N_3258);
xor U3579 (N_3579,N_3467,N_3328);
or U3580 (N_3580,N_3273,N_3482);
and U3581 (N_3581,N_3303,N_3174);
or U3582 (N_3582,N_3193,N_3276);
nor U3583 (N_3583,N_3289,N_3309);
nand U3584 (N_3584,N_3261,N_3409);
and U3585 (N_3585,N_3080,N_3324);
xnor U3586 (N_3586,N_3379,N_3345);
and U3587 (N_3587,N_3005,N_3043);
nand U3588 (N_3588,N_3081,N_3236);
nand U3589 (N_3589,N_3472,N_3334);
xor U3590 (N_3590,N_3373,N_3439);
and U3591 (N_3591,N_3357,N_3018);
or U3592 (N_3592,N_3454,N_3041);
xnor U3593 (N_3593,N_3169,N_3238);
or U3594 (N_3594,N_3230,N_3383);
and U3595 (N_3595,N_3413,N_3410);
nor U3596 (N_3596,N_3388,N_3248);
nand U3597 (N_3597,N_3115,N_3109);
nand U3598 (N_3598,N_3447,N_3480);
nand U3599 (N_3599,N_3394,N_3189);
and U3600 (N_3600,N_3263,N_3188);
nor U3601 (N_3601,N_3491,N_3246);
nand U3602 (N_3602,N_3396,N_3255);
or U3603 (N_3603,N_3397,N_3191);
and U3604 (N_3604,N_3231,N_3479);
or U3605 (N_3605,N_3160,N_3332);
or U3606 (N_3606,N_3234,N_3265);
and U3607 (N_3607,N_3438,N_3060);
nand U3608 (N_3608,N_3423,N_3119);
nor U3609 (N_3609,N_3251,N_3215);
and U3610 (N_3610,N_3034,N_3428);
nor U3611 (N_3611,N_3031,N_3219);
nand U3612 (N_3612,N_3290,N_3016);
and U3613 (N_3613,N_3093,N_3126);
and U3614 (N_3614,N_3176,N_3199);
nand U3615 (N_3615,N_3054,N_3227);
and U3616 (N_3616,N_3178,N_3008);
nand U3617 (N_3617,N_3250,N_3367);
nor U3618 (N_3618,N_3146,N_3390);
nor U3619 (N_3619,N_3020,N_3315);
xnor U3620 (N_3620,N_3025,N_3061);
xnor U3621 (N_3621,N_3127,N_3444);
or U3622 (N_3622,N_3430,N_3463);
xnor U3623 (N_3623,N_3110,N_3460);
xnor U3624 (N_3624,N_3292,N_3461);
and U3625 (N_3625,N_3414,N_3097);
or U3626 (N_3626,N_3496,N_3200);
nor U3627 (N_3627,N_3205,N_3435);
and U3628 (N_3628,N_3442,N_3464);
and U3629 (N_3629,N_3312,N_3229);
and U3630 (N_3630,N_3445,N_3003);
and U3631 (N_3631,N_3089,N_3492);
nand U3632 (N_3632,N_3343,N_3116);
nand U3633 (N_3633,N_3067,N_3340);
nor U3634 (N_3634,N_3149,N_3190);
xor U3635 (N_3635,N_3100,N_3304);
nand U3636 (N_3636,N_3001,N_3253);
nor U3637 (N_3637,N_3481,N_3135);
xnor U3638 (N_3638,N_3141,N_3049);
or U3639 (N_3639,N_3162,N_3164);
nor U3640 (N_3640,N_3136,N_3076);
nor U3641 (N_3641,N_3044,N_3412);
and U3642 (N_3642,N_3257,N_3245);
and U3643 (N_3643,N_3440,N_3052);
and U3644 (N_3644,N_3195,N_3028);
nand U3645 (N_3645,N_3055,N_3351);
or U3646 (N_3646,N_3092,N_3449);
and U3647 (N_3647,N_3356,N_3474);
and U3648 (N_3648,N_3498,N_3314);
nand U3649 (N_3649,N_3056,N_3237);
xor U3650 (N_3650,N_3477,N_3036);
or U3651 (N_3651,N_3202,N_3166);
nor U3652 (N_3652,N_3073,N_3330);
xor U3653 (N_3653,N_3322,N_3368);
nor U3654 (N_3654,N_3009,N_3451);
nand U3655 (N_3655,N_3032,N_3220);
xnor U3656 (N_3656,N_3279,N_3348);
nand U3657 (N_3657,N_3051,N_3476);
nand U3658 (N_3658,N_3117,N_3282);
nor U3659 (N_3659,N_3456,N_3068);
nand U3660 (N_3660,N_3082,N_3323);
nor U3661 (N_3661,N_3125,N_3077);
xnor U3662 (N_3662,N_3264,N_3186);
xor U3663 (N_3663,N_3118,N_3059);
and U3664 (N_3664,N_3180,N_3150);
nand U3665 (N_3665,N_3353,N_3208);
xor U3666 (N_3666,N_3375,N_3391);
and U3667 (N_3667,N_3085,N_3295);
xor U3668 (N_3668,N_3000,N_3158);
nor U3669 (N_3669,N_3404,N_3139);
or U3670 (N_3670,N_3046,N_3014);
xnor U3671 (N_3671,N_3421,N_3443);
xnor U3672 (N_3672,N_3310,N_3487);
or U3673 (N_3673,N_3241,N_3341);
xnor U3674 (N_3674,N_3224,N_3161);
nand U3675 (N_3675,N_3172,N_3347);
and U3676 (N_3676,N_3272,N_3284);
nand U3677 (N_3677,N_3256,N_3453);
nand U3678 (N_3678,N_3038,N_3360);
xor U3679 (N_3679,N_3071,N_3401);
and U3680 (N_3680,N_3319,N_3424);
or U3681 (N_3681,N_3021,N_3103);
or U3682 (N_3682,N_3434,N_3266);
nor U3683 (N_3683,N_3301,N_3385);
and U3684 (N_3684,N_3106,N_3201);
nand U3685 (N_3685,N_3156,N_3173);
or U3686 (N_3686,N_3342,N_3361);
nand U3687 (N_3687,N_3030,N_3197);
or U3688 (N_3688,N_3002,N_3362);
or U3689 (N_3689,N_3129,N_3239);
or U3690 (N_3690,N_3214,N_3393);
nand U3691 (N_3691,N_3493,N_3198);
xnor U3692 (N_3692,N_3131,N_3235);
xnor U3693 (N_3693,N_3218,N_3308);
or U3694 (N_3694,N_3426,N_3192);
xnor U3695 (N_3695,N_3349,N_3457);
xnor U3696 (N_3696,N_3431,N_3179);
xor U3697 (N_3697,N_3140,N_3037);
xor U3698 (N_3698,N_3483,N_3217);
nand U3699 (N_3699,N_3168,N_3094);
and U3700 (N_3700,N_3416,N_3079);
xor U3701 (N_3701,N_3207,N_3455);
xnor U3702 (N_3702,N_3074,N_3050);
xnor U3703 (N_3703,N_3137,N_3069);
or U3704 (N_3704,N_3157,N_3244);
or U3705 (N_3705,N_3159,N_3254);
nand U3706 (N_3706,N_3147,N_3377);
nor U3707 (N_3707,N_3365,N_3363);
nand U3708 (N_3708,N_3183,N_3299);
or U3709 (N_3709,N_3386,N_3321);
xor U3710 (N_3710,N_3063,N_3222);
nor U3711 (N_3711,N_3271,N_3114);
or U3712 (N_3712,N_3378,N_3039);
xor U3713 (N_3713,N_3194,N_3023);
or U3714 (N_3714,N_3181,N_3142);
nor U3715 (N_3715,N_3111,N_3405);
nor U3716 (N_3716,N_3288,N_3305);
xnor U3717 (N_3717,N_3267,N_3145);
nor U3718 (N_3718,N_3108,N_3427);
nor U3719 (N_3719,N_3144,N_3163);
or U3720 (N_3720,N_3458,N_3064);
or U3721 (N_3721,N_3317,N_3133);
nand U3722 (N_3722,N_3337,N_3182);
nor U3723 (N_3723,N_3336,N_3494);
and U3724 (N_3724,N_3465,N_3499);
or U3725 (N_3725,N_3088,N_3242);
xnor U3726 (N_3726,N_3024,N_3283);
nand U3727 (N_3727,N_3048,N_3425);
xnor U3728 (N_3728,N_3096,N_3381);
and U3729 (N_3729,N_3495,N_3387);
xor U3730 (N_3730,N_3053,N_3286);
nor U3731 (N_3731,N_3471,N_3485);
and U3732 (N_3732,N_3084,N_3128);
nand U3733 (N_3733,N_3042,N_3380);
or U3734 (N_3734,N_3325,N_3099);
and U3735 (N_3735,N_3045,N_3210);
and U3736 (N_3736,N_3029,N_3211);
xnor U3737 (N_3737,N_3113,N_3228);
and U3738 (N_3738,N_3132,N_3019);
xor U3739 (N_3739,N_3155,N_3403);
or U3740 (N_3740,N_3316,N_3065);
nor U3741 (N_3741,N_3296,N_3102);
nor U3742 (N_3742,N_3090,N_3070);
or U3743 (N_3743,N_3369,N_3320);
xor U3744 (N_3744,N_3095,N_3154);
nand U3745 (N_3745,N_3411,N_3259);
xor U3746 (N_3746,N_3293,N_3419);
and U3747 (N_3747,N_3004,N_3475);
nand U3748 (N_3748,N_3040,N_3112);
xnor U3749 (N_3749,N_3130,N_3206);
or U3750 (N_3750,N_3170,N_3013);
or U3751 (N_3751,N_3192,N_3206);
and U3752 (N_3752,N_3219,N_3044);
xnor U3753 (N_3753,N_3454,N_3386);
nor U3754 (N_3754,N_3220,N_3404);
nor U3755 (N_3755,N_3178,N_3449);
and U3756 (N_3756,N_3358,N_3396);
nand U3757 (N_3757,N_3396,N_3406);
nand U3758 (N_3758,N_3133,N_3391);
and U3759 (N_3759,N_3298,N_3291);
or U3760 (N_3760,N_3390,N_3268);
nor U3761 (N_3761,N_3136,N_3306);
nor U3762 (N_3762,N_3435,N_3208);
and U3763 (N_3763,N_3398,N_3035);
nor U3764 (N_3764,N_3088,N_3136);
nor U3765 (N_3765,N_3392,N_3090);
nand U3766 (N_3766,N_3403,N_3023);
or U3767 (N_3767,N_3493,N_3181);
and U3768 (N_3768,N_3462,N_3145);
or U3769 (N_3769,N_3356,N_3334);
or U3770 (N_3770,N_3099,N_3339);
nand U3771 (N_3771,N_3329,N_3078);
nand U3772 (N_3772,N_3005,N_3275);
nand U3773 (N_3773,N_3436,N_3419);
nor U3774 (N_3774,N_3317,N_3364);
xor U3775 (N_3775,N_3370,N_3025);
nor U3776 (N_3776,N_3265,N_3196);
nand U3777 (N_3777,N_3285,N_3360);
xor U3778 (N_3778,N_3177,N_3285);
nor U3779 (N_3779,N_3125,N_3479);
nand U3780 (N_3780,N_3052,N_3431);
nor U3781 (N_3781,N_3051,N_3154);
or U3782 (N_3782,N_3285,N_3394);
and U3783 (N_3783,N_3432,N_3135);
nand U3784 (N_3784,N_3043,N_3369);
or U3785 (N_3785,N_3472,N_3474);
xor U3786 (N_3786,N_3134,N_3152);
nor U3787 (N_3787,N_3134,N_3200);
xor U3788 (N_3788,N_3244,N_3206);
nand U3789 (N_3789,N_3062,N_3420);
and U3790 (N_3790,N_3308,N_3000);
nor U3791 (N_3791,N_3308,N_3474);
or U3792 (N_3792,N_3123,N_3126);
and U3793 (N_3793,N_3199,N_3450);
or U3794 (N_3794,N_3348,N_3261);
xnor U3795 (N_3795,N_3331,N_3074);
or U3796 (N_3796,N_3443,N_3417);
or U3797 (N_3797,N_3275,N_3381);
nand U3798 (N_3798,N_3186,N_3228);
and U3799 (N_3799,N_3046,N_3055);
nand U3800 (N_3800,N_3228,N_3339);
nand U3801 (N_3801,N_3378,N_3452);
or U3802 (N_3802,N_3409,N_3313);
xor U3803 (N_3803,N_3364,N_3191);
and U3804 (N_3804,N_3275,N_3233);
nand U3805 (N_3805,N_3225,N_3395);
and U3806 (N_3806,N_3255,N_3120);
nor U3807 (N_3807,N_3037,N_3007);
or U3808 (N_3808,N_3402,N_3096);
xor U3809 (N_3809,N_3150,N_3091);
or U3810 (N_3810,N_3156,N_3365);
xor U3811 (N_3811,N_3061,N_3423);
or U3812 (N_3812,N_3149,N_3419);
or U3813 (N_3813,N_3275,N_3201);
and U3814 (N_3814,N_3235,N_3307);
and U3815 (N_3815,N_3211,N_3045);
and U3816 (N_3816,N_3218,N_3489);
nand U3817 (N_3817,N_3195,N_3126);
xnor U3818 (N_3818,N_3077,N_3117);
or U3819 (N_3819,N_3380,N_3420);
and U3820 (N_3820,N_3434,N_3350);
and U3821 (N_3821,N_3025,N_3006);
or U3822 (N_3822,N_3324,N_3406);
or U3823 (N_3823,N_3070,N_3183);
or U3824 (N_3824,N_3021,N_3092);
nor U3825 (N_3825,N_3247,N_3264);
xor U3826 (N_3826,N_3422,N_3111);
nand U3827 (N_3827,N_3243,N_3436);
nor U3828 (N_3828,N_3025,N_3244);
nor U3829 (N_3829,N_3403,N_3284);
nor U3830 (N_3830,N_3310,N_3123);
nor U3831 (N_3831,N_3014,N_3438);
nand U3832 (N_3832,N_3469,N_3298);
nand U3833 (N_3833,N_3430,N_3294);
xnor U3834 (N_3834,N_3111,N_3133);
or U3835 (N_3835,N_3106,N_3455);
and U3836 (N_3836,N_3383,N_3067);
xnor U3837 (N_3837,N_3038,N_3102);
nor U3838 (N_3838,N_3196,N_3231);
and U3839 (N_3839,N_3453,N_3222);
nand U3840 (N_3840,N_3056,N_3442);
nor U3841 (N_3841,N_3199,N_3042);
or U3842 (N_3842,N_3452,N_3246);
or U3843 (N_3843,N_3175,N_3267);
nor U3844 (N_3844,N_3489,N_3483);
and U3845 (N_3845,N_3119,N_3232);
nand U3846 (N_3846,N_3216,N_3288);
nor U3847 (N_3847,N_3332,N_3140);
or U3848 (N_3848,N_3214,N_3479);
nor U3849 (N_3849,N_3093,N_3139);
and U3850 (N_3850,N_3222,N_3302);
and U3851 (N_3851,N_3499,N_3328);
xor U3852 (N_3852,N_3485,N_3389);
nand U3853 (N_3853,N_3326,N_3072);
or U3854 (N_3854,N_3188,N_3142);
or U3855 (N_3855,N_3351,N_3110);
xnor U3856 (N_3856,N_3111,N_3155);
and U3857 (N_3857,N_3262,N_3132);
or U3858 (N_3858,N_3060,N_3084);
nand U3859 (N_3859,N_3425,N_3084);
nor U3860 (N_3860,N_3311,N_3175);
nor U3861 (N_3861,N_3383,N_3076);
nand U3862 (N_3862,N_3302,N_3308);
and U3863 (N_3863,N_3283,N_3368);
nand U3864 (N_3864,N_3049,N_3254);
nor U3865 (N_3865,N_3082,N_3378);
xor U3866 (N_3866,N_3451,N_3188);
xor U3867 (N_3867,N_3154,N_3060);
and U3868 (N_3868,N_3332,N_3397);
nor U3869 (N_3869,N_3492,N_3232);
or U3870 (N_3870,N_3048,N_3169);
xor U3871 (N_3871,N_3205,N_3098);
and U3872 (N_3872,N_3473,N_3436);
nor U3873 (N_3873,N_3095,N_3224);
or U3874 (N_3874,N_3313,N_3497);
and U3875 (N_3875,N_3375,N_3114);
nor U3876 (N_3876,N_3469,N_3406);
or U3877 (N_3877,N_3145,N_3211);
xor U3878 (N_3878,N_3396,N_3262);
or U3879 (N_3879,N_3196,N_3003);
and U3880 (N_3880,N_3393,N_3402);
xnor U3881 (N_3881,N_3332,N_3157);
or U3882 (N_3882,N_3099,N_3316);
nor U3883 (N_3883,N_3191,N_3452);
or U3884 (N_3884,N_3388,N_3364);
and U3885 (N_3885,N_3250,N_3131);
and U3886 (N_3886,N_3140,N_3458);
and U3887 (N_3887,N_3063,N_3396);
or U3888 (N_3888,N_3378,N_3357);
and U3889 (N_3889,N_3297,N_3318);
nor U3890 (N_3890,N_3065,N_3338);
and U3891 (N_3891,N_3403,N_3177);
nand U3892 (N_3892,N_3015,N_3414);
nor U3893 (N_3893,N_3346,N_3109);
nor U3894 (N_3894,N_3040,N_3254);
nor U3895 (N_3895,N_3444,N_3462);
or U3896 (N_3896,N_3470,N_3475);
or U3897 (N_3897,N_3070,N_3497);
xor U3898 (N_3898,N_3052,N_3395);
nor U3899 (N_3899,N_3257,N_3357);
or U3900 (N_3900,N_3498,N_3201);
nor U3901 (N_3901,N_3219,N_3269);
nand U3902 (N_3902,N_3488,N_3250);
nor U3903 (N_3903,N_3308,N_3248);
nor U3904 (N_3904,N_3117,N_3127);
and U3905 (N_3905,N_3107,N_3329);
nor U3906 (N_3906,N_3408,N_3297);
nand U3907 (N_3907,N_3273,N_3304);
xor U3908 (N_3908,N_3260,N_3201);
nor U3909 (N_3909,N_3445,N_3268);
or U3910 (N_3910,N_3060,N_3470);
and U3911 (N_3911,N_3298,N_3475);
nand U3912 (N_3912,N_3407,N_3033);
and U3913 (N_3913,N_3375,N_3188);
xnor U3914 (N_3914,N_3179,N_3040);
and U3915 (N_3915,N_3322,N_3307);
or U3916 (N_3916,N_3255,N_3479);
or U3917 (N_3917,N_3025,N_3443);
nor U3918 (N_3918,N_3239,N_3329);
or U3919 (N_3919,N_3205,N_3280);
nand U3920 (N_3920,N_3295,N_3485);
or U3921 (N_3921,N_3144,N_3253);
nor U3922 (N_3922,N_3158,N_3300);
and U3923 (N_3923,N_3256,N_3205);
xor U3924 (N_3924,N_3184,N_3045);
and U3925 (N_3925,N_3477,N_3482);
and U3926 (N_3926,N_3153,N_3433);
and U3927 (N_3927,N_3397,N_3045);
nor U3928 (N_3928,N_3293,N_3400);
nor U3929 (N_3929,N_3350,N_3081);
and U3930 (N_3930,N_3155,N_3113);
and U3931 (N_3931,N_3473,N_3425);
and U3932 (N_3932,N_3422,N_3361);
xnor U3933 (N_3933,N_3350,N_3039);
and U3934 (N_3934,N_3104,N_3077);
nor U3935 (N_3935,N_3447,N_3034);
xnor U3936 (N_3936,N_3258,N_3151);
nor U3937 (N_3937,N_3165,N_3224);
xnor U3938 (N_3938,N_3135,N_3115);
xnor U3939 (N_3939,N_3008,N_3225);
xor U3940 (N_3940,N_3282,N_3173);
and U3941 (N_3941,N_3257,N_3392);
nand U3942 (N_3942,N_3107,N_3410);
or U3943 (N_3943,N_3473,N_3217);
and U3944 (N_3944,N_3154,N_3401);
xnor U3945 (N_3945,N_3141,N_3183);
nand U3946 (N_3946,N_3322,N_3152);
or U3947 (N_3947,N_3191,N_3430);
xnor U3948 (N_3948,N_3446,N_3020);
nand U3949 (N_3949,N_3098,N_3126);
or U3950 (N_3950,N_3372,N_3298);
and U3951 (N_3951,N_3281,N_3026);
and U3952 (N_3952,N_3171,N_3352);
nor U3953 (N_3953,N_3465,N_3002);
nand U3954 (N_3954,N_3193,N_3106);
nor U3955 (N_3955,N_3020,N_3408);
nor U3956 (N_3956,N_3291,N_3195);
xnor U3957 (N_3957,N_3448,N_3325);
nor U3958 (N_3958,N_3023,N_3172);
nor U3959 (N_3959,N_3062,N_3422);
or U3960 (N_3960,N_3463,N_3467);
and U3961 (N_3961,N_3264,N_3298);
nand U3962 (N_3962,N_3440,N_3387);
and U3963 (N_3963,N_3264,N_3344);
nor U3964 (N_3964,N_3245,N_3137);
nor U3965 (N_3965,N_3183,N_3406);
xor U3966 (N_3966,N_3353,N_3447);
nand U3967 (N_3967,N_3195,N_3110);
nand U3968 (N_3968,N_3187,N_3128);
or U3969 (N_3969,N_3383,N_3153);
or U3970 (N_3970,N_3461,N_3346);
nand U3971 (N_3971,N_3106,N_3299);
or U3972 (N_3972,N_3288,N_3250);
and U3973 (N_3973,N_3080,N_3028);
and U3974 (N_3974,N_3322,N_3330);
or U3975 (N_3975,N_3312,N_3446);
nor U3976 (N_3976,N_3313,N_3281);
nand U3977 (N_3977,N_3128,N_3173);
nor U3978 (N_3978,N_3371,N_3403);
nor U3979 (N_3979,N_3364,N_3082);
nor U3980 (N_3980,N_3109,N_3399);
nand U3981 (N_3981,N_3389,N_3332);
and U3982 (N_3982,N_3120,N_3051);
or U3983 (N_3983,N_3091,N_3324);
xnor U3984 (N_3984,N_3014,N_3304);
nor U3985 (N_3985,N_3148,N_3085);
nor U3986 (N_3986,N_3115,N_3492);
xor U3987 (N_3987,N_3419,N_3484);
xnor U3988 (N_3988,N_3413,N_3084);
nor U3989 (N_3989,N_3498,N_3278);
or U3990 (N_3990,N_3321,N_3493);
xor U3991 (N_3991,N_3400,N_3230);
and U3992 (N_3992,N_3114,N_3100);
xor U3993 (N_3993,N_3060,N_3464);
nor U3994 (N_3994,N_3404,N_3108);
or U3995 (N_3995,N_3353,N_3463);
or U3996 (N_3996,N_3494,N_3199);
nand U3997 (N_3997,N_3450,N_3260);
and U3998 (N_3998,N_3152,N_3064);
or U3999 (N_3999,N_3205,N_3019);
nor U4000 (N_4000,N_3796,N_3829);
nand U4001 (N_4001,N_3566,N_3858);
xor U4002 (N_4002,N_3672,N_3572);
or U4003 (N_4003,N_3909,N_3710);
or U4004 (N_4004,N_3805,N_3747);
nor U4005 (N_4005,N_3703,N_3833);
nor U4006 (N_4006,N_3732,N_3719);
nand U4007 (N_4007,N_3507,N_3607);
nor U4008 (N_4008,N_3966,N_3897);
nand U4009 (N_4009,N_3871,N_3995);
nand U4010 (N_4010,N_3821,N_3576);
nand U4011 (N_4011,N_3724,N_3853);
and U4012 (N_4012,N_3979,N_3538);
nand U4013 (N_4013,N_3973,N_3891);
and U4014 (N_4014,N_3579,N_3911);
nor U4015 (N_4015,N_3661,N_3827);
or U4016 (N_4016,N_3881,N_3647);
nor U4017 (N_4017,N_3549,N_3770);
and U4018 (N_4018,N_3813,N_3842);
and U4019 (N_4019,N_3823,N_3761);
nor U4020 (N_4020,N_3716,N_3963);
or U4021 (N_4021,N_3508,N_3941);
and U4022 (N_4022,N_3830,N_3651);
xor U4023 (N_4023,N_3601,N_3534);
nand U4024 (N_4024,N_3967,N_3559);
and U4025 (N_4025,N_3928,N_3844);
xnor U4026 (N_4026,N_3779,N_3933);
nor U4027 (N_4027,N_3650,N_3916);
xor U4028 (N_4028,N_3504,N_3878);
or U4029 (N_4029,N_3575,N_3992);
and U4030 (N_4030,N_3637,N_3804);
or U4031 (N_4031,N_3634,N_3937);
nor U4032 (N_4032,N_3723,N_3692);
and U4033 (N_4033,N_3910,N_3729);
nand U4034 (N_4034,N_3521,N_3654);
xor U4035 (N_4035,N_3797,N_3686);
nor U4036 (N_4036,N_3894,N_3629);
nor U4037 (N_4037,N_3569,N_3548);
and U4038 (N_4038,N_3552,N_3763);
and U4039 (N_4039,N_3644,N_3917);
or U4040 (N_4040,N_3513,N_3918);
and U4041 (N_4041,N_3617,N_3915);
xnor U4042 (N_4042,N_3595,N_3817);
xnor U4043 (N_4043,N_3746,N_3989);
or U4044 (N_4044,N_3743,N_3808);
or U4045 (N_4045,N_3608,N_3996);
and U4046 (N_4046,N_3599,N_3795);
xnor U4047 (N_4047,N_3960,N_3877);
nand U4048 (N_4048,N_3848,N_3893);
xnor U4049 (N_4049,N_3852,N_3886);
nand U4050 (N_4050,N_3593,N_3955);
nand U4051 (N_4051,N_3828,N_3585);
nand U4052 (N_4052,N_3653,N_3982);
nor U4053 (N_4053,N_3621,N_3868);
or U4054 (N_4054,N_3988,N_3938);
and U4055 (N_4055,N_3857,N_3753);
and U4056 (N_4056,N_3624,N_3849);
and U4057 (N_4057,N_3768,N_3865);
and U4058 (N_4058,N_3684,N_3749);
nor U4059 (N_4059,N_3990,N_3819);
xor U4060 (N_4060,N_3929,N_3913);
nand U4061 (N_4061,N_3999,N_3978);
and U4062 (N_4062,N_3876,N_3643);
or U4063 (N_4063,N_3900,N_3883);
nand U4064 (N_4064,N_3954,N_3958);
nor U4065 (N_4065,N_3767,N_3616);
nand U4066 (N_4066,N_3528,N_3547);
nor U4067 (N_4067,N_3859,N_3649);
nor U4068 (N_4068,N_3976,N_3554);
or U4069 (N_4069,N_3862,N_3777);
nand U4070 (N_4070,N_3631,N_3623);
or U4071 (N_4071,N_3760,N_3720);
nor U4072 (N_4072,N_3591,N_3503);
xnor U4073 (N_4073,N_3984,N_3639);
xnor U4074 (N_4074,N_3731,N_3907);
or U4075 (N_4075,N_3951,N_3690);
nand U4076 (N_4076,N_3879,N_3974);
and U4077 (N_4077,N_3993,N_3789);
or U4078 (N_4078,N_3540,N_3884);
nor U4079 (N_4079,N_3807,N_3944);
xor U4080 (N_4080,N_3652,N_3970);
nand U4081 (N_4081,N_3632,N_3557);
xor U4082 (N_4082,N_3903,N_3959);
nor U4083 (N_4083,N_3711,N_3501);
nand U4084 (N_4084,N_3737,N_3772);
xor U4085 (N_4085,N_3679,N_3526);
and U4086 (N_4086,N_3541,N_3820);
or U4087 (N_4087,N_3529,N_3935);
and U4088 (N_4088,N_3843,N_3904);
nand U4089 (N_4089,N_3983,N_3590);
or U4090 (N_4090,N_3773,N_3571);
and U4091 (N_4091,N_3733,N_3535);
nand U4092 (N_4092,N_3872,N_3781);
nand U4093 (N_4093,N_3707,N_3751);
xor U4094 (N_4094,N_3588,N_3896);
and U4095 (N_4095,N_3555,N_3586);
xnor U4096 (N_4096,N_3721,N_3712);
and U4097 (N_4097,N_3536,N_3930);
nor U4098 (N_4098,N_3792,N_3565);
or U4099 (N_4099,N_3577,N_3834);
nor U4100 (N_4100,N_3664,N_3854);
and U4101 (N_4101,N_3934,N_3923);
xor U4102 (N_4102,N_3505,N_3546);
or U4103 (N_4103,N_3646,N_3597);
nand U4104 (N_4104,N_3835,N_3663);
and U4105 (N_4105,N_3674,N_3919);
nand U4106 (N_4106,N_3573,N_3961);
nor U4107 (N_4107,N_3932,N_3782);
nand U4108 (N_4108,N_3867,N_3510);
and U4109 (N_4109,N_3850,N_3880);
and U4110 (N_4110,N_3689,N_3682);
or U4111 (N_4111,N_3809,N_3515);
xor U4112 (N_4112,N_3525,N_3818);
nand U4113 (N_4113,N_3582,N_3619);
nand U4114 (N_4114,N_3625,N_3977);
nor U4115 (N_4115,N_3783,N_3965);
or U4116 (N_4116,N_3956,N_3776);
nand U4117 (N_4117,N_3740,N_3939);
xor U4118 (N_4118,N_3543,N_3801);
or U4119 (N_4119,N_3701,N_3936);
xnor U4120 (N_4120,N_3757,N_3764);
nand U4121 (N_4121,N_3635,N_3603);
or U4122 (N_4122,N_3660,N_3698);
nand U4123 (N_4123,N_3502,N_3892);
nand U4124 (N_4124,N_3785,N_3730);
xor U4125 (N_4125,N_3592,N_3864);
xor U4126 (N_4126,N_3980,N_3614);
xnor U4127 (N_4127,N_3532,N_3742);
and U4128 (N_4128,N_3618,N_3840);
and U4129 (N_4129,N_3622,N_3659);
nor U4130 (N_4130,N_3717,N_3855);
and U4131 (N_4131,N_3790,N_3671);
and U4132 (N_4132,N_3898,N_3885);
nor U4133 (N_4133,N_3931,N_3887);
xnor U4134 (N_4134,N_3756,N_3596);
and U4135 (N_4135,N_3519,N_3561);
and U4136 (N_4136,N_3836,N_3500);
and U4137 (N_4137,N_3545,N_3658);
xor U4138 (N_4138,N_3681,N_3926);
or U4139 (N_4139,N_3687,N_3645);
nand U4140 (N_4140,N_3627,N_3873);
or U4141 (N_4141,N_3824,N_3726);
nand U4142 (N_4142,N_3553,N_3722);
xnor U4143 (N_4143,N_3787,N_3986);
and U4144 (N_4144,N_3810,N_3762);
or U4145 (N_4145,N_3704,N_3816);
xnor U4146 (N_4146,N_3856,N_3814);
nand U4147 (N_4147,N_3673,N_3985);
nand U4148 (N_4148,N_3677,N_3826);
or U4149 (N_4149,N_3968,N_3564);
and U4150 (N_4150,N_3696,N_3902);
and U4151 (N_4151,N_3665,N_3517);
xnor U4152 (N_4152,N_3694,N_3791);
nor U4153 (N_4153,N_3612,N_3727);
or U4154 (N_4154,N_3949,N_3516);
and U4155 (N_4155,N_3981,N_3888);
xnor U4156 (N_4156,N_3560,N_3613);
and U4157 (N_4157,N_3793,N_3666);
xor U4158 (N_4158,N_3890,N_3551);
nor U4159 (N_4159,N_3562,N_3839);
xnor U4160 (N_4160,N_3802,N_3874);
nand U4161 (N_4161,N_3530,N_3863);
nor U4162 (N_4162,N_3655,N_3544);
or U4163 (N_4163,N_3765,N_3771);
nor U4164 (N_4164,N_3754,N_3927);
nor U4165 (N_4165,N_3539,N_3708);
and U4166 (N_4166,N_3583,N_3638);
and U4167 (N_4167,N_3558,N_3744);
or U4168 (N_4168,N_3943,N_3837);
xor U4169 (N_4169,N_3769,N_3506);
xnor U4170 (N_4170,N_3811,N_3861);
nor U4171 (N_4171,N_3914,N_3714);
and U4172 (N_4172,N_3523,N_3642);
nand U4173 (N_4173,N_3606,N_3870);
nor U4174 (N_4174,N_3522,N_3942);
or U4175 (N_4175,N_3825,N_3803);
and U4176 (N_4176,N_3832,N_3725);
and U4177 (N_4177,N_3718,N_3531);
nor U4178 (N_4178,N_3905,N_3574);
nand U4179 (N_4179,N_3901,N_3972);
xnor U4180 (N_4180,N_3568,N_3640);
nor U4181 (N_4181,N_3739,N_3581);
nand U4182 (N_4182,N_3563,N_3598);
nand U4183 (N_4183,N_3812,N_3699);
nor U4184 (N_4184,N_3620,N_3925);
xor U4185 (N_4185,N_3589,N_3994);
nor U4186 (N_4186,N_3688,N_3800);
and U4187 (N_4187,N_3678,N_3786);
and U4188 (N_4188,N_3997,N_3922);
and U4189 (N_4189,N_3969,N_3709);
or U4190 (N_4190,N_3778,N_3542);
xnor U4191 (N_4191,N_3831,N_3798);
or U4192 (N_4192,N_3602,N_3946);
and U4193 (N_4193,N_3615,N_3774);
and U4194 (N_4194,N_3752,N_3527);
or U4195 (N_4195,N_3657,N_3685);
xor U4196 (N_4196,N_3846,N_3587);
or U4197 (N_4197,N_3991,N_3706);
nand U4198 (N_4198,N_3509,N_3669);
xnor U4199 (N_4199,N_3630,N_3734);
and U4200 (N_4200,N_3741,N_3775);
or U4201 (N_4201,N_3860,N_3924);
nand U4202 (N_4202,N_3869,N_3697);
and U4203 (N_4203,N_3680,N_3676);
and U4204 (N_4204,N_3748,N_3950);
nor U4205 (N_4205,N_3847,N_3845);
nand U4206 (N_4206,N_3755,N_3512);
nand U4207 (N_4207,N_3567,N_3514);
and U4208 (N_4208,N_3524,N_3728);
xnor U4209 (N_4209,N_3838,N_3691);
nand U4210 (N_4210,N_3987,N_3636);
nor U4211 (N_4211,N_3683,N_3975);
nor U4212 (N_4212,N_3609,N_3906);
nor U4213 (N_4213,N_3715,N_3920);
or U4214 (N_4214,N_3784,N_3611);
and U4215 (N_4215,N_3964,N_3610);
nor U4216 (N_4216,N_3750,N_3866);
xnor U4217 (N_4217,N_3953,N_3735);
xor U4218 (N_4218,N_3895,N_3667);
and U4219 (N_4219,N_3641,N_3670);
xnor U4220 (N_4220,N_3948,N_3780);
nand U4221 (N_4221,N_3556,N_3520);
and U4222 (N_4222,N_3912,N_3537);
or U4223 (N_4223,N_3633,N_3693);
or U4224 (N_4224,N_3578,N_3626);
xnor U4225 (N_4225,N_3908,N_3584);
or U4226 (N_4226,N_3533,N_3700);
and U4227 (N_4227,N_3675,N_3947);
nor U4228 (N_4228,N_3962,N_3713);
or U4229 (N_4229,N_3759,N_3511);
and U4230 (N_4230,N_3921,N_3600);
nand U4231 (N_4231,N_3841,N_3604);
and U4232 (N_4232,N_3668,N_3656);
or U4233 (N_4233,N_3957,N_3875);
and U4234 (N_4234,N_3882,N_3695);
nand U4235 (N_4235,N_3851,N_3899);
nand U4236 (N_4236,N_3736,N_3952);
and U4237 (N_4237,N_3822,N_3788);
nand U4238 (N_4238,N_3570,N_3766);
and U4239 (N_4239,N_3758,N_3662);
or U4240 (N_4240,N_3889,N_3806);
nand U4241 (N_4241,N_3702,N_3738);
and U4242 (N_4242,N_3940,N_3648);
nand U4243 (N_4243,N_3518,N_3971);
xnor U4244 (N_4244,N_3998,N_3550);
or U4245 (N_4245,N_3745,N_3605);
and U4246 (N_4246,N_3945,N_3794);
nand U4247 (N_4247,N_3580,N_3628);
and U4248 (N_4248,N_3799,N_3594);
nand U4249 (N_4249,N_3705,N_3815);
nor U4250 (N_4250,N_3639,N_3913);
nor U4251 (N_4251,N_3566,N_3509);
and U4252 (N_4252,N_3587,N_3908);
and U4253 (N_4253,N_3964,N_3618);
and U4254 (N_4254,N_3922,N_3540);
nor U4255 (N_4255,N_3523,N_3808);
nor U4256 (N_4256,N_3805,N_3950);
or U4257 (N_4257,N_3769,N_3609);
or U4258 (N_4258,N_3676,N_3963);
nor U4259 (N_4259,N_3559,N_3804);
nor U4260 (N_4260,N_3729,N_3593);
xnor U4261 (N_4261,N_3678,N_3880);
nor U4262 (N_4262,N_3981,N_3571);
xor U4263 (N_4263,N_3516,N_3865);
or U4264 (N_4264,N_3792,N_3536);
and U4265 (N_4265,N_3688,N_3823);
xnor U4266 (N_4266,N_3914,N_3860);
or U4267 (N_4267,N_3525,N_3529);
nand U4268 (N_4268,N_3601,N_3502);
nand U4269 (N_4269,N_3839,N_3790);
or U4270 (N_4270,N_3839,N_3789);
nor U4271 (N_4271,N_3995,N_3632);
and U4272 (N_4272,N_3722,N_3789);
and U4273 (N_4273,N_3623,N_3975);
nor U4274 (N_4274,N_3634,N_3819);
xnor U4275 (N_4275,N_3592,N_3863);
or U4276 (N_4276,N_3717,N_3980);
and U4277 (N_4277,N_3994,N_3555);
nor U4278 (N_4278,N_3639,N_3972);
and U4279 (N_4279,N_3629,N_3948);
xnor U4280 (N_4280,N_3759,N_3614);
xnor U4281 (N_4281,N_3866,N_3610);
xnor U4282 (N_4282,N_3899,N_3661);
and U4283 (N_4283,N_3941,N_3840);
nor U4284 (N_4284,N_3989,N_3973);
and U4285 (N_4285,N_3530,N_3679);
or U4286 (N_4286,N_3535,N_3678);
or U4287 (N_4287,N_3753,N_3540);
xnor U4288 (N_4288,N_3544,N_3710);
or U4289 (N_4289,N_3627,N_3856);
xnor U4290 (N_4290,N_3780,N_3847);
nor U4291 (N_4291,N_3568,N_3671);
or U4292 (N_4292,N_3969,N_3971);
and U4293 (N_4293,N_3557,N_3595);
and U4294 (N_4294,N_3734,N_3676);
xor U4295 (N_4295,N_3635,N_3883);
or U4296 (N_4296,N_3666,N_3769);
and U4297 (N_4297,N_3638,N_3946);
and U4298 (N_4298,N_3814,N_3900);
or U4299 (N_4299,N_3966,N_3737);
nor U4300 (N_4300,N_3899,N_3987);
xnor U4301 (N_4301,N_3515,N_3846);
xor U4302 (N_4302,N_3978,N_3768);
and U4303 (N_4303,N_3657,N_3505);
nand U4304 (N_4304,N_3585,N_3793);
nor U4305 (N_4305,N_3593,N_3624);
nand U4306 (N_4306,N_3661,N_3742);
nor U4307 (N_4307,N_3860,N_3611);
nand U4308 (N_4308,N_3835,N_3830);
or U4309 (N_4309,N_3716,N_3547);
nand U4310 (N_4310,N_3805,N_3572);
nor U4311 (N_4311,N_3962,N_3823);
nor U4312 (N_4312,N_3690,N_3599);
xor U4313 (N_4313,N_3841,N_3989);
and U4314 (N_4314,N_3945,N_3918);
nand U4315 (N_4315,N_3736,N_3751);
nand U4316 (N_4316,N_3756,N_3643);
or U4317 (N_4317,N_3851,N_3864);
xor U4318 (N_4318,N_3511,N_3717);
and U4319 (N_4319,N_3996,N_3773);
nand U4320 (N_4320,N_3749,N_3588);
and U4321 (N_4321,N_3673,N_3519);
nor U4322 (N_4322,N_3970,N_3799);
nand U4323 (N_4323,N_3932,N_3873);
nand U4324 (N_4324,N_3727,N_3891);
or U4325 (N_4325,N_3622,N_3705);
xnor U4326 (N_4326,N_3617,N_3996);
nand U4327 (N_4327,N_3653,N_3650);
xnor U4328 (N_4328,N_3637,N_3914);
nor U4329 (N_4329,N_3803,N_3826);
xor U4330 (N_4330,N_3551,N_3881);
nor U4331 (N_4331,N_3999,N_3581);
xor U4332 (N_4332,N_3993,N_3670);
xor U4333 (N_4333,N_3587,N_3827);
and U4334 (N_4334,N_3843,N_3987);
nor U4335 (N_4335,N_3561,N_3719);
nor U4336 (N_4336,N_3515,N_3597);
or U4337 (N_4337,N_3647,N_3929);
and U4338 (N_4338,N_3828,N_3965);
nand U4339 (N_4339,N_3819,N_3742);
xor U4340 (N_4340,N_3884,N_3815);
and U4341 (N_4341,N_3971,N_3682);
nand U4342 (N_4342,N_3711,N_3549);
nor U4343 (N_4343,N_3595,N_3986);
and U4344 (N_4344,N_3658,N_3744);
nor U4345 (N_4345,N_3866,N_3533);
or U4346 (N_4346,N_3859,N_3788);
or U4347 (N_4347,N_3941,N_3808);
nand U4348 (N_4348,N_3565,N_3705);
or U4349 (N_4349,N_3846,N_3980);
nor U4350 (N_4350,N_3632,N_3534);
nand U4351 (N_4351,N_3901,N_3580);
nor U4352 (N_4352,N_3853,N_3701);
and U4353 (N_4353,N_3545,N_3727);
xor U4354 (N_4354,N_3784,N_3608);
and U4355 (N_4355,N_3644,N_3709);
xor U4356 (N_4356,N_3646,N_3566);
xor U4357 (N_4357,N_3983,N_3912);
xnor U4358 (N_4358,N_3669,N_3675);
nand U4359 (N_4359,N_3716,N_3965);
xnor U4360 (N_4360,N_3833,N_3942);
or U4361 (N_4361,N_3802,N_3610);
or U4362 (N_4362,N_3626,N_3766);
nor U4363 (N_4363,N_3938,N_3795);
or U4364 (N_4364,N_3823,N_3658);
nor U4365 (N_4365,N_3842,N_3720);
or U4366 (N_4366,N_3685,N_3522);
nor U4367 (N_4367,N_3502,N_3997);
and U4368 (N_4368,N_3690,N_3906);
xnor U4369 (N_4369,N_3699,N_3741);
nor U4370 (N_4370,N_3775,N_3945);
nand U4371 (N_4371,N_3579,N_3613);
xor U4372 (N_4372,N_3633,N_3891);
xnor U4373 (N_4373,N_3862,N_3627);
xor U4374 (N_4374,N_3769,N_3626);
nor U4375 (N_4375,N_3693,N_3675);
and U4376 (N_4376,N_3708,N_3808);
nor U4377 (N_4377,N_3922,N_3637);
nor U4378 (N_4378,N_3659,N_3663);
or U4379 (N_4379,N_3580,N_3906);
or U4380 (N_4380,N_3919,N_3598);
or U4381 (N_4381,N_3708,N_3880);
and U4382 (N_4382,N_3906,N_3981);
nand U4383 (N_4383,N_3698,N_3828);
nor U4384 (N_4384,N_3782,N_3625);
xnor U4385 (N_4385,N_3699,N_3920);
or U4386 (N_4386,N_3508,N_3775);
and U4387 (N_4387,N_3516,N_3820);
nor U4388 (N_4388,N_3559,N_3884);
xnor U4389 (N_4389,N_3508,N_3513);
nand U4390 (N_4390,N_3836,N_3954);
nand U4391 (N_4391,N_3800,N_3641);
or U4392 (N_4392,N_3748,N_3537);
nand U4393 (N_4393,N_3501,N_3757);
nor U4394 (N_4394,N_3737,N_3647);
xnor U4395 (N_4395,N_3804,N_3698);
nand U4396 (N_4396,N_3825,N_3970);
nand U4397 (N_4397,N_3930,N_3769);
nand U4398 (N_4398,N_3916,N_3742);
xor U4399 (N_4399,N_3776,N_3600);
and U4400 (N_4400,N_3543,N_3857);
nor U4401 (N_4401,N_3665,N_3953);
and U4402 (N_4402,N_3772,N_3896);
nor U4403 (N_4403,N_3785,N_3841);
and U4404 (N_4404,N_3590,N_3703);
and U4405 (N_4405,N_3752,N_3762);
nor U4406 (N_4406,N_3503,N_3612);
or U4407 (N_4407,N_3594,N_3858);
and U4408 (N_4408,N_3579,N_3978);
or U4409 (N_4409,N_3814,N_3678);
xnor U4410 (N_4410,N_3899,N_3518);
xor U4411 (N_4411,N_3586,N_3574);
nand U4412 (N_4412,N_3734,N_3604);
or U4413 (N_4413,N_3606,N_3565);
or U4414 (N_4414,N_3669,N_3897);
xor U4415 (N_4415,N_3706,N_3993);
or U4416 (N_4416,N_3763,N_3654);
and U4417 (N_4417,N_3757,N_3799);
nor U4418 (N_4418,N_3655,N_3973);
xor U4419 (N_4419,N_3914,N_3507);
and U4420 (N_4420,N_3640,N_3996);
or U4421 (N_4421,N_3554,N_3821);
xnor U4422 (N_4422,N_3822,N_3665);
xnor U4423 (N_4423,N_3514,N_3588);
and U4424 (N_4424,N_3936,N_3914);
xor U4425 (N_4425,N_3551,N_3886);
xor U4426 (N_4426,N_3580,N_3947);
xnor U4427 (N_4427,N_3948,N_3715);
or U4428 (N_4428,N_3862,N_3772);
xnor U4429 (N_4429,N_3778,N_3833);
or U4430 (N_4430,N_3842,N_3887);
xor U4431 (N_4431,N_3740,N_3805);
and U4432 (N_4432,N_3841,N_3511);
and U4433 (N_4433,N_3796,N_3595);
nand U4434 (N_4434,N_3975,N_3932);
nor U4435 (N_4435,N_3696,N_3916);
nor U4436 (N_4436,N_3735,N_3703);
or U4437 (N_4437,N_3935,N_3688);
or U4438 (N_4438,N_3558,N_3806);
nand U4439 (N_4439,N_3884,N_3872);
xnor U4440 (N_4440,N_3554,N_3929);
nand U4441 (N_4441,N_3935,N_3771);
xor U4442 (N_4442,N_3995,N_3864);
xor U4443 (N_4443,N_3874,N_3895);
nor U4444 (N_4444,N_3754,N_3957);
nand U4445 (N_4445,N_3635,N_3517);
nand U4446 (N_4446,N_3608,N_3929);
nor U4447 (N_4447,N_3905,N_3820);
or U4448 (N_4448,N_3691,N_3656);
nor U4449 (N_4449,N_3724,N_3714);
nand U4450 (N_4450,N_3835,N_3956);
and U4451 (N_4451,N_3734,N_3567);
nor U4452 (N_4452,N_3646,N_3768);
or U4453 (N_4453,N_3738,N_3911);
or U4454 (N_4454,N_3860,N_3682);
nand U4455 (N_4455,N_3839,N_3720);
or U4456 (N_4456,N_3786,N_3542);
nor U4457 (N_4457,N_3539,N_3643);
nand U4458 (N_4458,N_3656,N_3905);
nand U4459 (N_4459,N_3739,N_3983);
or U4460 (N_4460,N_3925,N_3897);
nor U4461 (N_4461,N_3656,N_3703);
and U4462 (N_4462,N_3530,N_3924);
nand U4463 (N_4463,N_3617,N_3638);
xnor U4464 (N_4464,N_3557,N_3691);
and U4465 (N_4465,N_3510,N_3691);
xor U4466 (N_4466,N_3862,N_3653);
or U4467 (N_4467,N_3592,N_3556);
nor U4468 (N_4468,N_3716,N_3519);
nand U4469 (N_4469,N_3645,N_3989);
xor U4470 (N_4470,N_3730,N_3540);
and U4471 (N_4471,N_3825,N_3810);
nand U4472 (N_4472,N_3859,N_3912);
nor U4473 (N_4473,N_3913,N_3711);
xor U4474 (N_4474,N_3565,N_3866);
and U4475 (N_4475,N_3658,N_3930);
or U4476 (N_4476,N_3567,N_3603);
nand U4477 (N_4477,N_3706,N_3588);
nand U4478 (N_4478,N_3532,N_3954);
or U4479 (N_4479,N_3662,N_3790);
xnor U4480 (N_4480,N_3593,N_3594);
xor U4481 (N_4481,N_3892,N_3643);
or U4482 (N_4482,N_3727,N_3559);
xor U4483 (N_4483,N_3521,N_3633);
nor U4484 (N_4484,N_3755,N_3559);
xor U4485 (N_4485,N_3537,N_3875);
nor U4486 (N_4486,N_3539,N_3742);
or U4487 (N_4487,N_3759,N_3937);
and U4488 (N_4488,N_3534,N_3517);
nand U4489 (N_4489,N_3994,N_3903);
nand U4490 (N_4490,N_3851,N_3998);
nand U4491 (N_4491,N_3851,N_3984);
nor U4492 (N_4492,N_3621,N_3683);
or U4493 (N_4493,N_3680,N_3564);
and U4494 (N_4494,N_3781,N_3753);
and U4495 (N_4495,N_3911,N_3853);
and U4496 (N_4496,N_3874,N_3979);
or U4497 (N_4497,N_3613,N_3570);
or U4498 (N_4498,N_3859,N_3535);
and U4499 (N_4499,N_3694,N_3661);
nor U4500 (N_4500,N_4315,N_4195);
and U4501 (N_4501,N_4273,N_4251);
nor U4502 (N_4502,N_4083,N_4257);
or U4503 (N_4503,N_4067,N_4335);
and U4504 (N_4504,N_4129,N_4055);
and U4505 (N_4505,N_4248,N_4327);
or U4506 (N_4506,N_4252,N_4301);
nor U4507 (N_4507,N_4220,N_4143);
and U4508 (N_4508,N_4260,N_4425);
nor U4509 (N_4509,N_4118,N_4439);
xor U4510 (N_4510,N_4391,N_4107);
and U4511 (N_4511,N_4213,N_4087);
or U4512 (N_4512,N_4007,N_4111);
or U4513 (N_4513,N_4134,N_4006);
and U4514 (N_4514,N_4303,N_4126);
or U4515 (N_4515,N_4093,N_4194);
nand U4516 (N_4516,N_4418,N_4319);
nand U4517 (N_4517,N_4364,N_4215);
nor U4518 (N_4518,N_4116,N_4460);
or U4519 (N_4519,N_4230,N_4035);
nand U4520 (N_4520,N_4233,N_4001);
nor U4521 (N_4521,N_4125,N_4286);
nand U4522 (N_4522,N_4099,N_4472);
or U4523 (N_4523,N_4149,N_4376);
nand U4524 (N_4524,N_4312,N_4232);
nand U4525 (N_4525,N_4408,N_4467);
or U4526 (N_4526,N_4123,N_4333);
nor U4527 (N_4527,N_4407,N_4427);
nor U4528 (N_4528,N_4174,N_4110);
nor U4529 (N_4529,N_4234,N_4399);
or U4530 (N_4530,N_4245,N_4026);
xnor U4531 (N_4531,N_4019,N_4272);
nor U4532 (N_4532,N_4043,N_4189);
nor U4533 (N_4533,N_4314,N_4293);
or U4534 (N_4534,N_4361,N_4036);
xnor U4535 (N_4535,N_4112,N_4449);
or U4536 (N_4536,N_4255,N_4154);
nor U4537 (N_4537,N_4323,N_4414);
xnor U4538 (N_4538,N_4211,N_4253);
xnor U4539 (N_4539,N_4290,N_4150);
and U4540 (N_4540,N_4196,N_4104);
xnor U4541 (N_4541,N_4358,N_4404);
nand U4542 (N_4542,N_4012,N_4294);
or U4543 (N_4543,N_4121,N_4365);
and U4544 (N_4544,N_4038,N_4400);
nor U4545 (N_4545,N_4015,N_4127);
nand U4546 (N_4546,N_4002,N_4435);
and U4547 (N_4547,N_4451,N_4448);
and U4548 (N_4548,N_4155,N_4373);
nor U4549 (N_4549,N_4031,N_4113);
xnor U4550 (N_4550,N_4442,N_4170);
or U4551 (N_4551,N_4167,N_4218);
xnor U4552 (N_4552,N_4094,N_4160);
and U4553 (N_4553,N_4000,N_4354);
xor U4554 (N_4554,N_4275,N_4090);
nor U4555 (N_4555,N_4047,N_4324);
nor U4556 (N_4556,N_4056,N_4080);
xor U4557 (N_4557,N_4289,N_4428);
xor U4558 (N_4558,N_4464,N_4025);
xnor U4559 (N_4559,N_4236,N_4406);
or U4560 (N_4560,N_4142,N_4356);
xor U4561 (N_4561,N_4417,N_4276);
nor U4562 (N_4562,N_4095,N_4355);
and U4563 (N_4563,N_4059,N_4359);
xor U4564 (N_4564,N_4077,N_4393);
nand U4565 (N_4565,N_4326,N_4420);
or U4566 (N_4566,N_4225,N_4307);
nand U4567 (N_4567,N_4139,N_4309);
and U4568 (N_4568,N_4071,N_4483);
nand U4569 (N_4569,N_4302,N_4264);
xnor U4570 (N_4570,N_4222,N_4370);
nor U4571 (N_4571,N_4117,N_4197);
xor U4572 (N_4572,N_4362,N_4413);
and U4573 (N_4573,N_4488,N_4469);
or U4574 (N_4574,N_4453,N_4088);
or U4575 (N_4575,N_4279,N_4446);
or U4576 (N_4576,N_4369,N_4148);
or U4577 (N_4577,N_4239,N_4402);
nand U4578 (N_4578,N_4024,N_4168);
and U4579 (N_4579,N_4054,N_4203);
nor U4580 (N_4580,N_4396,N_4482);
nand U4581 (N_4581,N_4076,N_4032);
nor U4582 (N_4582,N_4023,N_4092);
nor U4583 (N_4583,N_4052,N_4045);
and U4584 (N_4584,N_4124,N_4228);
and U4585 (N_4585,N_4291,N_4422);
or U4586 (N_4586,N_4388,N_4351);
and U4587 (N_4587,N_4332,N_4183);
and U4588 (N_4588,N_4171,N_4336);
nand U4589 (N_4589,N_4454,N_4156);
or U4590 (N_4590,N_4141,N_4489);
nand U4591 (N_4591,N_4157,N_4325);
or U4592 (N_4592,N_4177,N_4034);
nor U4593 (N_4593,N_4205,N_4219);
and U4594 (N_4594,N_4295,N_4221);
or U4595 (N_4595,N_4473,N_4374);
and U4596 (N_4596,N_4386,N_4193);
xnor U4597 (N_4597,N_4444,N_4178);
xor U4598 (N_4598,N_4337,N_4072);
xor U4599 (N_4599,N_4062,N_4204);
nand U4600 (N_4600,N_4162,N_4310);
xor U4601 (N_4601,N_4341,N_4097);
nor U4602 (N_4602,N_4020,N_4456);
and U4603 (N_4603,N_4050,N_4046);
or U4604 (N_4604,N_4053,N_4186);
nand U4605 (N_4605,N_4210,N_4101);
xnor U4606 (N_4606,N_4223,N_4188);
or U4607 (N_4607,N_4438,N_4089);
nor U4608 (N_4608,N_4136,N_4411);
and U4609 (N_4609,N_4190,N_4287);
xnor U4610 (N_4610,N_4263,N_4037);
nand U4611 (N_4611,N_4468,N_4022);
xnor U4612 (N_4612,N_4209,N_4334);
or U4613 (N_4613,N_4200,N_4256);
nand U4614 (N_4614,N_4497,N_4165);
nand U4615 (N_4615,N_4330,N_4366);
nand U4616 (N_4616,N_4108,N_4119);
and U4617 (N_4617,N_4145,N_4202);
and U4618 (N_4618,N_4070,N_4246);
xor U4619 (N_4619,N_4383,N_4216);
nand U4620 (N_4620,N_4014,N_4135);
xor U4621 (N_4621,N_4360,N_4207);
nor U4622 (N_4622,N_4387,N_4426);
or U4623 (N_4623,N_4419,N_4100);
nand U4624 (N_4624,N_4085,N_4176);
or U4625 (N_4625,N_4440,N_4492);
and U4626 (N_4626,N_4231,N_4131);
nand U4627 (N_4627,N_4465,N_4086);
nor U4628 (N_4628,N_4328,N_4184);
xnor U4629 (N_4629,N_4380,N_4133);
nand U4630 (N_4630,N_4270,N_4470);
and U4631 (N_4631,N_4267,N_4033);
nand U4632 (N_4632,N_4172,N_4284);
or U4633 (N_4633,N_4159,N_4410);
or U4634 (N_4634,N_4152,N_4029);
or U4635 (N_4635,N_4227,N_4350);
nor U4636 (N_4636,N_4318,N_4068);
and U4637 (N_4637,N_4430,N_4181);
or U4638 (N_4638,N_4340,N_4283);
nor U4639 (N_4639,N_4058,N_4238);
xor U4640 (N_4640,N_4348,N_4079);
nor U4641 (N_4641,N_4028,N_4214);
or U4642 (N_4642,N_4229,N_4201);
xnor U4643 (N_4643,N_4182,N_4030);
or U4644 (N_4644,N_4173,N_4415);
and U4645 (N_4645,N_4445,N_4405);
or U4646 (N_4646,N_4421,N_4441);
and U4647 (N_4647,N_4300,N_4437);
nor U4648 (N_4648,N_4115,N_4353);
or U4649 (N_4649,N_4065,N_4049);
nor U4650 (N_4650,N_4423,N_4306);
xnor U4651 (N_4651,N_4192,N_4431);
and U4652 (N_4652,N_4485,N_4494);
nand U4653 (N_4653,N_4384,N_4109);
nand U4654 (N_4654,N_4144,N_4475);
xor U4655 (N_4655,N_4042,N_4471);
and U4656 (N_4656,N_4495,N_4243);
or U4657 (N_4657,N_4039,N_4329);
nand U4658 (N_4658,N_4061,N_4164);
and U4659 (N_4659,N_4098,N_4389);
xnor U4660 (N_4660,N_4169,N_4320);
nand U4661 (N_4661,N_4381,N_4122);
or U4662 (N_4662,N_4292,N_4249);
or U4663 (N_4663,N_4132,N_4392);
or U4664 (N_4664,N_4258,N_4147);
nand U4665 (N_4665,N_4371,N_4140);
or U4666 (N_4666,N_4322,N_4128);
nand U4667 (N_4667,N_4321,N_4259);
nor U4668 (N_4668,N_4463,N_4146);
nor U4669 (N_4669,N_4277,N_4208);
nand U4670 (N_4670,N_4297,N_4005);
xnor U4671 (N_4671,N_4048,N_4455);
or U4672 (N_4672,N_4349,N_4274);
nand U4673 (N_4673,N_4305,N_4352);
xor U4674 (N_4674,N_4345,N_4018);
xnor U4675 (N_4675,N_4447,N_4476);
nand U4676 (N_4676,N_4241,N_4308);
xnor U4677 (N_4677,N_4363,N_4479);
xnor U4678 (N_4678,N_4344,N_4016);
xnor U4679 (N_4679,N_4226,N_4316);
xor U4680 (N_4680,N_4271,N_4066);
and U4681 (N_4681,N_4382,N_4385);
xor U4682 (N_4682,N_4187,N_4106);
nand U4683 (N_4683,N_4161,N_4466);
or U4684 (N_4684,N_4429,N_4191);
nor U4685 (N_4685,N_4436,N_4212);
and U4686 (N_4686,N_4346,N_4397);
xor U4687 (N_4687,N_4285,N_4452);
or U4688 (N_4688,N_4368,N_4008);
and U4689 (N_4689,N_4158,N_4069);
nor U4690 (N_4690,N_4261,N_4247);
nand U4691 (N_4691,N_4013,N_4331);
and U4692 (N_4692,N_4102,N_4394);
and U4693 (N_4693,N_4011,N_4051);
nor U4694 (N_4694,N_4244,N_4130);
nor U4695 (N_4695,N_4199,N_4498);
or U4696 (N_4696,N_4487,N_4484);
or U4697 (N_4697,N_4317,N_4450);
nand U4698 (N_4698,N_4403,N_4462);
xnor U4699 (N_4699,N_4217,N_4338);
and U4700 (N_4700,N_4010,N_4237);
or U4701 (N_4701,N_4390,N_4278);
nor U4702 (N_4702,N_4457,N_4073);
xor U4703 (N_4703,N_4240,N_4235);
xor U4704 (N_4704,N_4490,N_4084);
and U4705 (N_4705,N_4416,N_4105);
xnor U4706 (N_4706,N_4311,N_4343);
or U4707 (N_4707,N_4281,N_4153);
nor U4708 (N_4708,N_4004,N_4224);
xnor U4709 (N_4709,N_4206,N_4091);
xnor U4710 (N_4710,N_4480,N_4461);
nor U4711 (N_4711,N_4040,N_4268);
xor U4712 (N_4712,N_4003,N_4296);
nand U4713 (N_4713,N_4474,N_4378);
xor U4714 (N_4714,N_4103,N_4009);
xnor U4715 (N_4715,N_4282,N_4313);
nor U4716 (N_4716,N_4075,N_4179);
nor U4717 (N_4717,N_4044,N_4262);
nor U4718 (N_4718,N_4180,N_4163);
xor U4719 (N_4719,N_4458,N_4078);
and U4720 (N_4720,N_4082,N_4481);
or U4721 (N_4721,N_4342,N_4432);
or U4722 (N_4722,N_4347,N_4138);
and U4723 (N_4723,N_4493,N_4063);
nor U4724 (N_4724,N_4096,N_4057);
nor U4725 (N_4725,N_4120,N_4434);
or U4726 (N_4726,N_4409,N_4372);
and U4727 (N_4727,N_4298,N_4041);
or U4728 (N_4728,N_4357,N_4242);
and U4729 (N_4729,N_4395,N_4250);
and U4730 (N_4730,N_4074,N_4269);
nor U4731 (N_4731,N_4175,N_4491);
and U4732 (N_4732,N_4114,N_4137);
and U4733 (N_4733,N_4401,N_4299);
xor U4734 (N_4734,N_4375,N_4443);
nand U4735 (N_4735,N_4254,N_4377);
nand U4736 (N_4736,N_4151,N_4304);
and U4737 (N_4737,N_4477,N_4265);
or U4738 (N_4738,N_4166,N_4185);
or U4739 (N_4739,N_4081,N_4060);
xnor U4740 (N_4740,N_4367,N_4379);
xnor U4741 (N_4741,N_4017,N_4288);
nand U4742 (N_4742,N_4280,N_4496);
nand U4743 (N_4743,N_4398,N_4266);
nand U4744 (N_4744,N_4021,N_4027);
xnor U4745 (N_4745,N_4412,N_4486);
nand U4746 (N_4746,N_4433,N_4339);
or U4747 (N_4747,N_4499,N_4424);
or U4748 (N_4748,N_4478,N_4198);
nor U4749 (N_4749,N_4459,N_4064);
xor U4750 (N_4750,N_4072,N_4344);
xor U4751 (N_4751,N_4152,N_4440);
or U4752 (N_4752,N_4329,N_4383);
nor U4753 (N_4753,N_4184,N_4401);
and U4754 (N_4754,N_4317,N_4420);
or U4755 (N_4755,N_4486,N_4297);
and U4756 (N_4756,N_4224,N_4205);
nor U4757 (N_4757,N_4197,N_4409);
nor U4758 (N_4758,N_4319,N_4044);
nand U4759 (N_4759,N_4204,N_4277);
xor U4760 (N_4760,N_4256,N_4039);
nand U4761 (N_4761,N_4145,N_4114);
nand U4762 (N_4762,N_4231,N_4155);
nand U4763 (N_4763,N_4249,N_4372);
or U4764 (N_4764,N_4230,N_4066);
nand U4765 (N_4765,N_4037,N_4228);
and U4766 (N_4766,N_4272,N_4309);
nand U4767 (N_4767,N_4379,N_4321);
xnor U4768 (N_4768,N_4152,N_4250);
nor U4769 (N_4769,N_4169,N_4001);
nor U4770 (N_4770,N_4457,N_4415);
or U4771 (N_4771,N_4346,N_4003);
nand U4772 (N_4772,N_4198,N_4255);
nor U4773 (N_4773,N_4119,N_4397);
nand U4774 (N_4774,N_4090,N_4420);
nand U4775 (N_4775,N_4398,N_4086);
and U4776 (N_4776,N_4200,N_4142);
or U4777 (N_4777,N_4451,N_4051);
nand U4778 (N_4778,N_4417,N_4168);
or U4779 (N_4779,N_4097,N_4194);
xor U4780 (N_4780,N_4029,N_4008);
xor U4781 (N_4781,N_4452,N_4492);
xor U4782 (N_4782,N_4168,N_4038);
or U4783 (N_4783,N_4328,N_4398);
and U4784 (N_4784,N_4007,N_4057);
nor U4785 (N_4785,N_4245,N_4136);
or U4786 (N_4786,N_4219,N_4095);
nand U4787 (N_4787,N_4125,N_4029);
nor U4788 (N_4788,N_4241,N_4089);
and U4789 (N_4789,N_4322,N_4089);
xnor U4790 (N_4790,N_4142,N_4129);
nand U4791 (N_4791,N_4346,N_4019);
xnor U4792 (N_4792,N_4320,N_4407);
nor U4793 (N_4793,N_4293,N_4331);
and U4794 (N_4794,N_4211,N_4304);
xor U4795 (N_4795,N_4109,N_4135);
nor U4796 (N_4796,N_4315,N_4057);
xnor U4797 (N_4797,N_4113,N_4218);
or U4798 (N_4798,N_4423,N_4157);
and U4799 (N_4799,N_4131,N_4055);
xor U4800 (N_4800,N_4425,N_4375);
nand U4801 (N_4801,N_4476,N_4029);
and U4802 (N_4802,N_4202,N_4050);
nand U4803 (N_4803,N_4142,N_4427);
xnor U4804 (N_4804,N_4032,N_4297);
and U4805 (N_4805,N_4075,N_4154);
and U4806 (N_4806,N_4273,N_4313);
and U4807 (N_4807,N_4179,N_4350);
nor U4808 (N_4808,N_4054,N_4023);
and U4809 (N_4809,N_4276,N_4080);
xor U4810 (N_4810,N_4136,N_4135);
and U4811 (N_4811,N_4459,N_4413);
nand U4812 (N_4812,N_4422,N_4031);
nor U4813 (N_4813,N_4193,N_4285);
or U4814 (N_4814,N_4218,N_4436);
xor U4815 (N_4815,N_4199,N_4453);
xor U4816 (N_4816,N_4435,N_4347);
xor U4817 (N_4817,N_4156,N_4054);
or U4818 (N_4818,N_4107,N_4201);
and U4819 (N_4819,N_4156,N_4341);
or U4820 (N_4820,N_4170,N_4490);
and U4821 (N_4821,N_4092,N_4356);
nand U4822 (N_4822,N_4031,N_4483);
xnor U4823 (N_4823,N_4066,N_4398);
or U4824 (N_4824,N_4310,N_4037);
or U4825 (N_4825,N_4411,N_4048);
nand U4826 (N_4826,N_4351,N_4374);
or U4827 (N_4827,N_4329,N_4402);
nor U4828 (N_4828,N_4370,N_4352);
nand U4829 (N_4829,N_4458,N_4225);
nor U4830 (N_4830,N_4317,N_4308);
nand U4831 (N_4831,N_4125,N_4445);
and U4832 (N_4832,N_4450,N_4175);
xnor U4833 (N_4833,N_4418,N_4093);
or U4834 (N_4834,N_4494,N_4419);
xnor U4835 (N_4835,N_4287,N_4202);
nor U4836 (N_4836,N_4128,N_4218);
nor U4837 (N_4837,N_4212,N_4013);
nor U4838 (N_4838,N_4280,N_4003);
xnor U4839 (N_4839,N_4340,N_4358);
nand U4840 (N_4840,N_4054,N_4043);
xor U4841 (N_4841,N_4498,N_4455);
and U4842 (N_4842,N_4000,N_4067);
and U4843 (N_4843,N_4408,N_4147);
and U4844 (N_4844,N_4417,N_4286);
xnor U4845 (N_4845,N_4025,N_4122);
nand U4846 (N_4846,N_4283,N_4094);
and U4847 (N_4847,N_4156,N_4267);
xor U4848 (N_4848,N_4382,N_4010);
or U4849 (N_4849,N_4490,N_4453);
or U4850 (N_4850,N_4139,N_4451);
nor U4851 (N_4851,N_4338,N_4362);
nand U4852 (N_4852,N_4314,N_4127);
nand U4853 (N_4853,N_4219,N_4073);
xor U4854 (N_4854,N_4060,N_4153);
nor U4855 (N_4855,N_4499,N_4053);
or U4856 (N_4856,N_4385,N_4272);
or U4857 (N_4857,N_4424,N_4239);
nand U4858 (N_4858,N_4249,N_4181);
xnor U4859 (N_4859,N_4358,N_4001);
and U4860 (N_4860,N_4157,N_4335);
nand U4861 (N_4861,N_4336,N_4005);
or U4862 (N_4862,N_4473,N_4062);
or U4863 (N_4863,N_4301,N_4458);
nand U4864 (N_4864,N_4152,N_4090);
and U4865 (N_4865,N_4196,N_4484);
nor U4866 (N_4866,N_4298,N_4240);
or U4867 (N_4867,N_4105,N_4384);
xor U4868 (N_4868,N_4043,N_4369);
and U4869 (N_4869,N_4241,N_4493);
xnor U4870 (N_4870,N_4482,N_4371);
xor U4871 (N_4871,N_4242,N_4018);
or U4872 (N_4872,N_4027,N_4324);
xnor U4873 (N_4873,N_4083,N_4301);
nor U4874 (N_4874,N_4162,N_4278);
or U4875 (N_4875,N_4381,N_4154);
and U4876 (N_4876,N_4111,N_4035);
nor U4877 (N_4877,N_4247,N_4025);
and U4878 (N_4878,N_4245,N_4392);
and U4879 (N_4879,N_4192,N_4168);
or U4880 (N_4880,N_4371,N_4336);
nand U4881 (N_4881,N_4113,N_4337);
nor U4882 (N_4882,N_4400,N_4371);
nor U4883 (N_4883,N_4362,N_4267);
and U4884 (N_4884,N_4300,N_4177);
or U4885 (N_4885,N_4395,N_4169);
or U4886 (N_4886,N_4432,N_4085);
xnor U4887 (N_4887,N_4464,N_4055);
nand U4888 (N_4888,N_4339,N_4224);
nor U4889 (N_4889,N_4111,N_4371);
or U4890 (N_4890,N_4146,N_4333);
xnor U4891 (N_4891,N_4304,N_4363);
or U4892 (N_4892,N_4189,N_4047);
nor U4893 (N_4893,N_4467,N_4184);
or U4894 (N_4894,N_4399,N_4473);
and U4895 (N_4895,N_4142,N_4034);
xnor U4896 (N_4896,N_4322,N_4260);
or U4897 (N_4897,N_4133,N_4021);
nor U4898 (N_4898,N_4248,N_4042);
and U4899 (N_4899,N_4482,N_4196);
nand U4900 (N_4900,N_4498,N_4346);
xor U4901 (N_4901,N_4132,N_4466);
xnor U4902 (N_4902,N_4031,N_4497);
and U4903 (N_4903,N_4383,N_4105);
nand U4904 (N_4904,N_4000,N_4372);
or U4905 (N_4905,N_4171,N_4495);
and U4906 (N_4906,N_4434,N_4327);
nor U4907 (N_4907,N_4413,N_4256);
and U4908 (N_4908,N_4281,N_4378);
and U4909 (N_4909,N_4145,N_4024);
or U4910 (N_4910,N_4419,N_4026);
nor U4911 (N_4911,N_4487,N_4002);
nand U4912 (N_4912,N_4236,N_4134);
nand U4913 (N_4913,N_4346,N_4171);
nor U4914 (N_4914,N_4265,N_4157);
xnor U4915 (N_4915,N_4071,N_4154);
or U4916 (N_4916,N_4051,N_4426);
xor U4917 (N_4917,N_4066,N_4323);
xor U4918 (N_4918,N_4060,N_4004);
and U4919 (N_4919,N_4367,N_4326);
nand U4920 (N_4920,N_4359,N_4397);
and U4921 (N_4921,N_4045,N_4491);
xnor U4922 (N_4922,N_4235,N_4136);
xnor U4923 (N_4923,N_4007,N_4054);
nand U4924 (N_4924,N_4495,N_4079);
nor U4925 (N_4925,N_4204,N_4245);
or U4926 (N_4926,N_4320,N_4345);
or U4927 (N_4927,N_4201,N_4046);
xor U4928 (N_4928,N_4356,N_4039);
and U4929 (N_4929,N_4056,N_4009);
nor U4930 (N_4930,N_4325,N_4326);
and U4931 (N_4931,N_4008,N_4198);
and U4932 (N_4932,N_4240,N_4075);
nor U4933 (N_4933,N_4257,N_4295);
nand U4934 (N_4934,N_4068,N_4418);
xor U4935 (N_4935,N_4175,N_4194);
nor U4936 (N_4936,N_4190,N_4397);
and U4937 (N_4937,N_4002,N_4341);
nand U4938 (N_4938,N_4309,N_4026);
or U4939 (N_4939,N_4381,N_4117);
xnor U4940 (N_4940,N_4127,N_4259);
and U4941 (N_4941,N_4119,N_4459);
nand U4942 (N_4942,N_4205,N_4372);
or U4943 (N_4943,N_4137,N_4351);
or U4944 (N_4944,N_4233,N_4223);
nor U4945 (N_4945,N_4212,N_4101);
nand U4946 (N_4946,N_4110,N_4487);
or U4947 (N_4947,N_4444,N_4009);
xnor U4948 (N_4948,N_4061,N_4297);
nand U4949 (N_4949,N_4274,N_4225);
xnor U4950 (N_4950,N_4490,N_4468);
nand U4951 (N_4951,N_4498,N_4073);
nand U4952 (N_4952,N_4015,N_4192);
xor U4953 (N_4953,N_4176,N_4427);
nand U4954 (N_4954,N_4266,N_4394);
or U4955 (N_4955,N_4154,N_4159);
nor U4956 (N_4956,N_4490,N_4287);
xnor U4957 (N_4957,N_4433,N_4471);
and U4958 (N_4958,N_4110,N_4172);
or U4959 (N_4959,N_4488,N_4418);
nor U4960 (N_4960,N_4406,N_4258);
or U4961 (N_4961,N_4498,N_4406);
or U4962 (N_4962,N_4464,N_4174);
and U4963 (N_4963,N_4489,N_4367);
xor U4964 (N_4964,N_4282,N_4302);
xor U4965 (N_4965,N_4005,N_4025);
xnor U4966 (N_4966,N_4259,N_4341);
nor U4967 (N_4967,N_4396,N_4041);
and U4968 (N_4968,N_4495,N_4343);
nor U4969 (N_4969,N_4370,N_4183);
nor U4970 (N_4970,N_4225,N_4198);
nand U4971 (N_4971,N_4131,N_4469);
nor U4972 (N_4972,N_4199,N_4292);
or U4973 (N_4973,N_4454,N_4088);
nand U4974 (N_4974,N_4143,N_4050);
or U4975 (N_4975,N_4337,N_4271);
xor U4976 (N_4976,N_4214,N_4382);
and U4977 (N_4977,N_4293,N_4332);
xor U4978 (N_4978,N_4370,N_4269);
and U4979 (N_4979,N_4486,N_4295);
nand U4980 (N_4980,N_4416,N_4037);
or U4981 (N_4981,N_4364,N_4311);
nor U4982 (N_4982,N_4362,N_4239);
or U4983 (N_4983,N_4008,N_4416);
or U4984 (N_4984,N_4248,N_4175);
xnor U4985 (N_4985,N_4351,N_4045);
nand U4986 (N_4986,N_4018,N_4112);
and U4987 (N_4987,N_4060,N_4427);
nor U4988 (N_4988,N_4062,N_4361);
and U4989 (N_4989,N_4485,N_4256);
and U4990 (N_4990,N_4028,N_4349);
nand U4991 (N_4991,N_4180,N_4009);
and U4992 (N_4992,N_4367,N_4350);
or U4993 (N_4993,N_4445,N_4490);
nor U4994 (N_4994,N_4288,N_4180);
xor U4995 (N_4995,N_4472,N_4020);
or U4996 (N_4996,N_4469,N_4338);
xor U4997 (N_4997,N_4268,N_4230);
nor U4998 (N_4998,N_4251,N_4215);
xnor U4999 (N_4999,N_4447,N_4481);
nand U5000 (N_5000,N_4573,N_4915);
xor U5001 (N_5001,N_4779,N_4791);
or U5002 (N_5002,N_4570,N_4877);
xnor U5003 (N_5003,N_4619,N_4898);
nand U5004 (N_5004,N_4902,N_4673);
nor U5005 (N_5005,N_4805,N_4895);
and U5006 (N_5006,N_4618,N_4714);
nand U5007 (N_5007,N_4996,N_4646);
nand U5008 (N_5008,N_4859,N_4800);
or U5009 (N_5009,N_4850,N_4732);
nand U5010 (N_5010,N_4807,N_4785);
and U5011 (N_5011,N_4706,N_4836);
nor U5012 (N_5012,N_4585,N_4775);
xor U5013 (N_5013,N_4802,N_4847);
xnor U5014 (N_5014,N_4599,N_4533);
nor U5015 (N_5015,N_4817,N_4739);
nor U5016 (N_5016,N_4955,N_4546);
nand U5017 (N_5017,N_4672,N_4645);
xnor U5018 (N_5018,N_4684,N_4629);
or U5019 (N_5019,N_4911,N_4989);
xnor U5020 (N_5020,N_4601,N_4505);
nand U5021 (N_5021,N_4889,N_4920);
xnor U5022 (N_5022,N_4951,N_4873);
and U5023 (N_5023,N_4874,N_4933);
xnor U5024 (N_5024,N_4880,N_4569);
nor U5025 (N_5025,N_4963,N_4829);
and U5026 (N_5026,N_4744,N_4832);
and U5027 (N_5027,N_4666,N_4509);
xnor U5028 (N_5028,N_4936,N_4690);
nor U5029 (N_5029,N_4658,N_4544);
and U5030 (N_5030,N_4980,N_4534);
and U5031 (N_5031,N_4710,N_4583);
xnor U5032 (N_5032,N_4649,N_4543);
or U5033 (N_5033,N_4537,N_4563);
or U5034 (N_5034,N_4592,N_4643);
nand U5035 (N_5035,N_4679,N_4532);
and U5036 (N_5036,N_4613,N_4598);
nor U5037 (N_5037,N_4635,N_4590);
and U5038 (N_5038,N_4753,N_4849);
nor U5039 (N_5039,N_4897,N_4667);
xnor U5040 (N_5040,N_4998,N_4747);
and U5041 (N_5041,N_4661,N_4787);
nand U5042 (N_5042,N_4610,N_4860);
nor U5043 (N_5043,N_4776,N_4677);
nor U5044 (N_5044,N_4741,N_4833);
xnor U5045 (N_5045,N_4934,N_4636);
xor U5046 (N_5046,N_4736,N_4865);
xnor U5047 (N_5047,N_4631,N_4514);
nor U5048 (N_5048,N_4788,N_4993);
and U5049 (N_5049,N_4841,N_4625);
and U5050 (N_5050,N_4918,N_4522);
nor U5051 (N_5051,N_4888,N_4864);
xnor U5052 (N_5052,N_4702,N_4948);
or U5053 (N_5053,N_4566,N_4759);
xnor U5054 (N_5054,N_4994,N_4502);
or U5055 (N_5055,N_4931,N_4905);
xnor U5056 (N_5056,N_4733,N_4735);
and U5057 (N_5057,N_4944,N_4781);
and U5058 (N_5058,N_4737,N_4561);
nor U5059 (N_5059,N_4565,N_4917);
nor U5060 (N_5060,N_4659,N_4571);
nor U5061 (N_5061,N_4754,N_4871);
nand U5062 (N_5062,N_4959,N_4899);
and U5063 (N_5063,N_4818,N_4508);
or U5064 (N_5064,N_4616,N_4878);
xnor U5065 (N_5065,N_4622,N_4538);
or U5066 (N_5066,N_4816,N_4988);
nor U5067 (N_5067,N_4912,N_4913);
nor U5068 (N_5068,N_4576,N_4579);
nand U5069 (N_5069,N_4801,N_4552);
nor U5070 (N_5070,N_4681,N_4794);
xor U5071 (N_5071,N_4831,N_4826);
or U5072 (N_5072,N_4995,N_4757);
nand U5073 (N_5073,N_4529,N_4891);
and U5074 (N_5074,N_4685,N_4966);
nor U5075 (N_5075,N_4881,N_4910);
or U5076 (N_5076,N_4740,N_4639);
nor U5077 (N_5077,N_4700,N_4624);
xor U5078 (N_5078,N_4630,N_4937);
nor U5079 (N_5079,N_4734,N_4678);
xor U5080 (N_5080,N_4548,N_4974);
and U5081 (N_5081,N_4970,N_4844);
xnor U5082 (N_5082,N_4526,N_4992);
nand U5083 (N_5083,N_4721,N_4729);
nand U5084 (N_5084,N_4553,N_4761);
xnor U5085 (N_5085,N_4773,N_4900);
or U5086 (N_5086,N_4506,N_4638);
or U5087 (N_5087,N_4572,N_4790);
xnor U5088 (N_5088,N_4550,N_4632);
nor U5089 (N_5089,N_4669,N_4595);
nor U5090 (N_5090,N_4965,N_4586);
xnor U5091 (N_5091,N_4614,N_4908);
nor U5092 (N_5092,N_4834,N_4676);
and U5093 (N_5093,N_4600,N_4777);
and U5094 (N_5094,N_4824,N_4708);
and U5095 (N_5095,N_4644,N_4535);
xnor U5096 (N_5096,N_4967,N_4882);
nor U5097 (N_5097,N_4683,N_4730);
xor U5098 (N_5098,N_4999,N_4503);
xor U5099 (N_5099,N_4767,N_4545);
or U5100 (N_5100,N_4766,N_4524);
nor U5101 (N_5101,N_4623,N_4555);
xnor U5102 (N_5102,N_4990,N_4940);
xor U5103 (N_5103,N_4928,N_4863);
nand U5104 (N_5104,N_4519,N_4774);
xor U5105 (N_5105,N_4954,N_4507);
nor U5106 (N_5106,N_4820,N_4605);
and U5107 (N_5107,N_4728,N_4770);
and U5108 (N_5108,N_4982,N_4694);
nand U5109 (N_5109,N_4609,N_4839);
and U5110 (N_5110,N_4972,N_4607);
nand U5111 (N_5111,N_4828,N_4782);
xnor U5112 (N_5112,N_4709,N_4591);
nand U5113 (N_5113,N_4830,N_4745);
nand U5114 (N_5114,N_4927,N_4977);
nand U5115 (N_5115,N_4577,N_4764);
or U5116 (N_5116,N_4870,N_4642);
and U5117 (N_5117,N_4652,N_4680);
or U5118 (N_5118,N_4789,N_4703);
nor U5119 (N_5119,N_4719,N_4528);
and U5120 (N_5120,N_4693,N_4808);
nand U5121 (N_5121,N_4711,N_4516);
xor U5122 (N_5122,N_4688,N_4896);
or U5123 (N_5123,N_4606,N_4979);
and U5124 (N_5124,N_4751,N_4884);
and U5125 (N_5125,N_4907,N_4671);
nand U5126 (N_5126,N_4866,N_4953);
nand U5127 (N_5127,N_4772,N_4584);
and U5128 (N_5128,N_4848,N_4938);
or U5129 (N_5129,N_4633,N_4810);
nand U5130 (N_5130,N_4564,N_4890);
nor U5131 (N_5131,N_4821,N_4675);
nor U5132 (N_5132,N_4815,N_4842);
xor U5133 (N_5133,N_4961,N_4562);
or U5134 (N_5134,N_4946,N_4947);
nor U5135 (N_5135,N_4872,N_4804);
and U5136 (N_5136,N_4755,N_4717);
or U5137 (N_5137,N_4660,N_4769);
xnor U5138 (N_5138,N_4501,N_4827);
or U5139 (N_5139,N_4715,N_4887);
nor U5140 (N_5140,N_4670,N_4922);
and U5141 (N_5141,N_4523,N_4760);
nand U5142 (N_5142,N_4530,N_4853);
or U5143 (N_5143,N_4540,N_4943);
nor U5144 (N_5144,N_4527,N_4875);
nand U5145 (N_5145,N_4783,N_4861);
or U5146 (N_5146,N_4554,N_4975);
nand U5147 (N_5147,N_4698,N_4855);
nor U5148 (N_5148,N_4539,N_4581);
xor U5149 (N_5149,N_4976,N_4867);
nand U5150 (N_5150,N_4726,N_4603);
nand U5151 (N_5151,N_4981,N_4626);
xor U5152 (N_5152,N_4727,N_4608);
xor U5153 (N_5153,N_4687,N_4686);
or U5154 (N_5154,N_4738,N_4691);
or U5155 (N_5155,N_4518,N_4634);
xnor U5156 (N_5156,N_4916,N_4695);
or U5157 (N_5157,N_4809,N_4615);
nand U5158 (N_5158,N_4750,N_4968);
and U5159 (N_5159,N_4587,N_4512);
and U5160 (N_5160,N_4582,N_4731);
and U5161 (N_5161,N_4851,N_4923);
xnor U5162 (N_5162,N_4707,N_4997);
xnor U5163 (N_5163,N_4664,N_4722);
nor U5164 (N_5164,N_4596,N_4892);
and U5165 (N_5165,N_4984,N_4696);
xnor U5166 (N_5166,N_4662,N_4748);
or U5167 (N_5167,N_4856,N_4558);
xnor U5168 (N_5168,N_4991,N_4654);
or U5169 (N_5169,N_4712,N_4604);
xor U5170 (N_5170,N_4799,N_4704);
nand U5171 (N_5171,N_4909,N_4868);
xnor U5172 (N_5172,N_4956,N_4960);
or U5173 (N_5173,N_4813,N_4511);
nand U5174 (N_5174,N_4743,N_4894);
xnor U5175 (N_5175,N_4521,N_4746);
nand U5176 (N_5176,N_4627,N_4567);
or U5177 (N_5177,N_4837,N_4987);
xor U5178 (N_5178,N_4846,N_4825);
nand U5179 (N_5179,N_4925,N_4893);
nor U5180 (N_5180,N_4797,N_4551);
nand U5181 (N_5181,N_4723,N_4513);
nand U5182 (N_5182,N_4803,N_4500);
and U5183 (N_5183,N_4958,N_4904);
and U5184 (N_5184,N_4611,N_4725);
or U5185 (N_5185,N_4510,N_4692);
and U5186 (N_5186,N_4932,N_4921);
or U5187 (N_5187,N_4793,N_4983);
xnor U5188 (N_5188,N_4612,N_4641);
or U5189 (N_5189,N_4640,N_4556);
and U5190 (N_5190,N_4559,N_4950);
nor U5191 (N_5191,N_4903,N_4857);
and U5192 (N_5192,N_4752,N_4765);
xor U5193 (N_5193,N_4574,N_4941);
and U5194 (N_5194,N_4531,N_4674);
or U5195 (N_5195,N_4762,N_4648);
nor U5196 (N_5196,N_4945,N_4978);
and U5197 (N_5197,N_4964,N_4758);
nand U5198 (N_5198,N_4542,N_4568);
xor U5199 (N_5199,N_4557,N_4699);
and U5200 (N_5200,N_4838,N_4926);
xnor U5201 (N_5201,N_4520,N_4780);
nor U5202 (N_5202,N_4786,N_4575);
nor U5203 (N_5203,N_4935,N_4742);
xnor U5204 (N_5204,N_4869,N_4578);
xnor U5205 (N_5205,N_4939,N_4806);
nor U5206 (N_5206,N_4653,N_4756);
and U5207 (N_5207,N_4823,N_4822);
or U5208 (N_5208,N_4814,N_4525);
nor U5209 (N_5209,N_4930,N_4986);
xnor U5210 (N_5210,N_4883,N_4549);
nor U5211 (N_5211,N_4914,N_4720);
nor U5212 (N_5212,N_4929,N_4840);
nand U5213 (N_5213,N_4843,N_4656);
nand U5214 (N_5214,N_4650,N_4778);
xnor U5215 (N_5215,N_4724,N_4628);
xor U5216 (N_5216,N_4515,N_4705);
nand U5217 (N_5217,N_4845,N_4547);
and U5218 (N_5218,N_4798,N_4580);
and U5219 (N_5219,N_4594,N_4617);
nand U5220 (N_5220,N_4885,N_4796);
xnor U5221 (N_5221,N_4763,N_4795);
or U5222 (N_5222,N_4854,N_4621);
nor U5223 (N_5223,N_4697,N_4589);
or U5224 (N_5224,N_4957,N_4665);
xnor U5225 (N_5225,N_4637,N_4906);
xor U5226 (N_5226,N_4812,N_4597);
or U5227 (N_5227,N_4971,N_4718);
or U5228 (N_5228,N_4862,N_4602);
xnor U5229 (N_5229,N_4952,N_4536);
nor U5230 (N_5230,N_4768,N_4541);
nor U5231 (N_5231,N_4663,N_4784);
nand U5232 (N_5232,N_4588,N_4713);
nand U5233 (N_5233,N_4886,N_4771);
and U5234 (N_5234,N_4949,N_4749);
xnor U5235 (N_5235,N_4835,N_4657);
xnor U5236 (N_5236,N_4969,N_4701);
or U5237 (N_5237,N_4517,N_4560);
or U5238 (N_5238,N_4620,N_4901);
nand U5239 (N_5239,N_4593,N_4792);
nor U5240 (N_5240,N_4985,N_4504);
and U5241 (N_5241,N_4876,N_4716);
and U5242 (N_5242,N_4682,N_4973);
nand U5243 (N_5243,N_4689,N_4655);
or U5244 (N_5244,N_4919,N_4852);
or U5245 (N_5245,N_4962,N_4879);
nor U5246 (N_5246,N_4668,N_4858);
or U5247 (N_5247,N_4942,N_4651);
xor U5248 (N_5248,N_4811,N_4924);
nand U5249 (N_5249,N_4647,N_4819);
xnor U5250 (N_5250,N_4907,N_4512);
or U5251 (N_5251,N_4698,N_4647);
or U5252 (N_5252,N_4658,N_4853);
nand U5253 (N_5253,N_4768,N_4599);
nor U5254 (N_5254,N_4939,N_4750);
and U5255 (N_5255,N_4767,N_4953);
xnor U5256 (N_5256,N_4709,N_4577);
nor U5257 (N_5257,N_4625,N_4530);
nor U5258 (N_5258,N_4931,N_4594);
and U5259 (N_5259,N_4703,N_4810);
nor U5260 (N_5260,N_4544,N_4621);
nor U5261 (N_5261,N_4929,N_4842);
xnor U5262 (N_5262,N_4746,N_4903);
xor U5263 (N_5263,N_4796,N_4784);
nand U5264 (N_5264,N_4641,N_4574);
nand U5265 (N_5265,N_4719,N_4832);
nand U5266 (N_5266,N_4589,N_4869);
nor U5267 (N_5267,N_4676,N_4955);
xnor U5268 (N_5268,N_4741,N_4809);
nand U5269 (N_5269,N_4985,N_4568);
nand U5270 (N_5270,N_4677,N_4718);
nor U5271 (N_5271,N_4676,N_4864);
nand U5272 (N_5272,N_4513,N_4501);
and U5273 (N_5273,N_4694,N_4782);
nand U5274 (N_5274,N_4934,N_4605);
xnor U5275 (N_5275,N_4790,N_4966);
and U5276 (N_5276,N_4578,N_4849);
or U5277 (N_5277,N_4660,N_4915);
and U5278 (N_5278,N_4862,N_4605);
nor U5279 (N_5279,N_4690,N_4739);
or U5280 (N_5280,N_4892,N_4991);
nor U5281 (N_5281,N_4616,N_4526);
and U5282 (N_5282,N_4797,N_4642);
nor U5283 (N_5283,N_4531,N_4509);
nor U5284 (N_5284,N_4964,N_4889);
and U5285 (N_5285,N_4671,N_4683);
or U5286 (N_5286,N_4678,N_4851);
nand U5287 (N_5287,N_4523,N_4908);
or U5288 (N_5288,N_4988,N_4532);
and U5289 (N_5289,N_4977,N_4710);
or U5290 (N_5290,N_4518,N_4695);
xnor U5291 (N_5291,N_4749,N_4906);
xor U5292 (N_5292,N_4614,N_4688);
or U5293 (N_5293,N_4964,N_4522);
nor U5294 (N_5294,N_4806,N_4507);
or U5295 (N_5295,N_4975,N_4711);
nand U5296 (N_5296,N_4913,N_4611);
and U5297 (N_5297,N_4779,N_4931);
nor U5298 (N_5298,N_4627,N_4999);
or U5299 (N_5299,N_4755,N_4754);
xor U5300 (N_5300,N_4866,N_4763);
xnor U5301 (N_5301,N_4592,N_4737);
xnor U5302 (N_5302,N_4821,N_4580);
and U5303 (N_5303,N_4853,N_4957);
and U5304 (N_5304,N_4629,N_4571);
nand U5305 (N_5305,N_4680,N_4857);
nor U5306 (N_5306,N_4501,N_4800);
xnor U5307 (N_5307,N_4772,N_4838);
nand U5308 (N_5308,N_4933,N_4771);
and U5309 (N_5309,N_4516,N_4852);
and U5310 (N_5310,N_4615,N_4504);
nor U5311 (N_5311,N_4541,N_4850);
xnor U5312 (N_5312,N_4959,N_4875);
or U5313 (N_5313,N_4614,N_4795);
xor U5314 (N_5314,N_4607,N_4910);
and U5315 (N_5315,N_4725,N_4946);
and U5316 (N_5316,N_4734,N_4835);
nor U5317 (N_5317,N_4633,N_4850);
xnor U5318 (N_5318,N_4771,N_4538);
nor U5319 (N_5319,N_4638,N_4673);
and U5320 (N_5320,N_4779,N_4541);
and U5321 (N_5321,N_4551,N_4521);
and U5322 (N_5322,N_4770,N_4542);
or U5323 (N_5323,N_4806,N_4914);
nor U5324 (N_5324,N_4622,N_4748);
and U5325 (N_5325,N_4593,N_4967);
or U5326 (N_5326,N_4646,N_4983);
or U5327 (N_5327,N_4883,N_4801);
and U5328 (N_5328,N_4912,N_4819);
xnor U5329 (N_5329,N_4961,N_4842);
xor U5330 (N_5330,N_4967,N_4503);
and U5331 (N_5331,N_4540,N_4794);
or U5332 (N_5332,N_4962,N_4847);
or U5333 (N_5333,N_4876,N_4941);
nand U5334 (N_5334,N_4500,N_4539);
nand U5335 (N_5335,N_4981,N_4596);
nor U5336 (N_5336,N_4901,N_4728);
xnor U5337 (N_5337,N_4993,N_4537);
nand U5338 (N_5338,N_4813,N_4858);
xor U5339 (N_5339,N_4525,N_4819);
xnor U5340 (N_5340,N_4609,N_4757);
nor U5341 (N_5341,N_4516,N_4937);
nand U5342 (N_5342,N_4914,N_4668);
and U5343 (N_5343,N_4636,N_4830);
xor U5344 (N_5344,N_4655,N_4775);
or U5345 (N_5345,N_4998,N_4893);
or U5346 (N_5346,N_4511,N_4564);
and U5347 (N_5347,N_4552,N_4648);
xnor U5348 (N_5348,N_4760,N_4900);
xor U5349 (N_5349,N_4577,N_4826);
or U5350 (N_5350,N_4706,N_4947);
nand U5351 (N_5351,N_4591,N_4577);
nand U5352 (N_5352,N_4991,N_4970);
or U5353 (N_5353,N_4581,N_4686);
nand U5354 (N_5354,N_4533,N_4983);
and U5355 (N_5355,N_4733,N_4995);
and U5356 (N_5356,N_4796,N_4572);
xnor U5357 (N_5357,N_4599,N_4990);
nand U5358 (N_5358,N_4925,N_4794);
xor U5359 (N_5359,N_4614,N_4911);
nand U5360 (N_5360,N_4532,N_4708);
and U5361 (N_5361,N_4700,N_4907);
nand U5362 (N_5362,N_4978,N_4916);
and U5363 (N_5363,N_4619,N_4757);
xnor U5364 (N_5364,N_4526,N_4869);
nand U5365 (N_5365,N_4519,N_4665);
or U5366 (N_5366,N_4893,N_4573);
or U5367 (N_5367,N_4776,N_4589);
and U5368 (N_5368,N_4651,N_4811);
or U5369 (N_5369,N_4801,N_4858);
xnor U5370 (N_5370,N_4565,N_4845);
and U5371 (N_5371,N_4992,N_4816);
or U5372 (N_5372,N_4882,N_4527);
or U5373 (N_5373,N_4960,N_4918);
nor U5374 (N_5374,N_4998,N_4745);
nor U5375 (N_5375,N_4779,N_4658);
nand U5376 (N_5376,N_4782,N_4901);
and U5377 (N_5377,N_4565,N_4911);
nand U5378 (N_5378,N_4585,N_4615);
nor U5379 (N_5379,N_4668,N_4802);
xor U5380 (N_5380,N_4577,N_4556);
and U5381 (N_5381,N_4629,N_4943);
nor U5382 (N_5382,N_4923,N_4728);
nor U5383 (N_5383,N_4964,N_4538);
or U5384 (N_5384,N_4808,N_4738);
xor U5385 (N_5385,N_4979,N_4628);
or U5386 (N_5386,N_4887,N_4536);
nor U5387 (N_5387,N_4992,N_4500);
xnor U5388 (N_5388,N_4668,N_4955);
xnor U5389 (N_5389,N_4539,N_4697);
or U5390 (N_5390,N_4620,N_4680);
nor U5391 (N_5391,N_4964,N_4675);
nor U5392 (N_5392,N_4938,N_4528);
xor U5393 (N_5393,N_4836,N_4779);
nor U5394 (N_5394,N_4647,N_4625);
nor U5395 (N_5395,N_4931,N_4817);
xor U5396 (N_5396,N_4576,N_4853);
and U5397 (N_5397,N_4786,N_4630);
xnor U5398 (N_5398,N_4506,N_4545);
nand U5399 (N_5399,N_4955,N_4554);
or U5400 (N_5400,N_4873,N_4590);
or U5401 (N_5401,N_4618,N_4787);
or U5402 (N_5402,N_4800,N_4785);
nor U5403 (N_5403,N_4824,N_4514);
xor U5404 (N_5404,N_4878,N_4944);
or U5405 (N_5405,N_4500,N_4953);
nor U5406 (N_5406,N_4696,N_4638);
or U5407 (N_5407,N_4620,N_4681);
xor U5408 (N_5408,N_4894,N_4860);
nor U5409 (N_5409,N_4709,N_4714);
xnor U5410 (N_5410,N_4889,N_4923);
xnor U5411 (N_5411,N_4838,N_4517);
xnor U5412 (N_5412,N_4950,N_4547);
or U5413 (N_5413,N_4871,N_4661);
xor U5414 (N_5414,N_4531,N_4827);
nand U5415 (N_5415,N_4800,N_4926);
xnor U5416 (N_5416,N_4845,N_4580);
xnor U5417 (N_5417,N_4763,N_4737);
or U5418 (N_5418,N_4968,N_4578);
xnor U5419 (N_5419,N_4674,N_4768);
nor U5420 (N_5420,N_4771,N_4734);
or U5421 (N_5421,N_4541,N_4766);
nor U5422 (N_5422,N_4773,N_4648);
or U5423 (N_5423,N_4881,N_4737);
nand U5424 (N_5424,N_4718,N_4591);
nand U5425 (N_5425,N_4556,N_4777);
xor U5426 (N_5426,N_4583,N_4637);
nor U5427 (N_5427,N_4973,N_4823);
nand U5428 (N_5428,N_4759,N_4752);
nand U5429 (N_5429,N_4990,N_4559);
or U5430 (N_5430,N_4831,N_4757);
nand U5431 (N_5431,N_4650,N_4769);
xnor U5432 (N_5432,N_4667,N_4972);
xor U5433 (N_5433,N_4627,N_4924);
or U5434 (N_5434,N_4899,N_4933);
xor U5435 (N_5435,N_4531,N_4996);
nand U5436 (N_5436,N_4804,N_4888);
nor U5437 (N_5437,N_4732,N_4996);
nor U5438 (N_5438,N_4746,N_4896);
or U5439 (N_5439,N_4668,N_4512);
and U5440 (N_5440,N_4580,N_4804);
nor U5441 (N_5441,N_4542,N_4516);
and U5442 (N_5442,N_4641,N_4963);
xnor U5443 (N_5443,N_4808,N_4641);
nor U5444 (N_5444,N_4863,N_4886);
or U5445 (N_5445,N_4732,N_4603);
nand U5446 (N_5446,N_4971,N_4672);
nand U5447 (N_5447,N_4888,N_4981);
and U5448 (N_5448,N_4501,N_4805);
and U5449 (N_5449,N_4860,N_4634);
and U5450 (N_5450,N_4681,N_4785);
xor U5451 (N_5451,N_4565,N_4506);
xnor U5452 (N_5452,N_4815,N_4604);
and U5453 (N_5453,N_4971,N_4646);
and U5454 (N_5454,N_4745,N_4662);
and U5455 (N_5455,N_4814,N_4797);
nor U5456 (N_5456,N_4986,N_4730);
nand U5457 (N_5457,N_4810,N_4529);
and U5458 (N_5458,N_4886,N_4597);
nor U5459 (N_5459,N_4834,N_4771);
nand U5460 (N_5460,N_4835,N_4799);
or U5461 (N_5461,N_4914,N_4649);
or U5462 (N_5462,N_4723,N_4895);
nor U5463 (N_5463,N_4954,N_4723);
and U5464 (N_5464,N_4628,N_4897);
xor U5465 (N_5465,N_4651,N_4884);
nor U5466 (N_5466,N_4839,N_4517);
xor U5467 (N_5467,N_4725,N_4865);
or U5468 (N_5468,N_4522,N_4544);
nor U5469 (N_5469,N_4793,N_4707);
or U5470 (N_5470,N_4944,N_4518);
or U5471 (N_5471,N_4524,N_4576);
nand U5472 (N_5472,N_4929,N_4566);
and U5473 (N_5473,N_4766,N_4986);
nor U5474 (N_5474,N_4656,N_4600);
or U5475 (N_5475,N_4800,N_4992);
nor U5476 (N_5476,N_4807,N_4769);
and U5477 (N_5477,N_4589,N_4762);
nand U5478 (N_5478,N_4793,N_4668);
xnor U5479 (N_5479,N_4603,N_4698);
xnor U5480 (N_5480,N_4797,N_4744);
nand U5481 (N_5481,N_4989,N_4997);
or U5482 (N_5482,N_4661,N_4844);
and U5483 (N_5483,N_4755,N_4892);
and U5484 (N_5484,N_4600,N_4940);
nor U5485 (N_5485,N_4969,N_4530);
nor U5486 (N_5486,N_4650,N_4749);
nor U5487 (N_5487,N_4942,N_4583);
or U5488 (N_5488,N_4905,N_4544);
or U5489 (N_5489,N_4632,N_4883);
xor U5490 (N_5490,N_4983,N_4886);
xnor U5491 (N_5491,N_4611,N_4556);
nand U5492 (N_5492,N_4951,N_4519);
or U5493 (N_5493,N_4926,N_4982);
or U5494 (N_5494,N_4865,N_4776);
xor U5495 (N_5495,N_4602,N_4795);
nand U5496 (N_5496,N_4909,N_4555);
nor U5497 (N_5497,N_4972,N_4747);
or U5498 (N_5498,N_4572,N_4706);
and U5499 (N_5499,N_4762,N_4726);
or U5500 (N_5500,N_5136,N_5105);
xnor U5501 (N_5501,N_5326,N_5214);
or U5502 (N_5502,N_5457,N_5365);
and U5503 (N_5503,N_5201,N_5167);
nor U5504 (N_5504,N_5343,N_5195);
nor U5505 (N_5505,N_5333,N_5254);
and U5506 (N_5506,N_5093,N_5434);
nand U5507 (N_5507,N_5020,N_5150);
xor U5508 (N_5508,N_5471,N_5194);
or U5509 (N_5509,N_5244,N_5320);
and U5510 (N_5510,N_5168,N_5347);
and U5511 (N_5511,N_5344,N_5369);
nand U5512 (N_5512,N_5275,N_5403);
xor U5513 (N_5513,N_5228,N_5239);
or U5514 (N_5514,N_5430,N_5406);
nand U5515 (N_5515,N_5265,N_5145);
or U5516 (N_5516,N_5138,N_5428);
xnor U5517 (N_5517,N_5459,N_5063);
or U5518 (N_5518,N_5114,N_5321);
nand U5519 (N_5519,N_5018,N_5031);
nor U5520 (N_5520,N_5454,N_5221);
or U5521 (N_5521,N_5090,N_5449);
xor U5522 (N_5522,N_5157,N_5006);
xnor U5523 (N_5523,N_5460,N_5215);
xnor U5524 (N_5524,N_5081,N_5355);
nor U5525 (N_5525,N_5234,N_5147);
xnor U5526 (N_5526,N_5183,N_5266);
nand U5527 (N_5527,N_5062,N_5376);
nor U5528 (N_5528,N_5352,N_5435);
nand U5529 (N_5529,N_5422,N_5156);
nor U5530 (N_5530,N_5046,N_5452);
and U5531 (N_5531,N_5137,N_5241);
nand U5532 (N_5532,N_5058,N_5324);
nor U5533 (N_5533,N_5419,N_5338);
or U5534 (N_5534,N_5287,N_5129);
xor U5535 (N_5535,N_5359,N_5330);
and U5536 (N_5536,N_5488,N_5117);
and U5537 (N_5537,N_5209,N_5124);
nor U5538 (N_5538,N_5380,N_5305);
nor U5539 (N_5539,N_5311,N_5075);
nand U5540 (N_5540,N_5251,N_5108);
nor U5541 (N_5541,N_5059,N_5178);
and U5542 (N_5542,N_5379,N_5323);
or U5543 (N_5543,N_5414,N_5104);
xnor U5544 (N_5544,N_5162,N_5101);
nand U5545 (N_5545,N_5440,N_5052);
nor U5546 (N_5546,N_5298,N_5328);
and U5547 (N_5547,N_5022,N_5021);
xor U5548 (N_5548,N_5140,N_5177);
nor U5549 (N_5549,N_5413,N_5198);
or U5550 (N_5550,N_5470,N_5426);
xnor U5551 (N_5551,N_5350,N_5030);
nand U5552 (N_5552,N_5128,N_5362);
nor U5553 (N_5553,N_5103,N_5396);
nor U5554 (N_5554,N_5279,N_5123);
and U5555 (N_5555,N_5047,N_5385);
and U5556 (N_5556,N_5013,N_5441);
and U5557 (N_5557,N_5354,N_5409);
or U5558 (N_5558,N_5076,N_5122);
nor U5559 (N_5559,N_5407,N_5249);
and U5560 (N_5560,N_5257,N_5002);
xor U5561 (N_5561,N_5278,N_5318);
xnor U5562 (N_5562,N_5392,N_5349);
or U5563 (N_5563,N_5481,N_5408);
and U5564 (N_5564,N_5023,N_5283);
and U5565 (N_5565,N_5447,N_5267);
nor U5566 (N_5566,N_5233,N_5292);
or U5567 (N_5567,N_5250,N_5367);
and U5568 (N_5568,N_5378,N_5065);
and U5569 (N_5569,N_5109,N_5039);
nor U5570 (N_5570,N_5444,N_5293);
or U5571 (N_5571,N_5374,N_5300);
or U5572 (N_5572,N_5258,N_5088);
xor U5573 (N_5573,N_5322,N_5256);
and U5574 (N_5574,N_5041,N_5325);
or U5575 (N_5575,N_5469,N_5486);
nor U5576 (N_5576,N_5053,N_5364);
xnor U5577 (N_5577,N_5061,N_5126);
or U5578 (N_5578,N_5288,N_5277);
nor U5579 (N_5579,N_5207,N_5084);
or U5580 (N_5580,N_5337,N_5000);
nand U5581 (N_5581,N_5184,N_5383);
nand U5582 (N_5582,N_5164,N_5433);
nor U5583 (N_5583,N_5432,N_5087);
nand U5584 (N_5584,N_5404,N_5410);
nor U5585 (N_5585,N_5237,N_5405);
nand U5586 (N_5586,N_5227,N_5095);
nor U5587 (N_5587,N_5232,N_5285);
or U5588 (N_5588,N_5313,N_5478);
and U5589 (N_5589,N_5210,N_5319);
nand U5590 (N_5590,N_5262,N_5218);
or U5591 (N_5591,N_5196,N_5371);
or U5592 (N_5592,N_5246,N_5295);
xnor U5593 (N_5593,N_5331,N_5094);
xnor U5594 (N_5594,N_5074,N_5357);
xnor U5595 (N_5595,N_5148,N_5049);
or U5596 (N_5596,N_5165,N_5025);
or U5597 (N_5597,N_5048,N_5353);
xor U5598 (N_5598,N_5118,N_5040);
nand U5599 (N_5599,N_5425,N_5180);
or U5600 (N_5600,N_5050,N_5391);
nor U5601 (N_5601,N_5327,N_5173);
and U5602 (N_5602,N_5092,N_5390);
nand U5603 (N_5603,N_5386,N_5034);
nor U5604 (N_5604,N_5045,N_5255);
xor U5605 (N_5605,N_5242,N_5436);
or U5606 (N_5606,N_5051,N_5336);
xor U5607 (N_5607,N_5315,N_5297);
or U5608 (N_5608,N_5202,N_5493);
xnor U5609 (N_5609,N_5247,N_5363);
and U5610 (N_5610,N_5192,N_5465);
or U5611 (N_5611,N_5420,N_5366);
and U5612 (N_5612,N_5453,N_5149);
xor U5613 (N_5613,N_5071,N_5252);
or U5614 (N_5614,N_5008,N_5270);
nor U5615 (N_5615,N_5189,N_5417);
nor U5616 (N_5616,N_5231,N_5400);
or U5617 (N_5617,N_5042,N_5370);
or U5618 (N_5618,N_5004,N_5368);
nor U5619 (N_5619,N_5271,N_5276);
or U5620 (N_5620,N_5290,N_5038);
nor U5621 (N_5621,N_5375,N_5001);
xnor U5622 (N_5622,N_5468,N_5424);
and U5623 (N_5623,N_5450,N_5015);
xnor U5624 (N_5624,N_5272,N_5455);
nor U5625 (N_5625,N_5448,N_5463);
xnor U5626 (N_5626,N_5462,N_5443);
xor U5627 (N_5627,N_5439,N_5029);
xor U5628 (N_5628,N_5066,N_5116);
nand U5629 (N_5629,N_5097,N_5203);
nand U5630 (N_5630,N_5281,N_5100);
and U5631 (N_5631,N_5190,N_5497);
and U5632 (N_5632,N_5382,N_5482);
or U5633 (N_5633,N_5024,N_5043);
and U5634 (N_5634,N_5153,N_5172);
and U5635 (N_5635,N_5308,N_5416);
and U5636 (N_5636,N_5102,N_5341);
nand U5637 (N_5637,N_5070,N_5208);
or U5638 (N_5638,N_5119,N_5476);
xnor U5639 (N_5639,N_5213,N_5037);
or U5640 (N_5640,N_5054,N_5402);
or U5641 (N_5641,N_5394,N_5146);
nor U5642 (N_5642,N_5229,N_5431);
and U5643 (N_5643,N_5446,N_5226);
and U5644 (N_5644,N_5003,N_5314);
or U5645 (N_5645,N_5223,N_5474);
and U5646 (N_5646,N_5268,N_5269);
or U5647 (N_5647,N_5389,N_5495);
or U5648 (N_5648,N_5211,N_5317);
nor U5649 (N_5649,N_5316,N_5115);
or U5650 (N_5650,N_5260,N_5423);
or U5651 (N_5651,N_5304,N_5345);
and U5652 (N_5652,N_5222,N_5132);
or U5653 (N_5653,N_5473,N_5259);
or U5654 (N_5654,N_5384,N_5358);
and U5655 (N_5655,N_5067,N_5301);
and U5656 (N_5656,N_5225,N_5158);
xnor U5657 (N_5657,N_5381,N_5296);
and U5658 (N_5658,N_5335,N_5479);
xnor U5659 (N_5659,N_5373,N_5193);
xor U5660 (N_5660,N_5219,N_5306);
or U5661 (N_5661,N_5206,N_5127);
nand U5662 (N_5662,N_5334,N_5028);
or U5663 (N_5663,N_5078,N_5134);
xor U5664 (N_5664,N_5346,N_5197);
or U5665 (N_5665,N_5361,N_5253);
nor U5666 (N_5666,N_5133,N_5032);
nand U5667 (N_5667,N_5429,N_5451);
nor U5668 (N_5668,N_5360,N_5397);
and U5669 (N_5669,N_5204,N_5498);
xor U5670 (N_5670,N_5125,N_5467);
xor U5671 (N_5671,N_5007,N_5289);
xnor U5672 (N_5672,N_5332,N_5069);
and U5673 (N_5673,N_5264,N_5351);
xnor U5674 (N_5674,N_5027,N_5477);
nor U5675 (N_5675,N_5174,N_5163);
and U5676 (N_5676,N_5171,N_5487);
and U5677 (N_5677,N_5142,N_5057);
nand U5678 (N_5678,N_5235,N_5388);
xnor U5679 (N_5679,N_5154,N_5496);
xnor U5680 (N_5680,N_5079,N_5035);
nor U5681 (N_5681,N_5160,N_5348);
and U5682 (N_5682,N_5169,N_5155);
or U5683 (N_5683,N_5291,N_5110);
nor U5684 (N_5684,N_5280,N_5484);
xnor U5685 (N_5685,N_5185,N_5036);
xor U5686 (N_5686,N_5438,N_5099);
and U5687 (N_5687,N_5161,N_5096);
or U5688 (N_5688,N_5098,N_5238);
xor U5689 (N_5689,N_5026,N_5236);
nor U5690 (N_5690,N_5068,N_5135);
xor U5691 (N_5691,N_5340,N_5060);
nand U5692 (N_5692,N_5217,N_5286);
nand U5693 (N_5693,N_5274,N_5339);
or U5694 (N_5694,N_5387,N_5212);
nand U5695 (N_5695,N_5010,N_5307);
or U5696 (N_5696,N_5490,N_5187);
nor U5697 (N_5697,N_5299,N_5205);
nor U5698 (N_5698,N_5056,N_5216);
and U5699 (N_5699,N_5393,N_5303);
xor U5700 (N_5700,N_5458,N_5072);
xor U5701 (N_5701,N_5411,N_5113);
xor U5702 (N_5702,N_5199,N_5442);
nand U5703 (N_5703,N_5055,N_5427);
or U5704 (N_5704,N_5398,N_5492);
xor U5705 (N_5705,N_5377,N_5245);
nand U5706 (N_5706,N_5263,N_5499);
or U5707 (N_5707,N_5273,N_5106);
nor U5708 (N_5708,N_5073,N_5086);
nand U5709 (N_5709,N_5188,N_5091);
nor U5710 (N_5710,N_5412,N_5395);
or U5711 (N_5711,N_5302,N_5342);
xor U5712 (N_5712,N_5489,N_5143);
nor U5713 (N_5713,N_5437,N_5312);
nand U5714 (N_5714,N_5082,N_5480);
or U5715 (N_5715,N_5151,N_5141);
nand U5716 (N_5716,N_5220,N_5005);
nor U5717 (N_5717,N_5310,N_5139);
xnor U5718 (N_5718,N_5472,N_5243);
xnor U5719 (N_5719,N_5080,N_5294);
nor U5720 (N_5720,N_5475,N_5356);
nand U5721 (N_5721,N_5170,N_5329);
and U5722 (N_5722,N_5077,N_5466);
or U5723 (N_5723,N_5200,N_5224);
nand U5724 (N_5724,N_5089,N_5012);
and U5725 (N_5725,N_5014,N_5445);
or U5726 (N_5726,N_5152,N_5011);
xnor U5727 (N_5727,N_5240,N_5120);
xnor U5728 (N_5728,N_5399,N_5186);
or U5729 (N_5729,N_5016,N_5483);
or U5730 (N_5730,N_5461,N_5111);
nand U5731 (N_5731,N_5159,N_5019);
and U5732 (N_5732,N_5121,N_5083);
nand U5733 (N_5733,N_5085,N_5107);
nand U5734 (N_5734,N_5166,N_5131);
or U5735 (N_5735,N_5494,N_5284);
xor U5736 (N_5736,N_5491,N_5009);
nand U5737 (N_5737,N_5230,N_5182);
and U5738 (N_5738,N_5418,N_5464);
xor U5739 (N_5739,N_5421,N_5401);
nand U5740 (N_5740,N_5176,N_5456);
nand U5741 (N_5741,N_5033,N_5282);
and U5742 (N_5742,N_5485,N_5181);
nor U5743 (N_5743,N_5175,N_5064);
nor U5744 (N_5744,N_5261,N_5112);
xnor U5745 (N_5745,N_5044,N_5309);
nor U5746 (N_5746,N_5248,N_5179);
nand U5747 (N_5747,N_5415,N_5191);
and U5748 (N_5748,N_5130,N_5372);
or U5749 (N_5749,N_5144,N_5017);
and U5750 (N_5750,N_5294,N_5370);
xor U5751 (N_5751,N_5239,N_5053);
and U5752 (N_5752,N_5238,N_5480);
nor U5753 (N_5753,N_5061,N_5437);
nand U5754 (N_5754,N_5453,N_5140);
nor U5755 (N_5755,N_5127,N_5023);
or U5756 (N_5756,N_5282,N_5010);
nand U5757 (N_5757,N_5415,N_5188);
xnor U5758 (N_5758,N_5235,N_5233);
and U5759 (N_5759,N_5247,N_5062);
xor U5760 (N_5760,N_5071,N_5243);
or U5761 (N_5761,N_5057,N_5441);
or U5762 (N_5762,N_5112,N_5141);
or U5763 (N_5763,N_5022,N_5426);
and U5764 (N_5764,N_5197,N_5401);
xor U5765 (N_5765,N_5380,N_5393);
xnor U5766 (N_5766,N_5231,N_5063);
and U5767 (N_5767,N_5137,N_5227);
or U5768 (N_5768,N_5291,N_5053);
or U5769 (N_5769,N_5030,N_5210);
nor U5770 (N_5770,N_5283,N_5355);
and U5771 (N_5771,N_5114,N_5183);
nor U5772 (N_5772,N_5340,N_5235);
or U5773 (N_5773,N_5265,N_5054);
nand U5774 (N_5774,N_5132,N_5390);
or U5775 (N_5775,N_5344,N_5208);
xnor U5776 (N_5776,N_5000,N_5049);
or U5777 (N_5777,N_5429,N_5401);
and U5778 (N_5778,N_5279,N_5339);
nand U5779 (N_5779,N_5187,N_5090);
and U5780 (N_5780,N_5269,N_5134);
nand U5781 (N_5781,N_5394,N_5207);
nand U5782 (N_5782,N_5356,N_5289);
nand U5783 (N_5783,N_5099,N_5177);
xnor U5784 (N_5784,N_5343,N_5209);
or U5785 (N_5785,N_5189,N_5140);
and U5786 (N_5786,N_5112,N_5408);
xnor U5787 (N_5787,N_5368,N_5347);
or U5788 (N_5788,N_5253,N_5047);
and U5789 (N_5789,N_5116,N_5498);
and U5790 (N_5790,N_5196,N_5314);
nor U5791 (N_5791,N_5123,N_5234);
or U5792 (N_5792,N_5153,N_5198);
and U5793 (N_5793,N_5285,N_5484);
and U5794 (N_5794,N_5113,N_5059);
nor U5795 (N_5795,N_5362,N_5251);
nor U5796 (N_5796,N_5356,N_5369);
nand U5797 (N_5797,N_5079,N_5294);
or U5798 (N_5798,N_5371,N_5435);
or U5799 (N_5799,N_5245,N_5247);
xnor U5800 (N_5800,N_5226,N_5227);
xor U5801 (N_5801,N_5137,N_5064);
nand U5802 (N_5802,N_5268,N_5283);
or U5803 (N_5803,N_5347,N_5106);
nor U5804 (N_5804,N_5038,N_5096);
and U5805 (N_5805,N_5362,N_5199);
nand U5806 (N_5806,N_5486,N_5239);
nor U5807 (N_5807,N_5337,N_5433);
nor U5808 (N_5808,N_5333,N_5123);
and U5809 (N_5809,N_5039,N_5331);
or U5810 (N_5810,N_5040,N_5241);
nand U5811 (N_5811,N_5444,N_5138);
and U5812 (N_5812,N_5452,N_5367);
or U5813 (N_5813,N_5286,N_5198);
xnor U5814 (N_5814,N_5341,N_5293);
nor U5815 (N_5815,N_5483,N_5295);
and U5816 (N_5816,N_5417,N_5083);
and U5817 (N_5817,N_5145,N_5292);
nor U5818 (N_5818,N_5045,N_5144);
or U5819 (N_5819,N_5000,N_5263);
nand U5820 (N_5820,N_5207,N_5035);
nand U5821 (N_5821,N_5305,N_5404);
nand U5822 (N_5822,N_5321,N_5308);
nand U5823 (N_5823,N_5410,N_5131);
and U5824 (N_5824,N_5231,N_5132);
nor U5825 (N_5825,N_5147,N_5455);
and U5826 (N_5826,N_5276,N_5096);
and U5827 (N_5827,N_5113,N_5211);
nor U5828 (N_5828,N_5114,N_5161);
nor U5829 (N_5829,N_5023,N_5194);
nor U5830 (N_5830,N_5497,N_5364);
and U5831 (N_5831,N_5109,N_5346);
nand U5832 (N_5832,N_5499,N_5452);
or U5833 (N_5833,N_5458,N_5198);
nand U5834 (N_5834,N_5121,N_5284);
nand U5835 (N_5835,N_5340,N_5126);
xnor U5836 (N_5836,N_5418,N_5424);
nand U5837 (N_5837,N_5223,N_5471);
nor U5838 (N_5838,N_5132,N_5244);
or U5839 (N_5839,N_5169,N_5114);
and U5840 (N_5840,N_5301,N_5453);
or U5841 (N_5841,N_5258,N_5376);
and U5842 (N_5842,N_5478,N_5435);
and U5843 (N_5843,N_5191,N_5464);
nand U5844 (N_5844,N_5286,N_5297);
nor U5845 (N_5845,N_5440,N_5383);
or U5846 (N_5846,N_5404,N_5330);
or U5847 (N_5847,N_5070,N_5096);
or U5848 (N_5848,N_5190,N_5076);
and U5849 (N_5849,N_5129,N_5209);
and U5850 (N_5850,N_5256,N_5492);
xor U5851 (N_5851,N_5091,N_5078);
nand U5852 (N_5852,N_5289,N_5040);
nor U5853 (N_5853,N_5078,N_5267);
or U5854 (N_5854,N_5343,N_5434);
or U5855 (N_5855,N_5447,N_5295);
or U5856 (N_5856,N_5254,N_5324);
nor U5857 (N_5857,N_5275,N_5287);
nor U5858 (N_5858,N_5018,N_5148);
nor U5859 (N_5859,N_5094,N_5348);
nand U5860 (N_5860,N_5390,N_5259);
nand U5861 (N_5861,N_5139,N_5134);
or U5862 (N_5862,N_5099,N_5499);
xor U5863 (N_5863,N_5428,N_5347);
nand U5864 (N_5864,N_5155,N_5454);
xor U5865 (N_5865,N_5196,N_5266);
or U5866 (N_5866,N_5454,N_5093);
or U5867 (N_5867,N_5348,N_5395);
nand U5868 (N_5868,N_5394,N_5102);
nand U5869 (N_5869,N_5148,N_5212);
nand U5870 (N_5870,N_5432,N_5489);
nand U5871 (N_5871,N_5025,N_5012);
nor U5872 (N_5872,N_5115,N_5286);
and U5873 (N_5873,N_5394,N_5335);
and U5874 (N_5874,N_5065,N_5228);
nand U5875 (N_5875,N_5239,N_5425);
xnor U5876 (N_5876,N_5434,N_5062);
and U5877 (N_5877,N_5379,N_5425);
xnor U5878 (N_5878,N_5309,N_5310);
nor U5879 (N_5879,N_5041,N_5388);
or U5880 (N_5880,N_5309,N_5234);
nand U5881 (N_5881,N_5372,N_5124);
or U5882 (N_5882,N_5057,N_5062);
nand U5883 (N_5883,N_5411,N_5202);
nand U5884 (N_5884,N_5066,N_5362);
nor U5885 (N_5885,N_5039,N_5389);
or U5886 (N_5886,N_5463,N_5279);
nand U5887 (N_5887,N_5357,N_5248);
and U5888 (N_5888,N_5285,N_5251);
nand U5889 (N_5889,N_5450,N_5028);
xor U5890 (N_5890,N_5449,N_5155);
nand U5891 (N_5891,N_5290,N_5367);
nor U5892 (N_5892,N_5236,N_5118);
or U5893 (N_5893,N_5461,N_5312);
nand U5894 (N_5894,N_5238,N_5333);
or U5895 (N_5895,N_5273,N_5263);
nor U5896 (N_5896,N_5150,N_5332);
xor U5897 (N_5897,N_5247,N_5457);
or U5898 (N_5898,N_5169,N_5120);
xnor U5899 (N_5899,N_5489,N_5405);
or U5900 (N_5900,N_5423,N_5414);
or U5901 (N_5901,N_5065,N_5037);
and U5902 (N_5902,N_5300,N_5337);
and U5903 (N_5903,N_5442,N_5493);
and U5904 (N_5904,N_5090,N_5207);
xnor U5905 (N_5905,N_5145,N_5211);
nand U5906 (N_5906,N_5448,N_5147);
and U5907 (N_5907,N_5314,N_5458);
nand U5908 (N_5908,N_5425,N_5490);
and U5909 (N_5909,N_5381,N_5405);
nand U5910 (N_5910,N_5472,N_5045);
nand U5911 (N_5911,N_5146,N_5188);
nor U5912 (N_5912,N_5489,N_5327);
nand U5913 (N_5913,N_5319,N_5378);
and U5914 (N_5914,N_5029,N_5312);
nor U5915 (N_5915,N_5146,N_5037);
nand U5916 (N_5916,N_5298,N_5211);
nor U5917 (N_5917,N_5489,N_5429);
nor U5918 (N_5918,N_5386,N_5343);
xor U5919 (N_5919,N_5047,N_5331);
or U5920 (N_5920,N_5234,N_5416);
and U5921 (N_5921,N_5224,N_5141);
or U5922 (N_5922,N_5081,N_5352);
nor U5923 (N_5923,N_5398,N_5057);
nand U5924 (N_5924,N_5401,N_5061);
nor U5925 (N_5925,N_5320,N_5003);
xor U5926 (N_5926,N_5381,N_5362);
nand U5927 (N_5927,N_5178,N_5140);
nor U5928 (N_5928,N_5096,N_5424);
nand U5929 (N_5929,N_5439,N_5203);
and U5930 (N_5930,N_5322,N_5264);
xor U5931 (N_5931,N_5075,N_5307);
and U5932 (N_5932,N_5001,N_5177);
nor U5933 (N_5933,N_5483,N_5155);
xnor U5934 (N_5934,N_5176,N_5301);
or U5935 (N_5935,N_5431,N_5293);
nor U5936 (N_5936,N_5365,N_5497);
nor U5937 (N_5937,N_5173,N_5319);
xor U5938 (N_5938,N_5497,N_5382);
or U5939 (N_5939,N_5367,N_5205);
nand U5940 (N_5940,N_5232,N_5070);
nand U5941 (N_5941,N_5128,N_5010);
and U5942 (N_5942,N_5412,N_5009);
or U5943 (N_5943,N_5237,N_5026);
nand U5944 (N_5944,N_5281,N_5480);
or U5945 (N_5945,N_5186,N_5021);
xor U5946 (N_5946,N_5148,N_5358);
and U5947 (N_5947,N_5129,N_5031);
xor U5948 (N_5948,N_5331,N_5169);
or U5949 (N_5949,N_5241,N_5096);
nor U5950 (N_5950,N_5248,N_5112);
xor U5951 (N_5951,N_5408,N_5290);
nor U5952 (N_5952,N_5083,N_5223);
or U5953 (N_5953,N_5055,N_5087);
nand U5954 (N_5954,N_5474,N_5184);
nand U5955 (N_5955,N_5342,N_5139);
nand U5956 (N_5956,N_5310,N_5447);
nor U5957 (N_5957,N_5360,N_5089);
nor U5958 (N_5958,N_5347,N_5459);
and U5959 (N_5959,N_5376,N_5083);
or U5960 (N_5960,N_5319,N_5325);
nor U5961 (N_5961,N_5114,N_5145);
or U5962 (N_5962,N_5346,N_5300);
and U5963 (N_5963,N_5398,N_5450);
and U5964 (N_5964,N_5133,N_5394);
xor U5965 (N_5965,N_5282,N_5075);
and U5966 (N_5966,N_5364,N_5152);
xor U5967 (N_5967,N_5075,N_5334);
and U5968 (N_5968,N_5333,N_5216);
nor U5969 (N_5969,N_5397,N_5341);
and U5970 (N_5970,N_5388,N_5240);
or U5971 (N_5971,N_5160,N_5459);
nor U5972 (N_5972,N_5248,N_5152);
nand U5973 (N_5973,N_5065,N_5110);
and U5974 (N_5974,N_5338,N_5273);
or U5975 (N_5975,N_5068,N_5396);
and U5976 (N_5976,N_5477,N_5434);
or U5977 (N_5977,N_5412,N_5154);
and U5978 (N_5978,N_5422,N_5389);
nor U5979 (N_5979,N_5192,N_5257);
nor U5980 (N_5980,N_5423,N_5186);
xnor U5981 (N_5981,N_5320,N_5343);
and U5982 (N_5982,N_5419,N_5035);
nor U5983 (N_5983,N_5448,N_5456);
nor U5984 (N_5984,N_5435,N_5201);
nor U5985 (N_5985,N_5251,N_5142);
nor U5986 (N_5986,N_5007,N_5336);
nor U5987 (N_5987,N_5370,N_5201);
xor U5988 (N_5988,N_5331,N_5072);
and U5989 (N_5989,N_5301,N_5276);
nor U5990 (N_5990,N_5150,N_5459);
xor U5991 (N_5991,N_5481,N_5093);
and U5992 (N_5992,N_5370,N_5393);
nor U5993 (N_5993,N_5215,N_5174);
or U5994 (N_5994,N_5022,N_5468);
nand U5995 (N_5995,N_5462,N_5342);
or U5996 (N_5996,N_5400,N_5112);
or U5997 (N_5997,N_5289,N_5435);
nor U5998 (N_5998,N_5407,N_5348);
and U5999 (N_5999,N_5095,N_5192);
nor U6000 (N_6000,N_5711,N_5817);
or U6001 (N_6001,N_5686,N_5973);
or U6002 (N_6002,N_5753,N_5909);
or U6003 (N_6003,N_5810,N_5510);
and U6004 (N_6004,N_5934,N_5698);
and U6005 (N_6005,N_5960,N_5693);
nor U6006 (N_6006,N_5680,N_5583);
and U6007 (N_6007,N_5563,N_5928);
xnor U6008 (N_6008,N_5559,N_5835);
xor U6009 (N_6009,N_5502,N_5856);
nand U6010 (N_6010,N_5906,N_5690);
xor U6011 (N_6011,N_5629,N_5791);
xnor U6012 (N_6012,N_5966,N_5819);
xor U6013 (N_6013,N_5780,N_5695);
nor U6014 (N_6014,N_5886,N_5815);
and U6015 (N_6015,N_5912,N_5808);
or U6016 (N_6016,N_5518,N_5859);
or U6017 (N_6017,N_5715,N_5801);
nor U6018 (N_6018,N_5950,N_5861);
nand U6019 (N_6019,N_5806,N_5643);
or U6020 (N_6020,N_5977,N_5972);
or U6021 (N_6021,N_5607,N_5903);
and U6022 (N_6022,N_5628,N_5752);
or U6023 (N_6023,N_5758,N_5764);
and U6024 (N_6024,N_5713,N_5888);
nor U6025 (N_6025,N_5831,N_5581);
xnor U6026 (N_6026,N_5814,N_5905);
or U6027 (N_6027,N_5595,N_5641);
nor U6028 (N_6028,N_5706,N_5805);
xnor U6029 (N_6029,N_5736,N_5959);
xnor U6030 (N_6030,N_5942,N_5967);
nand U6031 (N_6031,N_5738,N_5956);
and U6032 (N_6032,N_5996,N_5517);
and U6033 (N_6033,N_5847,N_5885);
xnor U6034 (N_6034,N_5919,N_5832);
nand U6035 (N_6035,N_5779,N_5900);
and U6036 (N_6036,N_5789,N_5932);
or U6037 (N_6037,N_5633,N_5917);
nand U6038 (N_6038,N_5655,N_5676);
and U6039 (N_6039,N_5648,N_5702);
and U6040 (N_6040,N_5634,N_5840);
or U6041 (N_6041,N_5936,N_5735);
xor U6042 (N_6042,N_5566,N_5976);
xor U6043 (N_6043,N_5908,N_5665);
and U6044 (N_6044,N_5710,N_5759);
xnor U6045 (N_6045,N_5747,N_5520);
and U6046 (N_6046,N_5845,N_5724);
and U6047 (N_6047,N_5667,N_5523);
nor U6048 (N_6048,N_5684,N_5569);
and U6049 (N_6049,N_5926,N_5534);
xor U6050 (N_6050,N_5714,N_5868);
nor U6051 (N_6051,N_5865,N_5874);
nor U6052 (N_6052,N_5842,N_5731);
nor U6053 (N_6053,N_5701,N_5526);
and U6054 (N_6054,N_5763,N_5744);
nand U6055 (N_6055,N_5683,N_5775);
nand U6056 (N_6056,N_5575,N_5866);
nand U6057 (N_6057,N_5631,N_5986);
xnor U6058 (N_6058,N_5708,N_5611);
nor U6059 (N_6059,N_5992,N_5915);
nor U6060 (N_6060,N_5864,N_5953);
and U6061 (N_6061,N_5982,N_5965);
and U6062 (N_6062,N_5538,N_5849);
nand U6063 (N_6063,N_5506,N_5687);
nand U6064 (N_6064,N_5910,N_5685);
or U6065 (N_6065,N_5688,N_5930);
or U6066 (N_6066,N_5567,N_5657);
nor U6067 (N_6067,N_5653,N_5732);
nand U6068 (N_6068,N_5858,N_5652);
xor U6069 (N_6069,N_5541,N_5841);
nor U6070 (N_6070,N_5991,N_5528);
nor U6071 (N_6071,N_5782,N_5556);
xnor U6072 (N_6072,N_5636,N_5597);
nor U6073 (N_6073,N_5794,N_5781);
nand U6074 (N_6074,N_5826,N_5830);
or U6075 (N_6075,N_5907,N_5968);
nand U6076 (N_6076,N_5659,N_5627);
nand U6077 (N_6077,N_5963,N_5602);
or U6078 (N_6078,N_5505,N_5621);
and U6079 (N_6079,N_5612,N_5703);
xnor U6080 (N_6080,N_5637,N_5700);
and U6081 (N_6081,N_5694,N_5516);
xnor U6082 (N_6082,N_5725,N_5705);
xor U6083 (N_6083,N_5639,N_5875);
nor U6084 (N_6084,N_5914,N_5925);
and U6085 (N_6085,N_5755,N_5591);
xnor U6086 (N_6086,N_5881,N_5798);
or U6087 (N_6087,N_5860,N_5571);
nor U6088 (N_6088,N_5589,N_5922);
or U6089 (N_6089,N_5560,N_5656);
xnor U6090 (N_6090,N_5924,N_5734);
xor U6091 (N_6091,N_5669,N_5957);
and U6092 (N_6092,N_5985,N_5843);
or U6093 (N_6093,N_5757,N_5943);
or U6094 (N_6094,N_5660,N_5890);
or U6095 (N_6095,N_5613,N_5527);
xnor U6096 (N_6096,N_5971,N_5696);
nor U6097 (N_6097,N_5772,N_5614);
or U6098 (N_6098,N_5618,N_5770);
xor U6099 (N_6099,N_5564,N_5557);
nor U6100 (N_6100,N_5709,N_5579);
nor U6101 (N_6101,N_5786,N_5941);
nor U6102 (N_6102,N_5540,N_5681);
nor U6103 (N_6103,N_5827,N_5729);
and U6104 (N_6104,N_5857,N_5978);
nor U6105 (N_6105,N_5813,N_5853);
nor U6106 (N_6106,N_5554,N_5839);
or U6107 (N_6107,N_5784,N_5716);
xor U6108 (N_6108,N_5501,N_5749);
and U6109 (N_6109,N_5604,N_5949);
xor U6110 (N_6110,N_5679,N_5773);
and U6111 (N_6111,N_5970,N_5507);
nand U6112 (N_6112,N_5938,N_5837);
xor U6113 (N_6113,N_5704,N_5783);
nor U6114 (N_6114,N_5542,N_5673);
or U6115 (N_6115,N_5593,N_5975);
or U6116 (N_6116,N_5882,N_5692);
xnor U6117 (N_6117,N_5848,N_5756);
xnor U6118 (N_6118,N_5532,N_5804);
and U6119 (N_6119,N_5997,N_5913);
or U6120 (N_6120,N_5987,N_5525);
xor U6121 (N_6121,N_5529,N_5577);
xnor U6122 (N_6122,N_5988,N_5619);
nor U6123 (N_6123,N_5879,N_5787);
nor U6124 (N_6124,N_5644,N_5568);
nand U6125 (N_6125,N_5661,N_5946);
nor U6126 (N_6126,N_5844,N_5598);
and U6127 (N_6127,N_5851,N_5723);
and U6128 (N_6128,N_5574,N_5902);
nand U6129 (N_6129,N_5767,N_5600);
nor U6130 (N_6130,N_5760,N_5741);
nor U6131 (N_6131,N_5547,N_5883);
xor U6132 (N_6132,N_5776,N_5682);
xor U6133 (N_6133,N_5521,N_5512);
nand U6134 (N_6134,N_5873,N_5620);
xor U6135 (N_6135,N_5699,N_5635);
and U6136 (N_6136,N_5592,N_5846);
xor U6137 (N_6137,N_5792,N_5552);
xor U6138 (N_6138,N_5573,N_5642);
xor U6139 (N_6139,N_5536,N_5964);
nor U6140 (N_6140,N_5901,N_5821);
nor U6141 (N_6141,N_5558,N_5720);
xnor U6142 (N_6142,N_5979,N_5766);
nand U6143 (N_6143,N_5721,N_5626);
xor U6144 (N_6144,N_5625,N_5834);
xnor U6145 (N_6145,N_5603,N_5609);
or U6146 (N_6146,N_5588,N_5855);
and U6147 (N_6147,N_5869,N_5954);
nand U6148 (N_6148,N_5630,N_5742);
and U6149 (N_6149,N_5722,N_5551);
nand U6150 (N_6150,N_5663,N_5990);
and U6151 (N_6151,N_5658,N_5668);
nor U6152 (N_6152,N_5500,N_5876);
xor U6153 (N_6153,N_5596,N_5546);
nand U6154 (N_6154,N_5646,N_5675);
and U6155 (N_6155,N_5825,N_5823);
or U6156 (N_6156,N_5727,N_5531);
nand U6157 (N_6157,N_5530,N_5923);
xnor U6158 (N_6158,N_5511,N_5945);
nor U6159 (N_6159,N_5891,N_5952);
or U6160 (N_6160,N_5896,N_5889);
and U6161 (N_6161,N_5691,N_5998);
or U6162 (N_6162,N_5993,N_5707);
xnor U6163 (N_6163,N_5862,N_5894);
or U6164 (N_6164,N_5533,N_5739);
and U6165 (N_6165,N_5820,N_5809);
nor U6166 (N_6166,N_5994,N_5623);
xnor U6167 (N_6167,N_5933,N_5553);
and U6168 (N_6168,N_5871,N_5615);
and U6169 (N_6169,N_5562,N_5867);
xor U6170 (N_6170,N_5638,N_5664);
and U6171 (N_6171,N_5921,N_5576);
and U6172 (N_6172,N_5584,N_5795);
nor U6173 (N_6173,N_5771,N_5748);
nand U6174 (N_6174,N_5649,N_5989);
nand U6175 (N_6175,N_5617,N_5899);
or U6176 (N_6176,N_5872,N_5951);
nand U6177 (N_6177,N_5544,N_5697);
or U6178 (N_6178,N_5980,N_5793);
and U6179 (N_6179,N_5537,N_5622);
xor U6180 (N_6180,N_5594,N_5800);
nand U6181 (N_6181,N_5565,N_5601);
nor U6182 (N_6182,N_5969,N_5790);
nand U6183 (N_6183,N_5895,N_5522);
nand U6184 (N_6184,N_5503,N_5893);
and U6185 (N_6185,N_5935,N_5981);
nor U6186 (N_6186,N_5671,N_5828);
xor U6187 (N_6187,N_5605,N_5666);
or U6188 (N_6188,N_5535,N_5816);
and U6189 (N_6189,N_5590,N_5898);
nand U6190 (N_6190,N_5931,N_5929);
nand U6191 (N_6191,N_5765,N_5911);
xnor U6192 (N_6192,N_5892,N_5740);
or U6193 (N_6193,N_5984,N_5927);
and U6194 (N_6194,N_5519,N_5587);
or U6195 (N_6195,N_5545,N_5948);
and U6196 (N_6196,N_5904,N_5548);
or U6197 (N_6197,N_5916,N_5730);
nor U6198 (N_6198,N_5983,N_5829);
or U6199 (N_6199,N_5778,N_5920);
nand U6200 (N_6200,N_5570,N_5797);
xor U6201 (N_6201,N_5572,N_5549);
nand U6202 (N_6202,N_5504,N_5513);
nand U6203 (N_6203,N_5751,N_5918);
nor U6204 (N_6204,N_5807,N_5754);
and U6205 (N_6205,N_5944,N_5750);
xnor U6206 (N_6206,N_5672,N_5677);
xnor U6207 (N_6207,N_5799,N_5958);
xnor U6208 (N_6208,N_5599,N_5774);
nor U6209 (N_6209,N_5850,N_5624);
and U6210 (N_6210,N_5647,N_5877);
and U6211 (N_6211,N_5650,N_5509);
nor U6212 (N_6212,N_5561,N_5818);
or U6213 (N_6213,N_5539,N_5670);
xor U6214 (N_6214,N_5822,N_5632);
nand U6215 (N_6215,N_5717,N_5796);
xor U6216 (N_6216,N_5610,N_5769);
xnor U6217 (N_6217,N_5974,N_5897);
nor U6218 (N_6218,N_5870,N_5838);
and U6219 (N_6219,N_5743,N_5728);
xor U6220 (N_6220,N_5550,N_5999);
or U6221 (N_6221,N_5863,N_5616);
and U6222 (N_6222,N_5947,N_5586);
nor U6223 (N_6223,N_5761,N_5645);
nand U6224 (N_6224,N_5606,N_5674);
xor U6225 (N_6225,N_5508,N_5737);
and U6226 (N_6226,N_5937,N_5961);
and U6227 (N_6227,N_5733,N_5803);
or U6228 (N_6228,N_5940,N_5662);
nor U6229 (N_6229,N_5580,N_5726);
nand U6230 (N_6230,N_5854,N_5651);
or U6231 (N_6231,N_5788,N_5719);
nand U6232 (N_6232,N_5811,N_5887);
nor U6233 (N_6233,N_5640,N_5824);
nand U6234 (N_6234,N_5878,N_5718);
nor U6235 (N_6235,N_5880,N_5762);
and U6236 (N_6236,N_5654,N_5582);
xor U6237 (N_6237,N_5852,N_5785);
nor U6238 (N_6238,N_5585,N_5777);
and U6239 (N_6239,N_5812,N_5746);
nor U6240 (N_6240,N_5962,N_5608);
and U6241 (N_6241,N_5833,N_5836);
xor U6242 (N_6242,N_5884,N_5689);
or U6243 (N_6243,N_5543,N_5678);
and U6244 (N_6244,N_5524,N_5802);
xor U6245 (N_6245,N_5578,N_5515);
and U6246 (N_6246,N_5995,N_5768);
xor U6247 (N_6247,N_5745,N_5514);
nor U6248 (N_6248,N_5955,N_5555);
and U6249 (N_6249,N_5712,N_5939);
nor U6250 (N_6250,N_5590,N_5505);
and U6251 (N_6251,N_5949,N_5947);
and U6252 (N_6252,N_5765,N_5771);
nor U6253 (N_6253,N_5642,N_5949);
or U6254 (N_6254,N_5877,N_5743);
and U6255 (N_6255,N_5725,N_5788);
nand U6256 (N_6256,N_5870,N_5796);
or U6257 (N_6257,N_5973,N_5735);
and U6258 (N_6258,N_5978,N_5684);
nor U6259 (N_6259,N_5635,N_5549);
nand U6260 (N_6260,N_5976,N_5512);
nand U6261 (N_6261,N_5682,N_5652);
or U6262 (N_6262,N_5562,N_5578);
or U6263 (N_6263,N_5626,N_5896);
nor U6264 (N_6264,N_5724,N_5977);
and U6265 (N_6265,N_5630,N_5522);
xnor U6266 (N_6266,N_5589,N_5746);
and U6267 (N_6267,N_5509,N_5685);
xnor U6268 (N_6268,N_5623,N_5515);
and U6269 (N_6269,N_5893,N_5660);
or U6270 (N_6270,N_5995,N_5537);
nor U6271 (N_6271,N_5692,N_5989);
nand U6272 (N_6272,N_5758,N_5557);
nor U6273 (N_6273,N_5718,N_5714);
and U6274 (N_6274,N_5741,N_5514);
nand U6275 (N_6275,N_5824,N_5687);
and U6276 (N_6276,N_5817,N_5890);
nor U6277 (N_6277,N_5999,N_5952);
and U6278 (N_6278,N_5709,N_5852);
nor U6279 (N_6279,N_5948,N_5720);
nand U6280 (N_6280,N_5907,N_5756);
or U6281 (N_6281,N_5517,N_5507);
and U6282 (N_6282,N_5703,N_5952);
or U6283 (N_6283,N_5989,N_5731);
nand U6284 (N_6284,N_5886,N_5872);
and U6285 (N_6285,N_5779,N_5951);
nor U6286 (N_6286,N_5556,N_5714);
nor U6287 (N_6287,N_5980,N_5932);
and U6288 (N_6288,N_5733,N_5706);
xnor U6289 (N_6289,N_5601,N_5542);
or U6290 (N_6290,N_5568,N_5897);
nor U6291 (N_6291,N_5883,N_5528);
nor U6292 (N_6292,N_5687,N_5567);
nand U6293 (N_6293,N_5765,N_5779);
nor U6294 (N_6294,N_5678,N_5505);
xor U6295 (N_6295,N_5701,N_5524);
and U6296 (N_6296,N_5798,N_5546);
nand U6297 (N_6297,N_5972,N_5854);
xor U6298 (N_6298,N_5696,N_5825);
xor U6299 (N_6299,N_5777,N_5644);
nor U6300 (N_6300,N_5785,N_5960);
nand U6301 (N_6301,N_5625,N_5998);
nor U6302 (N_6302,N_5920,N_5898);
xor U6303 (N_6303,N_5909,N_5846);
or U6304 (N_6304,N_5866,N_5770);
xor U6305 (N_6305,N_5673,N_5932);
nor U6306 (N_6306,N_5997,N_5985);
nor U6307 (N_6307,N_5987,N_5819);
or U6308 (N_6308,N_5720,N_5847);
nor U6309 (N_6309,N_5618,N_5775);
xnor U6310 (N_6310,N_5865,N_5990);
or U6311 (N_6311,N_5866,N_5989);
and U6312 (N_6312,N_5562,N_5963);
nor U6313 (N_6313,N_5979,N_5568);
nor U6314 (N_6314,N_5775,N_5773);
or U6315 (N_6315,N_5602,N_5654);
xnor U6316 (N_6316,N_5510,N_5993);
xnor U6317 (N_6317,N_5605,N_5723);
xnor U6318 (N_6318,N_5558,N_5962);
and U6319 (N_6319,N_5611,N_5657);
or U6320 (N_6320,N_5570,N_5941);
nor U6321 (N_6321,N_5722,N_5559);
xor U6322 (N_6322,N_5846,N_5508);
nor U6323 (N_6323,N_5508,N_5689);
nand U6324 (N_6324,N_5970,N_5855);
nor U6325 (N_6325,N_5524,N_5506);
nand U6326 (N_6326,N_5728,N_5597);
and U6327 (N_6327,N_5703,N_5508);
nor U6328 (N_6328,N_5896,N_5739);
nand U6329 (N_6329,N_5723,N_5996);
or U6330 (N_6330,N_5871,N_5964);
nand U6331 (N_6331,N_5959,N_5703);
or U6332 (N_6332,N_5854,N_5701);
and U6333 (N_6333,N_5837,N_5601);
and U6334 (N_6334,N_5673,N_5513);
and U6335 (N_6335,N_5710,N_5716);
or U6336 (N_6336,N_5523,N_5641);
xnor U6337 (N_6337,N_5899,N_5806);
nor U6338 (N_6338,N_5939,N_5719);
nand U6339 (N_6339,N_5910,N_5827);
nand U6340 (N_6340,N_5536,N_5563);
xor U6341 (N_6341,N_5793,N_5900);
and U6342 (N_6342,N_5539,N_5566);
nand U6343 (N_6343,N_5761,N_5756);
nand U6344 (N_6344,N_5894,N_5875);
and U6345 (N_6345,N_5690,N_5550);
nand U6346 (N_6346,N_5559,N_5687);
nor U6347 (N_6347,N_5847,N_5814);
or U6348 (N_6348,N_5951,N_5582);
or U6349 (N_6349,N_5969,N_5683);
or U6350 (N_6350,N_5545,N_5842);
or U6351 (N_6351,N_5719,N_5706);
nand U6352 (N_6352,N_5545,N_5931);
xor U6353 (N_6353,N_5699,N_5957);
nand U6354 (N_6354,N_5809,N_5845);
xor U6355 (N_6355,N_5889,N_5897);
and U6356 (N_6356,N_5708,N_5541);
and U6357 (N_6357,N_5602,N_5899);
xnor U6358 (N_6358,N_5544,N_5649);
nand U6359 (N_6359,N_5816,N_5836);
nand U6360 (N_6360,N_5574,N_5919);
and U6361 (N_6361,N_5807,N_5782);
or U6362 (N_6362,N_5838,N_5951);
and U6363 (N_6363,N_5717,N_5530);
xnor U6364 (N_6364,N_5805,N_5900);
xnor U6365 (N_6365,N_5837,N_5838);
and U6366 (N_6366,N_5596,N_5841);
and U6367 (N_6367,N_5987,N_5672);
or U6368 (N_6368,N_5739,N_5752);
nor U6369 (N_6369,N_5891,N_5875);
nand U6370 (N_6370,N_5661,N_5798);
or U6371 (N_6371,N_5908,N_5746);
nand U6372 (N_6372,N_5587,N_5590);
xnor U6373 (N_6373,N_5863,N_5748);
or U6374 (N_6374,N_5592,N_5591);
nor U6375 (N_6375,N_5820,N_5619);
nand U6376 (N_6376,N_5505,N_5902);
and U6377 (N_6377,N_5707,N_5866);
or U6378 (N_6378,N_5672,N_5897);
or U6379 (N_6379,N_5558,N_5745);
and U6380 (N_6380,N_5960,N_5527);
nor U6381 (N_6381,N_5685,N_5558);
and U6382 (N_6382,N_5776,N_5808);
nand U6383 (N_6383,N_5934,N_5800);
and U6384 (N_6384,N_5973,N_5527);
nor U6385 (N_6385,N_5856,N_5524);
nand U6386 (N_6386,N_5848,N_5866);
nor U6387 (N_6387,N_5987,N_5843);
xnor U6388 (N_6388,N_5954,N_5958);
or U6389 (N_6389,N_5915,N_5839);
and U6390 (N_6390,N_5980,N_5844);
or U6391 (N_6391,N_5656,N_5877);
nand U6392 (N_6392,N_5740,N_5613);
and U6393 (N_6393,N_5830,N_5586);
xnor U6394 (N_6394,N_5681,N_5967);
or U6395 (N_6395,N_5797,N_5739);
and U6396 (N_6396,N_5714,N_5735);
nand U6397 (N_6397,N_5812,N_5954);
and U6398 (N_6398,N_5916,N_5905);
or U6399 (N_6399,N_5815,N_5851);
nand U6400 (N_6400,N_5941,N_5848);
nand U6401 (N_6401,N_5871,N_5919);
or U6402 (N_6402,N_5686,N_5875);
xor U6403 (N_6403,N_5637,N_5582);
xor U6404 (N_6404,N_5533,N_5895);
or U6405 (N_6405,N_5864,N_5632);
nand U6406 (N_6406,N_5657,N_5780);
or U6407 (N_6407,N_5962,N_5967);
and U6408 (N_6408,N_5915,N_5700);
nand U6409 (N_6409,N_5652,N_5931);
and U6410 (N_6410,N_5562,N_5708);
nand U6411 (N_6411,N_5742,N_5924);
xor U6412 (N_6412,N_5568,N_5610);
nor U6413 (N_6413,N_5591,N_5657);
nor U6414 (N_6414,N_5588,N_5953);
nand U6415 (N_6415,N_5979,N_5755);
or U6416 (N_6416,N_5550,N_5972);
or U6417 (N_6417,N_5540,N_5815);
or U6418 (N_6418,N_5951,N_5523);
xor U6419 (N_6419,N_5676,N_5950);
and U6420 (N_6420,N_5625,N_5517);
and U6421 (N_6421,N_5536,N_5646);
and U6422 (N_6422,N_5957,N_5530);
xnor U6423 (N_6423,N_5528,N_5979);
nand U6424 (N_6424,N_5732,N_5684);
and U6425 (N_6425,N_5959,N_5726);
or U6426 (N_6426,N_5512,N_5886);
nor U6427 (N_6427,N_5873,N_5524);
or U6428 (N_6428,N_5620,N_5677);
nor U6429 (N_6429,N_5594,N_5988);
xor U6430 (N_6430,N_5522,N_5945);
and U6431 (N_6431,N_5795,N_5674);
or U6432 (N_6432,N_5764,N_5798);
or U6433 (N_6433,N_5596,N_5878);
or U6434 (N_6434,N_5999,N_5834);
nand U6435 (N_6435,N_5694,N_5902);
or U6436 (N_6436,N_5855,N_5683);
and U6437 (N_6437,N_5531,N_5660);
xor U6438 (N_6438,N_5628,N_5970);
and U6439 (N_6439,N_5755,N_5945);
nand U6440 (N_6440,N_5612,N_5536);
or U6441 (N_6441,N_5511,N_5646);
xor U6442 (N_6442,N_5860,N_5620);
and U6443 (N_6443,N_5873,N_5895);
and U6444 (N_6444,N_5826,N_5724);
xnor U6445 (N_6445,N_5622,N_5881);
or U6446 (N_6446,N_5703,N_5874);
xor U6447 (N_6447,N_5602,N_5558);
or U6448 (N_6448,N_5961,N_5896);
or U6449 (N_6449,N_5739,N_5826);
nand U6450 (N_6450,N_5710,N_5964);
xnor U6451 (N_6451,N_5970,N_5838);
xor U6452 (N_6452,N_5874,N_5636);
xor U6453 (N_6453,N_5823,N_5868);
xor U6454 (N_6454,N_5733,N_5540);
xor U6455 (N_6455,N_5770,N_5515);
and U6456 (N_6456,N_5700,N_5555);
xor U6457 (N_6457,N_5577,N_5641);
nand U6458 (N_6458,N_5705,N_5927);
nand U6459 (N_6459,N_5554,N_5661);
nand U6460 (N_6460,N_5688,N_5749);
nand U6461 (N_6461,N_5515,N_5576);
and U6462 (N_6462,N_5872,N_5916);
xor U6463 (N_6463,N_5956,N_5875);
nand U6464 (N_6464,N_5579,N_5674);
and U6465 (N_6465,N_5805,N_5573);
xnor U6466 (N_6466,N_5692,N_5945);
and U6467 (N_6467,N_5551,N_5553);
nand U6468 (N_6468,N_5575,N_5988);
and U6469 (N_6469,N_5987,N_5950);
or U6470 (N_6470,N_5502,N_5639);
nand U6471 (N_6471,N_5589,N_5891);
and U6472 (N_6472,N_5505,N_5771);
and U6473 (N_6473,N_5565,N_5901);
nor U6474 (N_6474,N_5999,N_5803);
xor U6475 (N_6475,N_5578,N_5703);
nand U6476 (N_6476,N_5598,N_5516);
xnor U6477 (N_6477,N_5897,N_5698);
nor U6478 (N_6478,N_5693,N_5953);
and U6479 (N_6479,N_5878,N_5999);
xnor U6480 (N_6480,N_5806,N_5938);
and U6481 (N_6481,N_5515,N_5647);
or U6482 (N_6482,N_5936,N_5979);
xnor U6483 (N_6483,N_5521,N_5510);
and U6484 (N_6484,N_5547,N_5885);
xor U6485 (N_6485,N_5815,N_5747);
xor U6486 (N_6486,N_5617,N_5556);
and U6487 (N_6487,N_5957,N_5800);
xnor U6488 (N_6488,N_5792,N_5932);
and U6489 (N_6489,N_5615,N_5570);
or U6490 (N_6490,N_5645,N_5852);
xnor U6491 (N_6491,N_5850,N_5562);
and U6492 (N_6492,N_5852,N_5511);
and U6493 (N_6493,N_5511,N_5529);
xor U6494 (N_6494,N_5891,N_5976);
xor U6495 (N_6495,N_5543,N_5627);
xnor U6496 (N_6496,N_5783,N_5804);
nor U6497 (N_6497,N_5583,N_5523);
or U6498 (N_6498,N_5687,N_5915);
xnor U6499 (N_6499,N_5869,N_5883);
or U6500 (N_6500,N_6032,N_6227);
xnor U6501 (N_6501,N_6479,N_6012);
nor U6502 (N_6502,N_6363,N_6486);
nand U6503 (N_6503,N_6317,N_6331);
xor U6504 (N_6504,N_6382,N_6308);
xor U6505 (N_6505,N_6006,N_6294);
nand U6506 (N_6506,N_6100,N_6403);
nand U6507 (N_6507,N_6328,N_6417);
or U6508 (N_6508,N_6264,N_6368);
or U6509 (N_6509,N_6322,N_6282);
nor U6510 (N_6510,N_6029,N_6082);
or U6511 (N_6511,N_6393,N_6121);
or U6512 (N_6512,N_6452,N_6267);
and U6513 (N_6513,N_6451,N_6206);
nor U6514 (N_6514,N_6341,N_6369);
nand U6515 (N_6515,N_6004,N_6350);
xnor U6516 (N_6516,N_6494,N_6216);
nor U6517 (N_6517,N_6288,N_6370);
nand U6518 (N_6518,N_6050,N_6063);
or U6519 (N_6519,N_6321,N_6318);
nand U6520 (N_6520,N_6073,N_6181);
and U6521 (N_6521,N_6477,N_6221);
nand U6522 (N_6522,N_6003,N_6296);
and U6523 (N_6523,N_6236,N_6078);
and U6524 (N_6524,N_6064,N_6258);
or U6525 (N_6525,N_6356,N_6414);
nand U6526 (N_6526,N_6239,N_6168);
and U6527 (N_6527,N_6250,N_6401);
and U6528 (N_6528,N_6231,N_6420);
xor U6529 (N_6529,N_6210,N_6375);
and U6530 (N_6530,N_6232,N_6223);
or U6531 (N_6531,N_6333,N_6085);
nand U6532 (N_6532,N_6238,N_6048);
nor U6533 (N_6533,N_6358,N_6315);
and U6534 (N_6534,N_6444,N_6243);
nand U6535 (N_6535,N_6274,N_6237);
nand U6536 (N_6536,N_6201,N_6017);
xor U6537 (N_6537,N_6482,N_6057);
or U6538 (N_6538,N_6359,N_6247);
or U6539 (N_6539,N_6449,N_6066);
nor U6540 (N_6540,N_6466,N_6304);
xnor U6541 (N_6541,N_6244,N_6240);
or U6542 (N_6542,N_6086,N_6139);
xnor U6543 (N_6543,N_6390,N_6122);
or U6544 (N_6544,N_6001,N_6007);
xor U6545 (N_6545,N_6203,N_6445);
nor U6546 (N_6546,N_6481,N_6079);
nor U6547 (N_6547,N_6010,N_6182);
nor U6548 (N_6548,N_6126,N_6355);
nand U6549 (N_6549,N_6438,N_6123);
nand U6550 (N_6550,N_6465,N_6125);
xor U6551 (N_6551,N_6097,N_6072);
nor U6552 (N_6552,N_6140,N_6141);
nand U6553 (N_6553,N_6474,N_6045);
or U6554 (N_6554,N_6406,N_6346);
or U6555 (N_6555,N_6084,N_6169);
nand U6556 (N_6556,N_6380,N_6415);
xor U6557 (N_6557,N_6177,N_6398);
nand U6558 (N_6558,N_6460,N_6497);
and U6559 (N_6559,N_6196,N_6259);
or U6560 (N_6560,N_6348,N_6336);
or U6561 (N_6561,N_6040,N_6150);
or U6562 (N_6562,N_6278,N_6291);
or U6563 (N_6563,N_6316,N_6428);
or U6564 (N_6564,N_6246,N_6448);
or U6565 (N_6565,N_6166,N_6133);
or U6566 (N_6566,N_6186,N_6446);
or U6567 (N_6567,N_6046,N_6260);
xor U6568 (N_6568,N_6340,N_6293);
nor U6569 (N_6569,N_6262,N_6491);
and U6570 (N_6570,N_6202,N_6018);
nor U6571 (N_6571,N_6156,N_6329);
and U6572 (N_6572,N_6307,N_6047);
xor U6573 (N_6573,N_6127,N_6495);
nand U6574 (N_6574,N_6049,N_6395);
nor U6575 (N_6575,N_6034,N_6372);
xnor U6576 (N_6576,N_6042,N_6379);
nand U6577 (N_6577,N_6480,N_6245);
nand U6578 (N_6578,N_6038,N_6263);
and U6579 (N_6579,N_6015,N_6478);
and U6580 (N_6580,N_6441,N_6151);
xnor U6581 (N_6581,N_6021,N_6374);
or U6582 (N_6582,N_6005,N_6373);
xnor U6583 (N_6583,N_6266,N_6104);
or U6584 (N_6584,N_6284,N_6213);
nor U6585 (N_6585,N_6404,N_6089);
nor U6586 (N_6586,N_6023,N_6002);
and U6587 (N_6587,N_6337,N_6458);
or U6588 (N_6588,N_6024,N_6187);
or U6589 (N_6589,N_6136,N_6043);
or U6590 (N_6590,N_6419,N_6191);
nor U6591 (N_6591,N_6060,N_6192);
xnor U6592 (N_6592,N_6114,N_6167);
nor U6593 (N_6593,N_6305,N_6366);
nor U6594 (N_6594,N_6313,N_6039);
and U6595 (N_6595,N_6378,N_6439);
nor U6596 (N_6596,N_6416,N_6459);
nor U6597 (N_6597,N_6146,N_6137);
and U6598 (N_6598,N_6334,N_6070);
nor U6599 (N_6599,N_6008,N_6099);
and U6600 (N_6600,N_6014,N_6352);
xnor U6601 (N_6601,N_6143,N_6484);
xnor U6602 (N_6602,N_6091,N_6455);
or U6603 (N_6603,N_6011,N_6389);
nand U6604 (N_6604,N_6179,N_6434);
or U6605 (N_6605,N_6306,N_6279);
or U6606 (N_6606,N_6364,N_6431);
and U6607 (N_6607,N_6440,N_6424);
xor U6608 (N_6608,N_6075,N_6295);
and U6609 (N_6609,N_6176,N_6081);
or U6610 (N_6610,N_6226,N_6098);
xnor U6611 (N_6611,N_6129,N_6092);
xnor U6612 (N_6612,N_6093,N_6160);
or U6613 (N_6613,N_6487,N_6178);
or U6614 (N_6614,N_6319,N_6116);
or U6615 (N_6615,N_6158,N_6432);
or U6616 (N_6616,N_6059,N_6095);
and U6617 (N_6617,N_6037,N_6138);
nor U6618 (N_6618,N_6184,N_6469);
or U6619 (N_6619,N_6430,N_6462);
and U6620 (N_6620,N_6426,N_6292);
and U6621 (N_6621,N_6286,N_6450);
nor U6622 (N_6622,N_6118,N_6120);
and U6623 (N_6623,N_6036,N_6147);
nor U6624 (N_6624,N_6498,N_6212);
xor U6625 (N_6625,N_6035,N_6344);
and U6626 (N_6626,N_6483,N_6130);
and U6627 (N_6627,N_6105,N_6367);
nor U6628 (N_6628,N_6219,N_6200);
and U6629 (N_6629,N_6400,N_6311);
xnor U6630 (N_6630,N_6000,N_6214);
or U6631 (N_6631,N_6044,N_6396);
nand U6632 (N_6632,N_6323,N_6392);
and U6633 (N_6633,N_6157,N_6290);
and U6634 (N_6634,N_6302,N_6220);
nor U6635 (N_6635,N_6327,N_6051);
and U6636 (N_6636,N_6019,N_6028);
xnor U6637 (N_6637,N_6235,N_6229);
xor U6638 (N_6638,N_6280,N_6111);
xnor U6639 (N_6639,N_6303,N_6471);
xnor U6640 (N_6640,N_6159,N_6224);
or U6641 (N_6641,N_6332,N_6496);
xor U6642 (N_6642,N_6467,N_6205);
nand U6643 (N_6643,N_6222,N_6463);
or U6644 (N_6644,N_6270,N_6488);
or U6645 (N_6645,N_6485,N_6300);
xor U6646 (N_6646,N_6054,N_6058);
nand U6647 (N_6647,N_6285,N_6476);
and U6648 (N_6648,N_6009,N_6189);
or U6649 (N_6649,N_6330,N_6335);
nor U6650 (N_6650,N_6065,N_6161);
or U6651 (N_6651,N_6371,N_6080);
nand U6652 (N_6652,N_6413,N_6094);
nor U6653 (N_6653,N_6277,N_6443);
nor U6654 (N_6654,N_6338,N_6387);
and U6655 (N_6655,N_6408,N_6394);
or U6656 (N_6656,N_6041,N_6257);
and U6657 (N_6657,N_6272,N_6310);
nor U6658 (N_6658,N_6088,N_6265);
or U6659 (N_6659,N_6261,N_6351);
xor U6660 (N_6660,N_6384,N_6436);
xor U6661 (N_6661,N_6271,N_6030);
and U6662 (N_6662,N_6197,N_6248);
or U6663 (N_6663,N_6254,N_6067);
nand U6664 (N_6664,N_6255,N_6405);
xor U6665 (N_6665,N_6230,N_6457);
nand U6666 (N_6666,N_6013,N_6171);
or U6667 (N_6667,N_6135,N_6437);
or U6668 (N_6668,N_6145,N_6252);
xor U6669 (N_6669,N_6362,N_6402);
or U6670 (N_6670,N_6134,N_6112);
nand U6671 (N_6671,N_6407,N_6052);
xnor U6672 (N_6672,N_6148,N_6218);
or U6673 (N_6673,N_6283,N_6102);
and U6674 (N_6674,N_6170,N_6251);
xor U6675 (N_6675,N_6386,N_6076);
nand U6676 (N_6676,N_6025,N_6115);
xnor U6677 (N_6677,N_6109,N_6031);
or U6678 (N_6678,N_6113,N_6193);
xnor U6679 (N_6679,N_6022,N_6108);
xor U6680 (N_6680,N_6273,N_6339);
nand U6681 (N_6681,N_6312,N_6198);
nor U6682 (N_6682,N_6175,N_6268);
nor U6683 (N_6683,N_6233,N_6183);
and U6684 (N_6684,N_6299,N_6298);
or U6685 (N_6685,N_6061,N_6360);
or U6686 (N_6686,N_6454,N_6103);
nor U6687 (N_6687,N_6020,N_6194);
and U6688 (N_6688,N_6074,N_6253);
nand U6689 (N_6689,N_6409,N_6204);
or U6690 (N_6690,N_6425,N_6256);
xor U6691 (N_6691,N_6185,N_6301);
xnor U6692 (N_6692,N_6472,N_6365);
xor U6693 (N_6693,N_6208,N_6132);
or U6694 (N_6694,N_6090,N_6033);
or U6695 (N_6695,N_6473,N_6199);
or U6696 (N_6696,N_6107,N_6418);
xnor U6697 (N_6697,N_6149,N_6096);
xnor U6698 (N_6698,N_6281,N_6016);
or U6699 (N_6699,N_6314,N_6433);
and U6700 (N_6700,N_6217,N_6297);
or U6701 (N_6701,N_6131,N_6453);
xnor U6702 (N_6702,N_6289,N_6153);
nor U6703 (N_6703,N_6228,N_6397);
or U6704 (N_6704,N_6381,N_6174);
xor U6705 (N_6705,N_6361,N_6275);
or U6706 (N_6706,N_6309,N_6461);
nor U6707 (N_6707,N_6056,N_6071);
nor U6708 (N_6708,N_6468,N_6209);
nand U6709 (N_6709,N_6357,N_6142);
nand U6710 (N_6710,N_6225,N_6412);
and U6711 (N_6711,N_6242,N_6195);
xnor U6712 (N_6712,N_6423,N_6053);
or U6713 (N_6713,N_6173,N_6421);
nand U6714 (N_6714,N_6342,N_6427);
xnor U6715 (N_6715,N_6101,N_6124);
and U6716 (N_6716,N_6087,N_6083);
nor U6717 (N_6717,N_6349,N_6026);
nand U6718 (N_6718,N_6347,N_6383);
and U6719 (N_6719,N_6027,N_6055);
xnor U6720 (N_6720,N_6207,N_6155);
xnor U6721 (N_6721,N_6276,N_6211);
and U6722 (N_6722,N_6429,N_6117);
and U6723 (N_6723,N_6470,N_6410);
or U6724 (N_6724,N_6106,N_6490);
xnor U6725 (N_6725,N_6377,N_6324);
xnor U6726 (N_6726,N_6345,N_6442);
nor U6727 (N_6727,N_6399,N_6287);
xnor U6728 (N_6728,N_6326,N_6391);
and U6729 (N_6729,N_6343,N_6215);
nand U6730 (N_6730,N_6110,N_6128);
nand U6731 (N_6731,N_6077,N_6456);
nand U6732 (N_6732,N_6154,N_6241);
nand U6733 (N_6733,N_6464,N_6234);
or U6734 (N_6734,N_6475,N_6489);
or U6735 (N_6735,N_6119,N_6188);
nor U6736 (N_6736,N_6144,N_6163);
or U6737 (N_6737,N_6411,N_6492);
and U6738 (N_6738,N_6062,N_6164);
xnor U6739 (N_6739,N_6499,N_6354);
or U6740 (N_6740,N_6152,N_6069);
and U6741 (N_6741,N_6376,N_6422);
and U6742 (N_6742,N_6180,N_6162);
nand U6743 (N_6743,N_6172,N_6493);
nor U6744 (N_6744,N_6249,N_6447);
xor U6745 (N_6745,N_6353,N_6190);
nand U6746 (N_6746,N_6165,N_6388);
and U6747 (N_6747,N_6385,N_6068);
nand U6748 (N_6748,N_6320,N_6325);
or U6749 (N_6749,N_6435,N_6269);
nand U6750 (N_6750,N_6383,N_6223);
xor U6751 (N_6751,N_6139,N_6071);
or U6752 (N_6752,N_6131,N_6084);
xnor U6753 (N_6753,N_6489,N_6212);
nor U6754 (N_6754,N_6462,N_6061);
and U6755 (N_6755,N_6288,N_6024);
and U6756 (N_6756,N_6468,N_6223);
xnor U6757 (N_6757,N_6008,N_6028);
xor U6758 (N_6758,N_6076,N_6353);
and U6759 (N_6759,N_6426,N_6109);
xor U6760 (N_6760,N_6225,N_6014);
xnor U6761 (N_6761,N_6229,N_6094);
and U6762 (N_6762,N_6108,N_6219);
nor U6763 (N_6763,N_6497,N_6194);
xnor U6764 (N_6764,N_6056,N_6091);
nand U6765 (N_6765,N_6088,N_6175);
and U6766 (N_6766,N_6009,N_6368);
or U6767 (N_6767,N_6337,N_6094);
nand U6768 (N_6768,N_6349,N_6327);
or U6769 (N_6769,N_6379,N_6483);
xor U6770 (N_6770,N_6423,N_6299);
xor U6771 (N_6771,N_6359,N_6099);
nor U6772 (N_6772,N_6067,N_6193);
and U6773 (N_6773,N_6458,N_6319);
nand U6774 (N_6774,N_6409,N_6161);
and U6775 (N_6775,N_6148,N_6321);
and U6776 (N_6776,N_6269,N_6265);
and U6777 (N_6777,N_6066,N_6023);
nor U6778 (N_6778,N_6452,N_6471);
and U6779 (N_6779,N_6212,N_6028);
xnor U6780 (N_6780,N_6188,N_6273);
or U6781 (N_6781,N_6273,N_6179);
nand U6782 (N_6782,N_6385,N_6245);
xor U6783 (N_6783,N_6440,N_6341);
nand U6784 (N_6784,N_6124,N_6087);
and U6785 (N_6785,N_6374,N_6318);
xnor U6786 (N_6786,N_6153,N_6168);
and U6787 (N_6787,N_6431,N_6403);
xor U6788 (N_6788,N_6136,N_6229);
or U6789 (N_6789,N_6481,N_6124);
or U6790 (N_6790,N_6242,N_6475);
or U6791 (N_6791,N_6098,N_6290);
nand U6792 (N_6792,N_6036,N_6345);
nor U6793 (N_6793,N_6257,N_6078);
nor U6794 (N_6794,N_6198,N_6017);
or U6795 (N_6795,N_6040,N_6256);
xor U6796 (N_6796,N_6134,N_6382);
nand U6797 (N_6797,N_6469,N_6172);
and U6798 (N_6798,N_6080,N_6177);
nor U6799 (N_6799,N_6200,N_6238);
nor U6800 (N_6800,N_6361,N_6120);
and U6801 (N_6801,N_6362,N_6071);
or U6802 (N_6802,N_6368,N_6375);
xor U6803 (N_6803,N_6385,N_6476);
nor U6804 (N_6804,N_6152,N_6314);
nand U6805 (N_6805,N_6303,N_6291);
xnor U6806 (N_6806,N_6032,N_6201);
nand U6807 (N_6807,N_6184,N_6315);
and U6808 (N_6808,N_6414,N_6089);
nand U6809 (N_6809,N_6018,N_6238);
nand U6810 (N_6810,N_6229,N_6035);
xor U6811 (N_6811,N_6175,N_6372);
xor U6812 (N_6812,N_6246,N_6164);
xor U6813 (N_6813,N_6056,N_6193);
nor U6814 (N_6814,N_6115,N_6380);
nor U6815 (N_6815,N_6036,N_6321);
nor U6816 (N_6816,N_6436,N_6320);
or U6817 (N_6817,N_6098,N_6159);
and U6818 (N_6818,N_6118,N_6200);
nand U6819 (N_6819,N_6344,N_6114);
or U6820 (N_6820,N_6080,N_6056);
xor U6821 (N_6821,N_6129,N_6376);
or U6822 (N_6822,N_6176,N_6446);
nor U6823 (N_6823,N_6249,N_6043);
or U6824 (N_6824,N_6053,N_6384);
nor U6825 (N_6825,N_6353,N_6388);
and U6826 (N_6826,N_6440,N_6347);
nor U6827 (N_6827,N_6490,N_6221);
or U6828 (N_6828,N_6212,N_6302);
and U6829 (N_6829,N_6210,N_6141);
and U6830 (N_6830,N_6348,N_6436);
nor U6831 (N_6831,N_6338,N_6498);
xor U6832 (N_6832,N_6040,N_6185);
or U6833 (N_6833,N_6484,N_6378);
xor U6834 (N_6834,N_6111,N_6029);
xnor U6835 (N_6835,N_6497,N_6155);
nand U6836 (N_6836,N_6313,N_6454);
nor U6837 (N_6837,N_6269,N_6258);
nor U6838 (N_6838,N_6267,N_6328);
or U6839 (N_6839,N_6268,N_6090);
nor U6840 (N_6840,N_6371,N_6030);
nor U6841 (N_6841,N_6169,N_6343);
and U6842 (N_6842,N_6465,N_6079);
nand U6843 (N_6843,N_6263,N_6278);
xnor U6844 (N_6844,N_6373,N_6394);
or U6845 (N_6845,N_6133,N_6386);
nor U6846 (N_6846,N_6403,N_6091);
nand U6847 (N_6847,N_6147,N_6260);
nor U6848 (N_6848,N_6277,N_6236);
nor U6849 (N_6849,N_6162,N_6233);
nand U6850 (N_6850,N_6039,N_6022);
and U6851 (N_6851,N_6425,N_6177);
and U6852 (N_6852,N_6280,N_6471);
nand U6853 (N_6853,N_6397,N_6167);
xnor U6854 (N_6854,N_6462,N_6248);
or U6855 (N_6855,N_6352,N_6495);
or U6856 (N_6856,N_6280,N_6053);
and U6857 (N_6857,N_6309,N_6142);
and U6858 (N_6858,N_6001,N_6222);
and U6859 (N_6859,N_6212,N_6400);
xor U6860 (N_6860,N_6008,N_6489);
or U6861 (N_6861,N_6109,N_6280);
xor U6862 (N_6862,N_6408,N_6386);
and U6863 (N_6863,N_6034,N_6047);
and U6864 (N_6864,N_6136,N_6406);
nand U6865 (N_6865,N_6120,N_6400);
xnor U6866 (N_6866,N_6267,N_6075);
nor U6867 (N_6867,N_6210,N_6098);
nor U6868 (N_6868,N_6204,N_6355);
nand U6869 (N_6869,N_6279,N_6439);
nor U6870 (N_6870,N_6025,N_6376);
nand U6871 (N_6871,N_6423,N_6369);
and U6872 (N_6872,N_6067,N_6326);
xnor U6873 (N_6873,N_6220,N_6241);
and U6874 (N_6874,N_6431,N_6169);
nor U6875 (N_6875,N_6445,N_6393);
xor U6876 (N_6876,N_6403,N_6098);
xor U6877 (N_6877,N_6094,N_6178);
nand U6878 (N_6878,N_6019,N_6187);
nand U6879 (N_6879,N_6204,N_6142);
nor U6880 (N_6880,N_6004,N_6301);
and U6881 (N_6881,N_6076,N_6461);
nand U6882 (N_6882,N_6347,N_6453);
or U6883 (N_6883,N_6392,N_6356);
nor U6884 (N_6884,N_6145,N_6305);
nand U6885 (N_6885,N_6222,N_6154);
or U6886 (N_6886,N_6288,N_6326);
nand U6887 (N_6887,N_6080,N_6044);
nand U6888 (N_6888,N_6465,N_6444);
and U6889 (N_6889,N_6200,N_6235);
or U6890 (N_6890,N_6307,N_6219);
or U6891 (N_6891,N_6249,N_6389);
or U6892 (N_6892,N_6415,N_6331);
or U6893 (N_6893,N_6194,N_6388);
and U6894 (N_6894,N_6471,N_6248);
nor U6895 (N_6895,N_6068,N_6496);
xor U6896 (N_6896,N_6393,N_6131);
nand U6897 (N_6897,N_6266,N_6154);
or U6898 (N_6898,N_6473,N_6397);
nand U6899 (N_6899,N_6388,N_6152);
or U6900 (N_6900,N_6442,N_6425);
nand U6901 (N_6901,N_6255,N_6061);
xor U6902 (N_6902,N_6173,N_6484);
nor U6903 (N_6903,N_6344,N_6305);
and U6904 (N_6904,N_6105,N_6143);
xor U6905 (N_6905,N_6205,N_6320);
nand U6906 (N_6906,N_6018,N_6258);
or U6907 (N_6907,N_6070,N_6363);
and U6908 (N_6908,N_6396,N_6286);
and U6909 (N_6909,N_6157,N_6215);
nand U6910 (N_6910,N_6034,N_6177);
nand U6911 (N_6911,N_6071,N_6094);
and U6912 (N_6912,N_6032,N_6221);
or U6913 (N_6913,N_6476,N_6137);
nor U6914 (N_6914,N_6043,N_6364);
nor U6915 (N_6915,N_6140,N_6033);
or U6916 (N_6916,N_6121,N_6201);
and U6917 (N_6917,N_6015,N_6339);
nand U6918 (N_6918,N_6390,N_6186);
nand U6919 (N_6919,N_6042,N_6262);
xnor U6920 (N_6920,N_6169,N_6290);
or U6921 (N_6921,N_6167,N_6195);
xnor U6922 (N_6922,N_6250,N_6272);
nand U6923 (N_6923,N_6277,N_6262);
and U6924 (N_6924,N_6264,N_6258);
or U6925 (N_6925,N_6384,N_6123);
nand U6926 (N_6926,N_6189,N_6255);
nor U6927 (N_6927,N_6379,N_6127);
xnor U6928 (N_6928,N_6026,N_6268);
nand U6929 (N_6929,N_6475,N_6027);
xnor U6930 (N_6930,N_6488,N_6053);
xnor U6931 (N_6931,N_6152,N_6471);
and U6932 (N_6932,N_6042,N_6361);
xnor U6933 (N_6933,N_6347,N_6442);
nand U6934 (N_6934,N_6250,N_6233);
nand U6935 (N_6935,N_6067,N_6458);
nand U6936 (N_6936,N_6482,N_6137);
nand U6937 (N_6937,N_6390,N_6054);
xnor U6938 (N_6938,N_6458,N_6422);
and U6939 (N_6939,N_6029,N_6489);
nand U6940 (N_6940,N_6489,N_6387);
or U6941 (N_6941,N_6310,N_6281);
xnor U6942 (N_6942,N_6307,N_6254);
nor U6943 (N_6943,N_6104,N_6154);
nand U6944 (N_6944,N_6124,N_6106);
nor U6945 (N_6945,N_6375,N_6211);
and U6946 (N_6946,N_6137,N_6033);
or U6947 (N_6947,N_6011,N_6366);
xnor U6948 (N_6948,N_6160,N_6306);
nor U6949 (N_6949,N_6064,N_6335);
nor U6950 (N_6950,N_6326,N_6460);
nor U6951 (N_6951,N_6210,N_6039);
and U6952 (N_6952,N_6268,N_6235);
or U6953 (N_6953,N_6042,N_6348);
xor U6954 (N_6954,N_6186,N_6449);
and U6955 (N_6955,N_6369,N_6060);
or U6956 (N_6956,N_6027,N_6497);
and U6957 (N_6957,N_6011,N_6433);
xor U6958 (N_6958,N_6142,N_6490);
or U6959 (N_6959,N_6366,N_6122);
xor U6960 (N_6960,N_6498,N_6181);
xnor U6961 (N_6961,N_6179,N_6209);
or U6962 (N_6962,N_6087,N_6230);
and U6963 (N_6963,N_6297,N_6065);
or U6964 (N_6964,N_6082,N_6361);
or U6965 (N_6965,N_6294,N_6199);
nand U6966 (N_6966,N_6112,N_6226);
nor U6967 (N_6967,N_6009,N_6496);
and U6968 (N_6968,N_6433,N_6025);
or U6969 (N_6969,N_6187,N_6274);
and U6970 (N_6970,N_6367,N_6458);
xor U6971 (N_6971,N_6044,N_6406);
xnor U6972 (N_6972,N_6152,N_6108);
or U6973 (N_6973,N_6367,N_6318);
nand U6974 (N_6974,N_6284,N_6107);
nor U6975 (N_6975,N_6010,N_6064);
and U6976 (N_6976,N_6493,N_6197);
or U6977 (N_6977,N_6080,N_6083);
nand U6978 (N_6978,N_6149,N_6354);
nor U6979 (N_6979,N_6042,N_6376);
nor U6980 (N_6980,N_6165,N_6110);
or U6981 (N_6981,N_6105,N_6216);
nor U6982 (N_6982,N_6162,N_6371);
nand U6983 (N_6983,N_6399,N_6473);
or U6984 (N_6984,N_6297,N_6102);
nor U6985 (N_6985,N_6108,N_6042);
or U6986 (N_6986,N_6346,N_6200);
and U6987 (N_6987,N_6043,N_6083);
nor U6988 (N_6988,N_6305,N_6490);
xor U6989 (N_6989,N_6104,N_6092);
xor U6990 (N_6990,N_6213,N_6365);
nand U6991 (N_6991,N_6093,N_6222);
or U6992 (N_6992,N_6078,N_6396);
xnor U6993 (N_6993,N_6116,N_6198);
nor U6994 (N_6994,N_6305,N_6409);
nor U6995 (N_6995,N_6287,N_6006);
or U6996 (N_6996,N_6030,N_6452);
and U6997 (N_6997,N_6427,N_6448);
and U6998 (N_6998,N_6249,N_6286);
nand U6999 (N_6999,N_6225,N_6125);
or U7000 (N_7000,N_6875,N_6751);
nor U7001 (N_7001,N_6781,N_6628);
or U7002 (N_7002,N_6704,N_6698);
xor U7003 (N_7003,N_6627,N_6907);
xor U7004 (N_7004,N_6942,N_6932);
or U7005 (N_7005,N_6763,N_6821);
xnor U7006 (N_7006,N_6707,N_6922);
or U7007 (N_7007,N_6984,N_6762);
and U7008 (N_7008,N_6888,N_6576);
nand U7009 (N_7009,N_6971,N_6752);
xnor U7010 (N_7010,N_6645,N_6826);
nand U7011 (N_7011,N_6766,N_6824);
and U7012 (N_7012,N_6609,N_6564);
nor U7013 (N_7013,N_6549,N_6745);
or U7014 (N_7014,N_6846,N_6709);
nor U7015 (N_7015,N_6644,N_6914);
or U7016 (N_7016,N_6519,N_6533);
nor U7017 (N_7017,N_6798,N_6748);
or U7018 (N_7018,N_6694,N_6795);
and U7019 (N_7019,N_6596,N_6518);
xnor U7020 (N_7020,N_6685,N_6960);
nor U7021 (N_7021,N_6854,N_6646);
and U7022 (N_7022,N_6584,N_6877);
or U7023 (N_7023,N_6775,N_6822);
or U7024 (N_7024,N_6892,N_6570);
or U7025 (N_7025,N_6970,N_6966);
or U7026 (N_7026,N_6565,N_6962);
xnor U7027 (N_7027,N_6989,N_6607);
xnor U7028 (N_7028,N_6626,N_6809);
nor U7029 (N_7029,N_6625,N_6567);
and U7030 (N_7030,N_6829,N_6827);
and U7031 (N_7031,N_6613,N_6948);
or U7032 (N_7032,N_6897,N_6818);
xnor U7033 (N_7033,N_6552,N_6718);
nor U7034 (N_7034,N_6623,N_6904);
or U7035 (N_7035,N_6872,N_6956);
nor U7036 (N_7036,N_6712,N_6783);
nand U7037 (N_7037,N_6873,N_6749);
or U7038 (N_7038,N_6771,N_6935);
or U7039 (N_7039,N_6589,N_6503);
xnor U7040 (N_7040,N_6890,N_6747);
or U7041 (N_7041,N_6514,N_6999);
or U7042 (N_7042,N_6760,N_6909);
or U7043 (N_7043,N_6993,N_6791);
nor U7044 (N_7044,N_6705,N_6719);
nand U7045 (N_7045,N_6841,N_6906);
nor U7046 (N_7046,N_6986,N_6515);
nand U7047 (N_7047,N_6582,N_6583);
nand U7048 (N_7048,N_6692,N_6544);
or U7049 (N_7049,N_6635,N_6615);
nand U7050 (N_7050,N_6742,N_6688);
nand U7051 (N_7051,N_6711,N_6592);
or U7052 (N_7052,N_6979,N_6900);
nor U7053 (N_7053,N_6658,N_6558);
nor U7054 (N_7054,N_6838,N_6949);
nor U7055 (N_7055,N_6996,N_6575);
and U7056 (N_7056,N_6980,N_6659);
and U7057 (N_7057,N_6974,N_6850);
nor U7058 (N_7058,N_6835,N_6786);
xor U7059 (N_7059,N_6664,N_6880);
and U7060 (N_7060,N_6637,N_6700);
and U7061 (N_7061,N_6563,N_6703);
xnor U7062 (N_7062,N_6797,N_6667);
or U7063 (N_7063,N_6785,N_6852);
xor U7064 (N_7064,N_6780,N_6530);
or U7065 (N_7065,N_6662,N_6656);
nor U7066 (N_7066,N_6642,N_6756);
xor U7067 (N_7067,N_6774,N_6605);
or U7068 (N_7068,N_6764,N_6950);
nor U7069 (N_7069,N_6777,N_6967);
nor U7070 (N_7070,N_6573,N_6758);
nand U7071 (N_7071,N_6863,N_6744);
or U7072 (N_7072,N_6677,N_6945);
xnor U7073 (N_7073,N_6968,N_6540);
xnor U7074 (N_7074,N_6679,N_6905);
or U7075 (N_7075,N_6696,N_6733);
nand U7076 (N_7076,N_6524,N_6663);
nand U7077 (N_7077,N_6923,N_6572);
nand U7078 (N_7078,N_6893,N_6640);
nor U7079 (N_7079,N_6591,N_6955);
xnor U7080 (N_7080,N_6988,N_6917);
or U7081 (N_7081,N_6976,N_6690);
nor U7082 (N_7082,N_6725,N_6604);
xor U7083 (N_7083,N_6687,N_6657);
nor U7084 (N_7084,N_6713,N_6648);
nand U7085 (N_7085,N_6750,N_6736);
nor U7086 (N_7086,N_6871,N_6896);
nand U7087 (N_7087,N_6804,N_6536);
xor U7088 (N_7088,N_6867,N_6855);
and U7089 (N_7089,N_6587,N_6969);
xnor U7090 (N_7090,N_6823,N_6860);
or U7091 (N_7091,N_6545,N_6702);
nor U7092 (N_7092,N_6884,N_6921);
or U7093 (N_7093,N_6620,N_6507);
nand U7094 (N_7094,N_6808,N_6669);
xnor U7095 (N_7095,N_6874,N_6913);
nor U7096 (N_7096,N_6761,N_6706);
nor U7097 (N_7097,N_6714,N_6856);
nand U7098 (N_7098,N_6882,N_6803);
nand U7099 (N_7099,N_6812,N_6738);
nor U7100 (N_7100,N_6721,N_6728);
and U7101 (N_7101,N_6580,N_6535);
xor U7102 (N_7102,N_6840,N_6528);
nor U7103 (N_7103,N_6831,N_6858);
xnor U7104 (N_7104,N_6502,N_6542);
and U7105 (N_7105,N_6836,N_6819);
xnor U7106 (N_7106,N_6772,N_6963);
nor U7107 (N_7107,N_6961,N_6708);
nor U7108 (N_7108,N_6666,N_6546);
xor U7109 (N_7109,N_6622,N_6633);
xnor U7110 (N_7110,N_6717,N_6992);
nand U7111 (N_7111,N_6911,N_6739);
or U7112 (N_7112,N_6610,N_6853);
or U7113 (N_7113,N_6652,N_6887);
nor U7114 (N_7114,N_6834,N_6539);
or U7115 (N_7115,N_6952,N_6522);
or U7116 (N_7116,N_6726,N_6765);
nor U7117 (N_7117,N_6941,N_6957);
and U7118 (N_7118,N_6683,N_6516);
or U7119 (N_7119,N_6878,N_6559);
nand U7120 (N_7120,N_6869,N_6767);
or U7121 (N_7121,N_6670,N_6531);
xnor U7122 (N_7122,N_6740,N_6947);
nand U7123 (N_7123,N_6870,N_6994);
xor U7124 (N_7124,N_6953,N_6543);
nand U7125 (N_7125,N_6634,N_6936);
and U7126 (N_7126,N_6534,N_6934);
or U7127 (N_7127,N_6825,N_6943);
nor U7128 (N_7128,N_6901,N_6828);
nor U7129 (N_7129,N_6569,N_6770);
xor U7130 (N_7130,N_6830,N_6886);
nand U7131 (N_7131,N_6987,N_6554);
nand U7132 (N_7132,N_6844,N_6602);
nor U7133 (N_7133,N_6513,N_6654);
and U7134 (N_7134,N_6930,N_6788);
xnor U7135 (N_7135,N_6595,N_6639);
nand U7136 (N_7136,N_6561,N_6735);
nand U7137 (N_7137,N_6729,N_6548);
and U7138 (N_7138,N_6837,N_6864);
and U7139 (N_7139,N_6940,N_6997);
nand U7140 (N_7140,N_6665,N_6682);
nor U7141 (N_7141,N_6865,N_6802);
and U7142 (N_7142,N_6693,N_6792);
xor U7143 (N_7143,N_6578,N_6972);
nand U7144 (N_7144,N_6510,N_6671);
xnor U7145 (N_7145,N_6814,N_6617);
or U7146 (N_7146,N_6927,N_6861);
and U7147 (N_7147,N_6807,N_6678);
xor U7148 (N_7148,N_6556,N_6796);
nand U7149 (N_7149,N_6898,N_6538);
nand U7150 (N_7150,N_6924,N_6789);
and U7151 (N_7151,N_6506,N_6649);
or U7152 (N_7152,N_6560,N_6737);
nor U7153 (N_7153,N_6551,N_6894);
nand U7154 (N_7154,N_6520,N_6632);
nand U7155 (N_7155,N_6574,N_6817);
or U7156 (N_7156,N_6883,N_6866);
and U7157 (N_7157,N_6973,N_6790);
xnor U7158 (N_7158,N_6910,N_6879);
nor U7159 (N_7159,N_6720,N_6915);
nand U7160 (N_7160,N_6689,N_6621);
xor U7161 (N_7161,N_6975,N_6612);
or U7162 (N_7162,N_6673,N_6650);
xnor U7163 (N_7163,N_6608,N_6724);
or U7164 (N_7164,N_6753,N_6815);
xor U7165 (N_7165,N_6833,N_6991);
nor U7166 (N_7166,N_6512,N_6523);
nand U7167 (N_7167,N_6810,N_6782);
xnor U7168 (N_7168,N_6964,N_6908);
nand U7169 (N_7169,N_6787,N_6876);
and U7170 (N_7170,N_6527,N_6759);
xor U7171 (N_7171,N_6746,N_6990);
nand U7172 (N_7172,N_6843,N_6547);
or U7173 (N_7173,N_6571,N_6902);
and U7174 (N_7174,N_6638,N_6614);
or U7175 (N_7175,N_6647,N_6616);
nand U7176 (N_7176,N_6641,N_6557);
xor U7177 (N_7177,N_6743,N_6768);
nand U7178 (N_7178,N_6918,N_6985);
nor U7179 (N_7179,N_6727,N_6937);
and U7180 (N_7180,N_6839,N_6889);
nor U7181 (N_7181,N_6920,N_6755);
nand U7182 (N_7182,N_6773,N_6508);
and U7183 (N_7183,N_6857,N_6568);
and U7184 (N_7184,N_6845,N_6715);
and U7185 (N_7185,N_6811,N_6723);
or U7186 (N_7186,N_6862,N_6562);
nand U7187 (N_7187,N_6699,N_6581);
and U7188 (N_7188,N_6599,N_6800);
or U7189 (N_7189,N_6776,N_6939);
nor U7190 (N_7190,N_6899,N_6660);
or U7191 (N_7191,N_6611,N_6805);
nand U7192 (N_7192,N_6550,N_6686);
and U7193 (N_7193,N_6944,N_6600);
xnor U7194 (N_7194,N_6500,N_6801);
and U7195 (N_7195,N_6849,N_6794);
and U7196 (N_7196,N_6653,N_6912);
nor U7197 (N_7197,N_6885,N_6606);
nand U7198 (N_7198,N_6594,N_6517);
nand U7199 (N_7199,N_6741,N_6806);
nor U7200 (N_7200,N_6691,N_6954);
nor U7201 (N_7201,N_6981,N_6619);
or U7202 (N_7202,N_6566,N_6925);
nand U7203 (N_7203,N_6778,N_6537);
or U7204 (N_7204,N_6842,N_6784);
and U7205 (N_7205,N_6680,N_6672);
nand U7206 (N_7206,N_6813,N_6848);
and U7207 (N_7207,N_6891,N_6732);
xor U7208 (N_7208,N_6668,N_6509);
nor U7209 (N_7209,N_6946,N_6730);
nand U7210 (N_7210,N_6529,N_6504);
nand U7211 (N_7211,N_6716,N_6995);
or U7212 (N_7212,N_6851,N_6701);
nand U7213 (N_7213,N_6521,N_6816);
xnor U7214 (N_7214,N_6590,N_6983);
nand U7215 (N_7215,N_6919,N_6881);
xor U7216 (N_7216,N_6618,N_6926);
or U7217 (N_7217,N_6631,N_6624);
and U7218 (N_7218,N_6933,N_6722);
nand U7219 (N_7219,N_6585,N_6916);
and U7220 (N_7220,N_6511,N_6799);
nor U7221 (N_7221,N_6977,N_6579);
and U7222 (N_7222,N_6998,N_6526);
or U7223 (N_7223,N_6674,N_6779);
xor U7224 (N_7224,N_6501,N_6958);
nand U7225 (N_7225,N_6731,N_6929);
or U7226 (N_7226,N_6675,N_6868);
and U7227 (N_7227,N_6697,N_6629);
nor U7228 (N_7228,N_6793,N_6553);
nor U7229 (N_7229,N_6959,N_6577);
nand U7230 (N_7230,N_6541,N_6661);
and U7231 (N_7231,N_6903,N_6655);
xor U7232 (N_7232,N_6982,N_6593);
or U7233 (N_7233,N_6710,N_6951);
nor U7234 (N_7234,N_6586,N_6603);
and U7235 (N_7235,N_6978,N_6681);
xnor U7236 (N_7236,N_6555,N_6630);
nor U7237 (N_7237,N_6769,N_6601);
nand U7238 (N_7238,N_6820,N_6643);
and U7239 (N_7239,N_6859,N_6588);
and U7240 (N_7240,N_6532,N_6931);
and U7241 (N_7241,N_6754,N_6598);
and U7242 (N_7242,N_6676,N_6847);
and U7243 (N_7243,N_6757,N_6651);
or U7244 (N_7244,N_6734,N_6938);
xnor U7245 (N_7245,N_6636,N_6965);
or U7246 (N_7246,N_6928,N_6597);
nand U7247 (N_7247,N_6832,N_6695);
nand U7248 (N_7248,N_6684,N_6895);
and U7249 (N_7249,N_6505,N_6525);
nor U7250 (N_7250,N_6786,N_6526);
nand U7251 (N_7251,N_6743,N_6584);
nor U7252 (N_7252,N_6907,N_6586);
nand U7253 (N_7253,N_6797,N_6881);
nand U7254 (N_7254,N_6565,N_6875);
nor U7255 (N_7255,N_6889,N_6992);
nand U7256 (N_7256,N_6607,N_6880);
nand U7257 (N_7257,N_6890,N_6741);
and U7258 (N_7258,N_6637,N_6555);
and U7259 (N_7259,N_6521,N_6598);
or U7260 (N_7260,N_6537,N_6840);
or U7261 (N_7261,N_6806,N_6548);
and U7262 (N_7262,N_6553,N_6782);
or U7263 (N_7263,N_6624,N_6939);
xnor U7264 (N_7264,N_6618,N_6722);
and U7265 (N_7265,N_6533,N_6776);
nand U7266 (N_7266,N_6504,N_6998);
nand U7267 (N_7267,N_6537,N_6598);
nand U7268 (N_7268,N_6976,N_6630);
or U7269 (N_7269,N_6596,N_6912);
nor U7270 (N_7270,N_6823,N_6648);
or U7271 (N_7271,N_6889,N_6735);
or U7272 (N_7272,N_6899,N_6523);
and U7273 (N_7273,N_6795,N_6984);
nand U7274 (N_7274,N_6792,N_6914);
xor U7275 (N_7275,N_6618,N_6780);
nand U7276 (N_7276,N_6879,N_6638);
nand U7277 (N_7277,N_6759,N_6581);
nand U7278 (N_7278,N_6654,N_6665);
and U7279 (N_7279,N_6665,N_6500);
or U7280 (N_7280,N_6519,N_6862);
xnor U7281 (N_7281,N_6997,N_6980);
nand U7282 (N_7282,N_6824,N_6624);
nand U7283 (N_7283,N_6737,N_6779);
nand U7284 (N_7284,N_6582,N_6757);
or U7285 (N_7285,N_6606,N_6869);
and U7286 (N_7286,N_6584,N_6508);
nand U7287 (N_7287,N_6891,N_6865);
or U7288 (N_7288,N_6558,N_6952);
nor U7289 (N_7289,N_6721,N_6772);
nand U7290 (N_7290,N_6615,N_6903);
or U7291 (N_7291,N_6890,N_6816);
or U7292 (N_7292,N_6776,N_6541);
or U7293 (N_7293,N_6840,N_6696);
nand U7294 (N_7294,N_6638,N_6954);
xnor U7295 (N_7295,N_6574,N_6924);
and U7296 (N_7296,N_6909,N_6574);
and U7297 (N_7297,N_6655,N_6953);
xnor U7298 (N_7298,N_6801,N_6638);
or U7299 (N_7299,N_6804,N_6761);
nand U7300 (N_7300,N_6723,N_6591);
nand U7301 (N_7301,N_6694,N_6628);
or U7302 (N_7302,N_6644,N_6827);
nor U7303 (N_7303,N_6572,N_6938);
or U7304 (N_7304,N_6519,N_6730);
xor U7305 (N_7305,N_6627,N_6898);
nor U7306 (N_7306,N_6909,N_6542);
nor U7307 (N_7307,N_6602,N_6583);
or U7308 (N_7308,N_6622,N_6508);
xnor U7309 (N_7309,N_6642,N_6958);
or U7310 (N_7310,N_6731,N_6590);
and U7311 (N_7311,N_6627,N_6902);
and U7312 (N_7312,N_6611,N_6845);
nor U7313 (N_7313,N_6504,N_6939);
or U7314 (N_7314,N_6949,N_6880);
or U7315 (N_7315,N_6873,N_6571);
nand U7316 (N_7316,N_6579,N_6870);
or U7317 (N_7317,N_6756,N_6879);
nand U7318 (N_7318,N_6973,N_6778);
or U7319 (N_7319,N_6824,N_6933);
and U7320 (N_7320,N_6729,N_6950);
nand U7321 (N_7321,N_6543,N_6732);
xor U7322 (N_7322,N_6741,N_6647);
or U7323 (N_7323,N_6720,N_6704);
nor U7324 (N_7324,N_6990,N_6888);
xnor U7325 (N_7325,N_6690,N_6956);
nor U7326 (N_7326,N_6526,N_6516);
xnor U7327 (N_7327,N_6961,N_6542);
or U7328 (N_7328,N_6794,N_6853);
and U7329 (N_7329,N_6968,N_6521);
or U7330 (N_7330,N_6722,N_6855);
nor U7331 (N_7331,N_6753,N_6893);
nor U7332 (N_7332,N_6766,N_6848);
xnor U7333 (N_7333,N_6694,N_6615);
xor U7334 (N_7334,N_6714,N_6523);
nor U7335 (N_7335,N_6549,N_6882);
and U7336 (N_7336,N_6511,N_6796);
or U7337 (N_7337,N_6646,N_6778);
and U7338 (N_7338,N_6576,N_6878);
or U7339 (N_7339,N_6635,N_6665);
xnor U7340 (N_7340,N_6875,N_6738);
xor U7341 (N_7341,N_6762,N_6638);
nand U7342 (N_7342,N_6858,N_6510);
or U7343 (N_7343,N_6552,N_6689);
xnor U7344 (N_7344,N_6596,N_6987);
and U7345 (N_7345,N_6634,N_6965);
or U7346 (N_7346,N_6869,N_6834);
xor U7347 (N_7347,N_6721,N_6848);
and U7348 (N_7348,N_6554,N_6652);
nor U7349 (N_7349,N_6823,N_6830);
nor U7350 (N_7350,N_6774,N_6586);
or U7351 (N_7351,N_6659,N_6581);
and U7352 (N_7352,N_6837,N_6977);
xnor U7353 (N_7353,N_6584,N_6923);
nand U7354 (N_7354,N_6931,N_6616);
or U7355 (N_7355,N_6856,N_6787);
nand U7356 (N_7356,N_6546,N_6928);
xnor U7357 (N_7357,N_6537,N_6508);
xor U7358 (N_7358,N_6665,N_6577);
and U7359 (N_7359,N_6680,N_6512);
nand U7360 (N_7360,N_6511,N_6828);
or U7361 (N_7361,N_6659,N_6564);
nand U7362 (N_7362,N_6870,N_6526);
or U7363 (N_7363,N_6746,N_6679);
nand U7364 (N_7364,N_6521,N_6583);
or U7365 (N_7365,N_6762,N_6847);
and U7366 (N_7366,N_6919,N_6846);
or U7367 (N_7367,N_6681,N_6799);
nor U7368 (N_7368,N_6951,N_6665);
xor U7369 (N_7369,N_6725,N_6692);
xor U7370 (N_7370,N_6997,N_6877);
xnor U7371 (N_7371,N_6587,N_6614);
nor U7372 (N_7372,N_6963,N_6998);
xnor U7373 (N_7373,N_6605,N_6780);
nand U7374 (N_7374,N_6788,N_6892);
nor U7375 (N_7375,N_6696,N_6940);
and U7376 (N_7376,N_6890,N_6596);
and U7377 (N_7377,N_6623,N_6894);
nand U7378 (N_7378,N_6553,N_6891);
and U7379 (N_7379,N_6833,N_6867);
nand U7380 (N_7380,N_6610,N_6947);
and U7381 (N_7381,N_6701,N_6628);
nor U7382 (N_7382,N_6600,N_6771);
or U7383 (N_7383,N_6840,N_6657);
and U7384 (N_7384,N_6839,N_6763);
nand U7385 (N_7385,N_6567,N_6896);
nor U7386 (N_7386,N_6972,N_6812);
and U7387 (N_7387,N_6933,N_6672);
or U7388 (N_7388,N_6705,N_6521);
or U7389 (N_7389,N_6785,N_6544);
nor U7390 (N_7390,N_6622,N_6578);
and U7391 (N_7391,N_6911,N_6741);
xnor U7392 (N_7392,N_6552,N_6784);
or U7393 (N_7393,N_6797,N_6744);
or U7394 (N_7394,N_6970,N_6971);
nand U7395 (N_7395,N_6888,N_6769);
and U7396 (N_7396,N_6562,N_6949);
nor U7397 (N_7397,N_6575,N_6808);
nand U7398 (N_7398,N_6651,N_6828);
nor U7399 (N_7399,N_6738,N_6937);
nand U7400 (N_7400,N_6514,N_6802);
xnor U7401 (N_7401,N_6505,N_6641);
nand U7402 (N_7402,N_6588,N_6884);
nor U7403 (N_7403,N_6951,N_6869);
nor U7404 (N_7404,N_6942,N_6661);
and U7405 (N_7405,N_6546,N_6949);
nand U7406 (N_7406,N_6997,N_6938);
nor U7407 (N_7407,N_6973,N_6974);
nor U7408 (N_7408,N_6819,N_6726);
and U7409 (N_7409,N_6517,N_6780);
or U7410 (N_7410,N_6872,N_6838);
nor U7411 (N_7411,N_6974,N_6569);
nand U7412 (N_7412,N_6667,N_6733);
and U7413 (N_7413,N_6754,N_6702);
nor U7414 (N_7414,N_6902,N_6638);
and U7415 (N_7415,N_6849,N_6696);
nand U7416 (N_7416,N_6931,N_6614);
and U7417 (N_7417,N_6643,N_6848);
xor U7418 (N_7418,N_6769,N_6537);
and U7419 (N_7419,N_6749,N_6783);
and U7420 (N_7420,N_6909,N_6658);
nor U7421 (N_7421,N_6620,N_6993);
xor U7422 (N_7422,N_6632,N_6990);
xor U7423 (N_7423,N_6906,N_6818);
xnor U7424 (N_7424,N_6882,N_6606);
or U7425 (N_7425,N_6750,N_6682);
xor U7426 (N_7426,N_6511,N_6588);
nand U7427 (N_7427,N_6925,N_6733);
nor U7428 (N_7428,N_6517,N_6766);
nand U7429 (N_7429,N_6764,N_6679);
or U7430 (N_7430,N_6664,N_6792);
or U7431 (N_7431,N_6749,N_6521);
and U7432 (N_7432,N_6625,N_6767);
and U7433 (N_7433,N_6892,N_6730);
nor U7434 (N_7434,N_6821,N_6650);
and U7435 (N_7435,N_6844,N_6731);
xor U7436 (N_7436,N_6567,N_6604);
nand U7437 (N_7437,N_6529,N_6896);
and U7438 (N_7438,N_6966,N_6558);
or U7439 (N_7439,N_6831,N_6747);
or U7440 (N_7440,N_6702,N_6597);
nor U7441 (N_7441,N_6537,N_6674);
nand U7442 (N_7442,N_6984,N_6662);
nor U7443 (N_7443,N_6669,N_6728);
nand U7444 (N_7444,N_6574,N_6694);
and U7445 (N_7445,N_6841,N_6677);
and U7446 (N_7446,N_6954,N_6537);
xor U7447 (N_7447,N_6709,N_6905);
nand U7448 (N_7448,N_6760,N_6596);
nand U7449 (N_7449,N_6503,N_6528);
nand U7450 (N_7450,N_6673,N_6656);
xor U7451 (N_7451,N_6526,N_6669);
nand U7452 (N_7452,N_6933,N_6811);
nor U7453 (N_7453,N_6742,N_6845);
nor U7454 (N_7454,N_6852,N_6730);
nand U7455 (N_7455,N_6543,N_6795);
and U7456 (N_7456,N_6523,N_6974);
and U7457 (N_7457,N_6548,N_6892);
and U7458 (N_7458,N_6624,N_6889);
nand U7459 (N_7459,N_6736,N_6839);
xor U7460 (N_7460,N_6571,N_6806);
nor U7461 (N_7461,N_6627,N_6600);
xnor U7462 (N_7462,N_6946,N_6505);
and U7463 (N_7463,N_6775,N_6507);
nand U7464 (N_7464,N_6623,N_6674);
or U7465 (N_7465,N_6544,N_6516);
or U7466 (N_7466,N_6936,N_6815);
and U7467 (N_7467,N_6519,N_6563);
nand U7468 (N_7468,N_6831,N_6925);
and U7469 (N_7469,N_6658,N_6565);
and U7470 (N_7470,N_6827,N_6588);
xnor U7471 (N_7471,N_6701,N_6922);
and U7472 (N_7472,N_6929,N_6727);
xnor U7473 (N_7473,N_6656,N_6700);
nand U7474 (N_7474,N_6986,N_6507);
or U7475 (N_7475,N_6884,N_6968);
nor U7476 (N_7476,N_6837,N_6735);
nor U7477 (N_7477,N_6515,N_6604);
xor U7478 (N_7478,N_6698,N_6753);
xnor U7479 (N_7479,N_6698,N_6627);
xor U7480 (N_7480,N_6911,N_6705);
or U7481 (N_7481,N_6663,N_6570);
xnor U7482 (N_7482,N_6879,N_6880);
nor U7483 (N_7483,N_6833,N_6967);
xnor U7484 (N_7484,N_6576,N_6996);
nor U7485 (N_7485,N_6910,N_6596);
and U7486 (N_7486,N_6531,N_6701);
nand U7487 (N_7487,N_6501,N_6760);
nor U7488 (N_7488,N_6838,N_6889);
nor U7489 (N_7489,N_6902,N_6883);
and U7490 (N_7490,N_6543,N_6725);
xnor U7491 (N_7491,N_6915,N_6714);
nand U7492 (N_7492,N_6620,N_6919);
xor U7493 (N_7493,N_6655,N_6927);
xor U7494 (N_7494,N_6841,N_6562);
nor U7495 (N_7495,N_6742,N_6662);
and U7496 (N_7496,N_6713,N_6798);
xor U7497 (N_7497,N_6971,N_6709);
nor U7498 (N_7498,N_6887,N_6739);
xnor U7499 (N_7499,N_6853,N_6688);
and U7500 (N_7500,N_7141,N_7210);
or U7501 (N_7501,N_7126,N_7058);
nand U7502 (N_7502,N_7226,N_7187);
xnor U7503 (N_7503,N_7160,N_7071);
or U7504 (N_7504,N_7108,N_7011);
nand U7505 (N_7505,N_7433,N_7315);
nand U7506 (N_7506,N_7239,N_7262);
nor U7507 (N_7507,N_7494,N_7134);
and U7508 (N_7508,N_7260,N_7478);
and U7509 (N_7509,N_7046,N_7458);
and U7510 (N_7510,N_7110,N_7174);
nand U7511 (N_7511,N_7432,N_7097);
nor U7512 (N_7512,N_7219,N_7124);
xor U7513 (N_7513,N_7419,N_7069);
nand U7514 (N_7514,N_7375,N_7183);
nand U7515 (N_7515,N_7332,N_7354);
nor U7516 (N_7516,N_7431,N_7122);
and U7517 (N_7517,N_7193,N_7257);
nor U7518 (N_7518,N_7161,N_7208);
xor U7519 (N_7519,N_7491,N_7218);
nor U7520 (N_7520,N_7337,N_7173);
nor U7521 (N_7521,N_7036,N_7255);
nand U7522 (N_7522,N_7280,N_7207);
nand U7523 (N_7523,N_7037,N_7310);
xor U7524 (N_7524,N_7103,N_7035);
or U7525 (N_7525,N_7383,N_7459);
nand U7526 (N_7526,N_7024,N_7231);
xor U7527 (N_7527,N_7001,N_7196);
nor U7528 (N_7528,N_7188,N_7087);
and U7529 (N_7529,N_7137,N_7059);
nor U7530 (N_7530,N_7055,N_7347);
xor U7531 (N_7531,N_7456,N_7406);
and U7532 (N_7532,N_7060,N_7291);
xor U7533 (N_7533,N_7129,N_7043);
nand U7534 (N_7534,N_7023,N_7083);
xor U7535 (N_7535,N_7009,N_7409);
xor U7536 (N_7536,N_7267,N_7412);
nand U7537 (N_7537,N_7440,N_7463);
nor U7538 (N_7538,N_7088,N_7364);
or U7539 (N_7539,N_7222,N_7002);
nand U7540 (N_7540,N_7057,N_7439);
and U7541 (N_7541,N_7109,N_7401);
xor U7542 (N_7542,N_7348,N_7446);
or U7543 (N_7543,N_7474,N_7086);
and U7544 (N_7544,N_7229,N_7042);
or U7545 (N_7545,N_7119,N_7167);
xor U7546 (N_7546,N_7212,N_7451);
xnor U7547 (N_7547,N_7471,N_7276);
and U7548 (N_7548,N_7013,N_7329);
nor U7549 (N_7549,N_7008,N_7151);
or U7550 (N_7550,N_7041,N_7068);
nand U7551 (N_7551,N_7465,N_7281);
xor U7552 (N_7552,N_7078,N_7470);
or U7553 (N_7553,N_7112,N_7007);
xor U7554 (N_7554,N_7472,N_7278);
nor U7555 (N_7555,N_7476,N_7095);
nand U7556 (N_7556,N_7085,N_7270);
or U7557 (N_7557,N_7405,N_7357);
nand U7558 (N_7558,N_7447,N_7289);
and U7559 (N_7559,N_7072,N_7436);
nor U7560 (N_7560,N_7148,N_7425);
nand U7561 (N_7561,N_7128,N_7185);
nand U7562 (N_7562,N_7344,N_7442);
nor U7563 (N_7563,N_7300,N_7441);
nand U7564 (N_7564,N_7101,N_7127);
xor U7565 (N_7565,N_7140,N_7396);
nor U7566 (N_7566,N_7313,N_7156);
nand U7567 (N_7567,N_7217,N_7341);
nand U7568 (N_7568,N_7482,N_7121);
nand U7569 (N_7569,N_7017,N_7469);
nor U7570 (N_7570,N_7150,N_7227);
xor U7571 (N_7571,N_7317,N_7498);
and U7572 (N_7572,N_7403,N_7374);
or U7573 (N_7573,N_7091,N_7273);
and U7574 (N_7574,N_7288,N_7154);
xnor U7575 (N_7575,N_7232,N_7152);
nor U7576 (N_7576,N_7343,N_7422);
nor U7577 (N_7577,N_7198,N_7445);
xnor U7578 (N_7578,N_7117,N_7307);
xnor U7579 (N_7579,N_7448,N_7319);
nand U7580 (N_7580,N_7455,N_7398);
nor U7581 (N_7581,N_7462,N_7336);
xor U7582 (N_7582,N_7428,N_7106);
or U7583 (N_7583,N_7022,N_7483);
nand U7584 (N_7584,N_7168,N_7430);
nor U7585 (N_7585,N_7388,N_7169);
nor U7586 (N_7586,N_7283,N_7053);
or U7587 (N_7587,N_7026,N_7203);
and U7588 (N_7588,N_7386,N_7242);
and U7589 (N_7589,N_7145,N_7179);
xnor U7590 (N_7590,N_7258,N_7484);
or U7591 (N_7591,N_7015,N_7486);
and U7592 (N_7592,N_7373,N_7468);
nand U7593 (N_7593,N_7186,N_7094);
xnor U7594 (N_7594,N_7067,N_7377);
and U7595 (N_7595,N_7118,N_7147);
or U7596 (N_7596,N_7382,N_7497);
and U7597 (N_7597,N_7453,N_7066);
xnor U7598 (N_7598,N_7261,N_7184);
nand U7599 (N_7599,N_7380,N_7163);
or U7600 (N_7600,N_7437,N_7178);
nand U7601 (N_7601,N_7292,N_7130);
nand U7602 (N_7602,N_7211,N_7221);
nor U7603 (N_7603,N_7166,N_7236);
nand U7604 (N_7604,N_7294,N_7414);
xor U7605 (N_7605,N_7296,N_7338);
and U7606 (N_7606,N_7321,N_7393);
nand U7607 (N_7607,N_7040,N_7423);
nor U7608 (N_7608,N_7157,N_7213);
or U7609 (N_7609,N_7075,N_7252);
nor U7610 (N_7610,N_7100,N_7215);
and U7611 (N_7611,N_7320,N_7492);
nand U7612 (N_7612,N_7133,N_7473);
or U7613 (N_7613,N_7352,N_7330);
or U7614 (N_7614,N_7084,N_7314);
or U7615 (N_7615,N_7480,N_7376);
and U7616 (N_7616,N_7065,N_7230);
xnor U7617 (N_7617,N_7390,N_7290);
nand U7618 (N_7618,N_7201,N_7367);
and U7619 (N_7619,N_7092,N_7302);
nand U7620 (N_7620,N_7254,N_7397);
and U7621 (N_7621,N_7062,N_7454);
or U7622 (N_7622,N_7420,N_7143);
nand U7623 (N_7623,N_7138,N_7131);
xnor U7624 (N_7624,N_7264,N_7499);
or U7625 (N_7625,N_7200,N_7256);
or U7626 (N_7626,N_7361,N_7146);
or U7627 (N_7627,N_7237,N_7204);
nor U7628 (N_7628,N_7263,N_7090);
or U7629 (N_7629,N_7172,N_7284);
nand U7630 (N_7630,N_7381,N_7391);
and U7631 (N_7631,N_7305,N_7177);
nand U7632 (N_7632,N_7113,N_7429);
nor U7633 (N_7633,N_7159,N_7030);
or U7634 (N_7634,N_7056,N_7410);
and U7635 (N_7635,N_7240,N_7489);
xnor U7636 (N_7636,N_7012,N_7387);
nor U7637 (N_7637,N_7358,N_7411);
nand U7638 (N_7638,N_7020,N_7250);
xnor U7639 (N_7639,N_7328,N_7404);
or U7640 (N_7640,N_7192,N_7351);
nand U7641 (N_7641,N_7334,N_7105);
xnor U7642 (N_7642,N_7050,N_7158);
and U7643 (N_7643,N_7327,N_7081);
xnor U7644 (N_7644,N_7228,N_7209);
or U7645 (N_7645,N_7238,N_7114);
nand U7646 (N_7646,N_7426,N_7182);
and U7647 (N_7647,N_7384,N_7438);
xnor U7648 (N_7648,N_7259,N_7049);
and U7649 (N_7649,N_7346,N_7413);
nand U7650 (N_7650,N_7076,N_7191);
and U7651 (N_7651,N_7444,N_7006);
or U7652 (N_7652,N_7467,N_7054);
and U7653 (N_7653,N_7171,N_7421);
nand U7654 (N_7654,N_7496,N_7312);
xor U7655 (N_7655,N_7039,N_7248);
and U7656 (N_7656,N_7490,N_7477);
nand U7657 (N_7657,N_7000,N_7111);
and U7658 (N_7658,N_7417,N_7326);
xor U7659 (N_7659,N_7019,N_7304);
and U7660 (N_7660,N_7450,N_7277);
or U7661 (N_7661,N_7457,N_7132);
xor U7662 (N_7662,N_7180,N_7322);
nor U7663 (N_7663,N_7268,N_7234);
xnor U7664 (N_7664,N_7416,N_7366);
nand U7665 (N_7665,N_7495,N_7355);
nand U7666 (N_7666,N_7034,N_7197);
nand U7667 (N_7667,N_7216,N_7339);
nor U7668 (N_7668,N_7360,N_7249);
nor U7669 (N_7669,N_7155,N_7335);
or U7670 (N_7670,N_7274,N_7125);
and U7671 (N_7671,N_7010,N_7162);
nand U7672 (N_7672,N_7074,N_7214);
nand U7673 (N_7673,N_7004,N_7402);
and U7674 (N_7674,N_7295,N_7029);
xor U7675 (N_7675,N_7123,N_7014);
and U7676 (N_7676,N_7120,N_7418);
or U7677 (N_7677,N_7139,N_7466);
nor U7678 (N_7678,N_7342,N_7176);
and U7679 (N_7679,N_7027,N_7251);
nor U7680 (N_7680,N_7485,N_7082);
and U7681 (N_7681,N_7362,N_7372);
nor U7682 (N_7682,N_7306,N_7356);
or U7683 (N_7683,N_7051,N_7311);
or U7684 (N_7684,N_7323,N_7205);
nand U7685 (N_7685,N_7224,N_7225);
nor U7686 (N_7686,N_7028,N_7247);
nor U7687 (N_7687,N_7149,N_7303);
and U7688 (N_7688,N_7135,N_7309);
nand U7689 (N_7689,N_7488,N_7044);
xnor U7690 (N_7690,N_7443,N_7297);
or U7691 (N_7691,N_7481,N_7153);
and U7692 (N_7692,N_7235,N_7385);
nor U7693 (N_7693,N_7025,N_7243);
nand U7694 (N_7694,N_7282,N_7116);
nand U7695 (N_7695,N_7245,N_7316);
nand U7696 (N_7696,N_7061,N_7093);
or U7697 (N_7697,N_7479,N_7223);
nor U7698 (N_7698,N_7233,N_7298);
nor U7699 (N_7699,N_7269,N_7005);
and U7700 (N_7700,N_7048,N_7031);
and U7701 (N_7701,N_7144,N_7102);
nand U7702 (N_7702,N_7340,N_7435);
xnor U7703 (N_7703,N_7331,N_7175);
xnor U7704 (N_7704,N_7368,N_7285);
xor U7705 (N_7705,N_7493,N_7370);
nand U7706 (N_7706,N_7038,N_7033);
xor U7707 (N_7707,N_7301,N_7080);
and U7708 (N_7708,N_7427,N_7275);
xor U7709 (N_7709,N_7392,N_7365);
xnor U7710 (N_7710,N_7202,N_7464);
and U7711 (N_7711,N_7206,N_7052);
or U7712 (N_7712,N_7181,N_7394);
and U7713 (N_7713,N_7308,N_7378);
xor U7714 (N_7714,N_7018,N_7333);
or U7715 (N_7715,N_7190,N_7244);
nand U7716 (N_7716,N_7099,N_7460);
or U7717 (N_7717,N_7064,N_7136);
and U7718 (N_7718,N_7089,N_7299);
xnor U7719 (N_7719,N_7359,N_7389);
xnor U7720 (N_7720,N_7271,N_7098);
xor U7721 (N_7721,N_7104,N_7079);
nand U7722 (N_7722,N_7142,N_7070);
or U7723 (N_7723,N_7003,N_7063);
xor U7724 (N_7724,N_7324,N_7318);
or U7725 (N_7725,N_7325,N_7369);
and U7726 (N_7726,N_7287,N_7241);
or U7727 (N_7727,N_7349,N_7415);
and U7728 (N_7728,N_7096,N_7253);
xor U7729 (N_7729,N_7353,N_7293);
xnor U7730 (N_7730,N_7272,N_7107);
or U7731 (N_7731,N_7461,N_7345);
and U7732 (N_7732,N_7189,N_7195);
nand U7733 (N_7733,N_7164,N_7266);
xor U7734 (N_7734,N_7194,N_7279);
nor U7735 (N_7735,N_7032,N_7363);
nor U7736 (N_7736,N_7408,N_7246);
nor U7737 (N_7737,N_7199,N_7016);
nand U7738 (N_7738,N_7286,N_7047);
xor U7739 (N_7739,N_7021,N_7475);
nor U7740 (N_7740,N_7449,N_7220);
xnor U7741 (N_7741,N_7395,N_7265);
or U7742 (N_7742,N_7407,N_7399);
nor U7743 (N_7743,N_7434,N_7424);
nand U7744 (N_7744,N_7400,N_7350);
and U7745 (N_7745,N_7073,N_7379);
xor U7746 (N_7746,N_7170,N_7165);
xnor U7747 (N_7747,N_7371,N_7115);
and U7748 (N_7748,N_7487,N_7452);
or U7749 (N_7749,N_7077,N_7045);
xnor U7750 (N_7750,N_7293,N_7390);
or U7751 (N_7751,N_7217,N_7247);
xnor U7752 (N_7752,N_7383,N_7303);
or U7753 (N_7753,N_7454,N_7366);
and U7754 (N_7754,N_7448,N_7135);
or U7755 (N_7755,N_7026,N_7380);
or U7756 (N_7756,N_7449,N_7363);
xor U7757 (N_7757,N_7118,N_7367);
and U7758 (N_7758,N_7021,N_7402);
xnor U7759 (N_7759,N_7426,N_7320);
xor U7760 (N_7760,N_7121,N_7206);
nand U7761 (N_7761,N_7075,N_7145);
xnor U7762 (N_7762,N_7108,N_7384);
or U7763 (N_7763,N_7449,N_7230);
and U7764 (N_7764,N_7495,N_7172);
xnor U7765 (N_7765,N_7446,N_7404);
xor U7766 (N_7766,N_7224,N_7168);
nor U7767 (N_7767,N_7405,N_7436);
xnor U7768 (N_7768,N_7044,N_7268);
and U7769 (N_7769,N_7449,N_7119);
xor U7770 (N_7770,N_7280,N_7418);
nand U7771 (N_7771,N_7152,N_7157);
and U7772 (N_7772,N_7101,N_7233);
or U7773 (N_7773,N_7214,N_7394);
nand U7774 (N_7774,N_7337,N_7101);
nand U7775 (N_7775,N_7234,N_7378);
xnor U7776 (N_7776,N_7123,N_7092);
nor U7777 (N_7777,N_7157,N_7216);
nor U7778 (N_7778,N_7260,N_7012);
nor U7779 (N_7779,N_7246,N_7095);
nand U7780 (N_7780,N_7486,N_7288);
and U7781 (N_7781,N_7064,N_7103);
xor U7782 (N_7782,N_7042,N_7003);
and U7783 (N_7783,N_7353,N_7056);
nor U7784 (N_7784,N_7009,N_7298);
and U7785 (N_7785,N_7306,N_7267);
nand U7786 (N_7786,N_7389,N_7161);
and U7787 (N_7787,N_7081,N_7338);
xnor U7788 (N_7788,N_7290,N_7294);
nand U7789 (N_7789,N_7443,N_7383);
nand U7790 (N_7790,N_7297,N_7253);
nor U7791 (N_7791,N_7040,N_7214);
or U7792 (N_7792,N_7326,N_7160);
or U7793 (N_7793,N_7107,N_7308);
nor U7794 (N_7794,N_7476,N_7091);
nand U7795 (N_7795,N_7333,N_7078);
nor U7796 (N_7796,N_7407,N_7020);
or U7797 (N_7797,N_7042,N_7461);
or U7798 (N_7798,N_7047,N_7453);
or U7799 (N_7799,N_7142,N_7450);
nor U7800 (N_7800,N_7342,N_7203);
xor U7801 (N_7801,N_7336,N_7353);
nor U7802 (N_7802,N_7232,N_7222);
or U7803 (N_7803,N_7016,N_7229);
xor U7804 (N_7804,N_7293,N_7283);
and U7805 (N_7805,N_7392,N_7112);
nand U7806 (N_7806,N_7364,N_7483);
nor U7807 (N_7807,N_7032,N_7472);
nand U7808 (N_7808,N_7302,N_7349);
xnor U7809 (N_7809,N_7067,N_7268);
or U7810 (N_7810,N_7488,N_7249);
xor U7811 (N_7811,N_7155,N_7395);
or U7812 (N_7812,N_7364,N_7498);
and U7813 (N_7813,N_7310,N_7306);
xor U7814 (N_7814,N_7416,N_7283);
nand U7815 (N_7815,N_7139,N_7207);
xor U7816 (N_7816,N_7308,N_7157);
and U7817 (N_7817,N_7237,N_7209);
or U7818 (N_7818,N_7034,N_7207);
or U7819 (N_7819,N_7222,N_7119);
and U7820 (N_7820,N_7492,N_7221);
and U7821 (N_7821,N_7399,N_7075);
xor U7822 (N_7822,N_7390,N_7349);
nand U7823 (N_7823,N_7368,N_7291);
xnor U7824 (N_7824,N_7012,N_7204);
nand U7825 (N_7825,N_7032,N_7245);
nor U7826 (N_7826,N_7404,N_7437);
nor U7827 (N_7827,N_7215,N_7253);
nand U7828 (N_7828,N_7251,N_7121);
and U7829 (N_7829,N_7159,N_7047);
nor U7830 (N_7830,N_7351,N_7281);
xnor U7831 (N_7831,N_7380,N_7483);
and U7832 (N_7832,N_7082,N_7162);
or U7833 (N_7833,N_7445,N_7087);
nand U7834 (N_7834,N_7310,N_7165);
xnor U7835 (N_7835,N_7488,N_7435);
or U7836 (N_7836,N_7168,N_7291);
nand U7837 (N_7837,N_7205,N_7490);
nand U7838 (N_7838,N_7294,N_7068);
and U7839 (N_7839,N_7173,N_7324);
or U7840 (N_7840,N_7453,N_7093);
or U7841 (N_7841,N_7294,N_7367);
nor U7842 (N_7842,N_7439,N_7079);
xor U7843 (N_7843,N_7100,N_7461);
nor U7844 (N_7844,N_7374,N_7063);
and U7845 (N_7845,N_7043,N_7480);
nand U7846 (N_7846,N_7100,N_7394);
nand U7847 (N_7847,N_7453,N_7416);
or U7848 (N_7848,N_7082,N_7114);
and U7849 (N_7849,N_7037,N_7007);
xor U7850 (N_7850,N_7349,N_7279);
or U7851 (N_7851,N_7097,N_7074);
or U7852 (N_7852,N_7114,N_7489);
xnor U7853 (N_7853,N_7440,N_7362);
and U7854 (N_7854,N_7310,N_7142);
or U7855 (N_7855,N_7206,N_7131);
xor U7856 (N_7856,N_7452,N_7198);
nand U7857 (N_7857,N_7228,N_7406);
nor U7858 (N_7858,N_7314,N_7300);
or U7859 (N_7859,N_7302,N_7165);
xnor U7860 (N_7860,N_7370,N_7053);
xor U7861 (N_7861,N_7454,N_7278);
nand U7862 (N_7862,N_7033,N_7021);
nand U7863 (N_7863,N_7091,N_7299);
nand U7864 (N_7864,N_7265,N_7145);
or U7865 (N_7865,N_7085,N_7436);
nand U7866 (N_7866,N_7498,N_7386);
xor U7867 (N_7867,N_7214,N_7324);
and U7868 (N_7868,N_7115,N_7135);
and U7869 (N_7869,N_7064,N_7330);
nand U7870 (N_7870,N_7085,N_7192);
or U7871 (N_7871,N_7432,N_7364);
and U7872 (N_7872,N_7440,N_7101);
and U7873 (N_7873,N_7299,N_7166);
xor U7874 (N_7874,N_7413,N_7172);
nor U7875 (N_7875,N_7086,N_7258);
or U7876 (N_7876,N_7390,N_7231);
xor U7877 (N_7877,N_7080,N_7126);
nor U7878 (N_7878,N_7188,N_7079);
and U7879 (N_7879,N_7431,N_7317);
and U7880 (N_7880,N_7449,N_7084);
xnor U7881 (N_7881,N_7201,N_7209);
xnor U7882 (N_7882,N_7269,N_7212);
xor U7883 (N_7883,N_7059,N_7273);
xnor U7884 (N_7884,N_7010,N_7219);
and U7885 (N_7885,N_7041,N_7012);
and U7886 (N_7886,N_7264,N_7273);
and U7887 (N_7887,N_7310,N_7437);
nor U7888 (N_7888,N_7197,N_7478);
nor U7889 (N_7889,N_7366,N_7346);
xnor U7890 (N_7890,N_7061,N_7230);
nand U7891 (N_7891,N_7172,N_7483);
nor U7892 (N_7892,N_7103,N_7332);
xnor U7893 (N_7893,N_7444,N_7090);
nand U7894 (N_7894,N_7127,N_7021);
nor U7895 (N_7895,N_7127,N_7180);
xnor U7896 (N_7896,N_7057,N_7260);
and U7897 (N_7897,N_7224,N_7286);
xor U7898 (N_7898,N_7464,N_7279);
xnor U7899 (N_7899,N_7086,N_7121);
and U7900 (N_7900,N_7194,N_7450);
xnor U7901 (N_7901,N_7125,N_7123);
nor U7902 (N_7902,N_7303,N_7350);
or U7903 (N_7903,N_7246,N_7139);
and U7904 (N_7904,N_7158,N_7044);
nand U7905 (N_7905,N_7499,N_7390);
or U7906 (N_7906,N_7273,N_7436);
nand U7907 (N_7907,N_7334,N_7139);
and U7908 (N_7908,N_7376,N_7406);
nor U7909 (N_7909,N_7151,N_7164);
and U7910 (N_7910,N_7021,N_7202);
or U7911 (N_7911,N_7375,N_7433);
xor U7912 (N_7912,N_7133,N_7325);
and U7913 (N_7913,N_7440,N_7469);
and U7914 (N_7914,N_7448,N_7154);
nor U7915 (N_7915,N_7402,N_7348);
xnor U7916 (N_7916,N_7062,N_7371);
xor U7917 (N_7917,N_7020,N_7306);
or U7918 (N_7918,N_7196,N_7190);
xnor U7919 (N_7919,N_7085,N_7098);
xor U7920 (N_7920,N_7076,N_7442);
and U7921 (N_7921,N_7226,N_7337);
or U7922 (N_7922,N_7008,N_7428);
or U7923 (N_7923,N_7142,N_7328);
nor U7924 (N_7924,N_7450,N_7172);
or U7925 (N_7925,N_7465,N_7314);
nor U7926 (N_7926,N_7318,N_7020);
nand U7927 (N_7927,N_7377,N_7251);
or U7928 (N_7928,N_7430,N_7164);
and U7929 (N_7929,N_7247,N_7278);
nand U7930 (N_7930,N_7295,N_7272);
and U7931 (N_7931,N_7023,N_7478);
nand U7932 (N_7932,N_7278,N_7367);
or U7933 (N_7933,N_7219,N_7434);
or U7934 (N_7934,N_7349,N_7268);
and U7935 (N_7935,N_7488,N_7127);
xor U7936 (N_7936,N_7420,N_7459);
xnor U7937 (N_7937,N_7069,N_7462);
nand U7938 (N_7938,N_7124,N_7340);
nor U7939 (N_7939,N_7351,N_7363);
xor U7940 (N_7940,N_7138,N_7214);
or U7941 (N_7941,N_7290,N_7354);
or U7942 (N_7942,N_7248,N_7069);
xnor U7943 (N_7943,N_7270,N_7264);
xnor U7944 (N_7944,N_7231,N_7262);
and U7945 (N_7945,N_7395,N_7196);
or U7946 (N_7946,N_7468,N_7280);
or U7947 (N_7947,N_7438,N_7471);
and U7948 (N_7948,N_7409,N_7359);
or U7949 (N_7949,N_7422,N_7345);
or U7950 (N_7950,N_7432,N_7044);
xor U7951 (N_7951,N_7449,N_7352);
nor U7952 (N_7952,N_7013,N_7430);
or U7953 (N_7953,N_7293,N_7499);
nand U7954 (N_7954,N_7370,N_7139);
xor U7955 (N_7955,N_7469,N_7063);
or U7956 (N_7956,N_7453,N_7139);
xnor U7957 (N_7957,N_7066,N_7462);
and U7958 (N_7958,N_7310,N_7350);
nand U7959 (N_7959,N_7320,N_7055);
nand U7960 (N_7960,N_7131,N_7217);
or U7961 (N_7961,N_7230,N_7300);
and U7962 (N_7962,N_7322,N_7328);
xor U7963 (N_7963,N_7427,N_7284);
or U7964 (N_7964,N_7031,N_7017);
xnor U7965 (N_7965,N_7213,N_7493);
and U7966 (N_7966,N_7010,N_7459);
xor U7967 (N_7967,N_7344,N_7375);
or U7968 (N_7968,N_7205,N_7191);
or U7969 (N_7969,N_7112,N_7374);
or U7970 (N_7970,N_7374,N_7318);
xor U7971 (N_7971,N_7109,N_7487);
nand U7972 (N_7972,N_7464,N_7206);
and U7973 (N_7973,N_7277,N_7172);
nor U7974 (N_7974,N_7430,N_7470);
xor U7975 (N_7975,N_7238,N_7081);
nor U7976 (N_7976,N_7127,N_7121);
and U7977 (N_7977,N_7426,N_7184);
xnor U7978 (N_7978,N_7055,N_7118);
nor U7979 (N_7979,N_7440,N_7437);
xnor U7980 (N_7980,N_7056,N_7473);
xnor U7981 (N_7981,N_7084,N_7221);
nor U7982 (N_7982,N_7454,N_7480);
nor U7983 (N_7983,N_7077,N_7466);
or U7984 (N_7984,N_7264,N_7454);
xor U7985 (N_7985,N_7357,N_7278);
nand U7986 (N_7986,N_7028,N_7393);
xnor U7987 (N_7987,N_7371,N_7253);
nand U7988 (N_7988,N_7219,N_7229);
or U7989 (N_7989,N_7058,N_7129);
xor U7990 (N_7990,N_7385,N_7154);
nand U7991 (N_7991,N_7462,N_7499);
nand U7992 (N_7992,N_7364,N_7092);
or U7993 (N_7993,N_7455,N_7320);
nand U7994 (N_7994,N_7270,N_7247);
xor U7995 (N_7995,N_7289,N_7483);
and U7996 (N_7996,N_7052,N_7040);
and U7997 (N_7997,N_7492,N_7094);
nor U7998 (N_7998,N_7316,N_7098);
nand U7999 (N_7999,N_7476,N_7088);
nor U8000 (N_8000,N_7926,N_7872);
or U8001 (N_8001,N_7618,N_7792);
nor U8002 (N_8002,N_7543,N_7973);
xor U8003 (N_8003,N_7550,N_7985);
nand U8004 (N_8004,N_7880,N_7750);
xor U8005 (N_8005,N_7732,N_7770);
or U8006 (N_8006,N_7947,N_7650);
or U8007 (N_8007,N_7779,N_7713);
xnor U8008 (N_8008,N_7517,N_7661);
and U8009 (N_8009,N_7606,N_7906);
or U8010 (N_8010,N_7610,N_7812);
nand U8011 (N_8011,N_7929,N_7678);
nand U8012 (N_8012,N_7931,N_7849);
xnor U8013 (N_8013,N_7876,N_7545);
nand U8014 (N_8014,N_7791,N_7911);
and U8015 (N_8015,N_7503,N_7711);
and U8016 (N_8016,N_7824,N_7832);
xnor U8017 (N_8017,N_7699,N_7975);
xnor U8018 (N_8018,N_7983,N_7687);
nor U8019 (N_8019,N_7788,N_7556);
nor U8020 (N_8020,N_7915,N_7706);
or U8021 (N_8021,N_7665,N_7596);
and U8022 (N_8022,N_7509,N_7857);
nand U8023 (N_8023,N_7619,N_7777);
xor U8024 (N_8024,N_7656,N_7666);
or U8025 (N_8025,N_7809,N_7978);
and U8026 (N_8026,N_7551,N_7722);
xor U8027 (N_8027,N_7840,N_7839);
xor U8028 (N_8028,N_7868,N_7755);
xnor U8029 (N_8029,N_7782,N_7982);
nor U8030 (N_8030,N_7515,N_7980);
and U8031 (N_8031,N_7932,N_7762);
nor U8032 (N_8032,N_7846,N_7505);
or U8033 (N_8033,N_7853,N_7753);
xnor U8034 (N_8034,N_7950,N_7508);
or U8035 (N_8035,N_7720,N_7647);
nand U8036 (N_8036,N_7574,N_7630);
and U8037 (N_8037,N_7524,N_7565);
or U8038 (N_8038,N_7916,N_7970);
or U8039 (N_8039,N_7953,N_7819);
nor U8040 (N_8040,N_7641,N_7771);
nand U8041 (N_8041,N_7654,N_7959);
xnor U8042 (N_8042,N_7585,N_7520);
nor U8043 (N_8043,N_7576,N_7512);
and U8044 (N_8044,N_7954,N_7579);
and U8045 (N_8045,N_7544,N_7659);
xor U8046 (N_8046,N_7958,N_7601);
nand U8047 (N_8047,N_7602,N_7967);
and U8048 (N_8048,N_7893,N_7935);
nand U8049 (N_8049,N_7856,N_7513);
xnor U8050 (N_8050,N_7940,N_7599);
or U8051 (N_8051,N_7859,N_7655);
xor U8052 (N_8052,N_7920,N_7588);
and U8053 (N_8053,N_7584,N_7575);
xor U8054 (N_8054,N_7863,N_7816);
nor U8055 (N_8055,N_7890,N_7884);
or U8056 (N_8056,N_7972,N_7651);
nor U8057 (N_8057,N_7761,N_7514);
nor U8058 (N_8058,N_7887,N_7541);
xor U8059 (N_8059,N_7608,N_7747);
xnor U8060 (N_8060,N_7852,N_7702);
xor U8061 (N_8061,N_7866,N_7718);
and U8062 (N_8062,N_7594,N_7673);
and U8063 (N_8063,N_7817,N_7581);
or U8064 (N_8064,N_7708,N_7552);
and U8065 (N_8065,N_7851,N_7997);
nor U8066 (N_8066,N_7578,N_7695);
or U8067 (N_8067,N_7729,N_7964);
nor U8068 (N_8068,N_7794,N_7639);
or U8069 (N_8069,N_7664,N_7912);
nor U8070 (N_8070,N_7539,N_7739);
xnor U8071 (N_8071,N_7583,N_7525);
or U8072 (N_8072,N_7765,N_7681);
nand U8073 (N_8073,N_7754,N_7534);
or U8074 (N_8074,N_7592,N_7790);
nor U8075 (N_8075,N_7821,N_7726);
and U8076 (N_8076,N_7632,N_7566);
or U8077 (N_8077,N_7614,N_7889);
nand U8078 (N_8078,N_7568,N_7527);
xor U8079 (N_8079,N_7553,N_7977);
xor U8080 (N_8080,N_7813,N_7921);
or U8081 (N_8081,N_7899,N_7786);
nor U8082 (N_8082,N_7784,N_7993);
and U8083 (N_8083,N_7591,N_7918);
nand U8084 (N_8084,N_7798,N_7757);
xnor U8085 (N_8085,N_7555,N_7700);
nand U8086 (N_8086,N_7617,N_7796);
xor U8087 (N_8087,N_7710,N_7737);
nor U8088 (N_8088,N_7774,N_7854);
xnor U8089 (N_8089,N_7598,N_7910);
nor U8090 (N_8090,N_7844,N_7586);
nor U8091 (N_8091,N_7537,N_7861);
xnor U8092 (N_8092,N_7989,N_7909);
or U8093 (N_8093,N_7806,N_7701);
nand U8094 (N_8094,N_7895,N_7956);
nand U8095 (N_8095,N_7728,N_7996);
nor U8096 (N_8096,N_7684,N_7736);
or U8097 (N_8097,N_7894,N_7628);
xnor U8098 (N_8098,N_7873,N_7886);
nand U8099 (N_8099,N_7607,N_7662);
nand U8100 (N_8100,N_7595,N_7669);
or U8101 (N_8101,N_7746,N_7690);
and U8102 (N_8102,N_7927,N_7877);
nor U8103 (N_8103,N_7674,N_7645);
nand U8104 (N_8104,N_7572,N_7529);
or U8105 (N_8105,N_7516,N_7671);
nor U8106 (N_8106,N_7905,N_7772);
nand U8107 (N_8107,N_7528,N_7526);
nand U8108 (N_8108,N_7917,N_7648);
xnor U8109 (N_8109,N_7871,N_7896);
nand U8110 (N_8110,N_7901,N_7810);
nor U8111 (N_8111,N_7533,N_7667);
xnor U8112 (N_8112,N_7941,N_7769);
nand U8113 (N_8113,N_7600,N_7603);
and U8114 (N_8114,N_7635,N_7763);
and U8115 (N_8115,N_7825,N_7837);
or U8116 (N_8116,N_7864,N_7914);
or U8117 (N_8117,N_7621,N_7587);
or U8118 (N_8118,N_7874,N_7968);
nor U8119 (N_8119,N_7963,N_7991);
nor U8120 (N_8120,N_7698,N_7760);
and U8121 (N_8121,N_7712,N_7878);
nand U8122 (N_8122,N_7974,N_7693);
nor U8123 (N_8123,N_7501,N_7580);
nand U8124 (N_8124,N_7843,N_7558);
and U8125 (N_8125,N_7946,N_7981);
and U8126 (N_8126,N_7797,N_7616);
xnor U8127 (N_8127,N_7676,N_7907);
nand U8128 (N_8128,N_7802,N_7631);
nand U8129 (N_8129,N_7738,N_7780);
nor U8130 (N_8130,N_7836,N_7823);
xor U8131 (N_8131,N_7721,N_7942);
or U8132 (N_8132,N_7875,N_7957);
xor U8133 (N_8133,N_7660,N_7948);
nor U8134 (N_8134,N_7742,N_7691);
or U8135 (N_8135,N_7766,N_7554);
nand U8136 (N_8136,N_7818,N_7745);
nor U8137 (N_8137,N_7799,N_7663);
or U8138 (N_8138,N_7727,N_7951);
nor U8139 (N_8139,N_7862,N_7506);
or U8140 (N_8140,N_7908,N_7749);
or U8141 (N_8141,N_7805,N_7923);
or U8142 (N_8142,N_7530,N_7775);
or U8143 (N_8143,N_7939,N_7623);
or U8144 (N_8144,N_7892,N_7891);
or U8145 (N_8145,N_7624,N_7627);
or U8146 (N_8146,N_7571,N_7507);
xnor U8147 (N_8147,N_7785,N_7783);
nand U8148 (N_8148,N_7882,N_7577);
nand U8149 (N_8149,N_7560,N_7930);
or U8150 (N_8150,N_7536,N_7789);
nand U8151 (N_8151,N_7962,N_7835);
nor U8152 (N_8152,N_7879,N_7865);
nand U8153 (N_8153,N_7833,N_7688);
and U8154 (N_8154,N_7697,N_7924);
nor U8155 (N_8155,N_7860,N_7960);
nand U8156 (N_8156,N_7820,N_7634);
and U8157 (N_8157,N_7764,N_7626);
nor U8158 (N_8158,N_7827,N_7987);
nor U8159 (N_8159,N_7888,N_7943);
and U8160 (N_8160,N_7900,N_7629);
nor U8161 (N_8161,N_7625,N_7547);
nor U8162 (N_8162,N_7672,N_7679);
nand U8163 (N_8163,N_7611,N_7692);
and U8164 (N_8164,N_7845,N_7999);
nand U8165 (N_8165,N_7500,N_7933);
nor U8166 (N_8166,N_7842,N_7850);
nor U8167 (N_8167,N_7620,N_7559);
xor U8168 (N_8168,N_7965,N_7613);
nand U8169 (N_8169,N_7609,N_7883);
or U8170 (N_8170,N_7535,N_7714);
nor U8171 (N_8171,N_7937,N_7969);
nor U8172 (N_8172,N_7546,N_7903);
and U8173 (N_8173,N_7604,N_7709);
nand U8174 (N_8174,N_7971,N_7828);
xnor U8175 (N_8175,N_7847,N_7740);
or U8176 (N_8176,N_7612,N_7694);
nand U8177 (N_8177,N_7902,N_7658);
nand U8178 (N_8178,N_7682,N_7961);
xnor U8179 (N_8179,N_7984,N_7640);
nor U8180 (N_8180,N_7925,N_7704);
nor U8181 (N_8181,N_7703,N_7653);
xnor U8182 (N_8182,N_7668,N_7756);
or U8183 (N_8183,N_7966,N_7787);
and U8184 (N_8184,N_7652,N_7689);
nor U8185 (N_8185,N_7815,N_7945);
or U8186 (N_8186,N_7686,N_7510);
or U8187 (N_8187,N_7938,N_7803);
and U8188 (N_8188,N_7758,N_7562);
nor U8189 (N_8189,N_7637,N_7502);
xor U8190 (N_8190,N_7646,N_7751);
and U8191 (N_8191,N_7622,N_7705);
or U8192 (N_8192,N_7724,N_7990);
and U8193 (N_8193,N_7532,N_7811);
or U8194 (N_8194,N_7743,N_7898);
nor U8195 (N_8195,N_7538,N_7934);
or U8196 (N_8196,N_7657,N_7913);
or U8197 (N_8197,N_7986,N_7573);
nand U8198 (N_8198,N_7944,N_7936);
and U8199 (N_8199,N_7597,N_7638);
or U8200 (N_8200,N_7952,N_7633);
nand U8201 (N_8201,N_7549,N_7519);
xor U8202 (N_8202,N_7838,N_7567);
and U8203 (N_8203,N_7593,N_7642);
xor U8204 (N_8204,N_7730,N_7735);
and U8205 (N_8205,N_7731,N_7670);
xnor U8206 (N_8206,N_7869,N_7522);
nor U8207 (N_8207,N_7707,N_7649);
nor U8208 (N_8208,N_7542,N_7570);
nor U8209 (N_8209,N_7808,N_7744);
xnor U8210 (N_8210,N_7870,N_7885);
xnor U8211 (N_8211,N_7561,N_7829);
or U8212 (N_8212,N_7826,N_7569);
and U8213 (N_8213,N_7680,N_7518);
nand U8214 (N_8214,N_7831,N_7848);
nor U8215 (N_8215,N_7855,N_7723);
nand U8216 (N_8216,N_7564,N_7976);
nand U8217 (N_8217,N_7685,N_7643);
nand U8218 (N_8218,N_7992,N_7834);
nand U8219 (N_8219,N_7725,N_7778);
and U8220 (N_8220,N_7841,N_7988);
and U8221 (N_8221,N_7800,N_7589);
nand U8222 (N_8222,N_7719,N_7677);
nand U8223 (N_8223,N_7949,N_7804);
xor U8224 (N_8224,N_7540,N_7904);
and U8225 (N_8225,N_7922,N_7858);
xnor U8226 (N_8226,N_7675,N_7683);
or U8227 (N_8227,N_7807,N_7897);
nand U8228 (N_8228,N_7557,N_7590);
xor U8229 (N_8229,N_7563,N_7773);
nor U8230 (N_8230,N_7995,N_7776);
and U8231 (N_8231,N_7795,N_7605);
xor U8232 (N_8232,N_7801,N_7994);
or U8233 (N_8233,N_7696,N_7523);
or U8234 (N_8234,N_7867,N_7781);
nand U8235 (N_8235,N_7615,N_7531);
nor U8236 (N_8236,N_7767,N_7881);
xnor U8237 (N_8237,N_7511,N_7830);
nand U8238 (N_8238,N_7955,N_7822);
or U8239 (N_8239,N_7717,N_7998);
nand U8240 (N_8240,N_7741,N_7644);
xnor U8241 (N_8241,N_7715,N_7636);
nand U8242 (N_8242,N_7548,N_7814);
xnor U8243 (N_8243,N_7752,N_7768);
nor U8244 (N_8244,N_7716,N_7979);
and U8245 (N_8245,N_7582,N_7733);
xor U8246 (N_8246,N_7748,N_7504);
or U8247 (N_8247,N_7759,N_7521);
nor U8248 (N_8248,N_7734,N_7928);
xnor U8249 (N_8249,N_7793,N_7919);
xor U8250 (N_8250,N_7818,N_7771);
nor U8251 (N_8251,N_7509,N_7808);
nor U8252 (N_8252,N_7846,N_7847);
nand U8253 (N_8253,N_7946,N_7869);
nand U8254 (N_8254,N_7606,N_7901);
xor U8255 (N_8255,N_7936,N_7778);
nor U8256 (N_8256,N_7694,N_7946);
nor U8257 (N_8257,N_7817,N_7935);
and U8258 (N_8258,N_7754,N_7755);
nor U8259 (N_8259,N_7542,N_7777);
nor U8260 (N_8260,N_7951,N_7763);
and U8261 (N_8261,N_7913,N_7699);
or U8262 (N_8262,N_7856,N_7787);
nor U8263 (N_8263,N_7982,N_7687);
xnor U8264 (N_8264,N_7798,N_7940);
nor U8265 (N_8265,N_7886,N_7618);
xor U8266 (N_8266,N_7928,N_7528);
or U8267 (N_8267,N_7599,N_7935);
and U8268 (N_8268,N_7795,N_7978);
or U8269 (N_8269,N_7906,N_7799);
nor U8270 (N_8270,N_7681,N_7861);
and U8271 (N_8271,N_7906,N_7905);
xnor U8272 (N_8272,N_7948,N_7932);
and U8273 (N_8273,N_7581,N_7593);
and U8274 (N_8274,N_7722,N_7987);
and U8275 (N_8275,N_7566,N_7558);
nor U8276 (N_8276,N_7508,N_7551);
nand U8277 (N_8277,N_7502,N_7538);
nor U8278 (N_8278,N_7710,N_7605);
and U8279 (N_8279,N_7503,N_7957);
nor U8280 (N_8280,N_7526,N_7938);
or U8281 (N_8281,N_7587,N_7838);
or U8282 (N_8282,N_7973,N_7734);
nand U8283 (N_8283,N_7957,N_7547);
nand U8284 (N_8284,N_7893,N_7777);
and U8285 (N_8285,N_7552,N_7778);
xnor U8286 (N_8286,N_7528,N_7779);
xnor U8287 (N_8287,N_7617,N_7962);
and U8288 (N_8288,N_7569,N_7864);
nand U8289 (N_8289,N_7911,N_7953);
xor U8290 (N_8290,N_7529,N_7801);
nand U8291 (N_8291,N_7856,N_7642);
nand U8292 (N_8292,N_7901,N_7799);
xor U8293 (N_8293,N_7554,N_7552);
nand U8294 (N_8294,N_7883,N_7732);
nor U8295 (N_8295,N_7961,N_7878);
or U8296 (N_8296,N_7523,N_7867);
or U8297 (N_8297,N_7773,N_7914);
xnor U8298 (N_8298,N_7782,N_7804);
nand U8299 (N_8299,N_7811,N_7714);
nand U8300 (N_8300,N_7982,N_7532);
or U8301 (N_8301,N_7977,N_7550);
nand U8302 (N_8302,N_7729,N_7555);
xor U8303 (N_8303,N_7597,N_7561);
nor U8304 (N_8304,N_7785,N_7503);
and U8305 (N_8305,N_7866,N_7838);
xor U8306 (N_8306,N_7545,N_7884);
or U8307 (N_8307,N_7932,N_7850);
nor U8308 (N_8308,N_7613,N_7959);
nand U8309 (N_8309,N_7881,N_7833);
and U8310 (N_8310,N_7723,N_7679);
nand U8311 (N_8311,N_7616,N_7622);
nand U8312 (N_8312,N_7706,N_7879);
nand U8313 (N_8313,N_7561,N_7846);
nand U8314 (N_8314,N_7626,N_7606);
and U8315 (N_8315,N_7978,N_7938);
nor U8316 (N_8316,N_7783,N_7588);
and U8317 (N_8317,N_7868,N_7606);
xnor U8318 (N_8318,N_7843,N_7531);
xor U8319 (N_8319,N_7645,N_7768);
xnor U8320 (N_8320,N_7847,N_7746);
xnor U8321 (N_8321,N_7975,N_7521);
xor U8322 (N_8322,N_7872,N_7511);
and U8323 (N_8323,N_7722,N_7751);
nand U8324 (N_8324,N_7991,N_7702);
and U8325 (N_8325,N_7663,N_7788);
nand U8326 (N_8326,N_7621,N_7899);
nor U8327 (N_8327,N_7997,N_7913);
and U8328 (N_8328,N_7911,N_7873);
nand U8329 (N_8329,N_7646,N_7554);
nor U8330 (N_8330,N_7864,N_7866);
and U8331 (N_8331,N_7976,N_7844);
xor U8332 (N_8332,N_7932,N_7740);
xor U8333 (N_8333,N_7674,N_7910);
or U8334 (N_8334,N_7738,N_7535);
and U8335 (N_8335,N_7651,N_7774);
nor U8336 (N_8336,N_7842,N_7747);
or U8337 (N_8337,N_7791,N_7859);
nand U8338 (N_8338,N_7685,N_7720);
and U8339 (N_8339,N_7575,N_7851);
nand U8340 (N_8340,N_7672,N_7531);
xnor U8341 (N_8341,N_7807,N_7556);
or U8342 (N_8342,N_7664,N_7941);
nand U8343 (N_8343,N_7967,N_7551);
or U8344 (N_8344,N_7919,N_7920);
and U8345 (N_8345,N_7595,N_7692);
nor U8346 (N_8346,N_7765,N_7512);
and U8347 (N_8347,N_7717,N_7805);
and U8348 (N_8348,N_7849,N_7692);
xnor U8349 (N_8349,N_7805,N_7681);
nor U8350 (N_8350,N_7884,N_7958);
or U8351 (N_8351,N_7879,N_7768);
nand U8352 (N_8352,N_7556,N_7565);
or U8353 (N_8353,N_7519,N_7802);
nand U8354 (N_8354,N_7722,N_7743);
and U8355 (N_8355,N_7872,N_7821);
nand U8356 (N_8356,N_7997,N_7734);
xnor U8357 (N_8357,N_7811,N_7949);
or U8358 (N_8358,N_7889,N_7866);
xnor U8359 (N_8359,N_7965,N_7954);
nand U8360 (N_8360,N_7780,N_7956);
nor U8361 (N_8361,N_7845,N_7595);
nand U8362 (N_8362,N_7919,N_7757);
nor U8363 (N_8363,N_7885,N_7722);
nand U8364 (N_8364,N_7801,N_7995);
or U8365 (N_8365,N_7867,N_7853);
nand U8366 (N_8366,N_7662,N_7738);
xor U8367 (N_8367,N_7776,N_7561);
xnor U8368 (N_8368,N_7897,N_7693);
nand U8369 (N_8369,N_7659,N_7793);
nor U8370 (N_8370,N_7583,N_7883);
and U8371 (N_8371,N_7972,N_7700);
nor U8372 (N_8372,N_7734,N_7604);
xor U8373 (N_8373,N_7613,N_7573);
nand U8374 (N_8374,N_7795,N_7732);
nand U8375 (N_8375,N_7646,N_7552);
nor U8376 (N_8376,N_7534,N_7810);
or U8377 (N_8377,N_7636,N_7644);
or U8378 (N_8378,N_7944,N_7836);
nor U8379 (N_8379,N_7649,N_7877);
xor U8380 (N_8380,N_7931,N_7834);
or U8381 (N_8381,N_7622,N_7637);
nor U8382 (N_8382,N_7531,N_7575);
nand U8383 (N_8383,N_7774,N_7556);
and U8384 (N_8384,N_7754,N_7616);
nand U8385 (N_8385,N_7914,N_7506);
nand U8386 (N_8386,N_7621,N_7960);
or U8387 (N_8387,N_7937,N_7691);
nor U8388 (N_8388,N_7902,N_7533);
nor U8389 (N_8389,N_7690,N_7885);
nor U8390 (N_8390,N_7951,N_7734);
or U8391 (N_8391,N_7828,N_7618);
and U8392 (N_8392,N_7673,N_7834);
or U8393 (N_8393,N_7599,N_7898);
xnor U8394 (N_8394,N_7912,N_7883);
and U8395 (N_8395,N_7766,N_7911);
nand U8396 (N_8396,N_7753,N_7509);
nand U8397 (N_8397,N_7731,N_7994);
or U8398 (N_8398,N_7632,N_7606);
and U8399 (N_8399,N_7710,N_7806);
or U8400 (N_8400,N_7862,N_7793);
nor U8401 (N_8401,N_7699,N_7599);
xnor U8402 (N_8402,N_7514,N_7772);
or U8403 (N_8403,N_7828,N_7794);
xnor U8404 (N_8404,N_7931,N_7613);
nand U8405 (N_8405,N_7995,N_7648);
or U8406 (N_8406,N_7658,N_7849);
nand U8407 (N_8407,N_7987,N_7571);
nand U8408 (N_8408,N_7800,N_7922);
and U8409 (N_8409,N_7649,N_7815);
nand U8410 (N_8410,N_7630,N_7928);
or U8411 (N_8411,N_7753,N_7959);
nand U8412 (N_8412,N_7879,N_7994);
nand U8413 (N_8413,N_7508,N_7704);
nor U8414 (N_8414,N_7600,N_7642);
xor U8415 (N_8415,N_7619,N_7549);
nand U8416 (N_8416,N_7915,N_7758);
xnor U8417 (N_8417,N_7788,N_7808);
nor U8418 (N_8418,N_7773,N_7540);
or U8419 (N_8419,N_7631,N_7958);
and U8420 (N_8420,N_7687,N_7580);
and U8421 (N_8421,N_7975,N_7764);
or U8422 (N_8422,N_7532,N_7757);
nand U8423 (N_8423,N_7816,N_7905);
xor U8424 (N_8424,N_7576,N_7752);
nor U8425 (N_8425,N_7900,N_7602);
or U8426 (N_8426,N_7726,N_7661);
and U8427 (N_8427,N_7686,N_7606);
and U8428 (N_8428,N_7685,N_7978);
xnor U8429 (N_8429,N_7627,N_7871);
and U8430 (N_8430,N_7788,N_7846);
nor U8431 (N_8431,N_7827,N_7865);
nand U8432 (N_8432,N_7849,N_7835);
nor U8433 (N_8433,N_7864,N_7872);
xnor U8434 (N_8434,N_7500,N_7795);
nand U8435 (N_8435,N_7719,N_7565);
nor U8436 (N_8436,N_7899,N_7930);
and U8437 (N_8437,N_7916,N_7831);
nor U8438 (N_8438,N_7703,N_7553);
and U8439 (N_8439,N_7812,N_7508);
nor U8440 (N_8440,N_7662,N_7521);
nor U8441 (N_8441,N_7500,N_7901);
nor U8442 (N_8442,N_7642,N_7805);
xor U8443 (N_8443,N_7533,N_7863);
nand U8444 (N_8444,N_7538,N_7790);
xor U8445 (N_8445,N_7562,N_7967);
xor U8446 (N_8446,N_7658,N_7836);
nor U8447 (N_8447,N_7762,N_7720);
xor U8448 (N_8448,N_7638,N_7608);
xor U8449 (N_8449,N_7630,N_7642);
nand U8450 (N_8450,N_7637,N_7508);
and U8451 (N_8451,N_7536,N_7849);
nand U8452 (N_8452,N_7774,N_7873);
nand U8453 (N_8453,N_7682,N_7773);
nor U8454 (N_8454,N_7957,N_7698);
nand U8455 (N_8455,N_7929,N_7542);
nor U8456 (N_8456,N_7609,N_7500);
nor U8457 (N_8457,N_7742,N_7583);
and U8458 (N_8458,N_7735,N_7715);
nand U8459 (N_8459,N_7580,N_7790);
nand U8460 (N_8460,N_7632,N_7997);
xnor U8461 (N_8461,N_7748,N_7518);
xor U8462 (N_8462,N_7610,N_7621);
and U8463 (N_8463,N_7584,N_7982);
nor U8464 (N_8464,N_7547,N_7793);
nor U8465 (N_8465,N_7604,N_7777);
nand U8466 (N_8466,N_7834,N_7716);
or U8467 (N_8467,N_7734,N_7975);
nand U8468 (N_8468,N_7702,N_7648);
xor U8469 (N_8469,N_7844,N_7705);
nor U8470 (N_8470,N_7752,N_7714);
and U8471 (N_8471,N_7641,N_7915);
and U8472 (N_8472,N_7639,N_7731);
xnor U8473 (N_8473,N_7976,N_7918);
nor U8474 (N_8474,N_7969,N_7520);
xor U8475 (N_8475,N_7930,N_7514);
nand U8476 (N_8476,N_7782,N_7607);
or U8477 (N_8477,N_7949,N_7847);
nor U8478 (N_8478,N_7643,N_7894);
nand U8479 (N_8479,N_7883,N_7779);
nor U8480 (N_8480,N_7576,N_7890);
nand U8481 (N_8481,N_7600,N_7546);
and U8482 (N_8482,N_7917,N_7974);
and U8483 (N_8483,N_7544,N_7668);
and U8484 (N_8484,N_7712,N_7530);
and U8485 (N_8485,N_7576,N_7957);
nand U8486 (N_8486,N_7964,N_7613);
xnor U8487 (N_8487,N_7741,N_7812);
and U8488 (N_8488,N_7710,N_7858);
nor U8489 (N_8489,N_7610,N_7802);
or U8490 (N_8490,N_7899,N_7763);
nor U8491 (N_8491,N_7521,N_7666);
nor U8492 (N_8492,N_7768,N_7769);
xnor U8493 (N_8493,N_7883,N_7909);
xor U8494 (N_8494,N_7678,N_7511);
nor U8495 (N_8495,N_7936,N_7605);
nor U8496 (N_8496,N_7543,N_7871);
or U8497 (N_8497,N_7586,N_7680);
and U8498 (N_8498,N_7730,N_7789);
nor U8499 (N_8499,N_7878,N_7944);
or U8500 (N_8500,N_8199,N_8238);
or U8501 (N_8501,N_8414,N_8221);
nor U8502 (N_8502,N_8269,N_8067);
nand U8503 (N_8503,N_8327,N_8307);
nand U8504 (N_8504,N_8422,N_8013);
or U8505 (N_8505,N_8407,N_8202);
nand U8506 (N_8506,N_8046,N_8039);
nor U8507 (N_8507,N_8137,N_8064);
xnor U8508 (N_8508,N_8430,N_8331);
xnor U8509 (N_8509,N_8127,N_8019);
nor U8510 (N_8510,N_8343,N_8033);
nor U8511 (N_8511,N_8465,N_8245);
and U8512 (N_8512,N_8399,N_8017);
xnor U8513 (N_8513,N_8003,N_8165);
and U8514 (N_8514,N_8442,N_8432);
or U8515 (N_8515,N_8295,N_8096);
or U8516 (N_8516,N_8333,N_8193);
or U8517 (N_8517,N_8301,N_8231);
nand U8518 (N_8518,N_8382,N_8380);
and U8519 (N_8519,N_8481,N_8479);
or U8520 (N_8520,N_8290,N_8337);
xnor U8521 (N_8521,N_8268,N_8120);
nand U8522 (N_8522,N_8248,N_8443);
nor U8523 (N_8523,N_8371,N_8330);
or U8524 (N_8524,N_8404,N_8474);
nand U8525 (N_8525,N_8392,N_8326);
xnor U8526 (N_8526,N_8411,N_8316);
and U8527 (N_8527,N_8104,N_8010);
nand U8528 (N_8528,N_8142,N_8183);
and U8529 (N_8529,N_8298,N_8354);
xor U8530 (N_8530,N_8053,N_8150);
nand U8531 (N_8531,N_8169,N_8141);
xor U8532 (N_8532,N_8418,N_8420);
or U8533 (N_8533,N_8243,N_8312);
nand U8534 (N_8534,N_8004,N_8396);
nor U8535 (N_8535,N_8031,N_8457);
nor U8536 (N_8536,N_8085,N_8112);
nand U8537 (N_8537,N_8216,N_8272);
and U8538 (N_8538,N_8277,N_8487);
nand U8539 (N_8539,N_8105,N_8296);
and U8540 (N_8540,N_8350,N_8223);
or U8541 (N_8541,N_8372,N_8473);
or U8542 (N_8542,N_8176,N_8138);
nand U8543 (N_8543,N_8357,N_8450);
xor U8544 (N_8544,N_8126,N_8251);
or U8545 (N_8545,N_8065,N_8449);
and U8546 (N_8546,N_8288,N_8116);
xor U8547 (N_8547,N_8247,N_8008);
xor U8548 (N_8548,N_8421,N_8304);
and U8549 (N_8549,N_8109,N_8149);
nand U8550 (N_8550,N_8032,N_8060);
nor U8551 (N_8551,N_8066,N_8082);
and U8552 (N_8552,N_8424,N_8070);
nand U8553 (N_8553,N_8485,N_8376);
nand U8554 (N_8554,N_8428,N_8208);
and U8555 (N_8555,N_8219,N_8419);
or U8556 (N_8556,N_8388,N_8348);
xnor U8557 (N_8557,N_8283,N_8262);
nor U8558 (N_8558,N_8101,N_8211);
and U8559 (N_8559,N_8029,N_8075);
xor U8560 (N_8560,N_8475,N_8198);
nand U8561 (N_8561,N_8106,N_8001);
nor U8562 (N_8562,N_8145,N_8117);
and U8563 (N_8563,N_8226,N_8488);
and U8564 (N_8564,N_8466,N_8284);
and U8565 (N_8565,N_8207,N_8427);
xnor U8566 (N_8566,N_8203,N_8244);
xnor U8567 (N_8567,N_8389,N_8016);
nand U8568 (N_8568,N_8214,N_8297);
or U8569 (N_8569,N_8002,N_8254);
nand U8570 (N_8570,N_8071,N_8072);
nor U8571 (N_8571,N_8306,N_8212);
nand U8572 (N_8572,N_8195,N_8115);
or U8573 (N_8573,N_8291,N_8433);
or U8574 (N_8574,N_8406,N_8157);
nand U8575 (N_8575,N_8246,N_8220);
and U8576 (N_8576,N_8040,N_8302);
xor U8577 (N_8577,N_8274,N_8186);
nor U8578 (N_8578,N_8081,N_8394);
nor U8579 (N_8579,N_8006,N_8403);
or U8580 (N_8580,N_8240,N_8287);
xnor U8581 (N_8581,N_8439,N_8477);
xor U8582 (N_8582,N_8147,N_8484);
xnor U8583 (N_8583,N_8467,N_8119);
nor U8584 (N_8584,N_8472,N_8448);
nor U8585 (N_8585,N_8218,N_8332);
or U8586 (N_8586,N_8061,N_8289);
or U8587 (N_8587,N_8197,N_8387);
nor U8588 (N_8588,N_8050,N_8471);
xor U8589 (N_8589,N_8148,N_8217);
and U8590 (N_8590,N_8166,N_8490);
and U8591 (N_8591,N_8163,N_8317);
nand U8592 (N_8592,N_8410,N_8063);
nand U8593 (N_8593,N_8400,N_8462);
or U8594 (N_8594,N_8324,N_8042);
xor U8595 (N_8595,N_8489,N_8021);
nor U8596 (N_8596,N_8267,N_8276);
nand U8597 (N_8597,N_8027,N_8305);
xnor U8598 (N_8598,N_8250,N_8131);
xor U8599 (N_8599,N_8275,N_8379);
nor U8600 (N_8600,N_8162,N_8359);
xnor U8601 (N_8601,N_8405,N_8413);
nor U8602 (N_8602,N_8018,N_8395);
nand U8603 (N_8603,N_8187,N_8076);
nor U8604 (N_8604,N_8089,N_8456);
and U8605 (N_8605,N_8177,N_8328);
nor U8606 (N_8606,N_8447,N_8007);
nand U8607 (N_8607,N_8415,N_8256);
and U8608 (N_8608,N_8113,N_8130);
nand U8609 (N_8609,N_8318,N_8263);
and U8610 (N_8610,N_8213,N_8300);
or U8611 (N_8611,N_8329,N_8340);
nor U8612 (N_8612,N_8498,N_8100);
xnor U8613 (N_8613,N_8239,N_8058);
or U8614 (N_8614,N_8125,N_8034);
nor U8615 (N_8615,N_8453,N_8230);
and U8616 (N_8616,N_8429,N_8325);
nand U8617 (N_8617,N_8286,N_8423);
xnor U8618 (N_8618,N_8228,N_8047);
nor U8619 (N_8619,N_8139,N_8092);
nor U8620 (N_8620,N_8152,N_8035);
or U8621 (N_8621,N_8417,N_8069);
and U8622 (N_8622,N_8043,N_8179);
nor U8623 (N_8623,N_8355,N_8270);
and U8624 (N_8624,N_8320,N_8074);
or U8625 (N_8625,N_8015,N_8486);
nor U8626 (N_8626,N_8215,N_8431);
or U8627 (N_8627,N_8049,N_8036);
xnor U8628 (N_8628,N_8401,N_8025);
xor U8629 (N_8629,N_8459,N_8279);
nor U8630 (N_8630,N_8129,N_8201);
and U8631 (N_8631,N_8460,N_8170);
xnor U8632 (N_8632,N_8103,N_8026);
nor U8633 (N_8633,N_8227,N_8482);
or U8634 (N_8634,N_8168,N_8383);
nand U8635 (N_8635,N_8178,N_8242);
nand U8636 (N_8636,N_8059,N_8237);
and U8637 (N_8637,N_8365,N_8140);
nor U8638 (N_8638,N_8252,N_8191);
nor U8639 (N_8639,N_8110,N_8153);
or U8640 (N_8640,N_8336,N_8342);
and U8641 (N_8641,N_8257,N_8079);
nand U8642 (N_8642,N_8345,N_8347);
and U8643 (N_8643,N_8133,N_8356);
xnor U8644 (N_8644,N_8483,N_8044);
and U8645 (N_8645,N_8224,N_8020);
and U8646 (N_8646,N_8155,N_8098);
nand U8647 (N_8647,N_8353,N_8088);
xnor U8648 (N_8648,N_8041,N_8366);
or U8649 (N_8649,N_8361,N_8122);
xor U8650 (N_8650,N_8206,N_8038);
and U8651 (N_8651,N_8167,N_8143);
or U8652 (N_8652,N_8095,N_8437);
nor U8653 (N_8653,N_8121,N_8260);
xnor U8654 (N_8654,N_8363,N_8196);
xnor U8655 (N_8655,N_8362,N_8144);
and U8656 (N_8656,N_8086,N_8154);
or U8657 (N_8657,N_8311,N_8390);
or U8658 (N_8658,N_8408,N_8077);
or U8659 (N_8659,N_8370,N_8232);
or U8660 (N_8660,N_8055,N_8452);
or U8661 (N_8661,N_8062,N_8194);
nand U8662 (N_8662,N_8210,N_8451);
nand U8663 (N_8663,N_8303,N_8334);
xor U8664 (N_8664,N_8159,N_8160);
xor U8665 (N_8665,N_8461,N_8023);
and U8666 (N_8666,N_8436,N_8346);
and U8667 (N_8667,N_8409,N_8377);
and U8668 (N_8668,N_8037,N_8273);
nand U8669 (N_8669,N_8315,N_8102);
nor U8670 (N_8670,N_8259,N_8083);
nand U8671 (N_8671,N_8281,N_8444);
nor U8672 (N_8672,N_8173,N_8135);
nor U8673 (N_8673,N_8124,N_8434);
or U8674 (N_8674,N_8373,N_8308);
xor U8675 (N_8675,N_8045,N_8011);
xnor U8676 (N_8676,N_8496,N_8146);
or U8677 (N_8677,N_8054,N_8381);
nand U8678 (N_8678,N_8181,N_8402);
nand U8679 (N_8679,N_8182,N_8294);
nand U8680 (N_8680,N_8398,N_8497);
xnor U8681 (N_8681,N_8323,N_8156);
or U8682 (N_8682,N_8374,N_8024);
and U8683 (N_8683,N_8249,N_8078);
xor U8684 (N_8684,N_8494,N_8292);
nand U8685 (N_8685,N_8087,N_8000);
xor U8686 (N_8686,N_8192,N_8090);
xnor U8687 (N_8687,N_8057,N_8200);
xor U8688 (N_8688,N_8368,N_8480);
nor U8689 (N_8689,N_8093,N_8378);
nand U8690 (N_8690,N_8299,N_8446);
and U8691 (N_8691,N_8118,N_8136);
nor U8692 (N_8692,N_8080,N_8493);
xor U8693 (N_8693,N_8180,N_8454);
xnor U8694 (N_8694,N_8385,N_8271);
nand U8695 (N_8695,N_8164,N_8158);
and U8696 (N_8696,N_8360,N_8364);
and U8697 (N_8697,N_8234,N_8123);
nand U8698 (N_8698,N_8204,N_8190);
and U8699 (N_8699,N_8222,N_8351);
xnor U8700 (N_8700,N_8293,N_8205);
nor U8701 (N_8701,N_8492,N_8416);
xor U8702 (N_8702,N_8012,N_8280);
or U8703 (N_8703,N_8335,N_8464);
or U8704 (N_8704,N_8491,N_8174);
xor U8705 (N_8705,N_8282,N_8229);
nor U8706 (N_8706,N_8175,N_8111);
nor U8707 (N_8707,N_8310,N_8352);
nand U8708 (N_8708,N_8476,N_8185);
nor U8709 (N_8709,N_8495,N_8313);
nor U8710 (N_8710,N_8233,N_8107);
xnor U8711 (N_8711,N_8309,N_8028);
nand U8712 (N_8712,N_8265,N_8261);
xor U8713 (N_8713,N_8397,N_8258);
and U8714 (N_8714,N_8068,N_8321);
nor U8715 (N_8715,N_8253,N_8266);
nor U8716 (N_8716,N_8009,N_8441);
or U8717 (N_8717,N_8225,N_8445);
nor U8718 (N_8718,N_8048,N_8369);
nor U8719 (N_8719,N_8458,N_8171);
nand U8720 (N_8720,N_8469,N_8285);
and U8721 (N_8721,N_8255,N_8438);
nor U8722 (N_8722,N_8114,N_8151);
nor U8723 (N_8723,N_8344,N_8188);
nor U8724 (N_8724,N_8052,N_8014);
xnor U8725 (N_8725,N_8278,N_8314);
nand U8726 (N_8726,N_8132,N_8264);
or U8727 (N_8727,N_8339,N_8499);
xor U8728 (N_8728,N_8235,N_8463);
nand U8729 (N_8729,N_8005,N_8241);
or U8730 (N_8730,N_8094,N_8056);
nand U8731 (N_8731,N_8051,N_8236);
and U8732 (N_8732,N_8128,N_8349);
xnor U8733 (N_8733,N_8468,N_8358);
or U8734 (N_8734,N_8099,N_8184);
or U8735 (N_8735,N_8426,N_8391);
xnor U8736 (N_8736,N_8367,N_8384);
and U8737 (N_8737,N_8386,N_8022);
nor U8738 (N_8738,N_8189,N_8341);
xnor U8739 (N_8739,N_8209,N_8030);
xnor U8740 (N_8740,N_8073,N_8172);
and U8741 (N_8741,N_8393,N_8412);
or U8742 (N_8742,N_8440,N_8478);
xnor U8743 (N_8743,N_8338,N_8134);
nor U8744 (N_8744,N_8470,N_8425);
nor U8745 (N_8745,N_8097,N_8375);
xor U8746 (N_8746,N_8435,N_8455);
nor U8747 (N_8747,N_8322,N_8161);
or U8748 (N_8748,N_8091,N_8319);
nand U8749 (N_8749,N_8084,N_8108);
or U8750 (N_8750,N_8284,N_8339);
nand U8751 (N_8751,N_8429,N_8180);
and U8752 (N_8752,N_8255,N_8131);
and U8753 (N_8753,N_8113,N_8339);
nor U8754 (N_8754,N_8100,N_8327);
xor U8755 (N_8755,N_8191,N_8276);
nand U8756 (N_8756,N_8441,N_8184);
nand U8757 (N_8757,N_8191,N_8133);
xor U8758 (N_8758,N_8376,N_8264);
or U8759 (N_8759,N_8435,N_8150);
nand U8760 (N_8760,N_8078,N_8302);
xnor U8761 (N_8761,N_8094,N_8011);
nand U8762 (N_8762,N_8088,N_8399);
or U8763 (N_8763,N_8105,N_8364);
nor U8764 (N_8764,N_8091,N_8080);
nor U8765 (N_8765,N_8385,N_8038);
xor U8766 (N_8766,N_8153,N_8338);
or U8767 (N_8767,N_8210,N_8458);
and U8768 (N_8768,N_8462,N_8382);
or U8769 (N_8769,N_8014,N_8087);
xor U8770 (N_8770,N_8167,N_8388);
and U8771 (N_8771,N_8306,N_8221);
nor U8772 (N_8772,N_8321,N_8367);
xnor U8773 (N_8773,N_8275,N_8189);
nor U8774 (N_8774,N_8154,N_8070);
nor U8775 (N_8775,N_8072,N_8035);
xnor U8776 (N_8776,N_8080,N_8281);
nor U8777 (N_8777,N_8479,N_8291);
xor U8778 (N_8778,N_8440,N_8082);
xor U8779 (N_8779,N_8053,N_8476);
xnor U8780 (N_8780,N_8108,N_8245);
xor U8781 (N_8781,N_8010,N_8459);
or U8782 (N_8782,N_8262,N_8142);
xnor U8783 (N_8783,N_8340,N_8261);
and U8784 (N_8784,N_8210,N_8416);
nand U8785 (N_8785,N_8331,N_8004);
nand U8786 (N_8786,N_8064,N_8348);
or U8787 (N_8787,N_8339,N_8158);
nor U8788 (N_8788,N_8369,N_8115);
nor U8789 (N_8789,N_8238,N_8333);
xnor U8790 (N_8790,N_8294,N_8168);
nand U8791 (N_8791,N_8100,N_8430);
nand U8792 (N_8792,N_8013,N_8327);
xor U8793 (N_8793,N_8100,N_8409);
xnor U8794 (N_8794,N_8401,N_8392);
and U8795 (N_8795,N_8428,N_8243);
xnor U8796 (N_8796,N_8288,N_8068);
xnor U8797 (N_8797,N_8429,N_8445);
nand U8798 (N_8798,N_8300,N_8407);
nor U8799 (N_8799,N_8373,N_8045);
nor U8800 (N_8800,N_8204,N_8093);
and U8801 (N_8801,N_8106,N_8360);
and U8802 (N_8802,N_8391,N_8133);
or U8803 (N_8803,N_8471,N_8105);
and U8804 (N_8804,N_8405,N_8364);
nor U8805 (N_8805,N_8317,N_8342);
nor U8806 (N_8806,N_8168,N_8267);
xor U8807 (N_8807,N_8097,N_8379);
and U8808 (N_8808,N_8448,N_8294);
xnor U8809 (N_8809,N_8193,N_8148);
or U8810 (N_8810,N_8359,N_8218);
or U8811 (N_8811,N_8106,N_8108);
or U8812 (N_8812,N_8329,N_8252);
or U8813 (N_8813,N_8329,N_8363);
nand U8814 (N_8814,N_8190,N_8125);
nor U8815 (N_8815,N_8264,N_8257);
nand U8816 (N_8816,N_8164,N_8132);
and U8817 (N_8817,N_8309,N_8030);
xnor U8818 (N_8818,N_8076,N_8059);
or U8819 (N_8819,N_8087,N_8250);
and U8820 (N_8820,N_8446,N_8329);
nor U8821 (N_8821,N_8233,N_8453);
or U8822 (N_8822,N_8283,N_8474);
nor U8823 (N_8823,N_8152,N_8014);
nand U8824 (N_8824,N_8055,N_8382);
or U8825 (N_8825,N_8344,N_8135);
and U8826 (N_8826,N_8277,N_8363);
and U8827 (N_8827,N_8028,N_8191);
nand U8828 (N_8828,N_8438,N_8451);
xnor U8829 (N_8829,N_8044,N_8489);
or U8830 (N_8830,N_8487,N_8058);
xnor U8831 (N_8831,N_8075,N_8180);
xor U8832 (N_8832,N_8124,N_8317);
nand U8833 (N_8833,N_8211,N_8337);
nor U8834 (N_8834,N_8012,N_8278);
or U8835 (N_8835,N_8469,N_8091);
and U8836 (N_8836,N_8301,N_8055);
nor U8837 (N_8837,N_8421,N_8054);
nand U8838 (N_8838,N_8060,N_8132);
or U8839 (N_8839,N_8036,N_8136);
nand U8840 (N_8840,N_8280,N_8499);
and U8841 (N_8841,N_8382,N_8476);
nand U8842 (N_8842,N_8028,N_8334);
xnor U8843 (N_8843,N_8301,N_8468);
or U8844 (N_8844,N_8232,N_8261);
nor U8845 (N_8845,N_8335,N_8185);
nand U8846 (N_8846,N_8000,N_8106);
and U8847 (N_8847,N_8409,N_8183);
and U8848 (N_8848,N_8297,N_8051);
xnor U8849 (N_8849,N_8331,N_8414);
xnor U8850 (N_8850,N_8352,N_8026);
or U8851 (N_8851,N_8433,N_8207);
or U8852 (N_8852,N_8077,N_8153);
and U8853 (N_8853,N_8014,N_8226);
xor U8854 (N_8854,N_8253,N_8173);
nor U8855 (N_8855,N_8468,N_8481);
xor U8856 (N_8856,N_8229,N_8324);
and U8857 (N_8857,N_8162,N_8227);
or U8858 (N_8858,N_8265,N_8461);
or U8859 (N_8859,N_8316,N_8375);
nand U8860 (N_8860,N_8251,N_8044);
xor U8861 (N_8861,N_8453,N_8301);
nand U8862 (N_8862,N_8413,N_8121);
nand U8863 (N_8863,N_8367,N_8320);
or U8864 (N_8864,N_8437,N_8077);
nor U8865 (N_8865,N_8478,N_8077);
nand U8866 (N_8866,N_8140,N_8006);
nand U8867 (N_8867,N_8356,N_8290);
and U8868 (N_8868,N_8397,N_8151);
or U8869 (N_8869,N_8179,N_8302);
and U8870 (N_8870,N_8086,N_8398);
nand U8871 (N_8871,N_8260,N_8382);
or U8872 (N_8872,N_8269,N_8145);
nand U8873 (N_8873,N_8282,N_8398);
xnor U8874 (N_8874,N_8432,N_8347);
or U8875 (N_8875,N_8201,N_8139);
or U8876 (N_8876,N_8355,N_8123);
nor U8877 (N_8877,N_8157,N_8062);
xnor U8878 (N_8878,N_8285,N_8069);
xnor U8879 (N_8879,N_8298,N_8246);
nor U8880 (N_8880,N_8196,N_8222);
or U8881 (N_8881,N_8065,N_8495);
nand U8882 (N_8882,N_8273,N_8417);
or U8883 (N_8883,N_8175,N_8117);
nand U8884 (N_8884,N_8418,N_8291);
xor U8885 (N_8885,N_8032,N_8199);
nor U8886 (N_8886,N_8023,N_8105);
and U8887 (N_8887,N_8300,N_8433);
xnor U8888 (N_8888,N_8016,N_8093);
and U8889 (N_8889,N_8227,N_8487);
or U8890 (N_8890,N_8424,N_8233);
or U8891 (N_8891,N_8415,N_8094);
xnor U8892 (N_8892,N_8350,N_8216);
or U8893 (N_8893,N_8311,N_8107);
or U8894 (N_8894,N_8342,N_8211);
nand U8895 (N_8895,N_8451,N_8263);
xor U8896 (N_8896,N_8026,N_8368);
xor U8897 (N_8897,N_8465,N_8058);
or U8898 (N_8898,N_8192,N_8149);
or U8899 (N_8899,N_8187,N_8361);
xor U8900 (N_8900,N_8357,N_8033);
nor U8901 (N_8901,N_8148,N_8466);
nand U8902 (N_8902,N_8185,N_8097);
nor U8903 (N_8903,N_8491,N_8251);
or U8904 (N_8904,N_8395,N_8409);
nand U8905 (N_8905,N_8143,N_8432);
nor U8906 (N_8906,N_8352,N_8202);
xor U8907 (N_8907,N_8014,N_8170);
nor U8908 (N_8908,N_8032,N_8066);
nor U8909 (N_8909,N_8442,N_8439);
or U8910 (N_8910,N_8130,N_8391);
nand U8911 (N_8911,N_8482,N_8167);
xor U8912 (N_8912,N_8274,N_8012);
and U8913 (N_8913,N_8158,N_8185);
xnor U8914 (N_8914,N_8446,N_8307);
nand U8915 (N_8915,N_8021,N_8193);
nand U8916 (N_8916,N_8046,N_8337);
nand U8917 (N_8917,N_8465,N_8228);
nand U8918 (N_8918,N_8213,N_8235);
or U8919 (N_8919,N_8270,N_8250);
xnor U8920 (N_8920,N_8342,N_8068);
and U8921 (N_8921,N_8487,N_8392);
xor U8922 (N_8922,N_8462,N_8130);
nand U8923 (N_8923,N_8385,N_8332);
nand U8924 (N_8924,N_8228,N_8149);
nand U8925 (N_8925,N_8023,N_8029);
nor U8926 (N_8926,N_8419,N_8005);
nand U8927 (N_8927,N_8185,N_8091);
and U8928 (N_8928,N_8455,N_8076);
or U8929 (N_8929,N_8494,N_8254);
and U8930 (N_8930,N_8253,N_8314);
nor U8931 (N_8931,N_8340,N_8035);
nand U8932 (N_8932,N_8131,N_8443);
and U8933 (N_8933,N_8102,N_8269);
and U8934 (N_8934,N_8257,N_8489);
xor U8935 (N_8935,N_8011,N_8329);
nor U8936 (N_8936,N_8409,N_8029);
nand U8937 (N_8937,N_8176,N_8395);
nand U8938 (N_8938,N_8010,N_8328);
and U8939 (N_8939,N_8352,N_8020);
nand U8940 (N_8940,N_8052,N_8275);
nor U8941 (N_8941,N_8490,N_8286);
and U8942 (N_8942,N_8406,N_8059);
xnor U8943 (N_8943,N_8052,N_8349);
xor U8944 (N_8944,N_8015,N_8004);
and U8945 (N_8945,N_8145,N_8440);
nand U8946 (N_8946,N_8357,N_8225);
nand U8947 (N_8947,N_8227,N_8270);
or U8948 (N_8948,N_8032,N_8361);
and U8949 (N_8949,N_8112,N_8042);
or U8950 (N_8950,N_8478,N_8268);
nand U8951 (N_8951,N_8276,N_8219);
or U8952 (N_8952,N_8464,N_8146);
nand U8953 (N_8953,N_8421,N_8370);
xnor U8954 (N_8954,N_8483,N_8203);
and U8955 (N_8955,N_8171,N_8239);
or U8956 (N_8956,N_8334,N_8393);
nand U8957 (N_8957,N_8462,N_8460);
nor U8958 (N_8958,N_8087,N_8273);
xor U8959 (N_8959,N_8094,N_8360);
xor U8960 (N_8960,N_8217,N_8388);
nor U8961 (N_8961,N_8118,N_8153);
and U8962 (N_8962,N_8442,N_8390);
and U8963 (N_8963,N_8000,N_8495);
and U8964 (N_8964,N_8229,N_8044);
nor U8965 (N_8965,N_8110,N_8401);
xnor U8966 (N_8966,N_8303,N_8350);
or U8967 (N_8967,N_8044,N_8190);
or U8968 (N_8968,N_8487,N_8337);
or U8969 (N_8969,N_8019,N_8112);
or U8970 (N_8970,N_8454,N_8437);
or U8971 (N_8971,N_8044,N_8025);
or U8972 (N_8972,N_8366,N_8193);
and U8973 (N_8973,N_8003,N_8055);
xor U8974 (N_8974,N_8426,N_8471);
xor U8975 (N_8975,N_8270,N_8173);
xnor U8976 (N_8976,N_8146,N_8024);
or U8977 (N_8977,N_8304,N_8236);
and U8978 (N_8978,N_8410,N_8372);
or U8979 (N_8979,N_8187,N_8011);
xor U8980 (N_8980,N_8018,N_8095);
and U8981 (N_8981,N_8222,N_8237);
nand U8982 (N_8982,N_8077,N_8419);
and U8983 (N_8983,N_8018,N_8290);
nand U8984 (N_8984,N_8427,N_8474);
nand U8985 (N_8985,N_8064,N_8393);
nor U8986 (N_8986,N_8040,N_8070);
xnor U8987 (N_8987,N_8277,N_8473);
and U8988 (N_8988,N_8234,N_8238);
and U8989 (N_8989,N_8318,N_8002);
or U8990 (N_8990,N_8092,N_8384);
xor U8991 (N_8991,N_8474,N_8385);
or U8992 (N_8992,N_8032,N_8413);
xor U8993 (N_8993,N_8412,N_8334);
or U8994 (N_8994,N_8082,N_8366);
or U8995 (N_8995,N_8439,N_8379);
and U8996 (N_8996,N_8183,N_8193);
nand U8997 (N_8997,N_8041,N_8432);
xor U8998 (N_8998,N_8030,N_8253);
or U8999 (N_8999,N_8168,N_8017);
or U9000 (N_9000,N_8686,N_8858);
nor U9001 (N_9001,N_8866,N_8553);
xor U9002 (N_9002,N_8533,N_8691);
nor U9003 (N_9003,N_8932,N_8685);
xor U9004 (N_9004,N_8623,N_8702);
or U9005 (N_9005,N_8895,N_8867);
xnor U9006 (N_9006,N_8819,N_8791);
xor U9007 (N_9007,N_8785,N_8899);
nand U9008 (N_9008,N_8645,N_8996);
and U9009 (N_9009,N_8667,N_8874);
xor U9010 (N_9010,N_8793,N_8949);
and U9011 (N_9011,N_8904,N_8954);
nor U9012 (N_9012,N_8711,N_8541);
or U9013 (N_9013,N_8739,N_8882);
nand U9014 (N_9014,N_8598,N_8896);
or U9015 (N_9015,N_8707,N_8901);
nor U9016 (N_9016,N_8751,N_8814);
nor U9017 (N_9017,N_8618,N_8688);
and U9018 (N_9018,N_8763,N_8734);
nor U9019 (N_9019,N_8738,N_8506);
nor U9020 (N_9020,N_8995,N_8872);
or U9021 (N_9021,N_8539,N_8526);
xor U9022 (N_9022,N_8997,N_8617);
nor U9023 (N_9023,N_8903,N_8717);
or U9024 (N_9024,N_8588,N_8730);
or U9025 (N_9025,N_8583,N_8608);
or U9026 (N_9026,N_8595,N_8562);
nand U9027 (N_9027,N_8829,N_8943);
or U9028 (N_9028,N_8891,N_8787);
nand U9029 (N_9029,N_8826,N_8985);
nor U9030 (N_9030,N_8663,N_8856);
nand U9031 (N_9031,N_8554,N_8710);
nor U9032 (N_9032,N_8646,N_8602);
or U9033 (N_9033,N_8757,N_8744);
nand U9034 (N_9034,N_8679,N_8536);
nor U9035 (N_9035,N_8655,N_8752);
nand U9036 (N_9036,N_8784,N_8596);
nor U9037 (N_9037,N_8869,N_8724);
nand U9038 (N_9038,N_8723,N_8687);
or U9039 (N_9039,N_8799,N_8962);
nor U9040 (N_9040,N_8756,N_8900);
and U9041 (N_9041,N_8511,N_8609);
nor U9042 (N_9042,N_8921,N_8574);
nand U9043 (N_9043,N_8518,N_8800);
nor U9044 (N_9044,N_8935,N_8589);
nand U9045 (N_9045,N_8516,N_8653);
or U9046 (N_9046,N_8525,N_8987);
and U9047 (N_9047,N_8853,N_8747);
or U9048 (N_9048,N_8925,N_8640);
nor U9049 (N_9049,N_8523,N_8778);
nor U9050 (N_9050,N_8549,N_8659);
nor U9051 (N_9051,N_8759,N_8825);
nor U9052 (N_9052,N_8934,N_8864);
and U9053 (N_9053,N_8822,N_8998);
or U9054 (N_9054,N_8887,N_8840);
or U9055 (N_9055,N_8704,N_8980);
nor U9056 (N_9056,N_8569,N_8681);
xor U9057 (N_9057,N_8776,N_8937);
and U9058 (N_9058,N_8851,N_8705);
xnor U9059 (N_9059,N_8753,N_8976);
nor U9060 (N_9060,N_8737,N_8794);
nor U9061 (N_9061,N_8818,N_8502);
xor U9062 (N_9062,N_8773,N_8999);
nor U9063 (N_9063,N_8931,N_8955);
nor U9064 (N_9064,N_8754,N_8939);
or U9065 (N_9065,N_8957,N_8764);
or U9066 (N_9066,N_8638,N_8585);
xnor U9067 (N_9067,N_8586,N_8577);
xor U9068 (N_9068,N_8918,N_8674);
or U9069 (N_9069,N_8876,N_8779);
xor U9070 (N_9070,N_8812,N_8917);
or U9071 (N_9071,N_8953,N_8660);
or U9072 (N_9072,N_8565,N_8593);
nor U9073 (N_9073,N_8571,N_8992);
nand U9074 (N_9074,N_8775,N_8677);
xor U9075 (N_9075,N_8678,N_8914);
xnor U9076 (N_9076,N_8733,N_8644);
xnor U9077 (N_9077,N_8969,N_8898);
and U9078 (N_9078,N_8993,N_8580);
xor U9079 (N_9079,N_8606,N_8546);
or U9080 (N_9080,N_8531,N_8944);
or U9081 (N_9081,N_8811,N_8718);
or U9082 (N_9082,N_8994,N_8620);
nor U9083 (N_9083,N_8802,N_8795);
nand U9084 (N_9084,N_8830,N_8971);
or U9085 (N_9085,N_8693,N_8855);
xnor U9086 (N_9086,N_8670,N_8651);
xnor U9087 (N_9087,N_8832,N_8634);
nand U9088 (N_9088,N_8770,N_8522);
xor U9089 (N_9089,N_8701,N_8766);
nor U9090 (N_9090,N_8948,N_8749);
and U9091 (N_9091,N_8888,N_8947);
or U9092 (N_9092,N_8956,N_8624);
xnor U9093 (N_9093,N_8870,N_8591);
or U9094 (N_9094,N_8871,N_8528);
xnor U9095 (N_9095,N_8614,N_8857);
and U9096 (N_9096,N_8719,N_8810);
and U9097 (N_9097,N_8605,N_8828);
xor U9098 (N_9098,N_8540,N_8792);
nor U9099 (N_9099,N_8515,N_8774);
or U9100 (N_9100,N_8748,N_8963);
nor U9101 (N_9101,N_8643,N_8781);
nand U9102 (N_9102,N_8862,N_8886);
nand U9103 (N_9103,N_8958,N_8804);
or U9104 (N_9104,N_8573,N_8849);
nor U9105 (N_9105,N_8637,N_8545);
nand U9106 (N_9106,N_8658,N_8767);
and U9107 (N_9107,N_8945,N_8988);
nand U9108 (N_9108,N_8788,N_8727);
or U9109 (N_9109,N_8661,N_8612);
and U9110 (N_9110,N_8893,N_8505);
or U9111 (N_9111,N_8880,N_8630);
or U9112 (N_9112,N_8669,N_8860);
and U9113 (N_9113,N_8504,N_8552);
or U9114 (N_9114,N_8649,N_8868);
nor U9115 (N_9115,N_8604,N_8510);
nor U9116 (N_9116,N_8514,N_8923);
nand U9117 (N_9117,N_8859,N_8885);
nand U9118 (N_9118,N_8557,N_8581);
and U9119 (N_9119,N_8501,N_8626);
xor U9120 (N_9120,N_8959,N_8877);
and U9121 (N_9121,N_8671,N_8991);
xnor U9122 (N_9122,N_8831,N_8902);
or U9123 (N_9123,N_8782,N_8594);
xor U9124 (N_9124,N_8534,N_8732);
and U9125 (N_9125,N_8797,N_8852);
xor U9126 (N_9126,N_8684,N_8507);
or U9127 (N_9127,N_8873,N_8850);
or U9128 (N_9128,N_8513,N_8970);
nor U9129 (N_9129,N_8524,N_8509);
or U9130 (N_9130,N_8750,N_8720);
or U9131 (N_9131,N_8879,N_8973);
nand U9132 (N_9132,N_8960,N_8807);
or U9133 (N_9133,N_8746,N_8911);
nor U9134 (N_9134,N_8913,N_8875);
or U9135 (N_9135,N_8616,N_8682);
and U9136 (N_9136,N_8735,N_8530);
xnor U9137 (N_9137,N_8535,N_8977);
nand U9138 (N_9138,N_8708,N_8668);
nor U9139 (N_9139,N_8548,N_8587);
nand U9140 (N_9140,N_8894,N_8713);
nor U9141 (N_9141,N_8647,N_8578);
or U9142 (N_9142,N_8865,N_8780);
nand U9143 (N_9143,N_8984,N_8847);
nand U9144 (N_9144,N_8582,N_8907);
xnor U9145 (N_9145,N_8758,N_8861);
xor U9146 (N_9146,N_8715,N_8599);
nand U9147 (N_9147,N_8801,N_8745);
nand U9148 (N_9148,N_8839,N_8783);
or U9149 (N_9149,N_8961,N_8611);
and U9150 (N_9150,N_8808,N_8560);
nor U9151 (N_9151,N_8619,N_8741);
xor U9152 (N_9152,N_8550,N_8521);
nand U9153 (N_9153,N_8978,N_8823);
xor U9154 (N_9154,N_8632,N_8680);
or U9155 (N_9155,N_8919,N_8964);
and U9156 (N_9156,N_8690,N_8639);
nand U9157 (N_9157,N_8817,N_8936);
nand U9158 (N_9158,N_8628,N_8940);
and U9159 (N_9159,N_8517,N_8706);
or U9160 (N_9160,N_8673,N_8728);
and U9161 (N_9161,N_8695,N_8740);
or U9162 (N_9162,N_8656,N_8665);
or U9163 (N_9163,N_8542,N_8983);
or U9164 (N_9164,N_8558,N_8743);
and U9165 (N_9165,N_8654,N_8790);
nor U9166 (N_9166,N_8567,N_8631);
xor U9167 (N_9167,N_8527,N_8884);
or U9168 (N_9168,N_8881,N_8897);
xor U9169 (N_9169,N_8846,N_8512);
xnor U9170 (N_9170,N_8863,N_8503);
or U9171 (N_9171,N_8555,N_8841);
and U9172 (N_9172,N_8716,N_8915);
and U9173 (N_9173,N_8538,N_8597);
xor U9174 (N_9174,N_8837,N_8974);
nor U9175 (N_9175,N_8508,N_8979);
xnor U9176 (N_9176,N_8803,N_8551);
nor U9177 (N_9177,N_8603,N_8777);
and U9178 (N_9178,N_8615,N_8951);
and U9179 (N_9179,N_8607,N_8579);
nor U9180 (N_9180,N_8700,N_8601);
or U9181 (N_9181,N_8543,N_8968);
and U9182 (N_9182,N_8889,N_8952);
or U9183 (N_9183,N_8666,N_8928);
or U9184 (N_9184,N_8664,N_8650);
xnor U9185 (N_9185,N_8835,N_8838);
or U9186 (N_9186,N_8786,N_8815);
xor U9187 (N_9187,N_8762,N_8627);
or U9188 (N_9188,N_8721,N_8547);
xnor U9189 (N_9189,N_8709,N_8692);
and U9190 (N_9190,N_8641,N_8566);
nand U9191 (N_9191,N_8683,N_8584);
nand U9192 (N_9192,N_8629,N_8848);
or U9193 (N_9193,N_8929,N_8648);
xor U9194 (N_9194,N_8910,N_8761);
or U9195 (N_9195,N_8712,N_8714);
nor U9196 (N_9196,N_8564,N_8878);
nor U9197 (N_9197,N_8845,N_8883);
nor U9198 (N_9198,N_8622,N_8676);
xnor U9199 (N_9199,N_8909,N_8689);
nand U9200 (N_9200,N_8729,N_8736);
nand U9201 (N_9201,N_8834,N_8742);
or U9202 (N_9202,N_8576,N_8570);
nand U9203 (N_9203,N_8559,N_8908);
nor U9204 (N_9204,N_8642,N_8854);
or U9205 (N_9205,N_8967,N_8771);
nor U9206 (N_9206,N_8575,N_8662);
nor U9207 (N_9207,N_8768,N_8906);
or U9208 (N_9208,N_8699,N_8916);
and U9209 (N_9209,N_8905,N_8697);
nand U9210 (N_9210,N_8544,N_8989);
xnor U9211 (N_9211,N_8942,N_8765);
nor U9212 (N_9212,N_8990,N_8590);
or U9213 (N_9213,N_8805,N_8563);
and U9214 (N_9214,N_8636,N_8813);
nor U9215 (N_9215,N_8843,N_8827);
or U9216 (N_9216,N_8625,N_8572);
xnor U9217 (N_9217,N_8927,N_8892);
nand U9218 (N_9218,N_8672,N_8966);
xor U9219 (N_9219,N_8796,N_8798);
xor U9220 (N_9220,N_8613,N_8890);
or U9221 (N_9221,N_8920,N_8789);
xor U9222 (N_9222,N_8696,N_8930);
and U9223 (N_9223,N_8760,N_8694);
and U9224 (N_9224,N_8657,N_8844);
nor U9225 (N_9225,N_8926,N_8982);
or U9226 (N_9226,N_8675,N_8772);
and U9227 (N_9227,N_8635,N_8769);
xnor U9228 (N_9228,N_8725,N_8698);
xor U9229 (N_9229,N_8529,N_8821);
xnor U9230 (N_9230,N_8731,N_8924);
or U9231 (N_9231,N_8520,N_8519);
and U9232 (N_9232,N_8532,N_8922);
or U9233 (N_9233,N_8633,N_8500);
or U9234 (N_9234,N_8975,N_8556);
nor U9235 (N_9235,N_8561,N_8703);
nor U9236 (N_9236,N_8972,N_8950);
or U9237 (N_9237,N_8965,N_8600);
nand U9238 (N_9238,N_8652,N_8592);
nor U9239 (N_9239,N_8537,N_8621);
or U9240 (N_9240,N_8824,N_8809);
and U9241 (N_9241,N_8820,N_8836);
nor U9242 (N_9242,N_8568,N_8842);
nand U9243 (N_9243,N_8833,N_8986);
and U9244 (N_9244,N_8941,N_8755);
or U9245 (N_9245,N_8726,N_8610);
nor U9246 (N_9246,N_8946,N_8912);
xor U9247 (N_9247,N_8981,N_8806);
nor U9248 (N_9248,N_8816,N_8938);
nor U9249 (N_9249,N_8933,N_8722);
nor U9250 (N_9250,N_8834,N_8877);
nand U9251 (N_9251,N_8868,N_8621);
nor U9252 (N_9252,N_8966,N_8571);
nor U9253 (N_9253,N_8542,N_8969);
and U9254 (N_9254,N_8724,N_8646);
xor U9255 (N_9255,N_8614,N_8680);
or U9256 (N_9256,N_8855,N_8902);
and U9257 (N_9257,N_8926,N_8653);
nand U9258 (N_9258,N_8730,N_8761);
nand U9259 (N_9259,N_8885,N_8557);
and U9260 (N_9260,N_8648,N_8844);
or U9261 (N_9261,N_8613,N_8757);
nand U9262 (N_9262,N_8882,N_8912);
nand U9263 (N_9263,N_8794,N_8875);
nor U9264 (N_9264,N_8901,N_8900);
and U9265 (N_9265,N_8771,N_8648);
nand U9266 (N_9266,N_8622,N_8860);
and U9267 (N_9267,N_8585,N_8827);
nor U9268 (N_9268,N_8987,N_8557);
or U9269 (N_9269,N_8733,N_8851);
xor U9270 (N_9270,N_8863,N_8805);
xor U9271 (N_9271,N_8624,N_8577);
xnor U9272 (N_9272,N_8568,N_8864);
or U9273 (N_9273,N_8906,N_8520);
xor U9274 (N_9274,N_8967,N_8910);
or U9275 (N_9275,N_8715,N_8511);
nor U9276 (N_9276,N_8506,N_8805);
nand U9277 (N_9277,N_8533,N_8948);
nand U9278 (N_9278,N_8884,N_8559);
nand U9279 (N_9279,N_8952,N_8687);
xnor U9280 (N_9280,N_8571,N_8844);
nor U9281 (N_9281,N_8854,N_8861);
or U9282 (N_9282,N_8505,N_8626);
xnor U9283 (N_9283,N_8998,N_8872);
nor U9284 (N_9284,N_8516,N_8915);
nor U9285 (N_9285,N_8963,N_8874);
xnor U9286 (N_9286,N_8826,N_8739);
nand U9287 (N_9287,N_8578,N_8742);
nor U9288 (N_9288,N_8925,N_8603);
or U9289 (N_9289,N_8657,N_8857);
xnor U9290 (N_9290,N_8870,N_8806);
nand U9291 (N_9291,N_8609,N_8809);
xor U9292 (N_9292,N_8726,N_8901);
and U9293 (N_9293,N_8796,N_8810);
nor U9294 (N_9294,N_8884,N_8724);
or U9295 (N_9295,N_8538,N_8887);
nor U9296 (N_9296,N_8691,N_8886);
xor U9297 (N_9297,N_8709,N_8929);
and U9298 (N_9298,N_8565,N_8850);
nor U9299 (N_9299,N_8554,N_8763);
xor U9300 (N_9300,N_8913,N_8567);
or U9301 (N_9301,N_8597,N_8537);
nor U9302 (N_9302,N_8538,N_8748);
and U9303 (N_9303,N_8682,N_8983);
or U9304 (N_9304,N_8796,N_8686);
nand U9305 (N_9305,N_8639,N_8623);
or U9306 (N_9306,N_8775,N_8792);
nand U9307 (N_9307,N_8972,N_8802);
nor U9308 (N_9308,N_8624,N_8873);
and U9309 (N_9309,N_8691,N_8831);
and U9310 (N_9310,N_8753,N_8522);
and U9311 (N_9311,N_8902,N_8593);
nand U9312 (N_9312,N_8798,N_8780);
nor U9313 (N_9313,N_8996,N_8823);
xor U9314 (N_9314,N_8566,N_8873);
xor U9315 (N_9315,N_8651,N_8709);
nand U9316 (N_9316,N_8734,N_8620);
nor U9317 (N_9317,N_8750,N_8600);
nor U9318 (N_9318,N_8789,N_8924);
or U9319 (N_9319,N_8681,N_8747);
nand U9320 (N_9320,N_8623,N_8937);
nor U9321 (N_9321,N_8804,N_8747);
nor U9322 (N_9322,N_8977,N_8529);
nor U9323 (N_9323,N_8911,N_8653);
nor U9324 (N_9324,N_8692,N_8787);
or U9325 (N_9325,N_8868,N_8808);
nand U9326 (N_9326,N_8927,N_8940);
nand U9327 (N_9327,N_8681,N_8955);
xnor U9328 (N_9328,N_8513,N_8521);
and U9329 (N_9329,N_8683,N_8563);
nand U9330 (N_9330,N_8860,N_8868);
nand U9331 (N_9331,N_8551,N_8720);
nor U9332 (N_9332,N_8643,N_8924);
or U9333 (N_9333,N_8671,N_8848);
or U9334 (N_9334,N_8960,N_8788);
nand U9335 (N_9335,N_8660,N_8514);
or U9336 (N_9336,N_8649,N_8516);
nor U9337 (N_9337,N_8932,N_8955);
and U9338 (N_9338,N_8558,N_8965);
or U9339 (N_9339,N_8529,N_8759);
nor U9340 (N_9340,N_8879,N_8963);
or U9341 (N_9341,N_8878,N_8932);
and U9342 (N_9342,N_8745,N_8864);
nor U9343 (N_9343,N_8839,N_8500);
xnor U9344 (N_9344,N_8929,N_8710);
nor U9345 (N_9345,N_8544,N_8889);
or U9346 (N_9346,N_8687,N_8680);
and U9347 (N_9347,N_8801,N_8655);
nor U9348 (N_9348,N_8704,N_8701);
and U9349 (N_9349,N_8550,N_8995);
nand U9350 (N_9350,N_8604,N_8621);
or U9351 (N_9351,N_8589,N_8607);
and U9352 (N_9352,N_8871,N_8706);
nor U9353 (N_9353,N_8714,N_8897);
xor U9354 (N_9354,N_8788,N_8984);
xor U9355 (N_9355,N_8678,N_8764);
nand U9356 (N_9356,N_8645,N_8934);
or U9357 (N_9357,N_8621,N_8609);
nor U9358 (N_9358,N_8668,N_8771);
xnor U9359 (N_9359,N_8999,N_8983);
nor U9360 (N_9360,N_8594,N_8995);
nand U9361 (N_9361,N_8680,N_8781);
and U9362 (N_9362,N_8722,N_8961);
nor U9363 (N_9363,N_8564,N_8735);
nor U9364 (N_9364,N_8996,N_8684);
nor U9365 (N_9365,N_8554,N_8917);
or U9366 (N_9366,N_8962,N_8501);
nand U9367 (N_9367,N_8933,N_8839);
nand U9368 (N_9368,N_8619,N_8902);
nor U9369 (N_9369,N_8860,N_8921);
nor U9370 (N_9370,N_8684,N_8665);
nand U9371 (N_9371,N_8831,N_8542);
nand U9372 (N_9372,N_8856,N_8684);
nor U9373 (N_9373,N_8650,N_8913);
and U9374 (N_9374,N_8738,N_8704);
xor U9375 (N_9375,N_8772,N_8868);
nand U9376 (N_9376,N_8569,N_8844);
nand U9377 (N_9377,N_8824,N_8855);
or U9378 (N_9378,N_8856,N_8816);
nand U9379 (N_9379,N_8659,N_8748);
nand U9380 (N_9380,N_8875,N_8788);
xnor U9381 (N_9381,N_8818,N_8519);
nor U9382 (N_9382,N_8629,N_8890);
nand U9383 (N_9383,N_8634,N_8899);
or U9384 (N_9384,N_8972,N_8821);
or U9385 (N_9385,N_8673,N_8830);
or U9386 (N_9386,N_8860,N_8832);
or U9387 (N_9387,N_8791,N_8661);
or U9388 (N_9388,N_8742,N_8822);
nor U9389 (N_9389,N_8500,N_8828);
and U9390 (N_9390,N_8612,N_8539);
xnor U9391 (N_9391,N_8611,N_8579);
or U9392 (N_9392,N_8686,N_8549);
nand U9393 (N_9393,N_8704,N_8877);
or U9394 (N_9394,N_8919,N_8552);
xor U9395 (N_9395,N_8622,N_8728);
or U9396 (N_9396,N_8566,N_8653);
xor U9397 (N_9397,N_8660,N_8523);
xor U9398 (N_9398,N_8722,N_8905);
nor U9399 (N_9399,N_8593,N_8520);
xnor U9400 (N_9400,N_8841,N_8540);
or U9401 (N_9401,N_8774,N_8500);
or U9402 (N_9402,N_8674,N_8801);
nor U9403 (N_9403,N_8648,N_8646);
nor U9404 (N_9404,N_8992,N_8706);
and U9405 (N_9405,N_8786,N_8930);
xnor U9406 (N_9406,N_8709,N_8525);
nor U9407 (N_9407,N_8575,N_8625);
xnor U9408 (N_9408,N_8536,N_8657);
xor U9409 (N_9409,N_8672,N_8905);
or U9410 (N_9410,N_8649,N_8976);
nand U9411 (N_9411,N_8517,N_8962);
nand U9412 (N_9412,N_8580,N_8682);
nand U9413 (N_9413,N_8990,N_8584);
or U9414 (N_9414,N_8778,N_8892);
xor U9415 (N_9415,N_8517,N_8653);
xor U9416 (N_9416,N_8852,N_8923);
nand U9417 (N_9417,N_8847,N_8889);
nand U9418 (N_9418,N_8801,N_8500);
or U9419 (N_9419,N_8864,N_8737);
nand U9420 (N_9420,N_8659,N_8506);
xor U9421 (N_9421,N_8744,N_8543);
nand U9422 (N_9422,N_8551,N_8728);
nand U9423 (N_9423,N_8791,N_8548);
xnor U9424 (N_9424,N_8661,N_8861);
and U9425 (N_9425,N_8950,N_8948);
nand U9426 (N_9426,N_8615,N_8691);
or U9427 (N_9427,N_8804,N_8765);
and U9428 (N_9428,N_8639,N_8763);
or U9429 (N_9429,N_8692,N_8888);
nor U9430 (N_9430,N_8541,N_8768);
and U9431 (N_9431,N_8502,N_8826);
xor U9432 (N_9432,N_8967,N_8693);
xor U9433 (N_9433,N_8595,N_8643);
or U9434 (N_9434,N_8686,N_8799);
nand U9435 (N_9435,N_8598,N_8532);
and U9436 (N_9436,N_8970,N_8980);
and U9437 (N_9437,N_8724,N_8726);
nor U9438 (N_9438,N_8647,N_8876);
and U9439 (N_9439,N_8770,N_8734);
nand U9440 (N_9440,N_8962,N_8665);
nand U9441 (N_9441,N_8564,N_8593);
xnor U9442 (N_9442,N_8960,N_8945);
or U9443 (N_9443,N_8743,N_8519);
or U9444 (N_9444,N_8836,N_8563);
or U9445 (N_9445,N_8951,N_8754);
and U9446 (N_9446,N_8879,N_8816);
nor U9447 (N_9447,N_8594,N_8870);
nand U9448 (N_9448,N_8518,N_8634);
or U9449 (N_9449,N_8979,N_8501);
nand U9450 (N_9450,N_8761,N_8736);
nor U9451 (N_9451,N_8962,N_8908);
or U9452 (N_9452,N_8722,N_8767);
nand U9453 (N_9453,N_8703,N_8850);
nor U9454 (N_9454,N_8761,N_8704);
or U9455 (N_9455,N_8926,N_8589);
xor U9456 (N_9456,N_8508,N_8924);
nand U9457 (N_9457,N_8991,N_8579);
nand U9458 (N_9458,N_8566,N_8703);
and U9459 (N_9459,N_8767,N_8696);
xnor U9460 (N_9460,N_8773,N_8890);
nor U9461 (N_9461,N_8859,N_8708);
xor U9462 (N_9462,N_8983,N_8926);
xnor U9463 (N_9463,N_8953,N_8781);
xor U9464 (N_9464,N_8535,N_8518);
or U9465 (N_9465,N_8503,N_8690);
nor U9466 (N_9466,N_8984,N_8590);
xor U9467 (N_9467,N_8560,N_8754);
and U9468 (N_9468,N_8685,N_8974);
or U9469 (N_9469,N_8580,N_8664);
nor U9470 (N_9470,N_8546,N_8927);
nor U9471 (N_9471,N_8973,N_8535);
xnor U9472 (N_9472,N_8575,N_8842);
or U9473 (N_9473,N_8608,N_8763);
or U9474 (N_9474,N_8781,N_8815);
xnor U9475 (N_9475,N_8766,N_8782);
or U9476 (N_9476,N_8891,N_8522);
or U9477 (N_9477,N_8922,N_8888);
and U9478 (N_9478,N_8634,N_8607);
xor U9479 (N_9479,N_8528,N_8800);
or U9480 (N_9480,N_8833,N_8624);
and U9481 (N_9481,N_8919,N_8740);
nor U9482 (N_9482,N_8601,N_8798);
nand U9483 (N_9483,N_8906,N_8516);
and U9484 (N_9484,N_8642,N_8518);
nor U9485 (N_9485,N_8509,N_8757);
or U9486 (N_9486,N_8846,N_8681);
nand U9487 (N_9487,N_8788,N_8822);
nor U9488 (N_9488,N_8680,N_8650);
and U9489 (N_9489,N_8978,N_8684);
and U9490 (N_9490,N_8961,N_8917);
nand U9491 (N_9491,N_8526,N_8802);
or U9492 (N_9492,N_8902,N_8865);
nand U9493 (N_9493,N_8583,N_8965);
xnor U9494 (N_9494,N_8705,N_8814);
nor U9495 (N_9495,N_8858,N_8890);
nand U9496 (N_9496,N_8679,N_8902);
nand U9497 (N_9497,N_8592,N_8710);
nor U9498 (N_9498,N_8736,N_8707);
nor U9499 (N_9499,N_8989,N_8820);
nor U9500 (N_9500,N_9407,N_9174);
xnor U9501 (N_9501,N_9498,N_9078);
nand U9502 (N_9502,N_9343,N_9454);
nand U9503 (N_9503,N_9120,N_9374);
xnor U9504 (N_9504,N_9182,N_9023);
and U9505 (N_9505,N_9497,N_9322);
and U9506 (N_9506,N_9496,N_9068);
nor U9507 (N_9507,N_9259,N_9226);
or U9508 (N_9508,N_9082,N_9196);
nor U9509 (N_9509,N_9117,N_9282);
or U9510 (N_9510,N_9064,N_9314);
or U9511 (N_9511,N_9048,N_9331);
xnor U9512 (N_9512,N_9440,N_9188);
nand U9513 (N_9513,N_9403,N_9281);
nand U9514 (N_9514,N_9084,N_9180);
nor U9515 (N_9515,N_9236,N_9336);
and U9516 (N_9516,N_9489,N_9161);
nor U9517 (N_9517,N_9195,N_9347);
or U9518 (N_9518,N_9304,N_9032);
nor U9519 (N_9519,N_9411,N_9003);
nor U9520 (N_9520,N_9235,N_9192);
and U9521 (N_9521,N_9387,N_9360);
xor U9522 (N_9522,N_9193,N_9044);
xor U9523 (N_9523,N_9391,N_9104);
and U9524 (N_9524,N_9455,N_9019);
and U9525 (N_9525,N_9465,N_9178);
nand U9526 (N_9526,N_9423,N_9184);
xor U9527 (N_9527,N_9299,N_9495);
nor U9528 (N_9528,N_9200,N_9037);
nand U9529 (N_9529,N_9397,N_9421);
xnor U9530 (N_9530,N_9324,N_9316);
xor U9531 (N_9531,N_9031,N_9116);
and U9532 (N_9532,N_9043,N_9434);
nor U9533 (N_9533,N_9464,N_9112);
nor U9534 (N_9534,N_9271,N_9400);
nand U9535 (N_9535,N_9306,N_9352);
xnor U9536 (N_9536,N_9435,N_9460);
xnor U9537 (N_9537,N_9227,N_9254);
or U9538 (N_9538,N_9444,N_9327);
nor U9539 (N_9539,N_9097,N_9144);
nor U9540 (N_9540,N_9012,N_9377);
xor U9541 (N_9541,N_9284,N_9127);
xnor U9542 (N_9542,N_9494,N_9008);
nand U9543 (N_9543,N_9147,N_9416);
or U9544 (N_9544,N_9344,N_9118);
nand U9545 (N_9545,N_9020,N_9279);
or U9546 (N_9546,N_9171,N_9207);
nand U9547 (N_9547,N_9109,N_9459);
nor U9548 (N_9548,N_9476,N_9475);
xor U9549 (N_9549,N_9402,N_9436);
nand U9550 (N_9550,N_9212,N_9057);
or U9551 (N_9551,N_9468,N_9348);
nand U9552 (N_9552,N_9208,N_9231);
or U9553 (N_9553,N_9055,N_9265);
nand U9554 (N_9554,N_9490,N_9315);
xnor U9555 (N_9555,N_9009,N_9292);
xnor U9556 (N_9556,N_9042,N_9443);
xor U9557 (N_9557,N_9240,N_9221);
xor U9558 (N_9558,N_9015,N_9309);
and U9559 (N_9559,N_9272,N_9007);
or U9560 (N_9560,N_9482,N_9145);
and U9561 (N_9561,N_9040,N_9075);
nand U9562 (N_9562,N_9228,N_9214);
nor U9563 (N_9563,N_9164,N_9383);
or U9564 (N_9564,N_9080,N_9130);
and U9565 (N_9565,N_9349,N_9312);
nor U9566 (N_9566,N_9341,N_9270);
nor U9567 (N_9567,N_9225,N_9237);
or U9568 (N_9568,N_9014,N_9373);
and U9569 (N_9569,N_9095,N_9318);
and U9570 (N_9570,N_9337,N_9473);
or U9571 (N_9571,N_9308,N_9026);
and U9572 (N_9572,N_9480,N_9293);
nand U9573 (N_9573,N_9388,N_9364);
or U9574 (N_9574,N_9217,N_9071);
xor U9575 (N_9575,N_9438,N_9142);
xnor U9576 (N_9576,N_9356,N_9307);
xnor U9577 (N_9577,N_9257,N_9245);
and U9578 (N_9578,N_9155,N_9431);
or U9579 (N_9579,N_9415,N_9456);
or U9580 (N_9580,N_9479,N_9437);
or U9581 (N_9581,N_9441,N_9050);
or U9582 (N_9582,N_9390,N_9338);
and U9583 (N_9583,N_9162,N_9099);
or U9584 (N_9584,N_9215,N_9005);
xor U9585 (N_9585,N_9041,N_9061);
nand U9586 (N_9586,N_9260,N_9385);
nor U9587 (N_9587,N_9426,N_9205);
or U9588 (N_9588,N_9133,N_9105);
and U9589 (N_9589,N_9072,N_9010);
nand U9590 (N_9590,N_9246,N_9034);
nor U9591 (N_9591,N_9286,N_9499);
xor U9592 (N_9592,N_9412,N_9076);
nor U9593 (N_9593,N_9179,N_9484);
xnor U9594 (N_9594,N_9273,N_9368);
xnor U9595 (N_9595,N_9362,N_9108);
and U9596 (N_9596,N_9168,N_9156);
nor U9597 (N_9597,N_9267,N_9425);
nor U9598 (N_9598,N_9128,N_9277);
nand U9599 (N_9599,N_9124,N_9285);
nor U9600 (N_9600,N_9485,N_9258);
xor U9601 (N_9601,N_9220,N_9126);
nor U9602 (N_9602,N_9107,N_9492);
and U9603 (N_9603,N_9319,N_9363);
or U9604 (N_9604,N_9021,N_9332);
nor U9605 (N_9605,N_9393,N_9091);
and U9606 (N_9606,N_9035,N_9414);
and U9607 (N_9607,N_9409,N_9086);
xor U9608 (N_9608,N_9030,N_9089);
xor U9609 (N_9609,N_9340,N_9289);
and U9610 (N_9610,N_9418,N_9298);
and U9611 (N_9611,N_9115,N_9244);
or U9612 (N_9612,N_9300,N_9189);
nand U9613 (N_9613,N_9102,N_9398);
xor U9614 (N_9614,N_9323,N_9313);
nor U9615 (N_9615,N_9394,N_9382);
xor U9616 (N_9616,N_9370,N_9052);
xnor U9617 (N_9617,N_9024,N_9269);
nor U9618 (N_9618,N_9125,N_9432);
xnor U9619 (N_9619,N_9039,N_9392);
nor U9620 (N_9620,N_9381,N_9063);
and U9621 (N_9621,N_9305,N_9478);
and U9622 (N_9622,N_9069,N_9384);
and U9623 (N_9623,N_9399,N_9266);
and U9624 (N_9624,N_9136,N_9185);
and U9625 (N_9625,N_9442,N_9430);
and U9626 (N_9626,N_9371,N_9458);
nand U9627 (N_9627,N_9051,N_9379);
nor U9628 (N_9628,N_9066,N_9328);
xnor U9629 (N_9629,N_9433,N_9467);
nand U9630 (N_9630,N_9049,N_9187);
or U9631 (N_9631,N_9481,N_9294);
nor U9632 (N_9632,N_9335,N_9198);
and U9633 (N_9633,N_9138,N_9181);
xor U9634 (N_9634,N_9297,N_9166);
nor U9635 (N_9635,N_9022,N_9210);
nand U9636 (N_9636,N_9167,N_9047);
nand U9637 (N_9637,N_9491,N_9346);
nor U9638 (N_9638,N_9074,N_9404);
and U9639 (N_9639,N_9038,N_9175);
xor U9640 (N_9640,N_9268,N_9204);
or U9641 (N_9641,N_9263,N_9280);
nand U9642 (N_9642,N_9369,N_9470);
nor U9643 (N_9643,N_9046,N_9229);
nor U9644 (N_9644,N_9083,N_9143);
and U9645 (N_9645,N_9165,N_9410);
and U9646 (N_9646,N_9354,N_9334);
or U9647 (N_9647,N_9296,N_9248);
nor U9648 (N_9648,N_9088,N_9422);
nor U9649 (N_9649,N_9222,N_9058);
nand U9650 (N_9650,N_9065,N_9123);
and U9651 (N_9651,N_9100,N_9113);
nor U9652 (N_9652,N_9350,N_9002);
and U9653 (N_9653,N_9070,N_9213);
nand U9654 (N_9654,N_9028,N_9081);
or U9655 (N_9655,N_9252,N_9001);
xor U9656 (N_9656,N_9311,N_9325);
or U9657 (N_9657,N_9018,N_9176);
xnor U9658 (N_9658,N_9408,N_9253);
and U9659 (N_9659,N_9446,N_9146);
nor U9660 (N_9660,N_9448,N_9357);
or U9661 (N_9661,N_9172,N_9461);
nand U9662 (N_9662,N_9288,N_9054);
nor U9663 (N_9663,N_9477,N_9199);
nor U9664 (N_9664,N_9139,N_9339);
xnor U9665 (N_9665,N_9211,N_9278);
nand U9666 (N_9666,N_9255,N_9276);
nand U9667 (N_9667,N_9420,N_9365);
nand U9668 (N_9668,N_9361,N_9085);
nor U9669 (N_9669,N_9098,N_9463);
or U9670 (N_9670,N_9209,N_9424);
or U9671 (N_9671,N_9110,N_9151);
nor U9672 (N_9672,N_9094,N_9449);
xnor U9673 (N_9673,N_9141,N_9380);
nand U9674 (N_9674,N_9186,N_9234);
nor U9675 (N_9675,N_9216,N_9000);
and U9676 (N_9676,N_9493,N_9367);
and U9677 (N_9677,N_9111,N_9129);
nor U9678 (N_9678,N_9487,N_9386);
xnor U9679 (N_9679,N_9247,N_9359);
xnor U9680 (N_9680,N_9376,N_9153);
xor U9681 (N_9681,N_9148,N_9004);
xnor U9682 (N_9682,N_9201,N_9079);
nand U9683 (N_9683,N_9450,N_9158);
xnor U9684 (N_9684,N_9342,N_9103);
nor U9685 (N_9685,N_9011,N_9087);
nand U9686 (N_9686,N_9053,N_9451);
and U9687 (N_9687,N_9017,N_9233);
and U9688 (N_9688,N_9378,N_9239);
nor U9689 (N_9689,N_9223,N_9483);
nor U9690 (N_9690,N_9372,N_9013);
xnor U9691 (N_9691,N_9466,N_9149);
nand U9692 (N_9692,N_9029,N_9194);
nand U9693 (N_9693,N_9036,N_9241);
or U9694 (N_9694,N_9238,N_9132);
nor U9695 (N_9695,N_9092,N_9206);
or U9696 (N_9696,N_9152,N_9474);
and U9697 (N_9697,N_9469,N_9366);
and U9698 (N_9698,N_9303,N_9405);
nand U9699 (N_9699,N_9067,N_9389);
and U9700 (N_9700,N_9106,N_9330);
nor U9701 (N_9701,N_9375,N_9261);
nand U9702 (N_9702,N_9159,N_9060);
or U9703 (N_9703,N_9163,N_9170);
nor U9704 (N_9704,N_9232,N_9096);
or U9705 (N_9705,N_9250,N_9025);
or U9706 (N_9706,N_9134,N_9452);
and U9707 (N_9707,N_9287,N_9290);
nor U9708 (N_9708,N_9256,N_9101);
xor U9709 (N_9709,N_9056,N_9471);
nand U9710 (N_9710,N_9321,N_9291);
or U9711 (N_9711,N_9150,N_9295);
nor U9712 (N_9712,N_9006,N_9242);
or U9713 (N_9713,N_9154,N_9413);
or U9714 (N_9714,N_9447,N_9401);
nor U9715 (N_9715,N_9251,N_9302);
xor U9716 (N_9716,N_9301,N_9355);
xnor U9717 (N_9717,N_9218,N_9027);
xnor U9718 (N_9718,N_9090,N_9274);
and U9719 (N_9719,N_9062,N_9077);
or U9720 (N_9720,N_9429,N_9283);
and U9721 (N_9721,N_9121,N_9173);
and U9722 (N_9722,N_9045,N_9457);
or U9723 (N_9723,N_9310,N_9395);
and U9724 (N_9724,N_9140,N_9243);
xnor U9725 (N_9725,N_9224,N_9275);
xnor U9726 (N_9726,N_9428,N_9329);
xnor U9727 (N_9727,N_9183,N_9135);
nor U9728 (N_9728,N_9445,N_9262);
xor U9729 (N_9729,N_9190,N_9326);
and U9730 (N_9730,N_9230,N_9093);
xor U9731 (N_9731,N_9320,N_9119);
nor U9732 (N_9732,N_9203,N_9333);
xor U9733 (N_9733,N_9317,N_9177);
nand U9734 (N_9734,N_9114,N_9345);
nand U9735 (N_9735,N_9358,N_9439);
nand U9736 (N_9736,N_9419,N_9249);
xor U9737 (N_9737,N_9202,N_9406);
xor U9738 (N_9738,N_9462,N_9488);
nand U9739 (N_9739,N_9122,N_9191);
and U9740 (N_9740,N_9157,N_9264);
or U9741 (N_9741,N_9453,N_9016);
and U9742 (N_9742,N_9197,N_9219);
nand U9743 (N_9743,N_9486,N_9353);
and U9744 (N_9744,N_9131,N_9137);
nor U9745 (N_9745,N_9427,N_9472);
nand U9746 (N_9746,N_9033,N_9059);
and U9747 (N_9747,N_9417,N_9169);
nand U9748 (N_9748,N_9073,N_9396);
nand U9749 (N_9749,N_9160,N_9351);
and U9750 (N_9750,N_9397,N_9193);
nand U9751 (N_9751,N_9482,N_9339);
nand U9752 (N_9752,N_9350,N_9481);
or U9753 (N_9753,N_9034,N_9256);
nor U9754 (N_9754,N_9069,N_9446);
xnor U9755 (N_9755,N_9031,N_9419);
nor U9756 (N_9756,N_9001,N_9040);
xnor U9757 (N_9757,N_9161,N_9201);
nor U9758 (N_9758,N_9240,N_9346);
and U9759 (N_9759,N_9275,N_9390);
nor U9760 (N_9760,N_9490,N_9332);
or U9761 (N_9761,N_9139,N_9248);
nand U9762 (N_9762,N_9183,N_9051);
or U9763 (N_9763,N_9142,N_9333);
nor U9764 (N_9764,N_9156,N_9466);
nor U9765 (N_9765,N_9267,N_9187);
nor U9766 (N_9766,N_9043,N_9373);
xnor U9767 (N_9767,N_9230,N_9205);
nand U9768 (N_9768,N_9340,N_9328);
xor U9769 (N_9769,N_9267,N_9089);
nand U9770 (N_9770,N_9180,N_9128);
xor U9771 (N_9771,N_9254,N_9114);
nand U9772 (N_9772,N_9455,N_9028);
nand U9773 (N_9773,N_9475,N_9298);
nor U9774 (N_9774,N_9143,N_9283);
or U9775 (N_9775,N_9013,N_9057);
and U9776 (N_9776,N_9005,N_9457);
xnor U9777 (N_9777,N_9389,N_9279);
nor U9778 (N_9778,N_9408,N_9031);
and U9779 (N_9779,N_9177,N_9008);
nand U9780 (N_9780,N_9312,N_9329);
nor U9781 (N_9781,N_9436,N_9478);
or U9782 (N_9782,N_9101,N_9234);
xnor U9783 (N_9783,N_9470,N_9297);
and U9784 (N_9784,N_9273,N_9098);
nand U9785 (N_9785,N_9444,N_9209);
xnor U9786 (N_9786,N_9361,N_9401);
nor U9787 (N_9787,N_9462,N_9458);
xor U9788 (N_9788,N_9482,N_9479);
nand U9789 (N_9789,N_9321,N_9246);
or U9790 (N_9790,N_9239,N_9284);
or U9791 (N_9791,N_9460,N_9088);
xnor U9792 (N_9792,N_9115,N_9438);
xnor U9793 (N_9793,N_9142,N_9362);
and U9794 (N_9794,N_9307,N_9054);
nor U9795 (N_9795,N_9201,N_9210);
or U9796 (N_9796,N_9021,N_9230);
or U9797 (N_9797,N_9233,N_9129);
and U9798 (N_9798,N_9474,N_9084);
nor U9799 (N_9799,N_9195,N_9488);
xnor U9800 (N_9800,N_9434,N_9288);
xor U9801 (N_9801,N_9413,N_9220);
nor U9802 (N_9802,N_9295,N_9170);
or U9803 (N_9803,N_9182,N_9383);
nand U9804 (N_9804,N_9373,N_9188);
or U9805 (N_9805,N_9488,N_9414);
nor U9806 (N_9806,N_9218,N_9115);
xnor U9807 (N_9807,N_9143,N_9432);
nand U9808 (N_9808,N_9226,N_9008);
xnor U9809 (N_9809,N_9224,N_9340);
and U9810 (N_9810,N_9323,N_9225);
nor U9811 (N_9811,N_9164,N_9460);
nand U9812 (N_9812,N_9344,N_9496);
and U9813 (N_9813,N_9368,N_9190);
xnor U9814 (N_9814,N_9318,N_9130);
and U9815 (N_9815,N_9473,N_9087);
xnor U9816 (N_9816,N_9054,N_9353);
or U9817 (N_9817,N_9423,N_9414);
or U9818 (N_9818,N_9419,N_9193);
nor U9819 (N_9819,N_9249,N_9038);
nand U9820 (N_9820,N_9017,N_9369);
nand U9821 (N_9821,N_9167,N_9316);
nor U9822 (N_9822,N_9086,N_9276);
or U9823 (N_9823,N_9024,N_9418);
xor U9824 (N_9824,N_9475,N_9082);
nor U9825 (N_9825,N_9145,N_9297);
or U9826 (N_9826,N_9060,N_9357);
xor U9827 (N_9827,N_9118,N_9311);
xnor U9828 (N_9828,N_9205,N_9074);
xor U9829 (N_9829,N_9197,N_9490);
and U9830 (N_9830,N_9136,N_9086);
or U9831 (N_9831,N_9223,N_9358);
nor U9832 (N_9832,N_9284,N_9426);
xnor U9833 (N_9833,N_9485,N_9174);
nand U9834 (N_9834,N_9137,N_9405);
or U9835 (N_9835,N_9044,N_9018);
nand U9836 (N_9836,N_9129,N_9406);
nand U9837 (N_9837,N_9270,N_9407);
or U9838 (N_9838,N_9395,N_9248);
or U9839 (N_9839,N_9217,N_9327);
nor U9840 (N_9840,N_9434,N_9362);
nand U9841 (N_9841,N_9244,N_9418);
nand U9842 (N_9842,N_9113,N_9436);
xor U9843 (N_9843,N_9499,N_9059);
nor U9844 (N_9844,N_9336,N_9135);
and U9845 (N_9845,N_9466,N_9025);
nor U9846 (N_9846,N_9443,N_9271);
and U9847 (N_9847,N_9473,N_9105);
xor U9848 (N_9848,N_9303,N_9121);
nand U9849 (N_9849,N_9192,N_9379);
xnor U9850 (N_9850,N_9404,N_9035);
xnor U9851 (N_9851,N_9065,N_9144);
and U9852 (N_9852,N_9020,N_9172);
nor U9853 (N_9853,N_9190,N_9045);
and U9854 (N_9854,N_9090,N_9341);
nand U9855 (N_9855,N_9314,N_9425);
or U9856 (N_9856,N_9195,N_9110);
nand U9857 (N_9857,N_9215,N_9320);
nor U9858 (N_9858,N_9482,N_9106);
xor U9859 (N_9859,N_9433,N_9491);
xnor U9860 (N_9860,N_9192,N_9437);
nand U9861 (N_9861,N_9364,N_9210);
nor U9862 (N_9862,N_9493,N_9198);
and U9863 (N_9863,N_9093,N_9162);
or U9864 (N_9864,N_9126,N_9071);
xnor U9865 (N_9865,N_9017,N_9031);
or U9866 (N_9866,N_9342,N_9043);
or U9867 (N_9867,N_9227,N_9055);
and U9868 (N_9868,N_9129,N_9391);
nor U9869 (N_9869,N_9170,N_9228);
nor U9870 (N_9870,N_9408,N_9272);
nand U9871 (N_9871,N_9000,N_9391);
or U9872 (N_9872,N_9096,N_9140);
nor U9873 (N_9873,N_9020,N_9082);
and U9874 (N_9874,N_9370,N_9496);
xor U9875 (N_9875,N_9493,N_9191);
and U9876 (N_9876,N_9383,N_9105);
or U9877 (N_9877,N_9430,N_9092);
or U9878 (N_9878,N_9237,N_9357);
nand U9879 (N_9879,N_9096,N_9379);
xor U9880 (N_9880,N_9283,N_9383);
xor U9881 (N_9881,N_9408,N_9271);
xor U9882 (N_9882,N_9444,N_9134);
or U9883 (N_9883,N_9283,N_9486);
nand U9884 (N_9884,N_9022,N_9025);
or U9885 (N_9885,N_9079,N_9262);
or U9886 (N_9886,N_9416,N_9146);
or U9887 (N_9887,N_9232,N_9055);
nand U9888 (N_9888,N_9007,N_9348);
and U9889 (N_9889,N_9380,N_9317);
or U9890 (N_9890,N_9409,N_9254);
and U9891 (N_9891,N_9164,N_9488);
and U9892 (N_9892,N_9246,N_9041);
and U9893 (N_9893,N_9144,N_9380);
nand U9894 (N_9894,N_9359,N_9023);
xnor U9895 (N_9895,N_9287,N_9221);
or U9896 (N_9896,N_9449,N_9118);
and U9897 (N_9897,N_9438,N_9377);
nand U9898 (N_9898,N_9121,N_9201);
nand U9899 (N_9899,N_9087,N_9225);
or U9900 (N_9900,N_9140,N_9436);
xnor U9901 (N_9901,N_9191,N_9101);
nor U9902 (N_9902,N_9413,N_9028);
xnor U9903 (N_9903,N_9192,N_9301);
nor U9904 (N_9904,N_9480,N_9216);
xor U9905 (N_9905,N_9302,N_9164);
nand U9906 (N_9906,N_9339,N_9028);
or U9907 (N_9907,N_9259,N_9292);
nor U9908 (N_9908,N_9277,N_9006);
xnor U9909 (N_9909,N_9265,N_9457);
xor U9910 (N_9910,N_9441,N_9439);
and U9911 (N_9911,N_9181,N_9217);
nand U9912 (N_9912,N_9322,N_9419);
or U9913 (N_9913,N_9081,N_9103);
nand U9914 (N_9914,N_9201,N_9297);
xnor U9915 (N_9915,N_9492,N_9464);
and U9916 (N_9916,N_9196,N_9025);
nand U9917 (N_9917,N_9073,N_9005);
or U9918 (N_9918,N_9297,N_9498);
or U9919 (N_9919,N_9258,N_9080);
nand U9920 (N_9920,N_9391,N_9191);
nor U9921 (N_9921,N_9057,N_9075);
nor U9922 (N_9922,N_9129,N_9417);
and U9923 (N_9923,N_9286,N_9161);
nand U9924 (N_9924,N_9307,N_9133);
nor U9925 (N_9925,N_9310,N_9443);
nand U9926 (N_9926,N_9466,N_9320);
xnor U9927 (N_9927,N_9411,N_9192);
nor U9928 (N_9928,N_9286,N_9448);
xor U9929 (N_9929,N_9418,N_9368);
and U9930 (N_9930,N_9491,N_9134);
nor U9931 (N_9931,N_9170,N_9373);
or U9932 (N_9932,N_9274,N_9001);
and U9933 (N_9933,N_9312,N_9100);
nor U9934 (N_9934,N_9059,N_9090);
nor U9935 (N_9935,N_9466,N_9409);
xor U9936 (N_9936,N_9177,N_9201);
or U9937 (N_9937,N_9226,N_9157);
nor U9938 (N_9938,N_9318,N_9366);
or U9939 (N_9939,N_9288,N_9155);
and U9940 (N_9940,N_9020,N_9123);
and U9941 (N_9941,N_9006,N_9249);
or U9942 (N_9942,N_9392,N_9063);
nor U9943 (N_9943,N_9383,N_9439);
xnor U9944 (N_9944,N_9044,N_9152);
nor U9945 (N_9945,N_9079,N_9049);
xor U9946 (N_9946,N_9227,N_9354);
and U9947 (N_9947,N_9172,N_9452);
nor U9948 (N_9948,N_9455,N_9349);
or U9949 (N_9949,N_9081,N_9237);
xnor U9950 (N_9950,N_9315,N_9209);
or U9951 (N_9951,N_9204,N_9056);
nand U9952 (N_9952,N_9412,N_9428);
xnor U9953 (N_9953,N_9039,N_9343);
nor U9954 (N_9954,N_9214,N_9451);
or U9955 (N_9955,N_9374,N_9088);
nor U9956 (N_9956,N_9465,N_9277);
nor U9957 (N_9957,N_9104,N_9296);
nand U9958 (N_9958,N_9299,N_9444);
nand U9959 (N_9959,N_9063,N_9084);
nand U9960 (N_9960,N_9135,N_9222);
nand U9961 (N_9961,N_9087,N_9434);
xnor U9962 (N_9962,N_9440,N_9319);
nor U9963 (N_9963,N_9445,N_9188);
or U9964 (N_9964,N_9250,N_9321);
and U9965 (N_9965,N_9241,N_9254);
xnor U9966 (N_9966,N_9029,N_9485);
nand U9967 (N_9967,N_9475,N_9471);
nand U9968 (N_9968,N_9412,N_9145);
xor U9969 (N_9969,N_9140,N_9105);
nand U9970 (N_9970,N_9473,N_9047);
or U9971 (N_9971,N_9187,N_9471);
nor U9972 (N_9972,N_9382,N_9004);
and U9973 (N_9973,N_9008,N_9133);
nor U9974 (N_9974,N_9254,N_9006);
and U9975 (N_9975,N_9230,N_9324);
xor U9976 (N_9976,N_9412,N_9179);
nand U9977 (N_9977,N_9126,N_9076);
nand U9978 (N_9978,N_9304,N_9079);
and U9979 (N_9979,N_9313,N_9314);
and U9980 (N_9980,N_9294,N_9276);
or U9981 (N_9981,N_9012,N_9325);
nor U9982 (N_9982,N_9322,N_9046);
nor U9983 (N_9983,N_9464,N_9289);
or U9984 (N_9984,N_9410,N_9129);
nand U9985 (N_9985,N_9271,N_9324);
nand U9986 (N_9986,N_9027,N_9196);
nor U9987 (N_9987,N_9151,N_9346);
and U9988 (N_9988,N_9336,N_9162);
or U9989 (N_9989,N_9392,N_9302);
and U9990 (N_9990,N_9324,N_9446);
nand U9991 (N_9991,N_9438,N_9263);
and U9992 (N_9992,N_9208,N_9114);
or U9993 (N_9993,N_9378,N_9054);
nor U9994 (N_9994,N_9128,N_9204);
and U9995 (N_9995,N_9318,N_9065);
and U9996 (N_9996,N_9428,N_9029);
nand U9997 (N_9997,N_9360,N_9424);
nand U9998 (N_9998,N_9028,N_9468);
xor U9999 (N_9999,N_9207,N_9361);
xor U10000 (N_10000,N_9787,N_9869);
nor U10001 (N_10001,N_9808,N_9587);
xnor U10002 (N_10002,N_9662,N_9954);
xor U10003 (N_10003,N_9677,N_9822);
nor U10004 (N_10004,N_9726,N_9760);
xnor U10005 (N_10005,N_9964,N_9674);
nor U10006 (N_10006,N_9518,N_9692);
nor U10007 (N_10007,N_9502,N_9871);
nor U10008 (N_10008,N_9565,N_9806);
nor U10009 (N_10009,N_9794,N_9588);
and U10010 (N_10010,N_9879,N_9872);
nor U10011 (N_10011,N_9881,N_9922);
nand U10012 (N_10012,N_9989,N_9977);
xor U10013 (N_10013,N_9702,N_9899);
xor U10014 (N_10014,N_9578,N_9573);
nor U10015 (N_10015,N_9915,N_9882);
nand U10016 (N_10016,N_9716,N_9558);
and U10017 (N_10017,N_9892,N_9925);
xnor U10018 (N_10018,N_9515,N_9812);
nand U10019 (N_10019,N_9975,N_9820);
nand U10020 (N_10020,N_9776,N_9870);
nand U10021 (N_10021,N_9624,N_9640);
or U10022 (N_10022,N_9765,N_9912);
and U10023 (N_10023,N_9982,N_9715);
nor U10024 (N_10024,N_9528,N_9681);
nor U10025 (N_10025,N_9804,N_9514);
nor U10026 (N_10026,N_9705,N_9958);
or U10027 (N_10027,N_9749,N_9685);
or U10028 (N_10028,N_9630,N_9920);
xor U10029 (N_10029,N_9534,N_9917);
or U10030 (N_10030,N_9967,N_9829);
and U10031 (N_10031,N_9670,N_9943);
nor U10032 (N_10032,N_9736,N_9696);
and U10033 (N_10033,N_9690,N_9947);
nor U10034 (N_10034,N_9704,N_9554);
or U10035 (N_10035,N_9768,N_9548);
xor U10036 (N_10036,N_9657,N_9933);
or U10037 (N_10037,N_9934,N_9599);
nor U10038 (N_10038,N_9613,N_9663);
and U10039 (N_10039,N_9672,N_9956);
and U10040 (N_10040,N_9836,N_9955);
nand U10041 (N_10041,N_9885,N_9873);
nand U10042 (N_10042,N_9896,N_9550);
nand U10043 (N_10043,N_9750,N_9532);
or U10044 (N_10044,N_9616,N_9942);
or U10045 (N_10045,N_9546,N_9751);
or U10046 (N_10046,N_9730,N_9997);
and U10047 (N_10047,N_9966,N_9762);
nor U10048 (N_10048,N_9608,N_9535);
nor U10049 (N_10049,N_9837,N_9887);
nand U10050 (N_10050,N_9553,N_9991);
nor U10051 (N_10051,N_9936,N_9543);
nor U10052 (N_10052,N_9615,N_9980);
and U10053 (N_10053,N_9684,N_9826);
xor U10054 (N_10054,N_9780,N_9676);
nor U10055 (N_10055,N_9522,N_9786);
xnor U10056 (N_10056,N_9619,N_9926);
nor U10057 (N_10057,N_9900,N_9863);
xor U10058 (N_10058,N_9503,N_9581);
or U10059 (N_10059,N_9665,N_9877);
nor U10060 (N_10060,N_9509,N_9907);
xnor U10061 (N_10061,N_9529,N_9905);
or U10062 (N_10062,N_9985,N_9513);
and U10063 (N_10063,N_9626,N_9713);
or U10064 (N_10064,N_9709,N_9678);
or U10065 (N_10065,N_9564,N_9718);
xnor U10066 (N_10066,N_9647,N_9970);
nand U10067 (N_10067,N_9703,N_9764);
and U10068 (N_10068,N_9830,N_9791);
and U10069 (N_10069,N_9590,N_9673);
or U10070 (N_10070,N_9719,N_9895);
nand U10071 (N_10071,N_9505,N_9853);
and U10072 (N_10072,N_9855,N_9792);
xor U10073 (N_10073,N_9723,N_9551);
or U10074 (N_10074,N_9720,N_9642);
and U10075 (N_10075,N_9567,N_9525);
and U10076 (N_10076,N_9852,N_9711);
nor U10077 (N_10077,N_9769,N_9913);
xnor U10078 (N_10078,N_9559,N_9914);
nand U10079 (N_10079,N_9854,N_9602);
nor U10080 (N_10080,N_9901,N_9748);
or U10081 (N_10081,N_9682,N_9686);
nand U10082 (N_10082,N_9841,N_9531);
nand U10083 (N_10083,N_9814,N_9618);
nor U10084 (N_10084,N_9628,N_9833);
and U10085 (N_10085,N_9617,N_9524);
nor U10086 (N_10086,N_9583,N_9941);
and U10087 (N_10087,N_9717,N_9990);
xnor U10088 (N_10088,N_9629,N_9517);
and U10089 (N_10089,N_9691,N_9566);
or U10090 (N_10090,N_9838,N_9951);
xor U10091 (N_10091,N_9862,N_9544);
and U10092 (N_10092,N_9880,N_9950);
nor U10093 (N_10093,N_9596,N_9731);
nand U10094 (N_10094,N_9798,N_9883);
and U10095 (N_10095,N_9533,N_9824);
xnor U10096 (N_10096,N_9577,N_9874);
nand U10097 (N_10097,N_9818,N_9664);
nor U10098 (N_10098,N_9957,N_9552);
nand U10099 (N_10099,N_9538,N_9738);
or U10100 (N_10100,N_9911,N_9530);
xor U10101 (N_10101,N_9646,N_9797);
or U10102 (N_10102,N_9969,N_9560);
nand U10103 (N_10103,N_9755,N_9927);
and U10104 (N_10104,N_9747,N_9600);
or U10105 (N_10105,N_9962,N_9779);
or U10106 (N_10106,N_9894,N_9699);
xor U10107 (N_10107,N_9821,N_9817);
nor U10108 (N_10108,N_9545,N_9807);
or U10109 (N_10109,N_9541,N_9952);
or U10110 (N_10110,N_9570,N_9849);
or U10111 (N_10111,N_9683,N_9784);
xor U10112 (N_10112,N_9953,N_9555);
and U10113 (N_10113,N_9631,N_9512);
nor U10114 (N_10114,N_9614,N_9557);
xor U10115 (N_10115,N_9754,N_9651);
or U10116 (N_10116,N_9766,N_9521);
nand U10117 (N_10117,N_9585,N_9639);
nand U10118 (N_10118,N_9921,N_9542);
and U10119 (N_10119,N_9501,N_9511);
xor U10120 (N_10120,N_9707,N_9793);
xnor U10121 (N_10121,N_9995,N_9732);
and U10122 (N_10122,N_9851,N_9759);
nor U10123 (N_10123,N_9661,N_9603);
or U10124 (N_10124,N_9993,N_9537);
xnor U10125 (N_10125,N_9612,N_9815);
or U10126 (N_10126,N_9697,N_9540);
and U10127 (N_10127,N_9782,N_9960);
xor U10128 (N_10128,N_9884,N_9984);
xnor U10129 (N_10129,N_9992,N_9799);
or U10130 (N_10130,N_9660,N_9777);
and U10131 (N_10131,N_9589,N_9781);
and U10132 (N_10132,N_9741,N_9520);
xnor U10133 (N_10133,N_9875,N_9737);
xnor U10134 (N_10134,N_9547,N_9916);
nand U10135 (N_10135,N_9563,N_9772);
or U10136 (N_10136,N_9591,N_9976);
xor U10137 (N_10137,N_9620,N_9734);
xor U10138 (N_10138,N_9625,N_9940);
or U10139 (N_10139,N_9756,N_9659);
and U10140 (N_10140,N_9667,N_9831);
or U10141 (N_10141,N_9606,N_9745);
and U10142 (N_10142,N_9842,N_9687);
nand U10143 (N_10143,N_9939,N_9740);
xnor U10144 (N_10144,N_9580,N_9773);
or U10145 (N_10145,N_9666,N_9832);
and U10146 (N_10146,N_9668,N_9593);
xor U10147 (N_10147,N_9770,N_9858);
or U10148 (N_10148,N_9857,N_9643);
or U10149 (N_10149,N_9839,N_9988);
nand U10150 (N_10150,N_9919,N_9742);
xor U10151 (N_10151,N_9778,N_9866);
and U10152 (N_10152,N_9519,N_9996);
and U10153 (N_10153,N_9706,N_9935);
and U10154 (N_10154,N_9979,N_9568);
xnor U10155 (N_10155,N_9847,N_9653);
nand U10156 (N_10156,N_9946,N_9825);
and U10157 (N_10157,N_9607,N_9861);
xor U10158 (N_10158,N_9819,N_9796);
xor U10159 (N_10159,N_9627,N_9767);
nor U10160 (N_10160,N_9635,N_9500);
xor U10161 (N_10161,N_9968,N_9802);
or U10162 (N_10162,N_9891,N_9827);
or U10163 (N_10163,N_9971,N_9889);
and U10164 (N_10164,N_9763,N_9611);
or U10165 (N_10165,N_9974,N_9910);
xnor U10166 (N_10166,N_9801,N_9843);
and U10167 (N_10167,N_9743,N_9986);
or U10168 (N_10168,N_9844,N_9850);
nor U10169 (N_10169,N_9721,N_9700);
xor U10170 (N_10170,N_9575,N_9902);
nand U10171 (N_10171,N_9865,N_9994);
nor U10172 (N_10172,N_9610,N_9680);
xor U10173 (N_10173,N_9930,N_9835);
or U10174 (N_10174,N_9908,N_9828);
or U10175 (N_10175,N_9576,N_9898);
nor U10176 (N_10176,N_9571,N_9928);
nand U10177 (N_10177,N_9810,N_9506);
xor U10178 (N_10178,N_9963,N_9688);
xor U10179 (N_10179,N_9972,N_9650);
xor U10180 (N_10180,N_9811,N_9886);
and U10181 (N_10181,N_9694,N_9998);
xnor U10182 (N_10182,N_9652,N_9539);
nand U10183 (N_10183,N_9638,N_9904);
xor U10184 (N_10184,N_9701,N_9549);
and U10185 (N_10185,N_9695,N_9728);
xnor U10186 (N_10186,N_9654,N_9675);
and U10187 (N_10187,N_9536,N_9710);
xnor U10188 (N_10188,N_9722,N_9597);
and U10189 (N_10189,N_9923,N_9803);
or U10190 (N_10190,N_9823,N_9800);
or U10191 (N_10191,N_9868,N_9733);
or U10192 (N_10192,N_9788,N_9679);
nand U10193 (N_10193,N_9816,N_9795);
or U10194 (N_10194,N_9595,N_9712);
nor U10195 (N_10195,N_9878,N_9859);
nor U10196 (N_10196,N_9689,N_9948);
or U10197 (N_10197,N_9937,N_9845);
nor U10198 (N_10198,N_9645,N_9648);
nor U10199 (N_10199,N_9725,N_9634);
and U10200 (N_10200,N_9938,N_9623);
xor U10201 (N_10201,N_9516,N_9724);
or U10202 (N_10202,N_9523,N_9785);
nor U10203 (N_10203,N_9698,N_9932);
nand U10204 (N_10204,N_9592,N_9961);
xor U10205 (N_10205,N_9708,N_9579);
nor U10206 (N_10206,N_9633,N_9918);
xnor U10207 (N_10207,N_9783,N_9508);
and U10208 (N_10208,N_9637,N_9999);
or U10209 (N_10209,N_9909,N_9757);
nand U10210 (N_10210,N_9658,N_9594);
nor U10211 (N_10211,N_9867,N_9805);
xnor U10212 (N_10212,N_9735,N_9890);
xnor U10213 (N_10213,N_9746,N_9632);
xor U10214 (N_10214,N_9604,N_9739);
or U10215 (N_10215,N_9965,N_9945);
xnor U10216 (N_10216,N_9561,N_9714);
or U10217 (N_10217,N_9876,N_9775);
nor U10218 (N_10218,N_9584,N_9601);
xnor U10219 (N_10219,N_9893,N_9774);
and U10220 (N_10220,N_9931,N_9507);
and U10221 (N_10221,N_9636,N_9983);
nand U10222 (N_10222,N_9813,N_9834);
nand U10223 (N_10223,N_9929,N_9510);
nor U10224 (N_10224,N_9641,N_9987);
and U10225 (N_10225,N_9973,N_9693);
nor U10226 (N_10226,N_9655,N_9744);
nor U10227 (N_10227,N_9649,N_9981);
and U10228 (N_10228,N_9903,N_9860);
xor U10229 (N_10229,N_9598,N_9864);
nor U10230 (N_10230,N_9758,N_9771);
nor U10231 (N_10231,N_9656,N_9727);
and U10232 (N_10232,N_9840,N_9924);
and U10233 (N_10233,N_9669,N_9621);
nand U10234 (N_10234,N_9944,N_9527);
xnor U10235 (N_10235,N_9888,N_9897);
or U10236 (N_10236,N_9586,N_9574);
nor U10237 (N_10237,N_9809,N_9609);
xnor U10238 (N_10238,N_9978,N_9504);
xnor U10239 (N_10239,N_9949,N_9761);
and U10240 (N_10240,N_9906,N_9671);
xor U10241 (N_10241,N_9572,N_9846);
nand U10242 (N_10242,N_9752,N_9644);
nand U10243 (N_10243,N_9753,N_9729);
nand U10244 (N_10244,N_9789,N_9556);
xor U10245 (N_10245,N_9562,N_9790);
nand U10246 (N_10246,N_9605,N_9622);
xnor U10247 (N_10247,N_9582,N_9856);
and U10248 (N_10248,N_9848,N_9959);
xor U10249 (N_10249,N_9526,N_9569);
nand U10250 (N_10250,N_9510,N_9912);
and U10251 (N_10251,N_9875,N_9929);
nand U10252 (N_10252,N_9759,N_9925);
or U10253 (N_10253,N_9614,N_9580);
and U10254 (N_10254,N_9840,N_9667);
xnor U10255 (N_10255,N_9656,N_9619);
and U10256 (N_10256,N_9532,N_9894);
or U10257 (N_10257,N_9903,N_9953);
xor U10258 (N_10258,N_9502,N_9776);
and U10259 (N_10259,N_9918,N_9600);
or U10260 (N_10260,N_9889,N_9706);
nand U10261 (N_10261,N_9955,N_9591);
or U10262 (N_10262,N_9872,N_9555);
nor U10263 (N_10263,N_9721,N_9854);
or U10264 (N_10264,N_9618,N_9776);
xnor U10265 (N_10265,N_9854,N_9514);
and U10266 (N_10266,N_9517,N_9684);
xnor U10267 (N_10267,N_9812,N_9838);
or U10268 (N_10268,N_9532,N_9551);
and U10269 (N_10269,N_9715,N_9899);
nand U10270 (N_10270,N_9994,N_9945);
nor U10271 (N_10271,N_9952,N_9624);
xnor U10272 (N_10272,N_9796,N_9731);
nand U10273 (N_10273,N_9881,N_9939);
nor U10274 (N_10274,N_9902,N_9725);
or U10275 (N_10275,N_9780,N_9880);
nand U10276 (N_10276,N_9629,N_9750);
and U10277 (N_10277,N_9803,N_9917);
or U10278 (N_10278,N_9973,N_9726);
nand U10279 (N_10279,N_9923,N_9660);
nor U10280 (N_10280,N_9950,N_9704);
nand U10281 (N_10281,N_9748,N_9971);
or U10282 (N_10282,N_9861,N_9817);
xor U10283 (N_10283,N_9529,N_9577);
xor U10284 (N_10284,N_9916,N_9806);
nand U10285 (N_10285,N_9950,N_9787);
or U10286 (N_10286,N_9929,N_9974);
and U10287 (N_10287,N_9671,N_9841);
xor U10288 (N_10288,N_9960,N_9704);
nand U10289 (N_10289,N_9825,N_9776);
or U10290 (N_10290,N_9882,N_9795);
or U10291 (N_10291,N_9657,N_9595);
or U10292 (N_10292,N_9760,N_9533);
xnor U10293 (N_10293,N_9744,N_9573);
or U10294 (N_10294,N_9871,N_9611);
xnor U10295 (N_10295,N_9671,N_9826);
xor U10296 (N_10296,N_9825,N_9527);
and U10297 (N_10297,N_9781,N_9709);
or U10298 (N_10298,N_9928,N_9882);
xnor U10299 (N_10299,N_9515,N_9824);
nor U10300 (N_10300,N_9542,N_9500);
nor U10301 (N_10301,N_9686,N_9766);
nor U10302 (N_10302,N_9576,N_9994);
and U10303 (N_10303,N_9635,N_9533);
nor U10304 (N_10304,N_9941,N_9901);
nor U10305 (N_10305,N_9742,N_9527);
nand U10306 (N_10306,N_9881,N_9956);
and U10307 (N_10307,N_9744,N_9629);
xnor U10308 (N_10308,N_9915,N_9722);
xnor U10309 (N_10309,N_9769,N_9757);
or U10310 (N_10310,N_9627,N_9541);
or U10311 (N_10311,N_9609,N_9566);
nand U10312 (N_10312,N_9576,N_9814);
or U10313 (N_10313,N_9700,N_9795);
and U10314 (N_10314,N_9708,N_9776);
xor U10315 (N_10315,N_9555,N_9559);
or U10316 (N_10316,N_9670,N_9812);
nand U10317 (N_10317,N_9827,N_9969);
or U10318 (N_10318,N_9610,N_9801);
xor U10319 (N_10319,N_9888,N_9895);
and U10320 (N_10320,N_9626,N_9717);
nand U10321 (N_10321,N_9594,N_9501);
or U10322 (N_10322,N_9544,N_9781);
or U10323 (N_10323,N_9775,N_9637);
or U10324 (N_10324,N_9878,N_9800);
xnor U10325 (N_10325,N_9946,N_9930);
or U10326 (N_10326,N_9816,N_9657);
nand U10327 (N_10327,N_9587,N_9697);
xor U10328 (N_10328,N_9689,N_9740);
or U10329 (N_10329,N_9716,N_9929);
nor U10330 (N_10330,N_9677,N_9630);
or U10331 (N_10331,N_9562,N_9934);
nand U10332 (N_10332,N_9655,N_9692);
nand U10333 (N_10333,N_9747,N_9766);
and U10334 (N_10334,N_9922,N_9785);
or U10335 (N_10335,N_9673,N_9529);
nor U10336 (N_10336,N_9524,N_9871);
nor U10337 (N_10337,N_9784,N_9689);
nand U10338 (N_10338,N_9730,N_9896);
or U10339 (N_10339,N_9989,N_9796);
xor U10340 (N_10340,N_9876,N_9989);
and U10341 (N_10341,N_9502,N_9927);
xor U10342 (N_10342,N_9531,N_9828);
xor U10343 (N_10343,N_9718,N_9751);
or U10344 (N_10344,N_9566,N_9701);
nand U10345 (N_10345,N_9501,N_9679);
nor U10346 (N_10346,N_9569,N_9938);
nor U10347 (N_10347,N_9984,N_9882);
and U10348 (N_10348,N_9984,N_9582);
or U10349 (N_10349,N_9976,N_9741);
or U10350 (N_10350,N_9894,N_9821);
and U10351 (N_10351,N_9888,N_9806);
and U10352 (N_10352,N_9638,N_9899);
or U10353 (N_10353,N_9730,N_9562);
nor U10354 (N_10354,N_9621,N_9929);
nand U10355 (N_10355,N_9676,N_9899);
xor U10356 (N_10356,N_9897,N_9734);
or U10357 (N_10357,N_9999,N_9697);
and U10358 (N_10358,N_9673,N_9645);
and U10359 (N_10359,N_9736,N_9608);
nor U10360 (N_10360,N_9615,N_9566);
nand U10361 (N_10361,N_9502,N_9766);
xnor U10362 (N_10362,N_9859,N_9548);
nand U10363 (N_10363,N_9573,N_9990);
or U10364 (N_10364,N_9679,N_9877);
and U10365 (N_10365,N_9559,N_9694);
or U10366 (N_10366,N_9860,N_9885);
nor U10367 (N_10367,N_9732,N_9859);
xor U10368 (N_10368,N_9660,N_9553);
xor U10369 (N_10369,N_9550,N_9855);
nand U10370 (N_10370,N_9630,N_9884);
nand U10371 (N_10371,N_9971,N_9577);
and U10372 (N_10372,N_9909,N_9931);
nor U10373 (N_10373,N_9575,N_9746);
nand U10374 (N_10374,N_9949,N_9787);
nand U10375 (N_10375,N_9978,N_9831);
and U10376 (N_10376,N_9552,N_9698);
xnor U10377 (N_10377,N_9608,N_9774);
nand U10378 (N_10378,N_9614,N_9927);
or U10379 (N_10379,N_9554,N_9635);
nor U10380 (N_10380,N_9876,N_9505);
nor U10381 (N_10381,N_9764,N_9903);
or U10382 (N_10382,N_9748,N_9507);
nor U10383 (N_10383,N_9758,N_9544);
or U10384 (N_10384,N_9583,N_9744);
nand U10385 (N_10385,N_9752,N_9599);
nand U10386 (N_10386,N_9798,N_9974);
or U10387 (N_10387,N_9646,N_9936);
nor U10388 (N_10388,N_9541,N_9518);
nor U10389 (N_10389,N_9655,N_9526);
or U10390 (N_10390,N_9706,N_9812);
xnor U10391 (N_10391,N_9990,N_9880);
or U10392 (N_10392,N_9785,N_9870);
nand U10393 (N_10393,N_9903,N_9940);
nor U10394 (N_10394,N_9958,N_9671);
nor U10395 (N_10395,N_9712,N_9947);
and U10396 (N_10396,N_9839,N_9735);
xnor U10397 (N_10397,N_9606,N_9996);
nor U10398 (N_10398,N_9990,N_9562);
xnor U10399 (N_10399,N_9942,N_9601);
xnor U10400 (N_10400,N_9950,N_9842);
and U10401 (N_10401,N_9578,N_9927);
nand U10402 (N_10402,N_9564,N_9721);
nand U10403 (N_10403,N_9534,N_9692);
nor U10404 (N_10404,N_9788,N_9627);
nor U10405 (N_10405,N_9557,N_9937);
or U10406 (N_10406,N_9974,N_9722);
or U10407 (N_10407,N_9939,N_9795);
or U10408 (N_10408,N_9587,N_9704);
nand U10409 (N_10409,N_9931,N_9854);
xor U10410 (N_10410,N_9583,N_9749);
or U10411 (N_10411,N_9511,N_9555);
and U10412 (N_10412,N_9849,N_9661);
nand U10413 (N_10413,N_9898,N_9791);
nor U10414 (N_10414,N_9593,N_9809);
xnor U10415 (N_10415,N_9536,N_9807);
nand U10416 (N_10416,N_9767,N_9803);
and U10417 (N_10417,N_9952,N_9529);
xor U10418 (N_10418,N_9884,N_9961);
or U10419 (N_10419,N_9814,N_9793);
or U10420 (N_10420,N_9675,N_9656);
or U10421 (N_10421,N_9573,N_9564);
nor U10422 (N_10422,N_9657,N_9887);
xor U10423 (N_10423,N_9580,N_9747);
nand U10424 (N_10424,N_9977,N_9963);
and U10425 (N_10425,N_9857,N_9615);
nand U10426 (N_10426,N_9801,N_9982);
or U10427 (N_10427,N_9602,N_9717);
nand U10428 (N_10428,N_9960,N_9757);
nand U10429 (N_10429,N_9526,N_9633);
and U10430 (N_10430,N_9875,N_9537);
xnor U10431 (N_10431,N_9738,N_9588);
nor U10432 (N_10432,N_9909,N_9601);
and U10433 (N_10433,N_9792,N_9977);
xor U10434 (N_10434,N_9619,N_9956);
and U10435 (N_10435,N_9545,N_9783);
or U10436 (N_10436,N_9865,N_9936);
nand U10437 (N_10437,N_9933,N_9882);
and U10438 (N_10438,N_9558,N_9544);
nand U10439 (N_10439,N_9752,N_9529);
or U10440 (N_10440,N_9877,N_9870);
nand U10441 (N_10441,N_9556,N_9532);
xor U10442 (N_10442,N_9508,N_9762);
nand U10443 (N_10443,N_9545,N_9649);
nor U10444 (N_10444,N_9642,N_9713);
and U10445 (N_10445,N_9755,N_9788);
or U10446 (N_10446,N_9567,N_9705);
or U10447 (N_10447,N_9923,N_9707);
nand U10448 (N_10448,N_9606,N_9629);
xor U10449 (N_10449,N_9692,N_9942);
nor U10450 (N_10450,N_9781,N_9802);
xnor U10451 (N_10451,N_9814,N_9561);
xnor U10452 (N_10452,N_9576,N_9569);
nand U10453 (N_10453,N_9572,N_9768);
or U10454 (N_10454,N_9820,N_9924);
xor U10455 (N_10455,N_9921,N_9546);
or U10456 (N_10456,N_9743,N_9960);
xor U10457 (N_10457,N_9547,N_9681);
nand U10458 (N_10458,N_9859,N_9871);
or U10459 (N_10459,N_9917,N_9634);
nand U10460 (N_10460,N_9916,N_9698);
or U10461 (N_10461,N_9626,N_9837);
nor U10462 (N_10462,N_9508,N_9510);
and U10463 (N_10463,N_9974,N_9928);
xnor U10464 (N_10464,N_9762,N_9906);
or U10465 (N_10465,N_9553,N_9541);
or U10466 (N_10466,N_9654,N_9891);
or U10467 (N_10467,N_9712,N_9585);
and U10468 (N_10468,N_9856,N_9665);
or U10469 (N_10469,N_9716,N_9705);
xnor U10470 (N_10470,N_9886,N_9953);
and U10471 (N_10471,N_9591,N_9505);
nor U10472 (N_10472,N_9872,N_9767);
or U10473 (N_10473,N_9600,N_9574);
and U10474 (N_10474,N_9519,N_9899);
nor U10475 (N_10475,N_9577,N_9990);
or U10476 (N_10476,N_9703,N_9709);
or U10477 (N_10477,N_9762,N_9554);
or U10478 (N_10478,N_9705,N_9856);
xnor U10479 (N_10479,N_9606,N_9995);
nand U10480 (N_10480,N_9922,N_9536);
and U10481 (N_10481,N_9723,N_9684);
and U10482 (N_10482,N_9795,N_9506);
or U10483 (N_10483,N_9654,N_9940);
nor U10484 (N_10484,N_9831,N_9940);
and U10485 (N_10485,N_9795,N_9611);
nand U10486 (N_10486,N_9959,N_9605);
nand U10487 (N_10487,N_9781,N_9683);
nor U10488 (N_10488,N_9795,N_9862);
or U10489 (N_10489,N_9501,N_9560);
xor U10490 (N_10490,N_9883,N_9817);
xor U10491 (N_10491,N_9701,N_9517);
nor U10492 (N_10492,N_9628,N_9730);
and U10493 (N_10493,N_9997,N_9500);
nand U10494 (N_10494,N_9911,N_9876);
xnor U10495 (N_10495,N_9678,N_9566);
xor U10496 (N_10496,N_9955,N_9547);
nor U10497 (N_10497,N_9747,N_9843);
xor U10498 (N_10498,N_9995,N_9800);
nand U10499 (N_10499,N_9991,N_9752);
nand U10500 (N_10500,N_10350,N_10468);
and U10501 (N_10501,N_10365,N_10269);
nand U10502 (N_10502,N_10218,N_10155);
or U10503 (N_10503,N_10368,N_10239);
nand U10504 (N_10504,N_10202,N_10276);
nand U10505 (N_10505,N_10119,N_10002);
nand U10506 (N_10506,N_10283,N_10219);
xnor U10507 (N_10507,N_10323,N_10179);
and U10508 (N_10508,N_10178,N_10253);
nor U10509 (N_10509,N_10160,N_10063);
nor U10510 (N_10510,N_10249,N_10245);
xor U10511 (N_10511,N_10047,N_10216);
nand U10512 (N_10512,N_10361,N_10366);
nand U10513 (N_10513,N_10125,N_10308);
nor U10514 (N_10514,N_10490,N_10076);
nand U10515 (N_10515,N_10317,N_10105);
xor U10516 (N_10516,N_10183,N_10459);
nor U10517 (N_10517,N_10142,N_10477);
nor U10518 (N_10518,N_10273,N_10093);
nor U10519 (N_10519,N_10133,N_10104);
xor U10520 (N_10520,N_10035,N_10338);
nand U10521 (N_10521,N_10400,N_10237);
nand U10522 (N_10522,N_10401,N_10187);
nand U10523 (N_10523,N_10347,N_10094);
nand U10524 (N_10524,N_10172,N_10058);
xnor U10525 (N_10525,N_10024,N_10146);
nor U10526 (N_10526,N_10443,N_10475);
and U10527 (N_10527,N_10255,N_10074);
xor U10528 (N_10528,N_10148,N_10286);
or U10529 (N_10529,N_10394,N_10268);
nor U10530 (N_10530,N_10422,N_10158);
or U10531 (N_10531,N_10083,N_10056);
and U10532 (N_10532,N_10441,N_10194);
nand U10533 (N_10533,N_10288,N_10207);
xnor U10534 (N_10534,N_10020,N_10407);
and U10535 (N_10535,N_10483,N_10021);
nor U10536 (N_10536,N_10306,N_10137);
nor U10537 (N_10537,N_10045,N_10185);
nand U10538 (N_10538,N_10033,N_10073);
nor U10539 (N_10539,N_10213,N_10162);
and U10540 (N_10540,N_10435,N_10373);
nand U10541 (N_10541,N_10437,N_10414);
nor U10542 (N_10542,N_10199,N_10360);
or U10543 (N_10543,N_10252,N_10208);
xnor U10544 (N_10544,N_10419,N_10188);
or U10545 (N_10545,N_10480,N_10244);
or U10546 (N_10546,N_10307,N_10032);
and U10547 (N_10547,N_10446,N_10295);
nor U10548 (N_10548,N_10092,N_10211);
and U10549 (N_10549,N_10271,N_10044);
or U10550 (N_10550,N_10221,N_10328);
nor U10551 (N_10551,N_10427,N_10432);
or U10552 (N_10552,N_10023,N_10018);
xor U10553 (N_10553,N_10467,N_10357);
nand U10554 (N_10554,N_10152,N_10242);
nand U10555 (N_10555,N_10327,N_10223);
nor U10556 (N_10556,N_10291,N_10462);
and U10557 (N_10557,N_10476,N_10111);
nand U10558 (N_10558,N_10456,N_10226);
or U10559 (N_10559,N_10012,N_10379);
nand U10560 (N_10560,N_10460,N_10377);
or U10561 (N_10561,N_10067,N_10272);
nand U10562 (N_10562,N_10120,N_10009);
or U10563 (N_10563,N_10465,N_10097);
xor U10564 (N_10564,N_10191,N_10210);
nor U10565 (N_10565,N_10329,N_10193);
xnor U10566 (N_10566,N_10485,N_10322);
or U10567 (N_10567,N_10197,N_10471);
nor U10568 (N_10568,N_10161,N_10220);
and U10569 (N_10569,N_10412,N_10367);
xor U10570 (N_10570,N_10371,N_10302);
or U10571 (N_10571,N_10209,N_10186);
nor U10572 (N_10572,N_10238,N_10054);
xnor U10573 (N_10573,N_10399,N_10167);
xnor U10574 (N_10574,N_10448,N_10095);
and U10575 (N_10575,N_10492,N_10413);
nor U10576 (N_10576,N_10000,N_10089);
xor U10577 (N_10577,N_10007,N_10037);
nor U10578 (N_10578,N_10318,N_10102);
nand U10579 (N_10579,N_10103,N_10233);
nand U10580 (N_10580,N_10433,N_10081);
nor U10581 (N_10581,N_10409,N_10229);
or U10582 (N_10582,N_10293,N_10128);
nand U10583 (N_10583,N_10326,N_10334);
and U10584 (N_10584,N_10248,N_10129);
or U10585 (N_10585,N_10052,N_10256);
nand U10586 (N_10586,N_10234,N_10404);
xnor U10587 (N_10587,N_10489,N_10333);
and U10588 (N_10588,N_10287,N_10236);
or U10589 (N_10589,N_10042,N_10461);
nor U10590 (N_10590,N_10402,N_10298);
or U10591 (N_10591,N_10396,N_10048);
xnor U10592 (N_10592,N_10030,N_10027);
nor U10593 (N_10593,N_10240,N_10494);
or U10594 (N_10594,N_10262,N_10098);
nor U10595 (N_10595,N_10168,N_10444);
or U10596 (N_10596,N_10359,N_10034);
and U10597 (N_10597,N_10484,N_10281);
or U10598 (N_10598,N_10458,N_10428);
xor U10599 (N_10599,N_10266,N_10270);
or U10600 (N_10600,N_10005,N_10082);
or U10601 (N_10601,N_10280,N_10116);
nor U10602 (N_10602,N_10043,N_10296);
nand U10603 (N_10603,N_10316,N_10393);
or U10604 (N_10604,N_10426,N_10455);
nand U10605 (N_10605,N_10397,N_10149);
nor U10606 (N_10606,N_10112,N_10062);
and U10607 (N_10607,N_10241,N_10079);
nor U10608 (N_10608,N_10292,N_10436);
or U10609 (N_10609,N_10060,N_10085);
and U10610 (N_10610,N_10006,N_10153);
nand U10611 (N_10611,N_10430,N_10297);
and U10612 (N_10612,N_10453,N_10294);
and U10613 (N_10613,N_10375,N_10040);
and U10614 (N_10614,N_10358,N_10343);
nor U10615 (N_10615,N_10154,N_10284);
or U10616 (N_10616,N_10450,N_10057);
nor U10617 (N_10617,N_10071,N_10055);
xnor U10618 (N_10618,N_10163,N_10046);
or U10619 (N_10619,N_10025,N_10001);
or U10620 (N_10620,N_10041,N_10277);
nor U10621 (N_10621,N_10051,N_10123);
or U10622 (N_10622,N_10201,N_10261);
nand U10623 (N_10623,N_10140,N_10145);
xnor U10624 (N_10624,N_10217,N_10066);
and U10625 (N_10625,N_10349,N_10439);
nor U10626 (N_10626,N_10447,N_10011);
xor U10627 (N_10627,N_10243,N_10049);
or U10628 (N_10628,N_10224,N_10132);
and U10629 (N_10629,N_10080,N_10362);
nor U10630 (N_10630,N_10247,N_10479);
or U10631 (N_10631,N_10110,N_10342);
nand U10632 (N_10632,N_10463,N_10088);
or U10633 (N_10633,N_10301,N_10144);
or U10634 (N_10634,N_10004,N_10114);
or U10635 (N_10635,N_10141,N_10225);
xor U10636 (N_10636,N_10127,N_10469);
or U10637 (N_10637,N_10330,N_10390);
nand U10638 (N_10638,N_10078,N_10230);
or U10639 (N_10639,N_10091,N_10068);
nand U10640 (N_10640,N_10053,N_10374);
xor U10641 (N_10641,N_10470,N_10304);
or U10642 (N_10642,N_10389,N_10382);
xor U10643 (N_10643,N_10231,N_10107);
and U10644 (N_10644,N_10171,N_10466);
and U10645 (N_10645,N_10335,N_10474);
nand U10646 (N_10646,N_10072,N_10337);
and U10647 (N_10647,N_10147,N_10332);
nor U10648 (N_10648,N_10438,N_10493);
xnor U10649 (N_10649,N_10320,N_10010);
xnor U10650 (N_10650,N_10309,N_10061);
xnor U10651 (N_10651,N_10391,N_10387);
xnor U10652 (N_10652,N_10384,N_10452);
nor U10653 (N_10653,N_10028,N_10014);
xor U10654 (N_10654,N_10015,N_10016);
or U10655 (N_10655,N_10312,N_10499);
and U10656 (N_10656,N_10369,N_10258);
and U10657 (N_10657,N_10165,N_10175);
xor U10658 (N_10658,N_10275,N_10143);
or U10659 (N_10659,N_10222,N_10086);
or U10660 (N_10660,N_10113,N_10008);
nand U10661 (N_10661,N_10192,N_10356);
and U10662 (N_10662,N_10313,N_10274);
or U10663 (N_10663,N_10099,N_10408);
nand U10664 (N_10664,N_10096,N_10036);
or U10665 (N_10665,N_10176,N_10124);
and U10666 (N_10666,N_10353,N_10077);
nand U10667 (N_10667,N_10232,N_10003);
and U10668 (N_10668,N_10454,N_10022);
and U10669 (N_10669,N_10370,N_10424);
xnor U10670 (N_10670,N_10331,N_10351);
nand U10671 (N_10671,N_10246,N_10355);
or U10672 (N_10672,N_10109,N_10200);
xnor U10673 (N_10673,N_10449,N_10101);
or U10674 (N_10674,N_10497,N_10206);
or U10675 (N_10675,N_10190,N_10265);
nor U10676 (N_10676,N_10300,N_10348);
nand U10677 (N_10677,N_10126,N_10013);
xnor U10678 (N_10678,N_10181,N_10108);
nor U10679 (N_10679,N_10038,N_10166);
nor U10680 (N_10680,N_10136,N_10457);
and U10681 (N_10681,N_10380,N_10403);
nand U10682 (N_10682,N_10118,N_10481);
xnor U10683 (N_10683,N_10406,N_10134);
nor U10684 (N_10684,N_10486,N_10180);
or U10685 (N_10685,N_10364,N_10344);
nand U10686 (N_10686,N_10189,N_10429);
nand U10687 (N_10687,N_10029,N_10423);
and U10688 (N_10688,N_10341,N_10420);
and U10689 (N_10689,N_10392,N_10064);
nor U10690 (N_10690,N_10346,N_10214);
nor U10691 (N_10691,N_10431,N_10445);
and U10692 (N_10692,N_10084,N_10372);
xnor U10693 (N_10693,N_10131,N_10121);
nor U10694 (N_10694,N_10196,N_10059);
and U10695 (N_10695,N_10299,N_10411);
and U10696 (N_10696,N_10264,N_10195);
and U10697 (N_10697,N_10050,N_10415);
nor U10698 (N_10698,N_10279,N_10405);
or U10699 (N_10699,N_10482,N_10498);
nor U10700 (N_10700,N_10017,N_10070);
nand U10701 (N_10701,N_10117,N_10340);
nand U10702 (N_10702,N_10352,N_10282);
and U10703 (N_10703,N_10257,N_10442);
or U10704 (N_10704,N_10325,N_10169);
nand U10705 (N_10705,N_10381,N_10410);
nand U10706 (N_10706,N_10026,N_10251);
nand U10707 (N_10707,N_10260,N_10130);
xor U10708 (N_10708,N_10363,N_10065);
and U10709 (N_10709,N_10151,N_10417);
xor U10710 (N_10710,N_10198,N_10321);
or U10711 (N_10711,N_10170,N_10069);
or U10712 (N_10712,N_10385,N_10090);
or U10713 (N_10713,N_10488,N_10164);
and U10714 (N_10714,N_10075,N_10157);
or U10715 (N_10715,N_10138,N_10182);
and U10716 (N_10716,N_10285,N_10354);
xor U10717 (N_10717,N_10339,N_10177);
and U10718 (N_10718,N_10203,N_10314);
or U10719 (N_10719,N_10386,N_10019);
or U10720 (N_10720,N_10336,N_10289);
and U10721 (N_10721,N_10106,N_10227);
xnor U10722 (N_10722,N_10115,N_10278);
and U10723 (N_10723,N_10345,N_10215);
or U10724 (N_10724,N_10303,N_10434);
xnor U10725 (N_10725,N_10388,N_10087);
nand U10726 (N_10726,N_10305,N_10156);
or U10727 (N_10727,N_10159,N_10324);
nand U10728 (N_10728,N_10440,N_10495);
xnor U10729 (N_10729,N_10376,N_10378);
nand U10730 (N_10730,N_10184,N_10267);
xor U10731 (N_10731,N_10395,N_10135);
and U10732 (N_10732,N_10290,N_10254);
and U10733 (N_10733,N_10259,N_10150);
xor U10734 (N_10734,N_10478,N_10263);
nor U10735 (N_10735,N_10451,N_10212);
nor U10736 (N_10736,N_10487,N_10205);
xor U10737 (N_10737,N_10228,N_10310);
nand U10738 (N_10738,N_10235,N_10122);
and U10739 (N_10739,N_10173,N_10472);
or U10740 (N_10740,N_10311,N_10464);
nand U10741 (N_10741,N_10204,N_10421);
xor U10742 (N_10742,N_10100,N_10319);
and U10743 (N_10743,N_10174,N_10139);
xnor U10744 (N_10744,N_10473,N_10383);
or U10745 (N_10745,N_10418,N_10425);
xor U10746 (N_10746,N_10250,N_10315);
and U10747 (N_10747,N_10496,N_10398);
and U10748 (N_10748,N_10031,N_10039);
nor U10749 (N_10749,N_10416,N_10491);
nor U10750 (N_10750,N_10409,N_10060);
and U10751 (N_10751,N_10403,N_10451);
and U10752 (N_10752,N_10224,N_10150);
nand U10753 (N_10753,N_10249,N_10079);
nand U10754 (N_10754,N_10496,N_10484);
and U10755 (N_10755,N_10471,N_10170);
xnor U10756 (N_10756,N_10242,N_10442);
and U10757 (N_10757,N_10417,N_10190);
and U10758 (N_10758,N_10401,N_10287);
or U10759 (N_10759,N_10108,N_10373);
and U10760 (N_10760,N_10152,N_10351);
xnor U10761 (N_10761,N_10230,N_10430);
and U10762 (N_10762,N_10029,N_10433);
nand U10763 (N_10763,N_10060,N_10016);
nor U10764 (N_10764,N_10415,N_10359);
nor U10765 (N_10765,N_10337,N_10272);
nor U10766 (N_10766,N_10367,N_10131);
and U10767 (N_10767,N_10432,N_10014);
nand U10768 (N_10768,N_10213,N_10208);
xor U10769 (N_10769,N_10498,N_10474);
nor U10770 (N_10770,N_10245,N_10498);
xnor U10771 (N_10771,N_10130,N_10049);
xnor U10772 (N_10772,N_10271,N_10158);
or U10773 (N_10773,N_10036,N_10455);
or U10774 (N_10774,N_10372,N_10366);
or U10775 (N_10775,N_10420,N_10077);
xnor U10776 (N_10776,N_10159,N_10068);
nor U10777 (N_10777,N_10327,N_10039);
or U10778 (N_10778,N_10305,N_10370);
and U10779 (N_10779,N_10491,N_10083);
xnor U10780 (N_10780,N_10071,N_10452);
xor U10781 (N_10781,N_10177,N_10336);
or U10782 (N_10782,N_10038,N_10000);
xnor U10783 (N_10783,N_10472,N_10057);
nor U10784 (N_10784,N_10090,N_10156);
and U10785 (N_10785,N_10104,N_10362);
and U10786 (N_10786,N_10058,N_10340);
nand U10787 (N_10787,N_10026,N_10387);
and U10788 (N_10788,N_10054,N_10115);
nor U10789 (N_10789,N_10238,N_10242);
or U10790 (N_10790,N_10290,N_10412);
nand U10791 (N_10791,N_10420,N_10129);
xnor U10792 (N_10792,N_10090,N_10086);
nand U10793 (N_10793,N_10151,N_10257);
nand U10794 (N_10794,N_10312,N_10498);
nor U10795 (N_10795,N_10434,N_10035);
or U10796 (N_10796,N_10008,N_10101);
xnor U10797 (N_10797,N_10381,N_10286);
or U10798 (N_10798,N_10227,N_10112);
xor U10799 (N_10799,N_10073,N_10454);
xnor U10800 (N_10800,N_10216,N_10077);
and U10801 (N_10801,N_10389,N_10341);
xor U10802 (N_10802,N_10414,N_10494);
nor U10803 (N_10803,N_10172,N_10428);
or U10804 (N_10804,N_10305,N_10076);
or U10805 (N_10805,N_10228,N_10036);
nand U10806 (N_10806,N_10014,N_10375);
nand U10807 (N_10807,N_10259,N_10375);
nor U10808 (N_10808,N_10447,N_10424);
or U10809 (N_10809,N_10481,N_10328);
nor U10810 (N_10810,N_10344,N_10055);
and U10811 (N_10811,N_10416,N_10287);
and U10812 (N_10812,N_10151,N_10150);
or U10813 (N_10813,N_10413,N_10205);
and U10814 (N_10814,N_10153,N_10272);
nor U10815 (N_10815,N_10326,N_10063);
nor U10816 (N_10816,N_10066,N_10397);
and U10817 (N_10817,N_10060,N_10431);
xor U10818 (N_10818,N_10015,N_10228);
nand U10819 (N_10819,N_10460,N_10370);
or U10820 (N_10820,N_10487,N_10039);
and U10821 (N_10821,N_10260,N_10326);
and U10822 (N_10822,N_10096,N_10155);
nand U10823 (N_10823,N_10125,N_10463);
or U10824 (N_10824,N_10001,N_10315);
xor U10825 (N_10825,N_10225,N_10464);
and U10826 (N_10826,N_10094,N_10375);
nor U10827 (N_10827,N_10286,N_10465);
nor U10828 (N_10828,N_10316,N_10383);
xnor U10829 (N_10829,N_10329,N_10119);
nor U10830 (N_10830,N_10259,N_10272);
or U10831 (N_10831,N_10188,N_10306);
and U10832 (N_10832,N_10162,N_10198);
and U10833 (N_10833,N_10327,N_10360);
and U10834 (N_10834,N_10490,N_10345);
nand U10835 (N_10835,N_10267,N_10452);
xnor U10836 (N_10836,N_10235,N_10309);
xnor U10837 (N_10837,N_10019,N_10394);
or U10838 (N_10838,N_10456,N_10073);
nor U10839 (N_10839,N_10375,N_10386);
and U10840 (N_10840,N_10308,N_10196);
or U10841 (N_10841,N_10276,N_10280);
and U10842 (N_10842,N_10435,N_10007);
and U10843 (N_10843,N_10092,N_10432);
and U10844 (N_10844,N_10113,N_10026);
nand U10845 (N_10845,N_10232,N_10445);
nand U10846 (N_10846,N_10422,N_10142);
and U10847 (N_10847,N_10247,N_10384);
nor U10848 (N_10848,N_10108,N_10286);
nand U10849 (N_10849,N_10050,N_10275);
xor U10850 (N_10850,N_10412,N_10488);
xnor U10851 (N_10851,N_10399,N_10300);
xor U10852 (N_10852,N_10144,N_10311);
xor U10853 (N_10853,N_10415,N_10068);
or U10854 (N_10854,N_10422,N_10480);
nand U10855 (N_10855,N_10496,N_10002);
nand U10856 (N_10856,N_10362,N_10303);
nor U10857 (N_10857,N_10019,N_10454);
xor U10858 (N_10858,N_10402,N_10383);
nor U10859 (N_10859,N_10150,N_10024);
xnor U10860 (N_10860,N_10130,N_10368);
xor U10861 (N_10861,N_10078,N_10051);
nor U10862 (N_10862,N_10279,N_10428);
nor U10863 (N_10863,N_10077,N_10335);
nand U10864 (N_10864,N_10224,N_10259);
or U10865 (N_10865,N_10173,N_10138);
nand U10866 (N_10866,N_10057,N_10329);
and U10867 (N_10867,N_10123,N_10104);
nor U10868 (N_10868,N_10007,N_10186);
and U10869 (N_10869,N_10088,N_10143);
or U10870 (N_10870,N_10313,N_10061);
nor U10871 (N_10871,N_10242,N_10308);
nand U10872 (N_10872,N_10242,N_10270);
xnor U10873 (N_10873,N_10013,N_10105);
nand U10874 (N_10874,N_10147,N_10004);
nor U10875 (N_10875,N_10425,N_10415);
and U10876 (N_10876,N_10047,N_10378);
nand U10877 (N_10877,N_10006,N_10327);
or U10878 (N_10878,N_10266,N_10459);
nor U10879 (N_10879,N_10484,N_10068);
nor U10880 (N_10880,N_10056,N_10298);
or U10881 (N_10881,N_10413,N_10487);
nand U10882 (N_10882,N_10438,N_10263);
nor U10883 (N_10883,N_10067,N_10136);
nor U10884 (N_10884,N_10072,N_10165);
xor U10885 (N_10885,N_10061,N_10240);
nand U10886 (N_10886,N_10206,N_10130);
nand U10887 (N_10887,N_10199,N_10135);
and U10888 (N_10888,N_10007,N_10415);
xor U10889 (N_10889,N_10222,N_10293);
xnor U10890 (N_10890,N_10347,N_10145);
xor U10891 (N_10891,N_10120,N_10269);
xor U10892 (N_10892,N_10301,N_10137);
and U10893 (N_10893,N_10211,N_10422);
or U10894 (N_10894,N_10405,N_10094);
or U10895 (N_10895,N_10387,N_10187);
nor U10896 (N_10896,N_10404,N_10169);
nor U10897 (N_10897,N_10058,N_10068);
xor U10898 (N_10898,N_10324,N_10354);
nand U10899 (N_10899,N_10362,N_10105);
nand U10900 (N_10900,N_10316,N_10095);
nor U10901 (N_10901,N_10393,N_10241);
or U10902 (N_10902,N_10012,N_10062);
or U10903 (N_10903,N_10476,N_10061);
nor U10904 (N_10904,N_10163,N_10169);
nor U10905 (N_10905,N_10309,N_10102);
nor U10906 (N_10906,N_10443,N_10275);
nand U10907 (N_10907,N_10422,N_10265);
xor U10908 (N_10908,N_10262,N_10441);
nand U10909 (N_10909,N_10474,N_10304);
nand U10910 (N_10910,N_10490,N_10200);
or U10911 (N_10911,N_10314,N_10382);
nand U10912 (N_10912,N_10112,N_10118);
or U10913 (N_10913,N_10344,N_10108);
and U10914 (N_10914,N_10458,N_10359);
nand U10915 (N_10915,N_10225,N_10369);
nand U10916 (N_10916,N_10043,N_10426);
nand U10917 (N_10917,N_10349,N_10479);
xor U10918 (N_10918,N_10390,N_10108);
and U10919 (N_10919,N_10083,N_10335);
or U10920 (N_10920,N_10256,N_10248);
and U10921 (N_10921,N_10069,N_10163);
or U10922 (N_10922,N_10142,N_10359);
nor U10923 (N_10923,N_10296,N_10125);
nand U10924 (N_10924,N_10164,N_10182);
or U10925 (N_10925,N_10318,N_10293);
nor U10926 (N_10926,N_10044,N_10028);
nor U10927 (N_10927,N_10411,N_10183);
nor U10928 (N_10928,N_10117,N_10422);
xnor U10929 (N_10929,N_10396,N_10193);
nor U10930 (N_10930,N_10082,N_10418);
and U10931 (N_10931,N_10029,N_10230);
nor U10932 (N_10932,N_10243,N_10417);
nand U10933 (N_10933,N_10091,N_10266);
nand U10934 (N_10934,N_10104,N_10120);
or U10935 (N_10935,N_10426,N_10428);
xnor U10936 (N_10936,N_10238,N_10231);
xor U10937 (N_10937,N_10371,N_10063);
or U10938 (N_10938,N_10186,N_10051);
nand U10939 (N_10939,N_10168,N_10482);
nand U10940 (N_10940,N_10280,N_10467);
and U10941 (N_10941,N_10243,N_10316);
or U10942 (N_10942,N_10416,N_10245);
or U10943 (N_10943,N_10329,N_10169);
or U10944 (N_10944,N_10010,N_10447);
and U10945 (N_10945,N_10329,N_10297);
nor U10946 (N_10946,N_10182,N_10372);
or U10947 (N_10947,N_10329,N_10160);
and U10948 (N_10948,N_10197,N_10006);
nand U10949 (N_10949,N_10225,N_10195);
and U10950 (N_10950,N_10442,N_10343);
nor U10951 (N_10951,N_10490,N_10212);
or U10952 (N_10952,N_10200,N_10418);
nor U10953 (N_10953,N_10488,N_10403);
or U10954 (N_10954,N_10366,N_10294);
or U10955 (N_10955,N_10449,N_10111);
or U10956 (N_10956,N_10172,N_10102);
xor U10957 (N_10957,N_10374,N_10108);
xnor U10958 (N_10958,N_10152,N_10277);
xor U10959 (N_10959,N_10173,N_10072);
nand U10960 (N_10960,N_10367,N_10446);
nand U10961 (N_10961,N_10072,N_10381);
nor U10962 (N_10962,N_10158,N_10345);
nand U10963 (N_10963,N_10307,N_10103);
xor U10964 (N_10964,N_10086,N_10159);
nand U10965 (N_10965,N_10014,N_10019);
and U10966 (N_10966,N_10082,N_10055);
nor U10967 (N_10967,N_10090,N_10046);
xnor U10968 (N_10968,N_10244,N_10344);
nand U10969 (N_10969,N_10141,N_10171);
nor U10970 (N_10970,N_10058,N_10038);
and U10971 (N_10971,N_10149,N_10369);
and U10972 (N_10972,N_10356,N_10487);
nor U10973 (N_10973,N_10263,N_10233);
and U10974 (N_10974,N_10305,N_10259);
and U10975 (N_10975,N_10002,N_10024);
nor U10976 (N_10976,N_10076,N_10078);
and U10977 (N_10977,N_10366,N_10133);
nand U10978 (N_10978,N_10101,N_10372);
xnor U10979 (N_10979,N_10132,N_10267);
xnor U10980 (N_10980,N_10252,N_10232);
xnor U10981 (N_10981,N_10349,N_10402);
and U10982 (N_10982,N_10318,N_10111);
nand U10983 (N_10983,N_10202,N_10402);
nand U10984 (N_10984,N_10215,N_10432);
xor U10985 (N_10985,N_10343,N_10063);
xnor U10986 (N_10986,N_10399,N_10481);
xor U10987 (N_10987,N_10372,N_10274);
nor U10988 (N_10988,N_10389,N_10419);
and U10989 (N_10989,N_10025,N_10290);
or U10990 (N_10990,N_10054,N_10472);
xor U10991 (N_10991,N_10310,N_10271);
or U10992 (N_10992,N_10300,N_10079);
nor U10993 (N_10993,N_10098,N_10471);
and U10994 (N_10994,N_10350,N_10124);
xnor U10995 (N_10995,N_10429,N_10046);
or U10996 (N_10996,N_10477,N_10445);
or U10997 (N_10997,N_10228,N_10214);
or U10998 (N_10998,N_10061,N_10222);
nor U10999 (N_10999,N_10204,N_10174);
or U11000 (N_11000,N_10723,N_10627);
xnor U11001 (N_11001,N_10527,N_10854);
and U11002 (N_11002,N_10639,N_10594);
or U11003 (N_11003,N_10550,N_10937);
xor U11004 (N_11004,N_10735,N_10941);
nor U11005 (N_11005,N_10544,N_10910);
nand U11006 (N_11006,N_10727,N_10912);
nor U11007 (N_11007,N_10645,N_10672);
and U11008 (N_11008,N_10537,N_10909);
nor U11009 (N_11009,N_10922,N_10644);
or U11010 (N_11010,N_10536,N_10541);
nor U11011 (N_11011,N_10923,N_10835);
or U11012 (N_11012,N_10695,N_10751);
nand U11013 (N_11013,N_10606,N_10888);
nand U11014 (N_11014,N_10913,N_10970);
nand U11015 (N_11015,N_10980,N_10688);
or U11016 (N_11016,N_10915,N_10685);
nand U11017 (N_11017,N_10809,N_10953);
xnor U11018 (N_11018,N_10858,N_10676);
nand U11019 (N_11019,N_10559,N_10729);
nand U11020 (N_11020,N_10956,N_10767);
nor U11021 (N_11021,N_10991,N_10518);
xor U11022 (N_11022,N_10692,N_10907);
nand U11023 (N_11023,N_10833,N_10571);
or U11024 (N_11024,N_10959,N_10505);
nor U11025 (N_11025,N_10648,N_10955);
xor U11026 (N_11026,N_10531,N_10696);
nor U11027 (N_11027,N_10812,N_10849);
or U11028 (N_11028,N_10581,N_10707);
nor U11029 (N_11029,N_10971,N_10660);
or U11030 (N_11030,N_10656,N_10629);
nor U11031 (N_11031,N_10958,N_10820);
nor U11032 (N_11032,N_10508,N_10891);
xnor U11033 (N_11033,N_10690,N_10788);
nor U11034 (N_11034,N_10616,N_10902);
nor U11035 (N_11035,N_10929,N_10947);
xor U11036 (N_11036,N_10700,N_10732);
and U11037 (N_11037,N_10600,N_10946);
nor U11038 (N_11038,N_10532,N_10609);
and U11039 (N_11039,N_10620,N_10617);
nand U11040 (N_11040,N_10844,N_10549);
xnor U11041 (N_11041,N_10869,N_10967);
and U11042 (N_11042,N_10733,N_10813);
xor U11043 (N_11043,N_10799,N_10899);
or U11044 (N_11044,N_10740,N_10882);
xnor U11045 (N_11045,N_10914,N_10574);
nand U11046 (N_11046,N_10597,N_10837);
nor U11047 (N_11047,N_10974,N_10989);
xor U11048 (N_11048,N_10784,N_10699);
nand U11049 (N_11049,N_10534,N_10624);
xnor U11050 (N_11050,N_10916,N_10755);
nand U11051 (N_11051,N_10719,N_10934);
nor U11052 (N_11052,N_10932,N_10528);
and U11053 (N_11053,N_10758,N_10502);
or U11054 (N_11054,N_10826,N_10779);
and U11055 (N_11055,N_10636,N_10730);
xor U11056 (N_11056,N_10984,N_10529);
nand U11057 (N_11057,N_10972,N_10569);
nor U11058 (N_11058,N_10840,N_10865);
nand U11059 (N_11059,N_10515,N_10674);
nor U11060 (N_11060,N_10710,N_10681);
nor U11061 (N_11061,N_10982,N_10880);
nor U11062 (N_11062,N_10641,N_10560);
xnor U11063 (N_11063,N_10774,N_10669);
nor U11064 (N_11064,N_10811,N_10592);
nand U11065 (N_11065,N_10966,N_10975);
xnor U11066 (N_11066,N_10708,N_10514);
and U11067 (N_11067,N_10583,N_10563);
xnor U11068 (N_11068,N_10731,N_10516);
nand U11069 (N_11069,N_10649,N_10717);
and U11070 (N_11070,N_10737,N_10501);
nor U11071 (N_11071,N_10872,N_10714);
and U11072 (N_11072,N_10679,N_10653);
nand U11073 (N_11073,N_10761,N_10911);
nand U11074 (N_11074,N_10698,N_10530);
or U11075 (N_11075,N_10783,N_10803);
xnor U11076 (N_11076,N_10513,N_10861);
and U11077 (N_11077,N_10847,N_10568);
or U11078 (N_11078,N_10703,N_10709);
nor U11079 (N_11079,N_10855,N_10757);
or U11080 (N_11080,N_10687,N_10931);
or U11081 (N_11081,N_10793,N_10866);
xor U11082 (N_11082,N_10603,N_10651);
nor U11083 (N_11083,N_10945,N_10743);
xnor U11084 (N_11084,N_10762,N_10851);
xor U11085 (N_11085,N_10815,N_10814);
nor U11086 (N_11086,N_10673,N_10852);
nor U11087 (N_11087,N_10924,N_10631);
nand U11088 (N_11088,N_10565,N_10765);
and U11089 (N_11089,N_10684,N_10566);
or U11090 (N_11090,N_10705,N_10990);
or U11091 (N_11091,N_10776,N_10864);
and U11092 (N_11092,N_10857,N_10867);
nand U11093 (N_11093,N_10800,N_10634);
nand U11094 (N_11094,N_10968,N_10877);
xor U11095 (N_11095,N_10570,N_10780);
or U11096 (N_11096,N_10768,N_10633);
nor U11097 (N_11097,N_10587,N_10547);
xor U11098 (N_11098,N_10591,N_10831);
or U11099 (N_11099,N_10667,N_10960);
or U11100 (N_11100,N_10706,N_10938);
nor U11101 (N_11101,N_10578,N_10944);
and U11102 (N_11102,N_10825,N_10658);
or U11103 (N_11103,N_10678,N_10846);
and U11104 (N_11104,N_10621,N_10903);
or U11105 (N_11105,N_10638,N_10567);
nand U11106 (N_11106,N_10610,N_10790);
nor U11107 (N_11107,N_10810,N_10662);
and U11108 (N_11108,N_10808,N_10954);
xor U11109 (N_11109,N_10511,N_10900);
nand U11110 (N_11110,N_10650,N_10716);
and U11111 (N_11111,N_10613,N_10963);
and U11112 (N_11112,N_10804,N_10786);
nor U11113 (N_11113,N_10670,N_10734);
and U11114 (N_11114,N_10775,N_10712);
xor U11115 (N_11115,N_10564,N_10794);
nand U11116 (N_11116,N_10618,N_10874);
xor U11117 (N_11117,N_10722,N_10890);
or U11118 (N_11118,N_10666,N_10647);
xnor U11119 (N_11119,N_10682,N_10871);
xnor U11120 (N_11120,N_10595,N_10576);
xor U11121 (N_11121,N_10646,N_10770);
or U11122 (N_11122,N_10976,N_10512);
and U11123 (N_11123,N_10680,N_10841);
and U11124 (N_11124,N_10842,N_10985);
nor U11125 (N_11125,N_10950,N_10961);
xor U11126 (N_11126,N_10773,N_10948);
nand U11127 (N_11127,N_10573,N_10893);
and U11128 (N_11128,N_10883,N_10701);
nor U11129 (N_11129,N_10589,N_10664);
and U11130 (N_11130,N_10500,N_10721);
nor U11131 (N_11131,N_10796,N_10885);
nor U11132 (N_11132,N_10523,N_10599);
or U11133 (N_11133,N_10720,N_10898);
or U11134 (N_11134,N_10821,N_10605);
nor U11135 (N_11135,N_10896,N_10818);
nor U11136 (N_11136,N_10764,N_10715);
nor U11137 (N_11137,N_10643,N_10601);
and U11138 (N_11138,N_10983,N_10817);
xor U11139 (N_11139,N_10632,N_10965);
and U11140 (N_11140,N_10894,N_10957);
xnor U11141 (N_11141,N_10797,N_10736);
nand U11142 (N_11142,N_10521,N_10901);
nand U11143 (N_11143,N_10718,N_10756);
nor U11144 (N_11144,N_10942,N_10819);
or U11145 (N_11145,N_10691,N_10824);
and U11146 (N_11146,N_10742,N_10652);
and U11147 (N_11147,N_10782,N_10747);
nor U11148 (N_11148,N_10791,N_10522);
and U11149 (N_11149,N_10711,N_10969);
or U11150 (N_11150,N_10943,N_10839);
or U11151 (N_11151,N_10655,N_10873);
and U11152 (N_11152,N_10580,N_10921);
nor U11153 (N_11153,N_10579,N_10752);
nor U11154 (N_11154,N_10848,N_10986);
xor U11155 (N_11155,N_10623,N_10952);
and U11156 (N_11156,N_10746,N_10769);
nor U11157 (N_11157,N_10551,N_10917);
nor U11158 (N_11158,N_10509,N_10807);
and U11159 (N_11159,N_10978,N_10889);
xor U11160 (N_11160,N_10642,N_10683);
xor U11161 (N_11161,N_10671,N_10798);
or U11162 (N_11162,N_10608,N_10895);
and U11163 (N_11163,N_10908,N_10507);
or U11164 (N_11164,N_10728,N_10704);
nand U11165 (N_11165,N_10850,N_10843);
xor U11166 (N_11166,N_10801,N_10859);
and U11167 (N_11167,N_10754,N_10926);
nand U11168 (N_11168,N_10881,N_10753);
and U11169 (N_11169,N_10677,N_10935);
nand U11170 (N_11170,N_10979,N_10879);
nand U11171 (N_11171,N_10602,N_10545);
xnor U11172 (N_11172,N_10919,N_10830);
or U11173 (N_11173,N_10654,N_10561);
nand U11174 (N_11174,N_10853,N_10862);
and U11175 (N_11175,N_10637,N_10834);
nor U11176 (N_11176,N_10822,N_10998);
and U11177 (N_11177,N_10665,N_10795);
nand U11178 (N_11178,N_10689,N_10539);
and U11179 (N_11179,N_10845,N_10738);
nor U11180 (N_11180,N_10763,N_10713);
or U11181 (N_11181,N_10994,N_10504);
or U11182 (N_11182,N_10556,N_10546);
nor U11183 (N_11183,N_10977,N_10607);
and U11184 (N_11184,N_10870,N_10816);
nor U11185 (N_11185,N_10925,N_10771);
or U11186 (N_11186,N_10598,N_10897);
nor U11187 (N_11187,N_10586,N_10951);
nand U11188 (N_11188,N_10535,N_10611);
nor U11189 (N_11189,N_10829,N_10884);
xnor U11190 (N_11190,N_10878,N_10694);
nor U11191 (N_11191,N_10787,N_10887);
nand U11192 (N_11192,N_10619,N_10973);
nand U11193 (N_11193,N_10554,N_10996);
and U11194 (N_11194,N_10558,N_10675);
nand U11195 (N_11195,N_10792,N_10918);
and U11196 (N_11196,N_10992,N_10823);
xor U11197 (N_11197,N_10997,N_10805);
and U11198 (N_11198,N_10772,N_10593);
nor U11199 (N_11199,N_10744,N_10749);
and U11200 (N_11200,N_10748,N_10868);
xnor U11201 (N_11201,N_10920,N_10590);
nand U11202 (N_11202,N_10741,N_10860);
nor U11203 (N_11203,N_10630,N_10588);
nor U11204 (N_11204,N_10614,N_10940);
nand U11205 (N_11205,N_10999,N_10572);
or U11206 (N_11206,N_10726,N_10828);
nand U11207 (N_11207,N_10936,N_10577);
nor U11208 (N_11208,N_10886,N_10856);
nand U11209 (N_11209,N_10686,N_10927);
xor U11210 (N_11210,N_10640,N_10585);
and U11211 (N_11211,N_10596,N_10553);
and U11212 (N_11212,N_10663,N_10557);
or U11213 (N_11213,N_10939,N_10766);
nor U11214 (N_11214,N_10933,N_10668);
or U11215 (N_11215,N_10949,N_10702);
nor U11216 (N_11216,N_10802,N_10785);
nor U11217 (N_11217,N_10838,N_10575);
nor U11218 (N_11218,N_10964,N_10836);
nand U11219 (N_11219,N_10993,N_10987);
or U11220 (N_11220,N_10533,N_10612);
nor U11221 (N_11221,N_10981,N_10777);
xnor U11222 (N_11222,N_10584,N_10930);
or U11223 (N_11223,N_10863,N_10506);
nand U11224 (N_11224,N_10759,N_10520);
and U11225 (N_11225,N_10626,N_10615);
xnor U11226 (N_11226,N_10745,N_10503);
or U11227 (N_11227,N_10739,N_10542);
and U11228 (N_11228,N_10995,N_10906);
or U11229 (N_11229,N_10517,N_10778);
nand U11230 (N_11230,N_10827,N_10832);
nor U11231 (N_11231,N_10693,N_10548);
and U11232 (N_11232,N_10635,N_10525);
or U11233 (N_11233,N_10806,N_10555);
xnor U11234 (N_11234,N_10582,N_10526);
nor U11235 (N_11235,N_10876,N_10519);
or U11236 (N_11236,N_10725,N_10928);
nand U11237 (N_11237,N_10750,N_10628);
or U11238 (N_11238,N_10697,N_10892);
xor U11239 (N_11239,N_10904,N_10604);
or U11240 (N_11240,N_10552,N_10657);
and U11241 (N_11241,N_10622,N_10724);
nor U11242 (N_11242,N_10538,N_10562);
xor U11243 (N_11243,N_10781,N_10875);
and U11244 (N_11244,N_10510,N_10905);
or U11245 (N_11245,N_10543,N_10524);
or U11246 (N_11246,N_10659,N_10540);
nor U11247 (N_11247,N_10760,N_10661);
nor U11248 (N_11248,N_10789,N_10625);
or U11249 (N_11249,N_10962,N_10988);
or U11250 (N_11250,N_10938,N_10953);
nand U11251 (N_11251,N_10716,N_10879);
and U11252 (N_11252,N_10564,N_10558);
xor U11253 (N_11253,N_10694,N_10917);
nor U11254 (N_11254,N_10528,N_10653);
and U11255 (N_11255,N_10775,N_10910);
nand U11256 (N_11256,N_10512,N_10803);
nor U11257 (N_11257,N_10551,N_10665);
or U11258 (N_11258,N_10665,N_10782);
xor U11259 (N_11259,N_10821,N_10918);
and U11260 (N_11260,N_10643,N_10852);
nor U11261 (N_11261,N_10576,N_10721);
or U11262 (N_11262,N_10514,N_10917);
nor U11263 (N_11263,N_10784,N_10635);
or U11264 (N_11264,N_10575,N_10501);
nand U11265 (N_11265,N_10549,N_10696);
nand U11266 (N_11266,N_10684,N_10673);
xnor U11267 (N_11267,N_10867,N_10676);
and U11268 (N_11268,N_10607,N_10881);
nor U11269 (N_11269,N_10740,N_10662);
nand U11270 (N_11270,N_10917,N_10563);
nand U11271 (N_11271,N_10696,N_10819);
xnor U11272 (N_11272,N_10769,N_10601);
xor U11273 (N_11273,N_10963,N_10628);
and U11274 (N_11274,N_10960,N_10673);
and U11275 (N_11275,N_10997,N_10598);
xor U11276 (N_11276,N_10730,N_10500);
or U11277 (N_11277,N_10791,N_10529);
and U11278 (N_11278,N_10501,N_10551);
nor U11279 (N_11279,N_10900,N_10877);
and U11280 (N_11280,N_10681,N_10777);
and U11281 (N_11281,N_10603,N_10768);
or U11282 (N_11282,N_10746,N_10890);
xnor U11283 (N_11283,N_10558,N_10695);
xor U11284 (N_11284,N_10734,N_10729);
nor U11285 (N_11285,N_10922,N_10666);
and U11286 (N_11286,N_10663,N_10543);
xor U11287 (N_11287,N_10727,N_10743);
and U11288 (N_11288,N_10818,N_10762);
nand U11289 (N_11289,N_10572,N_10588);
xnor U11290 (N_11290,N_10861,N_10818);
and U11291 (N_11291,N_10615,N_10788);
nor U11292 (N_11292,N_10644,N_10784);
nand U11293 (N_11293,N_10625,N_10861);
nand U11294 (N_11294,N_10558,N_10742);
nand U11295 (N_11295,N_10633,N_10524);
nand U11296 (N_11296,N_10709,N_10917);
xor U11297 (N_11297,N_10642,N_10860);
nor U11298 (N_11298,N_10696,N_10609);
and U11299 (N_11299,N_10683,N_10863);
xor U11300 (N_11300,N_10790,N_10827);
xor U11301 (N_11301,N_10958,N_10776);
nand U11302 (N_11302,N_10582,N_10782);
or U11303 (N_11303,N_10910,N_10932);
nand U11304 (N_11304,N_10766,N_10773);
nand U11305 (N_11305,N_10860,N_10995);
or U11306 (N_11306,N_10951,N_10718);
or U11307 (N_11307,N_10707,N_10679);
xor U11308 (N_11308,N_10945,N_10885);
nand U11309 (N_11309,N_10705,N_10929);
xnor U11310 (N_11310,N_10751,N_10569);
or U11311 (N_11311,N_10748,N_10955);
xor U11312 (N_11312,N_10555,N_10683);
or U11313 (N_11313,N_10617,N_10535);
xor U11314 (N_11314,N_10569,N_10694);
or U11315 (N_11315,N_10817,N_10866);
and U11316 (N_11316,N_10863,N_10571);
or U11317 (N_11317,N_10919,N_10573);
xnor U11318 (N_11318,N_10579,N_10743);
and U11319 (N_11319,N_10777,N_10970);
nand U11320 (N_11320,N_10771,N_10998);
nand U11321 (N_11321,N_10500,N_10719);
and U11322 (N_11322,N_10736,N_10908);
xor U11323 (N_11323,N_10923,N_10799);
nor U11324 (N_11324,N_10962,N_10558);
nand U11325 (N_11325,N_10901,N_10896);
and U11326 (N_11326,N_10545,N_10842);
xnor U11327 (N_11327,N_10766,N_10554);
or U11328 (N_11328,N_10764,N_10763);
and U11329 (N_11329,N_10605,N_10786);
or U11330 (N_11330,N_10765,N_10885);
or U11331 (N_11331,N_10986,N_10895);
and U11332 (N_11332,N_10753,N_10792);
nand U11333 (N_11333,N_10665,N_10873);
or U11334 (N_11334,N_10930,N_10705);
xor U11335 (N_11335,N_10734,N_10686);
and U11336 (N_11336,N_10778,N_10509);
xnor U11337 (N_11337,N_10777,N_10866);
and U11338 (N_11338,N_10707,N_10966);
nand U11339 (N_11339,N_10767,N_10691);
or U11340 (N_11340,N_10647,N_10577);
nand U11341 (N_11341,N_10902,N_10819);
nor U11342 (N_11342,N_10536,N_10731);
nand U11343 (N_11343,N_10912,N_10919);
nand U11344 (N_11344,N_10782,N_10911);
xnor U11345 (N_11345,N_10877,N_10944);
nand U11346 (N_11346,N_10915,N_10981);
nand U11347 (N_11347,N_10698,N_10856);
and U11348 (N_11348,N_10768,N_10924);
nor U11349 (N_11349,N_10597,N_10832);
nand U11350 (N_11350,N_10701,N_10924);
xor U11351 (N_11351,N_10552,N_10770);
xor U11352 (N_11352,N_10840,N_10777);
nand U11353 (N_11353,N_10710,N_10798);
xor U11354 (N_11354,N_10502,N_10619);
or U11355 (N_11355,N_10947,N_10823);
nor U11356 (N_11356,N_10879,N_10947);
nor U11357 (N_11357,N_10893,N_10708);
and U11358 (N_11358,N_10548,N_10731);
nand U11359 (N_11359,N_10648,N_10886);
nand U11360 (N_11360,N_10807,N_10815);
and U11361 (N_11361,N_10712,N_10840);
or U11362 (N_11362,N_10950,N_10838);
nand U11363 (N_11363,N_10871,N_10778);
nor U11364 (N_11364,N_10975,N_10742);
nor U11365 (N_11365,N_10581,N_10761);
nand U11366 (N_11366,N_10875,N_10900);
or U11367 (N_11367,N_10816,N_10616);
and U11368 (N_11368,N_10995,N_10677);
nand U11369 (N_11369,N_10983,N_10876);
xnor U11370 (N_11370,N_10689,N_10662);
or U11371 (N_11371,N_10818,N_10777);
xnor U11372 (N_11372,N_10546,N_10800);
xnor U11373 (N_11373,N_10624,N_10701);
xor U11374 (N_11374,N_10844,N_10829);
nor U11375 (N_11375,N_10786,N_10537);
nor U11376 (N_11376,N_10605,N_10973);
and U11377 (N_11377,N_10591,N_10847);
and U11378 (N_11378,N_10639,N_10999);
nor U11379 (N_11379,N_10807,N_10840);
or U11380 (N_11380,N_10597,N_10539);
nor U11381 (N_11381,N_10658,N_10982);
and U11382 (N_11382,N_10928,N_10558);
or U11383 (N_11383,N_10614,N_10627);
nor U11384 (N_11384,N_10888,N_10713);
xnor U11385 (N_11385,N_10604,N_10755);
and U11386 (N_11386,N_10742,N_10545);
xnor U11387 (N_11387,N_10833,N_10507);
and U11388 (N_11388,N_10831,N_10572);
or U11389 (N_11389,N_10654,N_10659);
and U11390 (N_11390,N_10878,N_10844);
xnor U11391 (N_11391,N_10567,N_10634);
nor U11392 (N_11392,N_10595,N_10837);
or U11393 (N_11393,N_10597,N_10972);
nand U11394 (N_11394,N_10712,N_10536);
and U11395 (N_11395,N_10578,N_10706);
nand U11396 (N_11396,N_10702,N_10844);
nand U11397 (N_11397,N_10798,N_10748);
or U11398 (N_11398,N_10768,N_10719);
and U11399 (N_11399,N_10945,N_10555);
or U11400 (N_11400,N_10926,N_10634);
and U11401 (N_11401,N_10968,N_10618);
and U11402 (N_11402,N_10764,N_10560);
nand U11403 (N_11403,N_10708,N_10540);
or U11404 (N_11404,N_10536,N_10555);
nor U11405 (N_11405,N_10664,N_10791);
or U11406 (N_11406,N_10750,N_10888);
nor U11407 (N_11407,N_10786,N_10597);
and U11408 (N_11408,N_10835,N_10530);
xor U11409 (N_11409,N_10705,N_10845);
nor U11410 (N_11410,N_10821,N_10743);
nor U11411 (N_11411,N_10831,N_10631);
xnor U11412 (N_11412,N_10706,N_10963);
nand U11413 (N_11413,N_10754,N_10947);
xnor U11414 (N_11414,N_10520,N_10548);
or U11415 (N_11415,N_10910,N_10969);
xnor U11416 (N_11416,N_10838,N_10609);
or U11417 (N_11417,N_10931,N_10541);
nand U11418 (N_11418,N_10895,N_10526);
nor U11419 (N_11419,N_10757,N_10847);
xnor U11420 (N_11420,N_10597,N_10925);
or U11421 (N_11421,N_10595,N_10624);
xor U11422 (N_11422,N_10581,N_10510);
and U11423 (N_11423,N_10882,N_10748);
and U11424 (N_11424,N_10953,N_10917);
or U11425 (N_11425,N_10527,N_10961);
xor U11426 (N_11426,N_10772,N_10920);
nand U11427 (N_11427,N_10975,N_10598);
nor U11428 (N_11428,N_10824,N_10794);
and U11429 (N_11429,N_10770,N_10796);
xor U11430 (N_11430,N_10518,N_10654);
nor U11431 (N_11431,N_10721,N_10718);
or U11432 (N_11432,N_10836,N_10586);
and U11433 (N_11433,N_10593,N_10807);
and U11434 (N_11434,N_10541,N_10937);
or U11435 (N_11435,N_10573,N_10900);
or U11436 (N_11436,N_10626,N_10588);
nor U11437 (N_11437,N_10915,N_10521);
nand U11438 (N_11438,N_10856,N_10647);
xor U11439 (N_11439,N_10611,N_10834);
nand U11440 (N_11440,N_10709,N_10860);
nor U11441 (N_11441,N_10728,N_10860);
xnor U11442 (N_11442,N_10542,N_10858);
nor U11443 (N_11443,N_10808,N_10827);
nand U11444 (N_11444,N_10532,N_10735);
nor U11445 (N_11445,N_10907,N_10628);
or U11446 (N_11446,N_10618,N_10522);
nand U11447 (N_11447,N_10696,N_10663);
xor U11448 (N_11448,N_10522,N_10923);
nor U11449 (N_11449,N_10978,N_10880);
and U11450 (N_11450,N_10502,N_10676);
and U11451 (N_11451,N_10558,N_10735);
nand U11452 (N_11452,N_10761,N_10696);
nand U11453 (N_11453,N_10838,N_10608);
or U11454 (N_11454,N_10678,N_10607);
xor U11455 (N_11455,N_10802,N_10584);
nand U11456 (N_11456,N_10951,N_10613);
xor U11457 (N_11457,N_10768,N_10630);
xnor U11458 (N_11458,N_10857,N_10749);
nand U11459 (N_11459,N_10940,N_10996);
nand U11460 (N_11460,N_10810,N_10829);
and U11461 (N_11461,N_10609,N_10957);
nor U11462 (N_11462,N_10611,N_10720);
and U11463 (N_11463,N_10917,N_10594);
nor U11464 (N_11464,N_10782,N_10542);
and U11465 (N_11465,N_10806,N_10621);
nor U11466 (N_11466,N_10501,N_10805);
nand U11467 (N_11467,N_10568,N_10806);
nor U11468 (N_11468,N_10674,N_10610);
nand U11469 (N_11469,N_10592,N_10667);
nand U11470 (N_11470,N_10832,N_10940);
xnor U11471 (N_11471,N_10907,N_10554);
xnor U11472 (N_11472,N_10671,N_10960);
and U11473 (N_11473,N_10534,N_10675);
nand U11474 (N_11474,N_10569,N_10560);
xor U11475 (N_11475,N_10562,N_10777);
or U11476 (N_11476,N_10755,N_10955);
or U11477 (N_11477,N_10504,N_10740);
or U11478 (N_11478,N_10718,N_10551);
nand U11479 (N_11479,N_10720,N_10818);
and U11480 (N_11480,N_10574,N_10866);
and U11481 (N_11481,N_10724,N_10709);
and U11482 (N_11482,N_10559,N_10546);
nor U11483 (N_11483,N_10503,N_10603);
nor U11484 (N_11484,N_10604,N_10817);
and U11485 (N_11485,N_10638,N_10771);
nand U11486 (N_11486,N_10587,N_10676);
xor U11487 (N_11487,N_10890,N_10806);
xnor U11488 (N_11488,N_10953,N_10513);
or U11489 (N_11489,N_10586,N_10915);
xor U11490 (N_11490,N_10700,N_10719);
or U11491 (N_11491,N_10947,N_10536);
and U11492 (N_11492,N_10714,N_10890);
nand U11493 (N_11493,N_10600,N_10632);
nor U11494 (N_11494,N_10984,N_10632);
xor U11495 (N_11495,N_10586,N_10551);
xnor U11496 (N_11496,N_10616,N_10642);
nand U11497 (N_11497,N_10759,N_10776);
nor U11498 (N_11498,N_10945,N_10924);
nand U11499 (N_11499,N_10666,N_10574);
and U11500 (N_11500,N_11457,N_11413);
and U11501 (N_11501,N_11022,N_11133);
and U11502 (N_11502,N_11425,N_11074);
nand U11503 (N_11503,N_11310,N_11161);
and U11504 (N_11504,N_11416,N_11339);
xor U11505 (N_11505,N_11323,N_11103);
and U11506 (N_11506,N_11344,N_11084);
nor U11507 (N_11507,N_11383,N_11153);
nor U11508 (N_11508,N_11246,N_11470);
xor U11509 (N_11509,N_11220,N_11405);
or U11510 (N_11510,N_11267,N_11298);
nor U11511 (N_11511,N_11156,N_11166);
nor U11512 (N_11512,N_11486,N_11420);
nand U11513 (N_11513,N_11483,N_11391);
nand U11514 (N_11514,N_11331,N_11001);
nand U11515 (N_11515,N_11168,N_11337);
or U11516 (N_11516,N_11287,N_11210);
nor U11517 (N_11517,N_11245,N_11414);
and U11518 (N_11518,N_11095,N_11055);
or U11519 (N_11519,N_11169,N_11113);
or U11520 (N_11520,N_11354,N_11250);
or U11521 (N_11521,N_11314,N_11367);
nand U11522 (N_11522,N_11300,N_11372);
xnor U11523 (N_11523,N_11116,N_11124);
nor U11524 (N_11524,N_11408,N_11481);
nand U11525 (N_11525,N_11307,N_11080);
or U11526 (N_11526,N_11233,N_11034);
nand U11527 (N_11527,N_11018,N_11479);
or U11528 (N_11528,N_11332,N_11375);
nor U11529 (N_11529,N_11217,N_11069);
nor U11530 (N_11530,N_11223,N_11144);
xnor U11531 (N_11531,N_11386,N_11378);
xnor U11532 (N_11532,N_11090,N_11057);
or U11533 (N_11533,N_11104,N_11087);
or U11534 (N_11534,N_11007,N_11061);
or U11535 (N_11535,N_11412,N_11119);
xnor U11536 (N_11536,N_11163,N_11361);
nand U11537 (N_11537,N_11053,N_11139);
nand U11538 (N_11538,N_11432,N_11443);
and U11539 (N_11539,N_11140,N_11454);
and U11540 (N_11540,N_11355,N_11302);
or U11541 (N_11541,N_11308,N_11187);
nand U11542 (N_11542,N_11376,N_11464);
or U11543 (N_11543,N_11142,N_11398);
xnor U11544 (N_11544,N_11494,N_11226);
or U11545 (N_11545,N_11474,N_11023);
or U11546 (N_11546,N_11205,N_11134);
or U11547 (N_11547,N_11261,N_11117);
nand U11548 (N_11548,N_11093,N_11241);
or U11549 (N_11549,N_11249,N_11222);
or U11550 (N_11550,N_11326,N_11437);
xnor U11551 (N_11551,N_11237,N_11199);
or U11552 (N_11552,N_11317,N_11050);
nand U11553 (N_11553,N_11268,N_11126);
or U11554 (N_11554,N_11114,N_11440);
or U11555 (N_11555,N_11350,N_11105);
and U11556 (N_11556,N_11145,N_11185);
nand U11557 (N_11557,N_11110,N_11316);
xnor U11558 (N_11558,N_11236,N_11136);
nand U11559 (N_11559,N_11219,N_11147);
or U11560 (N_11560,N_11004,N_11286);
or U11561 (N_11561,N_11348,N_11487);
and U11562 (N_11562,N_11384,N_11043);
nand U11563 (N_11563,N_11044,N_11397);
nor U11564 (N_11564,N_11496,N_11276);
nand U11565 (N_11565,N_11441,N_11107);
and U11566 (N_11566,N_11253,N_11306);
or U11567 (N_11567,N_11434,N_11466);
nor U11568 (N_11568,N_11186,N_11438);
or U11569 (N_11569,N_11002,N_11021);
nor U11570 (N_11570,N_11212,N_11473);
and U11571 (N_11571,N_11225,N_11291);
xnor U11572 (N_11572,N_11164,N_11356);
and U11573 (N_11573,N_11081,N_11431);
and U11574 (N_11574,N_11272,N_11465);
or U11575 (N_11575,N_11131,N_11277);
nor U11576 (N_11576,N_11035,N_11303);
nand U11577 (N_11577,N_11419,N_11146);
xor U11578 (N_11578,N_11099,N_11079);
xnor U11579 (N_11579,N_11138,N_11190);
nand U11580 (N_11580,N_11442,N_11330);
or U11581 (N_11581,N_11343,N_11446);
xor U11582 (N_11582,N_11489,N_11396);
nand U11583 (N_11583,N_11281,N_11058);
and U11584 (N_11584,N_11180,N_11070);
xor U11585 (N_11585,N_11029,N_11322);
or U11586 (N_11586,N_11135,N_11448);
nor U11587 (N_11587,N_11160,N_11294);
nor U11588 (N_11588,N_11423,N_11275);
or U11589 (N_11589,N_11215,N_11141);
nand U11590 (N_11590,N_11410,N_11313);
or U11591 (N_11591,N_11468,N_11014);
nand U11592 (N_11592,N_11013,N_11488);
xnor U11593 (N_11593,N_11255,N_11174);
and U11594 (N_11594,N_11240,N_11497);
or U11595 (N_11595,N_11498,N_11078);
and U11596 (N_11596,N_11439,N_11399);
xnor U11597 (N_11597,N_11201,N_11365);
nand U11598 (N_11598,N_11243,N_11274);
xnor U11599 (N_11599,N_11123,N_11336);
nor U11600 (N_11600,N_11094,N_11312);
or U11601 (N_11601,N_11183,N_11129);
and U11602 (N_11602,N_11400,N_11435);
or U11603 (N_11603,N_11216,N_11230);
or U11604 (N_11604,N_11289,N_11171);
and U11605 (N_11605,N_11132,N_11284);
nor U11606 (N_11606,N_11453,N_11430);
or U11607 (N_11607,N_11182,N_11092);
and U11608 (N_11608,N_11064,N_11460);
and U11609 (N_11609,N_11278,N_11211);
xor U11610 (N_11610,N_11292,N_11197);
nand U11611 (N_11611,N_11387,N_11444);
nor U11612 (N_11612,N_11328,N_11042);
or U11613 (N_11613,N_11194,N_11121);
xor U11614 (N_11614,N_11088,N_11297);
nand U11615 (N_11615,N_11020,N_11130);
or U11616 (N_11616,N_11478,N_11347);
or U11617 (N_11617,N_11491,N_11429);
nand U11618 (N_11618,N_11380,N_11385);
xnor U11619 (N_11619,N_11016,N_11056);
nor U11620 (N_11620,N_11046,N_11063);
xnor U11621 (N_11621,N_11327,N_11005);
or U11622 (N_11622,N_11177,N_11433);
nor U11623 (N_11623,N_11493,N_11279);
or U11624 (N_11624,N_11196,N_11159);
xor U11625 (N_11625,N_11207,N_11083);
and U11626 (N_11626,N_11321,N_11204);
nor U11627 (N_11627,N_11041,N_11009);
nor U11628 (N_11628,N_11340,N_11049);
nor U11629 (N_11629,N_11394,N_11024);
xor U11630 (N_11630,N_11106,N_11428);
or U11631 (N_11631,N_11127,N_11232);
nor U11632 (N_11632,N_11086,N_11172);
nor U11633 (N_11633,N_11052,N_11238);
nand U11634 (N_11634,N_11368,N_11477);
nand U11635 (N_11635,N_11112,N_11346);
nor U11636 (N_11636,N_11102,N_11319);
xnor U11637 (N_11637,N_11320,N_11381);
nand U11638 (N_11638,N_11451,N_11032);
and U11639 (N_11639,N_11234,N_11068);
or U11640 (N_11640,N_11198,N_11072);
nor U11641 (N_11641,N_11100,N_11262);
nand U11642 (N_11642,N_11341,N_11475);
and U11643 (N_11643,N_11436,N_11089);
xnor U11644 (N_11644,N_11170,N_11309);
nand U11645 (N_11645,N_11143,N_11445);
nand U11646 (N_11646,N_11158,N_11036);
nor U11647 (N_11647,N_11273,N_11244);
and U11648 (N_11648,N_11352,N_11388);
or U11649 (N_11649,N_11259,N_11415);
and U11650 (N_11650,N_11192,N_11155);
xor U11651 (N_11651,N_11299,N_11362);
or U11652 (N_11652,N_11040,N_11382);
and U11653 (N_11653,N_11150,N_11252);
xnor U11654 (N_11654,N_11333,N_11390);
xor U11655 (N_11655,N_11358,N_11345);
nand U11656 (N_11656,N_11426,N_11162);
nand U11657 (N_11657,N_11359,N_11165);
or U11658 (N_11658,N_11447,N_11045);
or U11659 (N_11659,N_11048,N_11221);
and U11660 (N_11660,N_11418,N_11173);
or U11661 (N_11661,N_11424,N_11176);
xor U11662 (N_11662,N_11097,N_11118);
nand U11663 (N_11663,N_11421,N_11269);
xnor U11664 (N_11664,N_11490,N_11366);
nand U11665 (N_11665,N_11265,N_11285);
or U11666 (N_11666,N_11349,N_11256);
nand U11667 (N_11667,N_11461,N_11282);
nand U11668 (N_11668,N_11293,N_11311);
or U11669 (N_11669,N_11015,N_11109);
xnor U11670 (N_11670,N_11059,N_11247);
xor U11671 (N_11671,N_11357,N_11266);
xor U11672 (N_11672,N_11037,N_11363);
nor U11673 (N_11673,N_11324,N_11301);
nor U11674 (N_11674,N_11377,N_11149);
nor U11675 (N_11675,N_11122,N_11373);
or U11676 (N_11676,N_11404,N_11334);
nor U11677 (N_11677,N_11427,N_11492);
or U11678 (N_11678,N_11148,N_11325);
nand U11679 (N_11679,N_11076,N_11101);
and U11680 (N_11680,N_11305,N_11054);
xnor U11681 (N_11681,N_11167,N_11495);
nand U11682 (N_11682,N_11030,N_11019);
nor U11683 (N_11683,N_11229,N_11364);
or U11684 (N_11684,N_11401,N_11304);
xnor U11685 (N_11685,N_11335,N_11038);
xor U11686 (N_11686,N_11315,N_11480);
nor U11687 (N_11687,N_11484,N_11389);
nor U11688 (N_11688,N_11290,N_11239);
xor U11689 (N_11689,N_11471,N_11189);
nor U11690 (N_11690,N_11264,N_11073);
nor U11691 (N_11691,N_11456,N_11027);
or U11692 (N_11692,N_11271,N_11066);
nand U11693 (N_11693,N_11422,N_11499);
or U11694 (N_11694,N_11369,N_11462);
or U11695 (N_11695,N_11096,N_11254);
xnor U11696 (N_11696,N_11000,N_11231);
or U11697 (N_11697,N_11224,N_11213);
xnor U11698 (N_11698,N_11179,N_11077);
and U11699 (N_11699,N_11111,N_11393);
nand U11700 (N_11700,N_11257,N_11353);
and U11701 (N_11701,N_11033,N_11258);
nand U11702 (N_11702,N_11338,N_11406);
or U11703 (N_11703,N_11051,N_11209);
nand U11704 (N_11704,N_11193,N_11214);
and U11705 (N_11705,N_11450,N_11200);
xnor U11706 (N_11706,N_11485,N_11008);
or U11707 (N_11707,N_11039,N_11178);
nand U11708 (N_11708,N_11260,N_11091);
nor U11709 (N_11709,N_11031,N_11012);
or U11710 (N_11710,N_11452,N_11270);
nand U11711 (N_11711,N_11288,N_11392);
nor U11712 (N_11712,N_11065,N_11047);
or U11713 (N_11713,N_11370,N_11025);
nand U11714 (N_11714,N_11060,N_11195);
or U11715 (N_11715,N_11151,N_11003);
and U11716 (N_11716,N_11071,N_11157);
xor U11717 (N_11717,N_11227,N_11191);
and U11718 (N_11718,N_11463,N_11010);
or U11719 (N_11719,N_11067,N_11459);
nor U11720 (N_11720,N_11125,N_11085);
nor U11721 (N_11721,N_11017,N_11469);
nand U11722 (N_11722,N_11098,N_11458);
nor U11723 (N_11723,N_11251,N_11154);
or U11724 (N_11724,N_11411,N_11360);
nor U11725 (N_11725,N_11318,N_11026);
and U11726 (N_11726,N_11482,N_11188);
and U11727 (N_11727,N_11407,N_11181);
or U11728 (N_11728,N_11011,N_11082);
nand U11729 (N_11729,N_11395,N_11108);
and U11730 (N_11730,N_11296,N_11184);
and U11731 (N_11731,N_11472,N_11075);
nand U11732 (N_11732,N_11283,N_11115);
xor U11733 (N_11733,N_11329,N_11403);
nor U11734 (N_11734,N_11218,N_11295);
and U11735 (N_11735,N_11263,N_11374);
xnor U11736 (N_11736,N_11128,N_11028);
and U11737 (N_11737,N_11206,N_11455);
nand U11738 (N_11738,N_11208,N_11242);
and U11739 (N_11739,N_11351,N_11280);
xor U11740 (N_11740,N_11137,N_11006);
xor U11741 (N_11741,N_11203,N_11175);
nand U11742 (N_11742,N_11417,N_11152);
xnor U11743 (N_11743,N_11228,N_11379);
nor U11744 (N_11744,N_11409,N_11120);
and U11745 (N_11745,N_11371,N_11248);
nor U11746 (N_11746,N_11449,N_11235);
or U11747 (N_11747,N_11402,N_11062);
nor U11748 (N_11748,N_11476,N_11202);
xnor U11749 (N_11749,N_11467,N_11342);
and U11750 (N_11750,N_11331,N_11228);
and U11751 (N_11751,N_11140,N_11464);
nand U11752 (N_11752,N_11422,N_11121);
xor U11753 (N_11753,N_11455,N_11417);
and U11754 (N_11754,N_11351,N_11010);
nand U11755 (N_11755,N_11465,N_11368);
or U11756 (N_11756,N_11303,N_11073);
xor U11757 (N_11757,N_11455,N_11274);
xnor U11758 (N_11758,N_11065,N_11458);
nor U11759 (N_11759,N_11070,N_11114);
nand U11760 (N_11760,N_11252,N_11373);
xor U11761 (N_11761,N_11026,N_11437);
and U11762 (N_11762,N_11141,N_11148);
or U11763 (N_11763,N_11426,N_11216);
or U11764 (N_11764,N_11123,N_11407);
or U11765 (N_11765,N_11440,N_11048);
nand U11766 (N_11766,N_11066,N_11265);
nor U11767 (N_11767,N_11147,N_11069);
nor U11768 (N_11768,N_11359,N_11352);
and U11769 (N_11769,N_11409,N_11112);
nand U11770 (N_11770,N_11476,N_11365);
nand U11771 (N_11771,N_11316,N_11179);
xnor U11772 (N_11772,N_11225,N_11076);
nor U11773 (N_11773,N_11102,N_11314);
xnor U11774 (N_11774,N_11150,N_11033);
nand U11775 (N_11775,N_11262,N_11111);
or U11776 (N_11776,N_11138,N_11328);
or U11777 (N_11777,N_11398,N_11459);
nor U11778 (N_11778,N_11030,N_11398);
xnor U11779 (N_11779,N_11439,N_11195);
xor U11780 (N_11780,N_11078,N_11440);
xnor U11781 (N_11781,N_11447,N_11160);
xnor U11782 (N_11782,N_11097,N_11091);
nor U11783 (N_11783,N_11080,N_11021);
nor U11784 (N_11784,N_11120,N_11200);
nand U11785 (N_11785,N_11200,N_11244);
xnor U11786 (N_11786,N_11289,N_11394);
nand U11787 (N_11787,N_11024,N_11352);
and U11788 (N_11788,N_11234,N_11297);
and U11789 (N_11789,N_11110,N_11282);
xor U11790 (N_11790,N_11194,N_11141);
nor U11791 (N_11791,N_11222,N_11107);
or U11792 (N_11792,N_11435,N_11227);
nand U11793 (N_11793,N_11375,N_11292);
or U11794 (N_11794,N_11426,N_11040);
nor U11795 (N_11795,N_11070,N_11160);
or U11796 (N_11796,N_11450,N_11382);
or U11797 (N_11797,N_11074,N_11360);
xnor U11798 (N_11798,N_11007,N_11295);
xnor U11799 (N_11799,N_11483,N_11340);
nand U11800 (N_11800,N_11148,N_11265);
and U11801 (N_11801,N_11284,N_11157);
nand U11802 (N_11802,N_11449,N_11372);
and U11803 (N_11803,N_11492,N_11486);
and U11804 (N_11804,N_11236,N_11474);
and U11805 (N_11805,N_11261,N_11493);
and U11806 (N_11806,N_11262,N_11324);
or U11807 (N_11807,N_11257,N_11123);
and U11808 (N_11808,N_11416,N_11331);
or U11809 (N_11809,N_11141,N_11181);
nor U11810 (N_11810,N_11043,N_11092);
nand U11811 (N_11811,N_11416,N_11370);
nor U11812 (N_11812,N_11031,N_11259);
xnor U11813 (N_11813,N_11161,N_11037);
xor U11814 (N_11814,N_11496,N_11264);
xnor U11815 (N_11815,N_11127,N_11271);
xnor U11816 (N_11816,N_11077,N_11117);
or U11817 (N_11817,N_11052,N_11275);
nor U11818 (N_11818,N_11199,N_11491);
nor U11819 (N_11819,N_11327,N_11244);
or U11820 (N_11820,N_11237,N_11221);
nor U11821 (N_11821,N_11237,N_11194);
and U11822 (N_11822,N_11175,N_11450);
or U11823 (N_11823,N_11392,N_11134);
and U11824 (N_11824,N_11149,N_11133);
xnor U11825 (N_11825,N_11095,N_11015);
nor U11826 (N_11826,N_11167,N_11288);
nand U11827 (N_11827,N_11499,N_11047);
xnor U11828 (N_11828,N_11249,N_11259);
or U11829 (N_11829,N_11321,N_11098);
nor U11830 (N_11830,N_11139,N_11352);
nand U11831 (N_11831,N_11417,N_11061);
and U11832 (N_11832,N_11350,N_11385);
nor U11833 (N_11833,N_11360,N_11446);
nand U11834 (N_11834,N_11394,N_11469);
nand U11835 (N_11835,N_11243,N_11085);
nand U11836 (N_11836,N_11491,N_11110);
and U11837 (N_11837,N_11268,N_11292);
nor U11838 (N_11838,N_11473,N_11347);
xnor U11839 (N_11839,N_11498,N_11090);
or U11840 (N_11840,N_11087,N_11022);
nand U11841 (N_11841,N_11313,N_11494);
nand U11842 (N_11842,N_11480,N_11209);
or U11843 (N_11843,N_11232,N_11196);
nand U11844 (N_11844,N_11252,N_11336);
and U11845 (N_11845,N_11452,N_11339);
or U11846 (N_11846,N_11037,N_11066);
and U11847 (N_11847,N_11042,N_11051);
xor U11848 (N_11848,N_11477,N_11076);
and U11849 (N_11849,N_11041,N_11269);
nand U11850 (N_11850,N_11328,N_11360);
nor U11851 (N_11851,N_11085,N_11248);
and U11852 (N_11852,N_11077,N_11206);
nand U11853 (N_11853,N_11265,N_11119);
and U11854 (N_11854,N_11350,N_11044);
nor U11855 (N_11855,N_11110,N_11263);
or U11856 (N_11856,N_11452,N_11312);
nand U11857 (N_11857,N_11459,N_11291);
nand U11858 (N_11858,N_11326,N_11035);
or U11859 (N_11859,N_11486,N_11023);
xor U11860 (N_11860,N_11106,N_11434);
xnor U11861 (N_11861,N_11096,N_11030);
and U11862 (N_11862,N_11483,N_11122);
nor U11863 (N_11863,N_11142,N_11048);
nor U11864 (N_11864,N_11440,N_11216);
or U11865 (N_11865,N_11135,N_11193);
and U11866 (N_11866,N_11160,N_11295);
and U11867 (N_11867,N_11011,N_11469);
or U11868 (N_11868,N_11471,N_11252);
nor U11869 (N_11869,N_11171,N_11366);
or U11870 (N_11870,N_11307,N_11483);
nand U11871 (N_11871,N_11302,N_11020);
nor U11872 (N_11872,N_11492,N_11156);
and U11873 (N_11873,N_11402,N_11397);
and U11874 (N_11874,N_11219,N_11405);
and U11875 (N_11875,N_11337,N_11441);
xor U11876 (N_11876,N_11294,N_11287);
xor U11877 (N_11877,N_11042,N_11435);
or U11878 (N_11878,N_11333,N_11298);
and U11879 (N_11879,N_11202,N_11136);
and U11880 (N_11880,N_11045,N_11037);
nand U11881 (N_11881,N_11311,N_11328);
nor U11882 (N_11882,N_11463,N_11394);
or U11883 (N_11883,N_11258,N_11443);
and U11884 (N_11884,N_11418,N_11027);
and U11885 (N_11885,N_11123,N_11488);
nand U11886 (N_11886,N_11454,N_11287);
and U11887 (N_11887,N_11255,N_11226);
or U11888 (N_11888,N_11184,N_11474);
nor U11889 (N_11889,N_11078,N_11194);
xor U11890 (N_11890,N_11311,N_11010);
and U11891 (N_11891,N_11142,N_11237);
or U11892 (N_11892,N_11036,N_11400);
nor U11893 (N_11893,N_11242,N_11194);
nor U11894 (N_11894,N_11075,N_11267);
xnor U11895 (N_11895,N_11176,N_11100);
nand U11896 (N_11896,N_11445,N_11103);
nor U11897 (N_11897,N_11076,N_11372);
or U11898 (N_11898,N_11200,N_11324);
nand U11899 (N_11899,N_11258,N_11304);
or U11900 (N_11900,N_11412,N_11202);
or U11901 (N_11901,N_11154,N_11130);
nor U11902 (N_11902,N_11011,N_11100);
xor U11903 (N_11903,N_11165,N_11302);
nor U11904 (N_11904,N_11391,N_11305);
xor U11905 (N_11905,N_11282,N_11475);
nor U11906 (N_11906,N_11403,N_11058);
nand U11907 (N_11907,N_11440,N_11328);
or U11908 (N_11908,N_11029,N_11364);
and U11909 (N_11909,N_11440,N_11455);
or U11910 (N_11910,N_11174,N_11077);
and U11911 (N_11911,N_11311,N_11449);
nor U11912 (N_11912,N_11003,N_11144);
or U11913 (N_11913,N_11468,N_11260);
nand U11914 (N_11914,N_11467,N_11418);
or U11915 (N_11915,N_11097,N_11152);
xnor U11916 (N_11916,N_11465,N_11143);
nor U11917 (N_11917,N_11354,N_11064);
and U11918 (N_11918,N_11361,N_11428);
or U11919 (N_11919,N_11195,N_11089);
and U11920 (N_11920,N_11267,N_11015);
xor U11921 (N_11921,N_11476,N_11408);
or U11922 (N_11922,N_11435,N_11443);
nor U11923 (N_11923,N_11301,N_11352);
nand U11924 (N_11924,N_11016,N_11316);
nand U11925 (N_11925,N_11243,N_11495);
nor U11926 (N_11926,N_11050,N_11302);
xor U11927 (N_11927,N_11051,N_11124);
nor U11928 (N_11928,N_11056,N_11346);
nor U11929 (N_11929,N_11226,N_11294);
or U11930 (N_11930,N_11388,N_11064);
and U11931 (N_11931,N_11210,N_11454);
nand U11932 (N_11932,N_11218,N_11167);
and U11933 (N_11933,N_11333,N_11198);
xor U11934 (N_11934,N_11391,N_11375);
and U11935 (N_11935,N_11029,N_11358);
nor U11936 (N_11936,N_11316,N_11022);
or U11937 (N_11937,N_11365,N_11013);
nor U11938 (N_11938,N_11330,N_11069);
nand U11939 (N_11939,N_11439,N_11345);
nand U11940 (N_11940,N_11006,N_11057);
xor U11941 (N_11941,N_11275,N_11166);
or U11942 (N_11942,N_11042,N_11221);
and U11943 (N_11943,N_11004,N_11414);
or U11944 (N_11944,N_11423,N_11310);
or U11945 (N_11945,N_11034,N_11318);
or U11946 (N_11946,N_11179,N_11233);
nor U11947 (N_11947,N_11211,N_11193);
or U11948 (N_11948,N_11433,N_11288);
xnor U11949 (N_11949,N_11041,N_11399);
and U11950 (N_11950,N_11002,N_11266);
nand U11951 (N_11951,N_11131,N_11040);
and U11952 (N_11952,N_11478,N_11443);
nor U11953 (N_11953,N_11033,N_11225);
and U11954 (N_11954,N_11499,N_11213);
nand U11955 (N_11955,N_11104,N_11487);
or U11956 (N_11956,N_11418,N_11129);
and U11957 (N_11957,N_11201,N_11044);
nor U11958 (N_11958,N_11328,N_11047);
xor U11959 (N_11959,N_11346,N_11136);
xor U11960 (N_11960,N_11411,N_11053);
or U11961 (N_11961,N_11381,N_11351);
or U11962 (N_11962,N_11422,N_11230);
and U11963 (N_11963,N_11439,N_11080);
nor U11964 (N_11964,N_11410,N_11422);
and U11965 (N_11965,N_11282,N_11212);
nor U11966 (N_11966,N_11001,N_11371);
xnor U11967 (N_11967,N_11288,N_11004);
or U11968 (N_11968,N_11432,N_11022);
and U11969 (N_11969,N_11041,N_11265);
xnor U11970 (N_11970,N_11011,N_11052);
or U11971 (N_11971,N_11255,N_11461);
or U11972 (N_11972,N_11123,N_11222);
nand U11973 (N_11973,N_11206,N_11071);
nor U11974 (N_11974,N_11356,N_11131);
or U11975 (N_11975,N_11144,N_11114);
and U11976 (N_11976,N_11381,N_11051);
or U11977 (N_11977,N_11046,N_11212);
or U11978 (N_11978,N_11237,N_11136);
nand U11979 (N_11979,N_11481,N_11245);
and U11980 (N_11980,N_11336,N_11346);
and U11981 (N_11981,N_11171,N_11042);
xor U11982 (N_11982,N_11123,N_11446);
xor U11983 (N_11983,N_11150,N_11453);
or U11984 (N_11984,N_11213,N_11294);
nor U11985 (N_11985,N_11253,N_11382);
and U11986 (N_11986,N_11394,N_11096);
and U11987 (N_11987,N_11108,N_11146);
xnor U11988 (N_11988,N_11439,N_11398);
or U11989 (N_11989,N_11440,N_11071);
or U11990 (N_11990,N_11283,N_11106);
or U11991 (N_11991,N_11022,N_11001);
nor U11992 (N_11992,N_11424,N_11492);
nor U11993 (N_11993,N_11436,N_11113);
and U11994 (N_11994,N_11234,N_11441);
or U11995 (N_11995,N_11070,N_11115);
xor U11996 (N_11996,N_11279,N_11357);
or U11997 (N_11997,N_11399,N_11326);
xor U11998 (N_11998,N_11232,N_11176);
xnor U11999 (N_11999,N_11377,N_11014);
or U12000 (N_12000,N_11599,N_11650);
xor U12001 (N_12001,N_11908,N_11807);
nor U12002 (N_12002,N_11765,N_11662);
nor U12003 (N_12003,N_11718,N_11685);
nand U12004 (N_12004,N_11999,N_11967);
nand U12005 (N_12005,N_11671,N_11538);
or U12006 (N_12006,N_11764,N_11531);
and U12007 (N_12007,N_11804,N_11966);
nor U12008 (N_12008,N_11851,N_11789);
nor U12009 (N_12009,N_11919,N_11895);
or U12010 (N_12010,N_11578,N_11547);
nor U12011 (N_12011,N_11680,N_11960);
xor U12012 (N_12012,N_11709,N_11517);
nor U12013 (N_12013,N_11643,N_11548);
nor U12014 (N_12014,N_11786,N_11897);
and U12015 (N_12015,N_11914,N_11752);
and U12016 (N_12016,N_11620,N_11901);
nand U12017 (N_12017,N_11596,N_11893);
and U12018 (N_12018,N_11781,N_11844);
and U12019 (N_12019,N_11744,N_11625);
or U12020 (N_12020,N_11637,N_11555);
xnor U12021 (N_12021,N_11911,N_11873);
xnor U12022 (N_12022,N_11597,N_11906);
xnor U12023 (N_12023,N_11820,N_11608);
xnor U12024 (N_12024,N_11552,N_11664);
nand U12025 (N_12025,N_11852,N_11594);
nand U12026 (N_12026,N_11834,N_11679);
nor U12027 (N_12027,N_11576,N_11611);
nand U12028 (N_12028,N_11891,N_11672);
and U12029 (N_12029,N_11649,N_11668);
xor U12030 (N_12030,N_11639,N_11924);
xor U12031 (N_12031,N_11708,N_11977);
xnor U12032 (N_12032,N_11926,N_11863);
nand U12033 (N_12033,N_11505,N_11582);
and U12034 (N_12034,N_11747,N_11678);
nor U12035 (N_12035,N_11721,N_11942);
nand U12036 (N_12036,N_11951,N_11722);
nor U12037 (N_12037,N_11806,N_11581);
nand U12038 (N_12038,N_11976,N_11824);
and U12039 (N_12039,N_11935,N_11841);
nand U12040 (N_12040,N_11887,N_11775);
nand U12041 (N_12041,N_11948,N_11588);
or U12042 (N_12042,N_11978,N_11601);
and U12043 (N_12043,N_11733,N_11669);
nor U12044 (N_12044,N_11575,N_11687);
nand U12045 (N_12045,N_11540,N_11802);
and U12046 (N_12046,N_11823,N_11683);
or U12047 (N_12047,N_11577,N_11882);
or U12048 (N_12048,N_11821,N_11715);
nand U12049 (N_12049,N_11598,N_11570);
or U12050 (N_12050,N_11516,N_11936);
or U12051 (N_12051,N_11616,N_11986);
nor U12052 (N_12052,N_11719,N_11512);
nand U12053 (N_12053,N_11970,N_11866);
nand U12054 (N_12054,N_11567,N_11988);
nand U12055 (N_12055,N_11626,N_11886);
or U12056 (N_12056,N_11542,N_11865);
nor U12057 (N_12057,N_11899,N_11544);
or U12058 (N_12058,N_11653,N_11571);
or U12059 (N_12059,N_11741,N_11840);
or U12060 (N_12060,N_11533,N_11583);
and U12061 (N_12061,N_11952,N_11956);
nand U12062 (N_12062,N_11749,N_11720);
nor U12063 (N_12063,N_11796,N_11586);
xor U12064 (N_12064,N_11798,N_11793);
nand U12065 (N_12065,N_11675,N_11883);
nor U12066 (N_12066,N_11788,N_11943);
nor U12067 (N_12067,N_11550,N_11892);
xnor U12068 (N_12068,N_11553,N_11572);
nor U12069 (N_12069,N_11562,N_11995);
xnor U12070 (N_12070,N_11869,N_11829);
xnor U12071 (N_12071,N_11545,N_11652);
xor U12072 (N_12072,N_11529,N_11716);
or U12073 (N_12073,N_11525,N_11723);
nor U12074 (N_12074,N_11923,N_11916);
nor U12075 (N_12075,N_11526,N_11808);
nand U12076 (N_12076,N_11871,N_11950);
nor U12077 (N_12077,N_11812,N_11580);
xor U12078 (N_12078,N_11930,N_11515);
nor U12079 (N_12079,N_11780,N_11946);
nor U12080 (N_12080,N_11993,N_11703);
or U12081 (N_12081,N_11697,N_11880);
nand U12082 (N_12082,N_11573,N_11772);
nor U12083 (N_12083,N_11758,N_11509);
xnor U12084 (N_12084,N_11565,N_11860);
xnor U12085 (N_12085,N_11830,N_11963);
or U12086 (N_12086,N_11667,N_11979);
and U12087 (N_12087,N_11508,N_11656);
and U12088 (N_12088,N_11640,N_11522);
nand U12089 (N_12089,N_11814,N_11759);
nand U12090 (N_12090,N_11927,N_11753);
nand U12091 (N_12091,N_11955,N_11827);
xor U12092 (N_12092,N_11913,N_11932);
nand U12093 (N_12093,N_11725,N_11607);
nor U12094 (N_12094,N_11700,N_11676);
xor U12095 (N_12095,N_11934,N_11707);
nand U12096 (N_12096,N_11785,N_11884);
xor U12097 (N_12097,N_11528,N_11809);
nor U12098 (N_12098,N_11568,N_11770);
xnor U12099 (N_12099,N_11595,N_11646);
and U12100 (N_12100,N_11504,N_11791);
nor U12101 (N_12101,N_11861,N_11973);
or U12102 (N_12102,N_11774,N_11638);
xnor U12103 (N_12103,N_11805,N_11511);
xor U12104 (N_12104,N_11954,N_11959);
and U12105 (N_12105,N_11881,N_11584);
and U12106 (N_12106,N_11610,N_11953);
nor U12107 (N_12107,N_11609,N_11694);
xnor U12108 (N_12108,N_11790,N_11831);
or U12109 (N_12109,N_11728,N_11842);
or U12110 (N_12110,N_11917,N_11879);
xnor U12111 (N_12111,N_11868,N_11704);
nor U12112 (N_12112,N_11876,N_11783);
nand U12113 (N_12113,N_11875,N_11998);
or U12114 (N_12114,N_11564,N_11604);
xor U12115 (N_12115,N_11739,N_11799);
nor U12116 (N_12116,N_11877,N_11519);
nand U12117 (N_12117,N_11856,N_11751);
xor U12118 (N_12118,N_11985,N_11848);
or U12119 (N_12119,N_11816,N_11849);
and U12120 (N_12120,N_11629,N_11845);
nor U12121 (N_12121,N_11712,N_11742);
nor U12122 (N_12122,N_11681,N_11592);
xor U12123 (N_12123,N_11850,N_11760);
nor U12124 (N_12124,N_11819,N_11510);
nor U12125 (N_12125,N_11524,N_11894);
nand U12126 (N_12126,N_11590,N_11717);
nand U12127 (N_12127,N_11624,N_11836);
nor U12128 (N_12128,N_11847,N_11925);
and U12129 (N_12129,N_11813,N_11904);
and U12130 (N_12130,N_11614,N_11619);
nor U12131 (N_12131,N_11506,N_11859);
and U12132 (N_12132,N_11644,N_11754);
nor U12133 (N_12133,N_11931,N_11928);
or U12134 (N_12134,N_11980,N_11556);
nor U12135 (N_12135,N_11815,N_11682);
or U12136 (N_12136,N_11561,N_11878);
or U12137 (N_12137,N_11623,N_11763);
xnor U12138 (N_12138,N_11787,N_11663);
xor U12139 (N_12139,N_11779,N_11989);
and U12140 (N_12140,N_11915,N_11982);
xnor U12141 (N_12141,N_11991,N_11628);
xor U12142 (N_12142,N_11705,N_11684);
nor U12143 (N_12143,N_11748,N_11794);
and U12144 (N_12144,N_11801,N_11501);
or U12145 (N_12145,N_11699,N_11541);
and U12146 (N_12146,N_11797,N_11536);
or U12147 (N_12147,N_11613,N_11941);
and U12148 (N_12148,N_11818,N_11910);
nand U12149 (N_12149,N_11958,N_11602);
nor U12150 (N_12150,N_11778,N_11714);
xor U12151 (N_12151,N_11903,N_11756);
nor U12152 (N_12152,N_11761,N_11566);
or U12153 (N_12153,N_11912,N_11557);
and U12154 (N_12154,N_11800,N_11846);
xor U12155 (N_12155,N_11855,N_11543);
and U12156 (N_12156,N_11621,N_11514);
xor U12157 (N_12157,N_11702,N_11937);
and U12158 (N_12158,N_11857,N_11726);
nand U12159 (N_12159,N_11691,N_11689);
and U12160 (N_12160,N_11658,N_11503);
and U12161 (N_12161,N_11922,N_11975);
and U12162 (N_12162,N_11838,N_11563);
or U12163 (N_12163,N_11773,N_11606);
xnor U12164 (N_12164,N_11826,N_11949);
nand U12165 (N_12165,N_11546,N_11898);
and U12166 (N_12166,N_11603,N_11974);
xor U12167 (N_12167,N_11835,N_11732);
and U12168 (N_12168,N_11502,N_11569);
and U12169 (N_12169,N_11858,N_11939);
nor U12170 (N_12170,N_11992,N_11768);
nand U12171 (N_12171,N_11521,N_11961);
xor U12172 (N_12172,N_11938,N_11535);
or U12173 (N_12173,N_11843,N_11659);
xor U12174 (N_12174,N_11729,N_11690);
or U12175 (N_12175,N_11929,N_11636);
and U12176 (N_12176,N_11810,N_11693);
and U12177 (N_12177,N_11641,N_11957);
xor U12178 (N_12178,N_11549,N_11771);
nor U12179 (N_12179,N_11647,N_11698);
nand U12180 (N_12180,N_11984,N_11853);
nor U12181 (N_12181,N_11987,N_11825);
nor U12182 (N_12182,N_11532,N_11635);
nor U12183 (N_12183,N_11634,N_11591);
and U12184 (N_12184,N_11981,N_11711);
xor U12185 (N_12185,N_11971,N_11520);
nor U12186 (N_12186,N_11735,N_11585);
and U12187 (N_12187,N_11888,N_11921);
and U12188 (N_12188,N_11657,N_11792);
nor U12189 (N_12189,N_11589,N_11885);
xor U12190 (N_12190,N_11507,N_11731);
xor U12191 (N_12191,N_11730,N_11688);
xor U12192 (N_12192,N_11554,N_11642);
xor U12193 (N_12193,N_11965,N_11666);
xor U12194 (N_12194,N_11902,N_11618);
xor U12195 (N_12195,N_11994,N_11933);
nand U12196 (N_12196,N_11837,N_11889);
and U12197 (N_12197,N_11944,N_11996);
or U12198 (N_12198,N_11560,N_11579);
and U12199 (N_12199,N_11655,N_11534);
nor U12200 (N_12200,N_11874,N_11947);
and U12201 (N_12201,N_11551,N_11832);
nand U12202 (N_12202,N_11500,N_11593);
and U12203 (N_12203,N_11918,N_11972);
nand U12204 (N_12204,N_11537,N_11817);
xor U12205 (N_12205,N_11962,N_11539);
or U12206 (N_12206,N_11734,N_11724);
nor U12207 (N_12207,N_11777,N_11632);
xnor U12208 (N_12208,N_11523,N_11661);
and U12209 (N_12209,N_11600,N_11612);
and U12210 (N_12210,N_11527,N_11896);
or U12211 (N_12211,N_11695,N_11530);
nand U12212 (N_12212,N_11518,N_11738);
nor U12213 (N_12213,N_11727,N_11762);
nand U12214 (N_12214,N_11605,N_11587);
or U12215 (N_12215,N_11648,N_11696);
nand U12216 (N_12216,N_11867,N_11674);
nand U12217 (N_12217,N_11558,N_11750);
or U12218 (N_12218,N_11782,N_11755);
or U12219 (N_12219,N_11651,N_11766);
nor U12220 (N_12220,N_11574,N_11745);
xnor U12221 (N_12221,N_11559,N_11900);
or U12222 (N_12222,N_11862,N_11990);
xor U12223 (N_12223,N_11890,N_11784);
nand U12224 (N_12224,N_11706,N_11692);
nand U12225 (N_12225,N_11665,N_11968);
xor U12226 (N_12226,N_11864,N_11713);
xor U12227 (N_12227,N_11633,N_11811);
nand U12228 (N_12228,N_11660,N_11854);
nand U12229 (N_12229,N_11627,N_11654);
xnor U12230 (N_12230,N_11645,N_11940);
xnor U12231 (N_12231,N_11872,N_11617);
xor U12232 (N_12232,N_11767,N_11769);
xnor U12233 (N_12233,N_11905,N_11746);
or U12234 (N_12234,N_11743,N_11615);
nand U12235 (N_12235,N_11776,N_11828);
nor U12236 (N_12236,N_11997,N_11670);
xor U12237 (N_12237,N_11757,N_11737);
xor U12238 (N_12238,N_11870,N_11920);
and U12239 (N_12239,N_11803,N_11686);
xnor U12240 (N_12240,N_11909,N_11622);
nor U12241 (N_12241,N_11677,N_11945);
nor U12242 (N_12242,N_11631,N_11513);
nor U12243 (N_12243,N_11964,N_11740);
xnor U12244 (N_12244,N_11710,N_11701);
and U12245 (N_12245,N_11907,N_11969);
xnor U12246 (N_12246,N_11673,N_11833);
nand U12247 (N_12247,N_11839,N_11822);
nor U12248 (N_12248,N_11630,N_11736);
and U12249 (N_12249,N_11983,N_11795);
nor U12250 (N_12250,N_11525,N_11983);
and U12251 (N_12251,N_11900,N_11636);
xnor U12252 (N_12252,N_11945,N_11972);
nor U12253 (N_12253,N_11503,N_11881);
xnor U12254 (N_12254,N_11817,N_11821);
nand U12255 (N_12255,N_11982,N_11812);
nor U12256 (N_12256,N_11728,N_11870);
nor U12257 (N_12257,N_11745,N_11658);
or U12258 (N_12258,N_11615,N_11854);
nand U12259 (N_12259,N_11910,N_11822);
xor U12260 (N_12260,N_11560,N_11804);
and U12261 (N_12261,N_11647,N_11749);
nor U12262 (N_12262,N_11994,N_11910);
nor U12263 (N_12263,N_11766,N_11827);
xor U12264 (N_12264,N_11974,N_11617);
or U12265 (N_12265,N_11546,N_11684);
xnor U12266 (N_12266,N_11696,N_11916);
nand U12267 (N_12267,N_11711,N_11829);
and U12268 (N_12268,N_11517,N_11965);
and U12269 (N_12269,N_11919,N_11717);
xnor U12270 (N_12270,N_11780,N_11537);
nor U12271 (N_12271,N_11597,N_11699);
xor U12272 (N_12272,N_11746,N_11556);
and U12273 (N_12273,N_11894,N_11842);
and U12274 (N_12274,N_11733,N_11833);
xnor U12275 (N_12275,N_11836,N_11882);
nand U12276 (N_12276,N_11600,N_11947);
or U12277 (N_12277,N_11835,N_11729);
or U12278 (N_12278,N_11848,N_11675);
or U12279 (N_12279,N_11867,N_11704);
nor U12280 (N_12280,N_11714,N_11869);
or U12281 (N_12281,N_11710,N_11640);
nor U12282 (N_12282,N_11654,N_11564);
or U12283 (N_12283,N_11550,N_11838);
or U12284 (N_12284,N_11595,N_11956);
nand U12285 (N_12285,N_11965,N_11970);
and U12286 (N_12286,N_11853,N_11594);
xor U12287 (N_12287,N_11613,N_11878);
and U12288 (N_12288,N_11555,N_11658);
and U12289 (N_12289,N_11914,N_11589);
xnor U12290 (N_12290,N_11858,N_11749);
xnor U12291 (N_12291,N_11540,N_11845);
or U12292 (N_12292,N_11564,N_11699);
xnor U12293 (N_12293,N_11967,N_11720);
and U12294 (N_12294,N_11809,N_11917);
nor U12295 (N_12295,N_11728,N_11543);
and U12296 (N_12296,N_11797,N_11591);
nor U12297 (N_12297,N_11683,N_11557);
nor U12298 (N_12298,N_11793,N_11919);
xor U12299 (N_12299,N_11897,N_11917);
or U12300 (N_12300,N_11835,N_11810);
xor U12301 (N_12301,N_11582,N_11584);
xnor U12302 (N_12302,N_11971,N_11799);
nor U12303 (N_12303,N_11588,N_11860);
nor U12304 (N_12304,N_11585,N_11854);
or U12305 (N_12305,N_11921,N_11974);
xnor U12306 (N_12306,N_11819,N_11954);
xnor U12307 (N_12307,N_11672,N_11572);
and U12308 (N_12308,N_11914,N_11631);
or U12309 (N_12309,N_11581,N_11530);
nor U12310 (N_12310,N_11686,N_11770);
and U12311 (N_12311,N_11737,N_11500);
or U12312 (N_12312,N_11898,N_11888);
or U12313 (N_12313,N_11565,N_11900);
nor U12314 (N_12314,N_11896,N_11888);
xor U12315 (N_12315,N_11839,N_11799);
nand U12316 (N_12316,N_11876,N_11772);
or U12317 (N_12317,N_11856,N_11501);
xnor U12318 (N_12318,N_11749,N_11561);
nor U12319 (N_12319,N_11749,N_11738);
or U12320 (N_12320,N_11767,N_11700);
nor U12321 (N_12321,N_11828,N_11690);
or U12322 (N_12322,N_11516,N_11761);
nand U12323 (N_12323,N_11710,N_11957);
xnor U12324 (N_12324,N_11738,N_11873);
or U12325 (N_12325,N_11799,N_11572);
and U12326 (N_12326,N_11923,N_11640);
nor U12327 (N_12327,N_11565,N_11734);
nor U12328 (N_12328,N_11675,N_11933);
xnor U12329 (N_12329,N_11564,N_11591);
and U12330 (N_12330,N_11514,N_11688);
or U12331 (N_12331,N_11770,N_11502);
and U12332 (N_12332,N_11663,N_11550);
nand U12333 (N_12333,N_11782,N_11605);
or U12334 (N_12334,N_11867,N_11745);
and U12335 (N_12335,N_11603,N_11980);
and U12336 (N_12336,N_11718,N_11836);
nand U12337 (N_12337,N_11971,N_11527);
nand U12338 (N_12338,N_11639,N_11925);
or U12339 (N_12339,N_11718,N_11665);
xnor U12340 (N_12340,N_11827,N_11763);
nor U12341 (N_12341,N_11928,N_11993);
nand U12342 (N_12342,N_11619,N_11597);
and U12343 (N_12343,N_11854,N_11735);
and U12344 (N_12344,N_11663,N_11665);
nor U12345 (N_12345,N_11744,N_11555);
and U12346 (N_12346,N_11964,N_11651);
xnor U12347 (N_12347,N_11778,N_11752);
or U12348 (N_12348,N_11559,N_11695);
and U12349 (N_12349,N_11748,N_11593);
nand U12350 (N_12350,N_11732,N_11780);
or U12351 (N_12351,N_11501,N_11531);
or U12352 (N_12352,N_11523,N_11672);
or U12353 (N_12353,N_11880,N_11970);
xor U12354 (N_12354,N_11809,N_11861);
or U12355 (N_12355,N_11765,N_11920);
nand U12356 (N_12356,N_11635,N_11845);
or U12357 (N_12357,N_11912,N_11863);
nor U12358 (N_12358,N_11900,N_11670);
and U12359 (N_12359,N_11536,N_11622);
and U12360 (N_12360,N_11927,N_11538);
xor U12361 (N_12361,N_11514,N_11634);
nand U12362 (N_12362,N_11797,N_11970);
and U12363 (N_12363,N_11788,N_11657);
nand U12364 (N_12364,N_11591,N_11747);
xor U12365 (N_12365,N_11766,N_11801);
xor U12366 (N_12366,N_11824,N_11706);
or U12367 (N_12367,N_11544,N_11705);
xor U12368 (N_12368,N_11655,N_11631);
or U12369 (N_12369,N_11652,N_11761);
nor U12370 (N_12370,N_11546,N_11737);
nor U12371 (N_12371,N_11646,N_11530);
nand U12372 (N_12372,N_11985,N_11763);
and U12373 (N_12373,N_11764,N_11859);
or U12374 (N_12374,N_11766,N_11710);
or U12375 (N_12375,N_11707,N_11721);
nand U12376 (N_12376,N_11696,N_11676);
and U12377 (N_12377,N_11758,N_11982);
nor U12378 (N_12378,N_11541,N_11750);
or U12379 (N_12379,N_11699,N_11899);
and U12380 (N_12380,N_11902,N_11602);
xor U12381 (N_12381,N_11878,N_11590);
nand U12382 (N_12382,N_11935,N_11628);
xnor U12383 (N_12383,N_11542,N_11839);
nor U12384 (N_12384,N_11543,N_11811);
nor U12385 (N_12385,N_11792,N_11779);
and U12386 (N_12386,N_11910,N_11588);
nand U12387 (N_12387,N_11781,N_11639);
nor U12388 (N_12388,N_11916,N_11905);
and U12389 (N_12389,N_11677,N_11565);
and U12390 (N_12390,N_11869,N_11805);
or U12391 (N_12391,N_11812,N_11600);
nand U12392 (N_12392,N_11534,N_11938);
nand U12393 (N_12393,N_11698,N_11848);
nand U12394 (N_12394,N_11631,N_11766);
or U12395 (N_12395,N_11523,N_11956);
nand U12396 (N_12396,N_11821,N_11855);
nor U12397 (N_12397,N_11948,N_11844);
nor U12398 (N_12398,N_11544,N_11715);
nand U12399 (N_12399,N_11666,N_11992);
and U12400 (N_12400,N_11918,N_11900);
and U12401 (N_12401,N_11577,N_11599);
or U12402 (N_12402,N_11972,N_11861);
or U12403 (N_12403,N_11967,N_11734);
and U12404 (N_12404,N_11683,N_11788);
or U12405 (N_12405,N_11847,N_11996);
xor U12406 (N_12406,N_11846,N_11939);
or U12407 (N_12407,N_11639,N_11876);
nand U12408 (N_12408,N_11519,N_11741);
nand U12409 (N_12409,N_11633,N_11855);
xnor U12410 (N_12410,N_11860,N_11946);
or U12411 (N_12411,N_11931,N_11514);
or U12412 (N_12412,N_11907,N_11586);
xnor U12413 (N_12413,N_11669,N_11517);
nand U12414 (N_12414,N_11836,N_11646);
and U12415 (N_12415,N_11681,N_11780);
xnor U12416 (N_12416,N_11759,N_11748);
or U12417 (N_12417,N_11591,N_11761);
nor U12418 (N_12418,N_11835,N_11596);
xnor U12419 (N_12419,N_11665,N_11955);
nand U12420 (N_12420,N_11577,N_11797);
xnor U12421 (N_12421,N_11643,N_11721);
nand U12422 (N_12422,N_11580,N_11788);
and U12423 (N_12423,N_11693,N_11759);
and U12424 (N_12424,N_11842,N_11646);
nor U12425 (N_12425,N_11763,N_11660);
or U12426 (N_12426,N_11970,N_11678);
and U12427 (N_12427,N_11573,N_11928);
xor U12428 (N_12428,N_11926,N_11601);
xnor U12429 (N_12429,N_11620,N_11597);
and U12430 (N_12430,N_11867,N_11758);
xor U12431 (N_12431,N_11901,N_11983);
nand U12432 (N_12432,N_11613,N_11936);
xor U12433 (N_12433,N_11506,N_11872);
and U12434 (N_12434,N_11616,N_11977);
or U12435 (N_12435,N_11695,N_11782);
and U12436 (N_12436,N_11976,N_11757);
or U12437 (N_12437,N_11806,N_11703);
xor U12438 (N_12438,N_11816,N_11916);
or U12439 (N_12439,N_11864,N_11688);
xor U12440 (N_12440,N_11777,N_11855);
nand U12441 (N_12441,N_11903,N_11621);
or U12442 (N_12442,N_11731,N_11594);
and U12443 (N_12443,N_11626,N_11652);
nor U12444 (N_12444,N_11826,N_11704);
and U12445 (N_12445,N_11673,N_11508);
nand U12446 (N_12446,N_11907,N_11732);
and U12447 (N_12447,N_11600,N_11743);
xnor U12448 (N_12448,N_11996,N_11787);
and U12449 (N_12449,N_11719,N_11555);
nand U12450 (N_12450,N_11747,N_11871);
xor U12451 (N_12451,N_11536,N_11561);
or U12452 (N_12452,N_11999,N_11906);
and U12453 (N_12453,N_11693,N_11597);
nand U12454 (N_12454,N_11645,N_11578);
or U12455 (N_12455,N_11754,N_11959);
or U12456 (N_12456,N_11556,N_11597);
nand U12457 (N_12457,N_11874,N_11600);
nand U12458 (N_12458,N_11553,N_11815);
or U12459 (N_12459,N_11598,N_11664);
xor U12460 (N_12460,N_11992,N_11894);
and U12461 (N_12461,N_11820,N_11526);
nand U12462 (N_12462,N_11592,N_11985);
and U12463 (N_12463,N_11641,N_11574);
or U12464 (N_12464,N_11708,N_11554);
nand U12465 (N_12465,N_11517,N_11573);
nand U12466 (N_12466,N_11951,N_11763);
and U12467 (N_12467,N_11643,N_11770);
nor U12468 (N_12468,N_11899,N_11551);
and U12469 (N_12469,N_11766,N_11729);
nand U12470 (N_12470,N_11716,N_11996);
or U12471 (N_12471,N_11883,N_11780);
or U12472 (N_12472,N_11507,N_11825);
and U12473 (N_12473,N_11656,N_11635);
xor U12474 (N_12474,N_11673,N_11909);
nor U12475 (N_12475,N_11568,N_11773);
xor U12476 (N_12476,N_11957,N_11575);
and U12477 (N_12477,N_11712,N_11959);
nand U12478 (N_12478,N_11820,N_11909);
nand U12479 (N_12479,N_11903,N_11942);
and U12480 (N_12480,N_11747,N_11578);
or U12481 (N_12481,N_11840,N_11577);
nor U12482 (N_12482,N_11844,N_11991);
or U12483 (N_12483,N_11730,N_11871);
and U12484 (N_12484,N_11685,N_11579);
or U12485 (N_12485,N_11870,N_11937);
nand U12486 (N_12486,N_11899,N_11814);
nor U12487 (N_12487,N_11736,N_11944);
xor U12488 (N_12488,N_11560,N_11796);
nand U12489 (N_12489,N_11549,N_11781);
nand U12490 (N_12490,N_11928,N_11794);
nand U12491 (N_12491,N_11951,N_11731);
and U12492 (N_12492,N_11852,N_11654);
nor U12493 (N_12493,N_11610,N_11692);
nor U12494 (N_12494,N_11585,N_11697);
nor U12495 (N_12495,N_11505,N_11762);
and U12496 (N_12496,N_11912,N_11570);
nor U12497 (N_12497,N_11923,N_11580);
nor U12498 (N_12498,N_11986,N_11578);
and U12499 (N_12499,N_11881,N_11607);
or U12500 (N_12500,N_12390,N_12278);
xnor U12501 (N_12501,N_12069,N_12244);
and U12502 (N_12502,N_12315,N_12030);
nor U12503 (N_12503,N_12024,N_12411);
nand U12504 (N_12504,N_12231,N_12361);
nor U12505 (N_12505,N_12393,N_12319);
or U12506 (N_12506,N_12182,N_12141);
nor U12507 (N_12507,N_12391,N_12345);
or U12508 (N_12508,N_12487,N_12386);
nor U12509 (N_12509,N_12392,N_12325);
xor U12510 (N_12510,N_12066,N_12300);
nor U12511 (N_12511,N_12305,N_12227);
and U12512 (N_12512,N_12236,N_12308);
nor U12513 (N_12513,N_12036,N_12034);
or U12514 (N_12514,N_12075,N_12173);
nand U12515 (N_12515,N_12493,N_12454);
or U12516 (N_12516,N_12372,N_12017);
and U12517 (N_12517,N_12062,N_12058);
xor U12518 (N_12518,N_12481,N_12329);
nand U12519 (N_12519,N_12047,N_12148);
xor U12520 (N_12520,N_12295,N_12020);
or U12521 (N_12521,N_12083,N_12450);
nand U12522 (N_12522,N_12344,N_12050);
or U12523 (N_12523,N_12277,N_12460);
or U12524 (N_12524,N_12002,N_12389);
or U12525 (N_12525,N_12137,N_12358);
and U12526 (N_12526,N_12230,N_12109);
nor U12527 (N_12527,N_12092,N_12202);
nor U12528 (N_12528,N_12216,N_12156);
or U12529 (N_12529,N_12165,N_12014);
or U12530 (N_12530,N_12312,N_12469);
nor U12531 (N_12531,N_12248,N_12441);
or U12532 (N_12532,N_12022,N_12354);
or U12533 (N_12533,N_12434,N_12387);
nor U12534 (N_12534,N_12416,N_12365);
nor U12535 (N_12535,N_12476,N_12417);
nand U12536 (N_12536,N_12268,N_12076);
xor U12537 (N_12537,N_12181,N_12394);
xnor U12538 (N_12538,N_12396,N_12471);
and U12539 (N_12539,N_12422,N_12294);
or U12540 (N_12540,N_12322,N_12483);
xnor U12541 (N_12541,N_12177,N_12335);
xor U12542 (N_12542,N_12215,N_12168);
and U12543 (N_12543,N_12346,N_12064);
and U12544 (N_12544,N_12174,N_12035);
xor U12545 (N_12545,N_12143,N_12149);
and U12546 (N_12546,N_12257,N_12081);
nor U12547 (N_12547,N_12249,N_12136);
xnor U12548 (N_12548,N_12042,N_12113);
and U12549 (N_12549,N_12170,N_12381);
or U12550 (N_12550,N_12179,N_12189);
nor U12551 (N_12551,N_12204,N_12104);
and U12552 (N_12552,N_12232,N_12028);
or U12553 (N_12553,N_12098,N_12280);
nor U12554 (N_12554,N_12160,N_12205);
nor U12555 (N_12555,N_12032,N_12110);
nand U12556 (N_12556,N_12453,N_12119);
nor U12557 (N_12557,N_12362,N_12135);
or U12558 (N_12558,N_12420,N_12371);
xor U12559 (N_12559,N_12192,N_12026);
xor U12560 (N_12560,N_12303,N_12423);
and U12561 (N_12561,N_12237,N_12171);
nand U12562 (N_12562,N_12432,N_12337);
or U12563 (N_12563,N_12251,N_12306);
nor U12564 (N_12564,N_12463,N_12053);
nor U12565 (N_12565,N_12061,N_12080);
or U12566 (N_12566,N_12485,N_12498);
xnor U12567 (N_12567,N_12128,N_12490);
nor U12568 (N_12568,N_12093,N_12304);
and U12569 (N_12569,N_12051,N_12163);
nor U12570 (N_12570,N_12054,N_12180);
and U12571 (N_12571,N_12224,N_12488);
nand U12572 (N_12572,N_12264,N_12027);
nand U12573 (N_12573,N_12044,N_12146);
xor U12574 (N_12574,N_12482,N_12222);
or U12575 (N_12575,N_12410,N_12497);
and U12576 (N_12576,N_12260,N_12433);
or U12577 (N_12577,N_12465,N_12031);
xor U12578 (N_12578,N_12099,N_12468);
and U12579 (N_12579,N_12238,N_12470);
and U12580 (N_12580,N_12087,N_12282);
nand U12581 (N_12581,N_12436,N_12261);
nand U12582 (N_12582,N_12349,N_12117);
or U12583 (N_12583,N_12382,N_12021);
xor U12584 (N_12584,N_12207,N_12091);
nor U12585 (N_12585,N_12052,N_12383);
xor U12586 (N_12586,N_12399,N_12364);
nand U12587 (N_12587,N_12183,N_12326);
xnor U12588 (N_12588,N_12293,N_12172);
xor U12589 (N_12589,N_12262,N_12112);
or U12590 (N_12590,N_12073,N_12418);
nand U12591 (N_12591,N_12287,N_12253);
xor U12592 (N_12592,N_12284,N_12254);
xor U12593 (N_12593,N_12437,N_12157);
nor U12594 (N_12594,N_12464,N_12342);
or U12595 (N_12595,N_12015,N_12195);
nor U12596 (N_12596,N_12140,N_12106);
nand U12597 (N_12597,N_12301,N_12255);
nand U12598 (N_12598,N_12286,N_12259);
nor U12599 (N_12599,N_12272,N_12245);
and U12600 (N_12600,N_12495,N_12153);
xor U12601 (N_12601,N_12025,N_12475);
xor U12602 (N_12602,N_12444,N_12200);
nor U12603 (N_12603,N_12199,N_12167);
nand U12604 (N_12604,N_12100,N_12378);
nor U12605 (N_12605,N_12296,N_12310);
nand U12606 (N_12606,N_12190,N_12404);
or U12607 (N_12607,N_12065,N_12122);
nor U12608 (N_12608,N_12428,N_12243);
xnor U12609 (N_12609,N_12492,N_12048);
nand U12610 (N_12610,N_12496,N_12366);
xor U12611 (N_12611,N_12445,N_12348);
and U12612 (N_12612,N_12413,N_12409);
nor U12613 (N_12613,N_12270,N_12321);
nor U12614 (N_12614,N_12016,N_12443);
and U12615 (N_12615,N_12265,N_12185);
nand U12616 (N_12616,N_12336,N_12363);
or U12617 (N_12617,N_12219,N_12247);
nand U12618 (N_12618,N_12159,N_12154);
nand U12619 (N_12619,N_12298,N_12400);
xnor U12620 (N_12620,N_12164,N_12467);
nor U12621 (N_12621,N_12339,N_12212);
or U12622 (N_12622,N_12068,N_12442);
nand U12623 (N_12623,N_12077,N_12127);
xor U12624 (N_12624,N_12375,N_12175);
and U12625 (N_12625,N_12045,N_12134);
nand U12626 (N_12626,N_12427,N_12331);
and U12627 (N_12627,N_12115,N_12431);
or U12628 (N_12628,N_12142,N_12290);
xnor U12629 (N_12629,N_12285,N_12279);
or U12630 (N_12630,N_12144,N_12479);
or U12631 (N_12631,N_12071,N_12228);
and U12632 (N_12632,N_12440,N_12407);
nor U12633 (N_12633,N_12191,N_12161);
or U12634 (N_12634,N_12456,N_12297);
xor U12635 (N_12635,N_12102,N_12357);
xnor U12636 (N_12636,N_12309,N_12395);
nor U12637 (N_12637,N_12033,N_12133);
or U12638 (N_12638,N_12352,N_12151);
nand U12639 (N_12639,N_12121,N_12446);
xnor U12640 (N_12640,N_12240,N_12088);
nor U12641 (N_12641,N_12435,N_12449);
or U12642 (N_12642,N_12461,N_12370);
xnor U12643 (N_12643,N_12341,N_12211);
and U12644 (N_12644,N_12320,N_12223);
nor U12645 (N_12645,N_12499,N_12038);
nand U12646 (N_12646,N_12203,N_12096);
nor U12647 (N_12647,N_12079,N_12108);
nand U12648 (N_12648,N_12425,N_12338);
xnor U12649 (N_12649,N_12457,N_12355);
xnor U12650 (N_12650,N_12006,N_12377);
nand U12651 (N_12651,N_12458,N_12063);
and U12652 (N_12652,N_12398,N_12367);
nand U12653 (N_12653,N_12274,N_12405);
or U12654 (N_12654,N_12334,N_12201);
and U12655 (N_12655,N_12059,N_12241);
nor U12656 (N_12656,N_12126,N_12007);
or U12657 (N_12657,N_12162,N_12406);
and U12658 (N_12658,N_12129,N_12474);
nand U12659 (N_12659,N_12340,N_12327);
nand U12660 (N_12660,N_12090,N_12131);
nor U12661 (N_12661,N_12343,N_12401);
or U12662 (N_12662,N_12328,N_12009);
nor U12663 (N_12663,N_12466,N_12473);
nor U12664 (N_12664,N_12289,N_12221);
and U12665 (N_12665,N_12239,N_12302);
and U12666 (N_12666,N_12250,N_12455);
nor U12667 (N_12667,N_12094,N_12424);
nand U12668 (N_12668,N_12374,N_12046);
nand U12669 (N_12669,N_12210,N_12004);
nor U12670 (N_12670,N_12246,N_12226);
and U12671 (N_12671,N_12451,N_12039);
xnor U12672 (N_12672,N_12056,N_12166);
and U12673 (N_12673,N_12214,N_12196);
xnor U12674 (N_12674,N_12040,N_12023);
nor U12675 (N_12675,N_12229,N_12187);
or U12676 (N_12676,N_12145,N_12206);
and U12677 (N_12677,N_12350,N_12123);
and U12678 (N_12678,N_12324,N_12356);
nand U12679 (N_12679,N_12447,N_12111);
nor U12680 (N_12680,N_12388,N_12208);
or U12681 (N_12681,N_12086,N_12147);
and U12682 (N_12682,N_12491,N_12256);
nand U12683 (N_12683,N_12266,N_12351);
nor U12684 (N_12684,N_12414,N_12218);
nor U12685 (N_12685,N_12072,N_12178);
or U12686 (N_12686,N_12484,N_12095);
nand U12687 (N_12687,N_12421,N_12318);
nor U12688 (N_12688,N_12176,N_12369);
or U12689 (N_12689,N_12438,N_12169);
xor U12690 (N_12690,N_12380,N_12130);
nor U12691 (N_12691,N_12292,N_12029);
xnor U12692 (N_12692,N_12258,N_12333);
nor U12693 (N_12693,N_12158,N_12008);
and U12694 (N_12694,N_12276,N_12220);
nor U12695 (N_12695,N_12385,N_12198);
or U12696 (N_12696,N_12311,N_12452);
xor U12697 (N_12697,N_12101,N_12184);
or U12698 (N_12698,N_12000,N_12118);
nor U12699 (N_12699,N_12299,N_12291);
xor U12700 (N_12700,N_12150,N_12011);
nand U12701 (N_12701,N_12448,N_12489);
or U12702 (N_12702,N_12057,N_12384);
and U12703 (N_12703,N_12107,N_12001);
nor U12704 (N_12704,N_12263,N_12415);
nand U12705 (N_12705,N_12273,N_12379);
or U12706 (N_12706,N_12041,N_12234);
or U12707 (N_12707,N_12013,N_12097);
and U12708 (N_12708,N_12478,N_12124);
or U12709 (N_12709,N_12459,N_12155);
nand U12710 (N_12710,N_12003,N_12402);
nand U12711 (N_12711,N_12271,N_12233);
nor U12712 (N_12712,N_12089,N_12267);
or U12713 (N_12713,N_12313,N_12314);
and U12714 (N_12714,N_12252,N_12439);
nand U12715 (N_12715,N_12116,N_12332);
nor U12716 (N_12716,N_12408,N_12103);
and U12717 (N_12717,N_12269,N_12472);
and U12718 (N_12718,N_12018,N_12359);
and U12719 (N_12719,N_12188,N_12412);
xor U12720 (N_12720,N_12307,N_12283);
nor U12721 (N_12721,N_12376,N_12403);
and U12722 (N_12722,N_12494,N_12281);
nand U12723 (N_12723,N_12084,N_12486);
and U12724 (N_12724,N_12209,N_12043);
xnor U12725 (N_12725,N_12235,N_12429);
nor U12726 (N_12726,N_12477,N_12074);
or U12727 (N_12727,N_12049,N_12347);
and U12728 (N_12728,N_12213,N_12085);
and U12729 (N_12729,N_12055,N_12082);
nand U12730 (N_12730,N_12019,N_12426);
or U12731 (N_12731,N_12225,N_12360);
and U12732 (N_12732,N_12275,N_12373);
nand U12733 (N_12733,N_12152,N_12330);
and U12734 (N_12734,N_12193,N_12105);
or U12735 (N_12735,N_12005,N_12480);
xnor U12736 (N_12736,N_12114,N_12288);
and U12737 (N_12737,N_12067,N_12430);
nor U12738 (N_12738,N_12012,N_12186);
or U12739 (N_12739,N_12078,N_12125);
xnor U12740 (N_12740,N_12139,N_12070);
xor U12741 (N_12741,N_12368,N_12037);
or U12742 (N_12742,N_12217,N_12353);
xnor U12743 (N_12743,N_12197,N_12194);
nand U12744 (N_12744,N_12462,N_12132);
and U12745 (N_12745,N_12242,N_12419);
and U12746 (N_12746,N_12138,N_12397);
nand U12747 (N_12747,N_12060,N_12323);
nor U12748 (N_12748,N_12010,N_12316);
and U12749 (N_12749,N_12120,N_12317);
nor U12750 (N_12750,N_12375,N_12014);
and U12751 (N_12751,N_12240,N_12486);
or U12752 (N_12752,N_12215,N_12269);
or U12753 (N_12753,N_12483,N_12150);
or U12754 (N_12754,N_12257,N_12347);
nand U12755 (N_12755,N_12438,N_12183);
xnor U12756 (N_12756,N_12076,N_12179);
nor U12757 (N_12757,N_12475,N_12252);
nor U12758 (N_12758,N_12195,N_12489);
and U12759 (N_12759,N_12463,N_12077);
xor U12760 (N_12760,N_12351,N_12247);
nand U12761 (N_12761,N_12140,N_12091);
xnor U12762 (N_12762,N_12373,N_12218);
nor U12763 (N_12763,N_12246,N_12432);
nand U12764 (N_12764,N_12397,N_12399);
and U12765 (N_12765,N_12167,N_12302);
xor U12766 (N_12766,N_12099,N_12200);
or U12767 (N_12767,N_12499,N_12043);
or U12768 (N_12768,N_12021,N_12445);
or U12769 (N_12769,N_12209,N_12356);
nor U12770 (N_12770,N_12274,N_12424);
nand U12771 (N_12771,N_12385,N_12191);
and U12772 (N_12772,N_12320,N_12418);
and U12773 (N_12773,N_12457,N_12495);
nand U12774 (N_12774,N_12469,N_12167);
and U12775 (N_12775,N_12370,N_12372);
or U12776 (N_12776,N_12273,N_12039);
or U12777 (N_12777,N_12274,N_12280);
nor U12778 (N_12778,N_12288,N_12305);
and U12779 (N_12779,N_12076,N_12424);
and U12780 (N_12780,N_12331,N_12394);
nor U12781 (N_12781,N_12216,N_12200);
xnor U12782 (N_12782,N_12304,N_12155);
nand U12783 (N_12783,N_12301,N_12466);
xnor U12784 (N_12784,N_12109,N_12062);
xnor U12785 (N_12785,N_12003,N_12067);
nand U12786 (N_12786,N_12161,N_12307);
or U12787 (N_12787,N_12433,N_12331);
or U12788 (N_12788,N_12044,N_12083);
and U12789 (N_12789,N_12452,N_12059);
xnor U12790 (N_12790,N_12225,N_12497);
nand U12791 (N_12791,N_12002,N_12127);
nand U12792 (N_12792,N_12063,N_12006);
nand U12793 (N_12793,N_12403,N_12078);
nand U12794 (N_12794,N_12232,N_12079);
nor U12795 (N_12795,N_12459,N_12411);
and U12796 (N_12796,N_12442,N_12159);
or U12797 (N_12797,N_12124,N_12339);
nor U12798 (N_12798,N_12407,N_12105);
or U12799 (N_12799,N_12211,N_12180);
and U12800 (N_12800,N_12264,N_12132);
nor U12801 (N_12801,N_12421,N_12352);
nand U12802 (N_12802,N_12161,N_12183);
and U12803 (N_12803,N_12494,N_12328);
nor U12804 (N_12804,N_12234,N_12028);
or U12805 (N_12805,N_12232,N_12213);
xnor U12806 (N_12806,N_12341,N_12063);
or U12807 (N_12807,N_12441,N_12426);
xor U12808 (N_12808,N_12064,N_12351);
nand U12809 (N_12809,N_12283,N_12018);
xor U12810 (N_12810,N_12366,N_12053);
or U12811 (N_12811,N_12009,N_12345);
or U12812 (N_12812,N_12121,N_12292);
and U12813 (N_12813,N_12148,N_12400);
or U12814 (N_12814,N_12421,N_12374);
xnor U12815 (N_12815,N_12335,N_12372);
and U12816 (N_12816,N_12454,N_12292);
nor U12817 (N_12817,N_12255,N_12187);
or U12818 (N_12818,N_12223,N_12209);
nor U12819 (N_12819,N_12436,N_12024);
or U12820 (N_12820,N_12261,N_12444);
or U12821 (N_12821,N_12433,N_12285);
nand U12822 (N_12822,N_12489,N_12086);
and U12823 (N_12823,N_12487,N_12397);
nand U12824 (N_12824,N_12069,N_12370);
and U12825 (N_12825,N_12304,N_12084);
nor U12826 (N_12826,N_12054,N_12395);
nor U12827 (N_12827,N_12456,N_12051);
nor U12828 (N_12828,N_12138,N_12385);
xnor U12829 (N_12829,N_12208,N_12463);
and U12830 (N_12830,N_12440,N_12145);
xor U12831 (N_12831,N_12115,N_12119);
xnor U12832 (N_12832,N_12346,N_12465);
or U12833 (N_12833,N_12247,N_12283);
nand U12834 (N_12834,N_12397,N_12285);
and U12835 (N_12835,N_12462,N_12317);
and U12836 (N_12836,N_12057,N_12164);
or U12837 (N_12837,N_12215,N_12046);
nor U12838 (N_12838,N_12389,N_12148);
xor U12839 (N_12839,N_12313,N_12104);
xnor U12840 (N_12840,N_12360,N_12468);
xnor U12841 (N_12841,N_12482,N_12142);
xor U12842 (N_12842,N_12238,N_12097);
and U12843 (N_12843,N_12220,N_12135);
and U12844 (N_12844,N_12356,N_12354);
and U12845 (N_12845,N_12164,N_12088);
or U12846 (N_12846,N_12185,N_12470);
xnor U12847 (N_12847,N_12181,N_12020);
nand U12848 (N_12848,N_12404,N_12156);
nand U12849 (N_12849,N_12252,N_12283);
or U12850 (N_12850,N_12124,N_12000);
nor U12851 (N_12851,N_12264,N_12387);
nand U12852 (N_12852,N_12255,N_12481);
xor U12853 (N_12853,N_12261,N_12287);
xnor U12854 (N_12854,N_12325,N_12409);
xor U12855 (N_12855,N_12290,N_12369);
nor U12856 (N_12856,N_12161,N_12401);
nand U12857 (N_12857,N_12287,N_12100);
nand U12858 (N_12858,N_12005,N_12474);
xnor U12859 (N_12859,N_12416,N_12105);
or U12860 (N_12860,N_12294,N_12259);
or U12861 (N_12861,N_12096,N_12359);
nand U12862 (N_12862,N_12349,N_12263);
and U12863 (N_12863,N_12351,N_12054);
nand U12864 (N_12864,N_12094,N_12423);
and U12865 (N_12865,N_12443,N_12460);
nor U12866 (N_12866,N_12328,N_12492);
nand U12867 (N_12867,N_12086,N_12289);
xor U12868 (N_12868,N_12203,N_12450);
and U12869 (N_12869,N_12174,N_12437);
nor U12870 (N_12870,N_12470,N_12353);
nand U12871 (N_12871,N_12124,N_12440);
and U12872 (N_12872,N_12300,N_12127);
and U12873 (N_12873,N_12307,N_12427);
or U12874 (N_12874,N_12212,N_12468);
and U12875 (N_12875,N_12084,N_12223);
and U12876 (N_12876,N_12229,N_12143);
and U12877 (N_12877,N_12012,N_12021);
or U12878 (N_12878,N_12231,N_12254);
and U12879 (N_12879,N_12326,N_12187);
nand U12880 (N_12880,N_12459,N_12267);
nand U12881 (N_12881,N_12244,N_12082);
and U12882 (N_12882,N_12368,N_12382);
and U12883 (N_12883,N_12475,N_12485);
nand U12884 (N_12884,N_12342,N_12184);
and U12885 (N_12885,N_12376,N_12281);
or U12886 (N_12886,N_12348,N_12471);
or U12887 (N_12887,N_12169,N_12333);
xor U12888 (N_12888,N_12145,N_12238);
xor U12889 (N_12889,N_12011,N_12086);
nand U12890 (N_12890,N_12193,N_12406);
nand U12891 (N_12891,N_12254,N_12433);
xor U12892 (N_12892,N_12357,N_12452);
nand U12893 (N_12893,N_12205,N_12013);
xor U12894 (N_12894,N_12271,N_12140);
and U12895 (N_12895,N_12219,N_12235);
nor U12896 (N_12896,N_12130,N_12076);
or U12897 (N_12897,N_12081,N_12266);
xor U12898 (N_12898,N_12043,N_12306);
or U12899 (N_12899,N_12489,N_12409);
and U12900 (N_12900,N_12477,N_12144);
or U12901 (N_12901,N_12454,N_12427);
xor U12902 (N_12902,N_12430,N_12226);
nor U12903 (N_12903,N_12389,N_12273);
nor U12904 (N_12904,N_12207,N_12474);
or U12905 (N_12905,N_12098,N_12431);
and U12906 (N_12906,N_12205,N_12262);
or U12907 (N_12907,N_12054,N_12469);
xnor U12908 (N_12908,N_12327,N_12043);
nor U12909 (N_12909,N_12137,N_12230);
xor U12910 (N_12910,N_12269,N_12234);
and U12911 (N_12911,N_12198,N_12328);
and U12912 (N_12912,N_12366,N_12004);
or U12913 (N_12913,N_12037,N_12385);
xor U12914 (N_12914,N_12470,N_12477);
or U12915 (N_12915,N_12172,N_12002);
or U12916 (N_12916,N_12270,N_12001);
and U12917 (N_12917,N_12435,N_12059);
xnor U12918 (N_12918,N_12247,N_12361);
nand U12919 (N_12919,N_12262,N_12195);
nand U12920 (N_12920,N_12354,N_12122);
and U12921 (N_12921,N_12148,N_12127);
nor U12922 (N_12922,N_12462,N_12420);
or U12923 (N_12923,N_12322,N_12255);
or U12924 (N_12924,N_12422,N_12445);
and U12925 (N_12925,N_12140,N_12284);
nand U12926 (N_12926,N_12101,N_12217);
or U12927 (N_12927,N_12226,N_12025);
or U12928 (N_12928,N_12125,N_12478);
nor U12929 (N_12929,N_12135,N_12023);
and U12930 (N_12930,N_12232,N_12207);
xor U12931 (N_12931,N_12382,N_12398);
or U12932 (N_12932,N_12459,N_12398);
nor U12933 (N_12933,N_12252,N_12432);
xnor U12934 (N_12934,N_12025,N_12351);
xnor U12935 (N_12935,N_12041,N_12425);
nand U12936 (N_12936,N_12013,N_12114);
or U12937 (N_12937,N_12447,N_12121);
or U12938 (N_12938,N_12236,N_12395);
or U12939 (N_12939,N_12301,N_12115);
or U12940 (N_12940,N_12041,N_12487);
nand U12941 (N_12941,N_12015,N_12189);
and U12942 (N_12942,N_12423,N_12120);
nand U12943 (N_12943,N_12293,N_12022);
and U12944 (N_12944,N_12489,N_12482);
and U12945 (N_12945,N_12442,N_12313);
and U12946 (N_12946,N_12144,N_12286);
xnor U12947 (N_12947,N_12459,N_12293);
or U12948 (N_12948,N_12069,N_12274);
or U12949 (N_12949,N_12233,N_12001);
and U12950 (N_12950,N_12353,N_12357);
nand U12951 (N_12951,N_12484,N_12169);
or U12952 (N_12952,N_12214,N_12473);
xor U12953 (N_12953,N_12042,N_12242);
xnor U12954 (N_12954,N_12445,N_12023);
nand U12955 (N_12955,N_12445,N_12434);
or U12956 (N_12956,N_12497,N_12499);
nand U12957 (N_12957,N_12481,N_12335);
xor U12958 (N_12958,N_12088,N_12132);
nor U12959 (N_12959,N_12452,N_12428);
xor U12960 (N_12960,N_12001,N_12071);
nand U12961 (N_12961,N_12274,N_12108);
nand U12962 (N_12962,N_12074,N_12421);
xor U12963 (N_12963,N_12160,N_12178);
nand U12964 (N_12964,N_12328,N_12428);
nand U12965 (N_12965,N_12168,N_12214);
and U12966 (N_12966,N_12463,N_12283);
xor U12967 (N_12967,N_12452,N_12048);
nor U12968 (N_12968,N_12252,N_12137);
nand U12969 (N_12969,N_12090,N_12493);
xor U12970 (N_12970,N_12451,N_12066);
or U12971 (N_12971,N_12115,N_12392);
and U12972 (N_12972,N_12275,N_12397);
nand U12973 (N_12973,N_12139,N_12449);
nor U12974 (N_12974,N_12356,N_12460);
nand U12975 (N_12975,N_12423,N_12136);
or U12976 (N_12976,N_12333,N_12329);
or U12977 (N_12977,N_12335,N_12117);
nand U12978 (N_12978,N_12016,N_12147);
or U12979 (N_12979,N_12310,N_12151);
or U12980 (N_12980,N_12136,N_12339);
or U12981 (N_12981,N_12141,N_12453);
or U12982 (N_12982,N_12414,N_12084);
and U12983 (N_12983,N_12258,N_12251);
or U12984 (N_12984,N_12046,N_12259);
and U12985 (N_12985,N_12384,N_12444);
nand U12986 (N_12986,N_12366,N_12163);
and U12987 (N_12987,N_12318,N_12131);
and U12988 (N_12988,N_12449,N_12297);
nor U12989 (N_12989,N_12049,N_12324);
xor U12990 (N_12990,N_12391,N_12379);
or U12991 (N_12991,N_12232,N_12344);
or U12992 (N_12992,N_12205,N_12018);
nand U12993 (N_12993,N_12018,N_12103);
xnor U12994 (N_12994,N_12479,N_12393);
or U12995 (N_12995,N_12357,N_12104);
or U12996 (N_12996,N_12494,N_12131);
nor U12997 (N_12997,N_12316,N_12263);
nor U12998 (N_12998,N_12312,N_12055);
xnor U12999 (N_12999,N_12425,N_12260);
nand U13000 (N_13000,N_12939,N_12922);
nor U13001 (N_13001,N_12887,N_12767);
nor U13002 (N_13002,N_12606,N_12885);
and U13003 (N_13003,N_12835,N_12982);
and U13004 (N_13004,N_12801,N_12799);
xor U13005 (N_13005,N_12914,N_12553);
nor U13006 (N_13006,N_12501,N_12664);
nor U13007 (N_13007,N_12540,N_12999);
or U13008 (N_13008,N_12564,N_12611);
xnor U13009 (N_13009,N_12884,N_12932);
xor U13010 (N_13010,N_12631,N_12906);
nand U13011 (N_13011,N_12772,N_12890);
nor U13012 (N_13012,N_12584,N_12855);
xor U13013 (N_13013,N_12850,N_12989);
nor U13014 (N_13014,N_12705,N_12945);
xnor U13015 (N_13015,N_12679,N_12597);
nand U13016 (N_13016,N_12810,N_12616);
xnor U13017 (N_13017,N_12919,N_12923);
and U13018 (N_13018,N_12693,N_12995);
xnor U13019 (N_13019,N_12665,N_12815);
xnor U13020 (N_13020,N_12949,N_12589);
and U13021 (N_13021,N_12676,N_12948);
xnor U13022 (N_13022,N_12940,N_12747);
nor U13023 (N_13023,N_12771,N_12613);
nor U13024 (N_13024,N_12714,N_12822);
nand U13025 (N_13025,N_12696,N_12870);
and U13026 (N_13026,N_12857,N_12785);
nor U13027 (N_13027,N_12987,N_12582);
xnor U13028 (N_13028,N_12637,N_12782);
or U13029 (N_13029,N_12554,N_12965);
and U13030 (N_13030,N_12831,N_12629);
nor U13031 (N_13031,N_12572,N_12826);
nor U13032 (N_13032,N_12626,N_12792);
xnor U13033 (N_13033,N_12682,N_12764);
nor U13034 (N_13034,N_12889,N_12548);
xor U13035 (N_13035,N_12773,N_12673);
nand U13036 (N_13036,N_12841,N_12909);
nand U13037 (N_13037,N_12655,N_12955);
nand U13038 (N_13038,N_12913,N_12701);
and U13039 (N_13039,N_12726,N_12837);
nor U13040 (N_13040,N_12690,N_12832);
nand U13041 (N_13041,N_12877,N_12866);
or U13042 (N_13042,N_12807,N_12619);
and U13043 (N_13043,N_12886,N_12508);
nand U13044 (N_13044,N_12901,N_12891);
and U13045 (N_13045,N_12615,N_12576);
and U13046 (N_13046,N_12650,N_12713);
nand U13047 (N_13047,N_12912,N_12678);
and U13048 (N_13048,N_12775,N_12507);
nor U13049 (N_13049,N_12961,N_12586);
or U13050 (N_13050,N_12527,N_12608);
nor U13051 (N_13051,N_12652,N_12738);
nor U13052 (N_13052,N_12844,N_12609);
nand U13053 (N_13053,N_12648,N_12607);
or U13054 (N_13054,N_12567,N_12969);
xnor U13055 (N_13055,N_12538,N_12575);
or U13056 (N_13056,N_12968,N_12902);
or U13057 (N_13057,N_12634,N_12854);
xnor U13058 (N_13058,N_12635,N_12531);
or U13059 (N_13059,N_12672,N_12743);
or U13060 (N_13060,N_12592,N_12896);
or U13061 (N_13061,N_12893,N_12994);
xnor U13062 (N_13062,N_12543,N_12763);
and U13063 (N_13063,N_12562,N_12636);
or U13064 (N_13064,N_12518,N_12649);
or U13065 (N_13065,N_12975,N_12544);
nor U13066 (N_13066,N_12873,N_12716);
or U13067 (N_13067,N_12529,N_12983);
or U13068 (N_13068,N_12514,N_12712);
nor U13069 (N_13069,N_12620,N_12596);
nand U13070 (N_13070,N_12722,N_12511);
nand U13071 (N_13071,N_12819,N_12604);
and U13072 (N_13072,N_12512,N_12700);
and U13073 (N_13073,N_12762,N_12779);
nor U13074 (N_13074,N_12859,N_12595);
xor U13075 (N_13075,N_12777,N_12744);
or U13076 (N_13076,N_12675,N_12663);
or U13077 (N_13077,N_12735,N_12504);
and U13078 (N_13078,N_12694,N_12746);
and U13079 (N_13079,N_12783,N_12521);
xor U13080 (N_13080,N_12823,N_12978);
xor U13081 (N_13081,N_12897,N_12996);
nand U13082 (N_13082,N_12852,N_12559);
nor U13083 (N_13083,N_12594,N_12555);
and U13084 (N_13084,N_12802,N_12814);
xnor U13085 (N_13085,N_12880,N_12733);
nand U13086 (N_13086,N_12520,N_12506);
or U13087 (N_13087,N_12711,N_12622);
nand U13088 (N_13088,N_12549,N_12769);
and U13089 (N_13089,N_12911,N_12936);
and U13090 (N_13090,N_12741,N_12537);
or U13091 (N_13091,N_12972,N_12643);
nor U13092 (N_13092,N_12900,N_12704);
nand U13093 (N_13093,N_12784,N_12661);
nor U13094 (N_13094,N_12917,N_12591);
and U13095 (N_13095,N_12723,N_12926);
and U13096 (N_13096,N_12551,N_12929);
xor U13097 (N_13097,N_12740,N_12780);
xnor U13098 (N_13098,N_12967,N_12730);
and U13099 (N_13099,N_12659,N_12976);
nand U13100 (N_13100,N_12944,N_12685);
or U13101 (N_13101,N_12985,N_12590);
or U13102 (N_13102,N_12980,N_12928);
and U13103 (N_13103,N_12959,N_12633);
nor U13104 (N_13104,N_12956,N_12882);
nand U13105 (N_13105,N_12724,N_12666);
and U13106 (N_13106,N_12581,N_12847);
and U13107 (N_13107,N_12848,N_12853);
and U13108 (N_13108,N_12786,N_12593);
and U13109 (N_13109,N_12825,N_12568);
and U13110 (N_13110,N_12556,N_12957);
nor U13111 (N_13111,N_12871,N_12503);
xnor U13112 (N_13112,N_12981,N_12702);
nor U13113 (N_13113,N_12789,N_12605);
xor U13114 (N_13114,N_12677,N_12578);
xnor U13115 (N_13115,N_12625,N_12753);
xnor U13116 (N_13116,N_12545,N_12715);
nor U13117 (N_13117,N_12888,N_12599);
or U13118 (N_13118,N_12588,N_12971);
xor U13119 (N_13119,N_12776,N_12680);
xor U13120 (N_13120,N_12770,N_12757);
nor U13121 (N_13121,N_12519,N_12800);
or U13122 (N_13122,N_12748,N_12951);
nor U13123 (N_13123,N_12931,N_12569);
and U13124 (N_13124,N_12861,N_12577);
xnor U13125 (N_13125,N_12573,N_12532);
nor U13126 (N_13126,N_12988,N_12563);
nor U13127 (N_13127,N_12541,N_12829);
nand U13128 (N_13128,N_12515,N_12865);
or U13129 (N_13129,N_12683,N_12974);
xnor U13130 (N_13130,N_12977,N_12918);
or U13131 (N_13131,N_12695,N_12565);
or U13132 (N_13132,N_12778,N_12522);
and U13133 (N_13133,N_12689,N_12874);
and U13134 (N_13134,N_12818,N_12752);
nor U13135 (N_13135,N_12739,N_12621);
xor U13136 (N_13136,N_12570,N_12674);
or U13137 (N_13137,N_12610,N_12845);
xor U13138 (N_13138,N_12804,N_12907);
and U13139 (N_13139,N_12526,N_12903);
nand U13140 (N_13140,N_12628,N_12642);
nor U13141 (N_13141,N_12546,N_12766);
nand U13142 (N_13142,N_12516,N_12530);
or U13143 (N_13143,N_12973,N_12646);
nand U13144 (N_13144,N_12760,N_12528);
nand U13145 (N_13145,N_12946,N_12915);
nand U13146 (N_13146,N_12813,N_12878);
nor U13147 (N_13147,N_12720,N_12547);
and U13148 (N_13148,N_12806,N_12930);
or U13149 (N_13149,N_12598,N_12579);
and U13150 (N_13150,N_12842,N_12964);
and U13151 (N_13151,N_12667,N_12979);
nor U13152 (N_13152,N_12600,N_12681);
nand U13153 (N_13153,N_12509,N_12805);
xnor U13154 (N_13154,N_12561,N_12524);
nand U13155 (N_13155,N_12552,N_12990);
xnor U13156 (N_13156,N_12699,N_12833);
nand U13157 (N_13157,N_12728,N_12754);
nor U13158 (N_13158,N_12653,N_12920);
xnor U13159 (N_13159,N_12585,N_12647);
nand U13160 (N_13160,N_12795,N_12881);
nand U13161 (N_13161,N_12703,N_12879);
or U13162 (N_13162,N_12533,N_12698);
nor U13163 (N_13163,N_12725,N_12898);
or U13164 (N_13164,N_12790,N_12808);
xnor U13165 (N_13165,N_12758,N_12717);
and U13166 (N_13166,N_12603,N_12614);
nand U13167 (N_13167,N_12617,N_12812);
and U13168 (N_13168,N_12560,N_12943);
or U13169 (N_13169,N_12793,N_12550);
nor U13170 (N_13170,N_12623,N_12856);
and U13171 (N_13171,N_12750,N_12719);
nor U13172 (N_13172,N_12883,N_12542);
nand U13173 (N_13173,N_12627,N_12638);
nand U13174 (N_13174,N_12759,N_12756);
nand U13175 (N_13175,N_12566,N_12787);
nand U13176 (N_13176,N_12868,N_12500);
nor U13177 (N_13177,N_12732,N_12872);
or U13178 (N_13178,N_12558,N_12954);
xnor U13179 (N_13179,N_12765,N_12927);
and U13180 (N_13180,N_12718,N_12505);
xor U13181 (N_13181,N_12539,N_12820);
nand U13182 (N_13182,N_12632,N_12618);
or U13183 (N_13183,N_12921,N_12953);
and U13184 (N_13184,N_12639,N_12669);
and U13185 (N_13185,N_12867,N_12966);
or U13186 (N_13186,N_12523,N_12580);
nor U13187 (N_13187,N_12688,N_12742);
nand U13188 (N_13188,N_12525,N_12710);
nor U13189 (N_13189,N_12602,N_12809);
xor U13190 (N_13190,N_12862,N_12630);
nor U13191 (N_13191,N_12654,N_12670);
nor U13192 (N_13192,N_12937,N_12601);
and U13193 (N_13193,N_12933,N_12640);
xnor U13194 (N_13194,N_12571,N_12788);
nand U13195 (N_13195,N_12816,N_12869);
nand U13196 (N_13196,N_12706,N_12827);
xor U13197 (N_13197,N_12904,N_12895);
and U13198 (N_13198,N_12997,N_12839);
xor U13199 (N_13199,N_12797,N_12941);
xnor U13200 (N_13200,N_12817,N_12657);
and U13201 (N_13201,N_12875,N_12745);
nor U13202 (N_13202,N_12849,N_12993);
and U13203 (N_13203,N_12645,N_12644);
xor U13204 (N_13204,N_12583,N_12924);
and U13205 (N_13205,N_12656,N_12935);
xor U13206 (N_13206,N_12899,N_12836);
or U13207 (N_13207,N_12824,N_12697);
xnor U13208 (N_13208,N_12751,N_12624);
nand U13209 (N_13209,N_12908,N_12938);
nor U13210 (N_13210,N_12796,N_12734);
nand U13211 (N_13211,N_12612,N_12651);
nor U13212 (N_13212,N_12557,N_12838);
xnor U13213 (N_13213,N_12536,N_12828);
nor U13214 (N_13214,N_12660,N_12641);
nor U13215 (N_13215,N_12892,N_12662);
nor U13216 (N_13216,N_12671,N_12830);
and U13217 (N_13217,N_12834,N_12876);
nor U13218 (N_13218,N_12840,N_12860);
xnor U13219 (N_13219,N_12950,N_12707);
nor U13220 (N_13220,N_12736,N_12942);
nand U13221 (N_13221,N_12947,N_12843);
or U13222 (N_13222,N_12761,N_12731);
nand U13223 (N_13223,N_12658,N_12984);
xor U13224 (N_13224,N_12749,N_12934);
or U13225 (N_13225,N_12986,N_12925);
and U13226 (N_13226,N_12510,N_12687);
or U13227 (N_13227,N_12692,N_12958);
nand U13228 (N_13228,N_12709,N_12721);
and U13229 (N_13229,N_12502,N_12894);
nor U13230 (N_13230,N_12534,N_12905);
nand U13231 (N_13231,N_12574,N_12684);
and U13232 (N_13232,N_12952,N_12535);
or U13233 (N_13233,N_12998,N_12774);
or U13234 (N_13234,N_12803,N_12513);
xnor U13235 (N_13235,N_12811,N_12864);
and U13236 (N_13236,N_12755,N_12863);
nand U13237 (N_13237,N_12798,N_12960);
and U13238 (N_13238,N_12686,N_12781);
xor U13239 (N_13239,N_12916,N_12992);
nor U13240 (N_13240,N_12768,N_12963);
nand U13241 (N_13241,N_12851,N_12791);
or U13242 (N_13242,N_12691,N_12991);
and U13243 (N_13243,N_12668,N_12858);
xor U13244 (N_13244,N_12846,N_12821);
xor U13245 (N_13245,N_12794,N_12737);
nor U13246 (N_13246,N_12962,N_12708);
xnor U13247 (N_13247,N_12970,N_12587);
nand U13248 (N_13248,N_12727,N_12910);
or U13249 (N_13249,N_12729,N_12517);
xnor U13250 (N_13250,N_12985,N_12851);
nand U13251 (N_13251,N_12681,N_12593);
nand U13252 (N_13252,N_12928,N_12647);
and U13253 (N_13253,N_12582,N_12526);
nor U13254 (N_13254,N_12513,N_12545);
nand U13255 (N_13255,N_12522,N_12959);
or U13256 (N_13256,N_12623,N_12931);
xnor U13257 (N_13257,N_12995,N_12571);
or U13258 (N_13258,N_12595,N_12995);
or U13259 (N_13259,N_12959,N_12801);
xor U13260 (N_13260,N_12966,N_12755);
nor U13261 (N_13261,N_12793,N_12583);
nand U13262 (N_13262,N_12631,N_12751);
nand U13263 (N_13263,N_12930,N_12964);
xnor U13264 (N_13264,N_12957,N_12951);
nor U13265 (N_13265,N_12563,N_12679);
nor U13266 (N_13266,N_12864,N_12897);
or U13267 (N_13267,N_12641,N_12633);
nand U13268 (N_13268,N_12724,N_12559);
xnor U13269 (N_13269,N_12993,N_12599);
nor U13270 (N_13270,N_12935,N_12632);
or U13271 (N_13271,N_12667,N_12737);
or U13272 (N_13272,N_12965,N_12883);
and U13273 (N_13273,N_12844,N_12827);
nor U13274 (N_13274,N_12970,N_12787);
nand U13275 (N_13275,N_12960,N_12895);
xor U13276 (N_13276,N_12745,N_12718);
xor U13277 (N_13277,N_12541,N_12630);
nand U13278 (N_13278,N_12542,N_12729);
nand U13279 (N_13279,N_12733,N_12662);
nand U13280 (N_13280,N_12691,N_12989);
nand U13281 (N_13281,N_12984,N_12696);
nor U13282 (N_13282,N_12994,N_12676);
and U13283 (N_13283,N_12966,N_12974);
or U13284 (N_13284,N_12889,N_12936);
nor U13285 (N_13285,N_12631,N_12943);
or U13286 (N_13286,N_12983,N_12725);
or U13287 (N_13287,N_12617,N_12833);
xor U13288 (N_13288,N_12502,N_12745);
xor U13289 (N_13289,N_12865,N_12667);
nor U13290 (N_13290,N_12591,N_12607);
nand U13291 (N_13291,N_12878,N_12820);
xor U13292 (N_13292,N_12601,N_12954);
xor U13293 (N_13293,N_12730,N_12652);
nor U13294 (N_13294,N_12609,N_12792);
and U13295 (N_13295,N_12936,N_12502);
nor U13296 (N_13296,N_12695,N_12797);
or U13297 (N_13297,N_12984,N_12966);
nand U13298 (N_13298,N_12574,N_12687);
nand U13299 (N_13299,N_12562,N_12901);
or U13300 (N_13300,N_12506,N_12860);
and U13301 (N_13301,N_12701,N_12676);
and U13302 (N_13302,N_12777,N_12722);
or U13303 (N_13303,N_12509,N_12564);
or U13304 (N_13304,N_12906,N_12720);
and U13305 (N_13305,N_12693,N_12745);
xor U13306 (N_13306,N_12589,N_12543);
or U13307 (N_13307,N_12861,N_12603);
and U13308 (N_13308,N_12923,N_12892);
nand U13309 (N_13309,N_12591,N_12727);
nor U13310 (N_13310,N_12578,N_12687);
nand U13311 (N_13311,N_12591,N_12979);
or U13312 (N_13312,N_12564,N_12738);
or U13313 (N_13313,N_12686,N_12966);
xnor U13314 (N_13314,N_12922,N_12850);
or U13315 (N_13315,N_12870,N_12571);
xor U13316 (N_13316,N_12829,N_12566);
or U13317 (N_13317,N_12536,N_12554);
and U13318 (N_13318,N_12657,N_12799);
nand U13319 (N_13319,N_12861,N_12816);
or U13320 (N_13320,N_12695,N_12629);
nor U13321 (N_13321,N_12895,N_12976);
nor U13322 (N_13322,N_12568,N_12860);
and U13323 (N_13323,N_12755,N_12794);
nor U13324 (N_13324,N_12554,N_12517);
or U13325 (N_13325,N_12987,N_12614);
nor U13326 (N_13326,N_12796,N_12991);
nand U13327 (N_13327,N_12687,N_12794);
nand U13328 (N_13328,N_12647,N_12977);
nor U13329 (N_13329,N_12900,N_12549);
nand U13330 (N_13330,N_12664,N_12978);
and U13331 (N_13331,N_12609,N_12587);
or U13332 (N_13332,N_12525,N_12766);
and U13333 (N_13333,N_12929,N_12941);
nand U13334 (N_13334,N_12526,N_12729);
and U13335 (N_13335,N_12708,N_12869);
or U13336 (N_13336,N_12688,N_12792);
or U13337 (N_13337,N_12594,N_12893);
nor U13338 (N_13338,N_12564,N_12961);
and U13339 (N_13339,N_12976,N_12705);
nand U13340 (N_13340,N_12584,N_12786);
or U13341 (N_13341,N_12675,N_12536);
or U13342 (N_13342,N_12735,N_12779);
or U13343 (N_13343,N_12717,N_12996);
nand U13344 (N_13344,N_12515,N_12538);
nor U13345 (N_13345,N_12921,N_12847);
nand U13346 (N_13346,N_12670,N_12505);
nand U13347 (N_13347,N_12695,N_12590);
or U13348 (N_13348,N_12874,N_12899);
or U13349 (N_13349,N_12522,N_12626);
nand U13350 (N_13350,N_12540,N_12675);
nor U13351 (N_13351,N_12955,N_12726);
and U13352 (N_13352,N_12805,N_12701);
xor U13353 (N_13353,N_12597,N_12631);
nand U13354 (N_13354,N_12624,N_12652);
nand U13355 (N_13355,N_12800,N_12857);
nor U13356 (N_13356,N_12713,N_12935);
and U13357 (N_13357,N_12998,N_12613);
nor U13358 (N_13358,N_12961,N_12541);
nor U13359 (N_13359,N_12784,N_12637);
nand U13360 (N_13360,N_12806,N_12535);
or U13361 (N_13361,N_12774,N_12550);
or U13362 (N_13362,N_12902,N_12749);
or U13363 (N_13363,N_12670,N_12703);
xor U13364 (N_13364,N_12664,N_12526);
nand U13365 (N_13365,N_12832,N_12530);
xnor U13366 (N_13366,N_12658,N_12879);
or U13367 (N_13367,N_12882,N_12681);
and U13368 (N_13368,N_12797,N_12804);
and U13369 (N_13369,N_12501,N_12767);
nand U13370 (N_13370,N_12726,N_12531);
nand U13371 (N_13371,N_12911,N_12668);
xnor U13372 (N_13372,N_12993,N_12534);
nor U13373 (N_13373,N_12872,N_12746);
nand U13374 (N_13374,N_12970,N_12754);
nand U13375 (N_13375,N_12787,N_12712);
nand U13376 (N_13376,N_12771,N_12783);
or U13377 (N_13377,N_12513,N_12770);
xor U13378 (N_13378,N_12607,N_12763);
xor U13379 (N_13379,N_12582,N_12969);
nor U13380 (N_13380,N_12594,N_12770);
and U13381 (N_13381,N_12947,N_12509);
xor U13382 (N_13382,N_12576,N_12847);
nor U13383 (N_13383,N_12746,N_12622);
xor U13384 (N_13384,N_12647,N_12765);
xor U13385 (N_13385,N_12803,N_12586);
xor U13386 (N_13386,N_12801,N_12711);
xnor U13387 (N_13387,N_12952,N_12725);
or U13388 (N_13388,N_12903,N_12753);
xor U13389 (N_13389,N_12562,N_12632);
nor U13390 (N_13390,N_12592,N_12570);
nor U13391 (N_13391,N_12707,N_12625);
and U13392 (N_13392,N_12607,N_12594);
and U13393 (N_13393,N_12629,N_12584);
xor U13394 (N_13394,N_12548,N_12840);
or U13395 (N_13395,N_12599,N_12926);
and U13396 (N_13396,N_12653,N_12936);
nand U13397 (N_13397,N_12842,N_12581);
or U13398 (N_13398,N_12551,N_12785);
xnor U13399 (N_13399,N_12718,N_12947);
xnor U13400 (N_13400,N_12998,N_12699);
nor U13401 (N_13401,N_12779,N_12625);
and U13402 (N_13402,N_12967,N_12921);
nand U13403 (N_13403,N_12532,N_12550);
nor U13404 (N_13404,N_12589,N_12907);
and U13405 (N_13405,N_12773,N_12745);
and U13406 (N_13406,N_12755,N_12547);
nand U13407 (N_13407,N_12958,N_12672);
and U13408 (N_13408,N_12758,N_12578);
and U13409 (N_13409,N_12666,N_12709);
xor U13410 (N_13410,N_12624,N_12682);
xor U13411 (N_13411,N_12987,N_12640);
or U13412 (N_13412,N_12759,N_12507);
or U13413 (N_13413,N_12956,N_12921);
xnor U13414 (N_13414,N_12544,N_12893);
and U13415 (N_13415,N_12767,N_12785);
nor U13416 (N_13416,N_12892,N_12575);
and U13417 (N_13417,N_12865,N_12763);
nor U13418 (N_13418,N_12884,N_12550);
xnor U13419 (N_13419,N_12830,N_12754);
xor U13420 (N_13420,N_12544,N_12831);
nand U13421 (N_13421,N_12898,N_12792);
xnor U13422 (N_13422,N_12773,N_12554);
xnor U13423 (N_13423,N_12617,N_12608);
and U13424 (N_13424,N_12618,N_12579);
nor U13425 (N_13425,N_12559,N_12963);
or U13426 (N_13426,N_12908,N_12700);
nor U13427 (N_13427,N_12751,N_12603);
xnor U13428 (N_13428,N_12521,N_12867);
xnor U13429 (N_13429,N_12714,N_12809);
nor U13430 (N_13430,N_12925,N_12510);
or U13431 (N_13431,N_12906,N_12698);
nand U13432 (N_13432,N_12796,N_12970);
nor U13433 (N_13433,N_12895,N_12818);
and U13434 (N_13434,N_12885,N_12782);
nand U13435 (N_13435,N_12977,N_12947);
xnor U13436 (N_13436,N_12517,N_12687);
or U13437 (N_13437,N_12993,N_12632);
xnor U13438 (N_13438,N_12607,N_12573);
nor U13439 (N_13439,N_12850,N_12938);
and U13440 (N_13440,N_12564,N_12638);
or U13441 (N_13441,N_12791,N_12682);
nand U13442 (N_13442,N_12845,N_12688);
nor U13443 (N_13443,N_12681,N_12667);
nand U13444 (N_13444,N_12874,N_12863);
nand U13445 (N_13445,N_12631,N_12539);
or U13446 (N_13446,N_12681,N_12640);
nor U13447 (N_13447,N_12759,N_12508);
and U13448 (N_13448,N_12976,N_12599);
xnor U13449 (N_13449,N_12677,N_12512);
and U13450 (N_13450,N_12683,N_12855);
or U13451 (N_13451,N_12805,N_12977);
and U13452 (N_13452,N_12558,N_12848);
or U13453 (N_13453,N_12505,N_12808);
xnor U13454 (N_13454,N_12680,N_12709);
nor U13455 (N_13455,N_12548,N_12682);
nor U13456 (N_13456,N_12920,N_12572);
and U13457 (N_13457,N_12923,N_12510);
xor U13458 (N_13458,N_12890,N_12668);
nand U13459 (N_13459,N_12629,N_12957);
xor U13460 (N_13460,N_12937,N_12904);
nand U13461 (N_13461,N_12569,N_12573);
or U13462 (N_13462,N_12620,N_12854);
and U13463 (N_13463,N_12997,N_12618);
nor U13464 (N_13464,N_12857,N_12812);
or U13465 (N_13465,N_12721,N_12658);
xnor U13466 (N_13466,N_12762,N_12928);
nand U13467 (N_13467,N_12914,N_12672);
xnor U13468 (N_13468,N_12911,N_12695);
nand U13469 (N_13469,N_12739,N_12929);
xnor U13470 (N_13470,N_12663,N_12699);
or U13471 (N_13471,N_12985,N_12537);
or U13472 (N_13472,N_12876,N_12961);
nor U13473 (N_13473,N_12619,N_12815);
nand U13474 (N_13474,N_12776,N_12975);
xnor U13475 (N_13475,N_12504,N_12612);
or U13476 (N_13476,N_12777,N_12775);
nand U13477 (N_13477,N_12509,N_12681);
and U13478 (N_13478,N_12878,N_12703);
nand U13479 (N_13479,N_12663,N_12689);
nor U13480 (N_13480,N_12553,N_12634);
xnor U13481 (N_13481,N_12944,N_12887);
nand U13482 (N_13482,N_12659,N_12810);
xnor U13483 (N_13483,N_12580,N_12911);
nand U13484 (N_13484,N_12688,N_12607);
xnor U13485 (N_13485,N_12726,N_12538);
nor U13486 (N_13486,N_12656,N_12783);
or U13487 (N_13487,N_12816,N_12642);
nand U13488 (N_13488,N_12685,N_12858);
nor U13489 (N_13489,N_12815,N_12898);
nand U13490 (N_13490,N_12691,N_12812);
nor U13491 (N_13491,N_12877,N_12589);
or U13492 (N_13492,N_12584,N_12717);
nand U13493 (N_13493,N_12714,N_12550);
or U13494 (N_13494,N_12697,N_12986);
nor U13495 (N_13495,N_12950,N_12745);
nor U13496 (N_13496,N_12664,N_12778);
xnor U13497 (N_13497,N_12853,N_12549);
nand U13498 (N_13498,N_12853,N_12636);
nor U13499 (N_13499,N_12518,N_12942);
or U13500 (N_13500,N_13147,N_13421);
nand U13501 (N_13501,N_13396,N_13217);
xor U13502 (N_13502,N_13032,N_13368);
xnor U13503 (N_13503,N_13313,N_13275);
xor U13504 (N_13504,N_13185,N_13168);
xnor U13505 (N_13505,N_13463,N_13143);
or U13506 (N_13506,N_13055,N_13346);
nor U13507 (N_13507,N_13027,N_13160);
nand U13508 (N_13508,N_13295,N_13362);
or U13509 (N_13509,N_13019,N_13023);
and U13510 (N_13510,N_13402,N_13215);
nand U13511 (N_13511,N_13468,N_13111);
xor U13512 (N_13512,N_13262,N_13239);
nor U13513 (N_13513,N_13198,N_13287);
xor U13514 (N_13514,N_13461,N_13149);
nand U13515 (N_13515,N_13114,N_13335);
xnor U13516 (N_13516,N_13497,N_13090);
nand U13517 (N_13517,N_13246,N_13271);
xnor U13518 (N_13518,N_13065,N_13151);
nand U13519 (N_13519,N_13124,N_13140);
xnor U13520 (N_13520,N_13203,N_13391);
nor U13521 (N_13521,N_13052,N_13058);
nand U13522 (N_13522,N_13233,N_13069);
nand U13523 (N_13523,N_13309,N_13486);
nor U13524 (N_13524,N_13355,N_13206);
nor U13525 (N_13525,N_13162,N_13455);
or U13526 (N_13526,N_13424,N_13181);
or U13527 (N_13527,N_13013,N_13130);
and U13528 (N_13528,N_13302,N_13199);
nor U13529 (N_13529,N_13393,N_13457);
xnor U13530 (N_13530,N_13093,N_13495);
or U13531 (N_13531,N_13125,N_13155);
and U13532 (N_13532,N_13316,N_13175);
xnor U13533 (N_13533,N_13172,N_13216);
nand U13534 (N_13534,N_13437,N_13242);
and U13535 (N_13535,N_13499,N_13282);
or U13536 (N_13536,N_13307,N_13045);
nor U13537 (N_13537,N_13317,N_13000);
xor U13538 (N_13538,N_13249,N_13112);
nor U13539 (N_13539,N_13253,N_13290);
nor U13540 (N_13540,N_13224,N_13076);
and U13541 (N_13541,N_13448,N_13191);
and U13542 (N_13542,N_13440,N_13494);
nor U13543 (N_13543,N_13025,N_13041);
and U13544 (N_13544,N_13277,N_13337);
nor U13545 (N_13545,N_13442,N_13481);
or U13546 (N_13546,N_13120,N_13414);
or U13547 (N_13547,N_13095,N_13356);
nand U13548 (N_13548,N_13301,N_13007);
or U13549 (N_13549,N_13129,N_13102);
and U13550 (N_13550,N_13070,N_13336);
or U13551 (N_13551,N_13431,N_13351);
nor U13552 (N_13552,N_13074,N_13116);
xnor U13553 (N_13553,N_13487,N_13326);
xnor U13554 (N_13554,N_13213,N_13009);
xnor U13555 (N_13555,N_13018,N_13022);
nor U13556 (N_13556,N_13108,N_13103);
or U13557 (N_13557,N_13423,N_13110);
or U13558 (N_13558,N_13458,N_13002);
xnor U13559 (N_13559,N_13491,N_13496);
and U13560 (N_13560,N_13445,N_13284);
nor U13561 (N_13561,N_13338,N_13148);
or U13562 (N_13562,N_13278,N_13433);
xor U13563 (N_13563,N_13375,N_13477);
nor U13564 (N_13564,N_13475,N_13352);
nor U13565 (N_13565,N_13240,N_13320);
nand U13566 (N_13566,N_13067,N_13011);
or U13567 (N_13567,N_13328,N_13480);
or U13568 (N_13568,N_13134,N_13082);
nor U13569 (N_13569,N_13286,N_13450);
xnor U13570 (N_13570,N_13042,N_13107);
or U13571 (N_13571,N_13408,N_13343);
xor U13572 (N_13572,N_13341,N_13306);
or U13573 (N_13573,N_13020,N_13285);
nand U13574 (N_13574,N_13441,N_13270);
and U13575 (N_13575,N_13451,N_13324);
xor U13576 (N_13576,N_13268,N_13254);
or U13577 (N_13577,N_13340,N_13398);
or U13578 (N_13578,N_13322,N_13484);
xor U13579 (N_13579,N_13383,N_13101);
or U13580 (N_13580,N_13482,N_13483);
xor U13581 (N_13581,N_13227,N_13017);
xnor U13582 (N_13582,N_13057,N_13312);
nand U13583 (N_13583,N_13071,N_13189);
nand U13584 (N_13584,N_13051,N_13293);
xnor U13585 (N_13585,N_13086,N_13193);
nand U13586 (N_13586,N_13347,N_13359);
xor U13587 (N_13587,N_13410,N_13364);
xnor U13588 (N_13588,N_13488,N_13209);
and U13589 (N_13589,N_13349,N_13182);
or U13590 (N_13590,N_13098,N_13026);
xor U13591 (N_13591,N_13136,N_13365);
nor U13592 (N_13592,N_13188,N_13409);
and U13593 (N_13593,N_13083,N_13050);
xnor U13594 (N_13594,N_13062,N_13138);
nand U13595 (N_13595,N_13367,N_13006);
or U13596 (N_13596,N_13106,N_13243);
and U13597 (N_13597,N_13248,N_13257);
nand U13598 (N_13598,N_13406,N_13190);
nor U13599 (N_13599,N_13272,N_13210);
xnor U13600 (N_13600,N_13161,N_13493);
nand U13601 (N_13601,N_13225,N_13259);
or U13602 (N_13602,N_13053,N_13049);
xor U13603 (N_13603,N_13121,N_13173);
xor U13604 (N_13604,N_13333,N_13256);
nand U13605 (N_13605,N_13374,N_13081);
nand U13606 (N_13606,N_13078,N_13251);
nand U13607 (N_13607,N_13449,N_13195);
nor U13608 (N_13608,N_13109,N_13135);
nor U13609 (N_13609,N_13178,N_13401);
or U13610 (N_13610,N_13310,N_13456);
xnor U13611 (N_13611,N_13382,N_13358);
xor U13612 (N_13612,N_13056,N_13229);
and U13613 (N_13613,N_13060,N_13003);
or U13614 (N_13614,N_13263,N_13258);
nand U13615 (N_13615,N_13250,N_13179);
or U13616 (N_13616,N_13184,N_13218);
nor U13617 (N_13617,N_13036,N_13092);
or U13618 (N_13618,N_13490,N_13476);
or U13619 (N_13619,N_13159,N_13321);
nor U13620 (N_13620,N_13465,N_13399);
nor U13621 (N_13621,N_13331,N_13460);
or U13622 (N_13622,N_13016,N_13154);
xor U13623 (N_13623,N_13418,N_13369);
xor U13624 (N_13624,N_13126,N_13381);
xnor U13625 (N_13625,N_13498,N_13299);
and U13626 (N_13626,N_13294,N_13370);
or U13627 (N_13627,N_13133,N_13446);
xor U13628 (N_13628,N_13222,N_13386);
or U13629 (N_13629,N_13139,N_13265);
and U13630 (N_13630,N_13360,N_13061);
nand U13631 (N_13631,N_13236,N_13459);
or U13632 (N_13632,N_13377,N_13466);
xnor U13633 (N_13633,N_13238,N_13376);
and U13634 (N_13634,N_13419,N_13066);
nor U13635 (N_13635,N_13366,N_13363);
nand U13636 (N_13636,N_13245,N_13400);
nor U13637 (N_13637,N_13084,N_13170);
and U13638 (N_13638,N_13244,N_13407);
xor U13639 (N_13639,N_13157,N_13261);
and U13640 (N_13640,N_13371,N_13046);
xor U13641 (N_13641,N_13059,N_13385);
nor U13642 (N_13642,N_13353,N_13231);
nand U13643 (N_13643,N_13273,N_13397);
xor U13644 (N_13644,N_13387,N_13415);
nand U13645 (N_13645,N_13208,N_13205);
nor U13646 (N_13646,N_13447,N_13165);
or U13647 (N_13647,N_13395,N_13392);
nor U13648 (N_13648,N_13378,N_13153);
xnor U13649 (N_13649,N_13033,N_13255);
nand U13650 (N_13650,N_13439,N_13472);
nor U13651 (N_13651,N_13150,N_13452);
nand U13652 (N_13652,N_13384,N_13174);
and U13653 (N_13653,N_13192,N_13436);
nor U13654 (N_13654,N_13202,N_13283);
and U13655 (N_13655,N_13068,N_13004);
and U13656 (N_13656,N_13241,N_13390);
and U13657 (N_13657,N_13156,N_13453);
xnor U13658 (N_13658,N_13204,N_13373);
nor U13659 (N_13659,N_13296,N_13144);
nor U13660 (N_13660,N_13350,N_13292);
nor U13661 (N_13661,N_13123,N_13064);
nor U13662 (N_13662,N_13088,N_13334);
nand U13663 (N_13663,N_13269,N_13425);
and U13664 (N_13664,N_13422,N_13276);
and U13665 (N_13665,N_13474,N_13237);
or U13666 (N_13666,N_13085,N_13211);
and U13667 (N_13667,N_13131,N_13274);
nand U13668 (N_13668,N_13075,N_13266);
xnor U13669 (N_13669,N_13300,N_13037);
and U13670 (N_13670,N_13438,N_13473);
and U13671 (N_13671,N_13411,N_13196);
xor U13672 (N_13672,N_13478,N_13394);
and U13673 (N_13673,N_13029,N_13247);
nor U13674 (N_13674,N_13080,N_13104);
nand U13675 (N_13675,N_13152,N_13389);
and U13676 (N_13676,N_13297,N_13339);
or U13677 (N_13677,N_13485,N_13289);
nor U13678 (N_13678,N_13344,N_13429);
nor U13679 (N_13679,N_13072,N_13420);
and U13680 (N_13680,N_13315,N_13176);
and U13681 (N_13681,N_13354,N_13047);
and U13682 (N_13682,N_13220,N_13403);
xnor U13683 (N_13683,N_13314,N_13180);
xnor U13684 (N_13684,N_13470,N_13318);
or U13685 (N_13685,N_13113,N_13122);
or U13686 (N_13686,N_13186,N_13212);
xor U13687 (N_13687,N_13094,N_13323);
and U13688 (N_13688,N_13279,N_13200);
and U13689 (N_13689,N_13388,N_13163);
xnor U13690 (N_13690,N_13345,N_13372);
nor U13691 (N_13691,N_13426,N_13311);
xor U13692 (N_13692,N_13031,N_13427);
nand U13693 (N_13693,N_13281,N_13197);
or U13694 (N_13694,N_13469,N_13444);
nor U13695 (N_13695,N_13038,N_13319);
xor U13696 (N_13696,N_13329,N_13119);
and U13697 (N_13697,N_13252,N_13361);
nand U13698 (N_13698,N_13308,N_13207);
nor U13699 (N_13699,N_13091,N_13280);
and U13700 (N_13700,N_13105,N_13332);
and U13701 (N_13701,N_13479,N_13226);
nand U13702 (N_13702,N_13303,N_13404);
xnor U13703 (N_13703,N_13291,N_13325);
nand U13704 (N_13704,N_13043,N_13330);
and U13705 (N_13705,N_13234,N_13063);
and U13706 (N_13706,N_13305,N_13379);
or U13707 (N_13707,N_13167,N_13288);
nor U13708 (N_13708,N_13137,N_13443);
nor U13709 (N_13709,N_13145,N_13171);
xnor U13710 (N_13710,N_13462,N_13435);
nor U13711 (N_13711,N_13228,N_13146);
and U13712 (N_13712,N_13267,N_13008);
nor U13713 (N_13713,N_13005,N_13010);
nand U13714 (N_13714,N_13132,N_13430);
nor U13715 (N_13715,N_13097,N_13235);
xor U13716 (N_13716,N_13021,N_13230);
or U13717 (N_13717,N_13183,N_13492);
or U13718 (N_13718,N_13223,N_13471);
nand U13719 (N_13719,N_13087,N_13035);
or U13720 (N_13720,N_13194,N_13489);
and U13721 (N_13721,N_13260,N_13089);
xor U13722 (N_13722,N_13030,N_13434);
nor U13723 (N_13723,N_13214,N_13298);
xnor U13724 (N_13724,N_13454,N_13128);
nor U13725 (N_13725,N_13467,N_13014);
nand U13726 (N_13726,N_13024,N_13380);
and U13727 (N_13727,N_13412,N_13012);
nor U13728 (N_13728,N_13039,N_13044);
nor U13729 (N_13729,N_13034,N_13100);
nand U13730 (N_13730,N_13221,N_13118);
nand U13731 (N_13731,N_13177,N_13264);
nand U13732 (N_13732,N_13015,N_13115);
nand U13733 (N_13733,N_13001,N_13464);
nor U13734 (N_13734,N_13079,N_13040);
or U13735 (N_13735,N_13417,N_13141);
nor U13736 (N_13736,N_13117,N_13348);
or U13737 (N_13737,N_13201,N_13127);
nand U13738 (N_13738,N_13342,N_13413);
nor U13739 (N_13739,N_13077,N_13073);
xnor U13740 (N_13740,N_13164,N_13219);
nand U13741 (N_13741,N_13166,N_13158);
and U13742 (N_13742,N_13096,N_13432);
xor U13743 (N_13743,N_13187,N_13054);
nand U13744 (N_13744,N_13028,N_13304);
nor U13745 (N_13745,N_13169,N_13327);
nor U13746 (N_13746,N_13428,N_13099);
or U13747 (N_13747,N_13416,N_13405);
or U13748 (N_13748,N_13142,N_13357);
nor U13749 (N_13749,N_13048,N_13232);
nor U13750 (N_13750,N_13393,N_13213);
nor U13751 (N_13751,N_13332,N_13226);
xnor U13752 (N_13752,N_13106,N_13262);
and U13753 (N_13753,N_13097,N_13132);
xor U13754 (N_13754,N_13302,N_13332);
and U13755 (N_13755,N_13381,N_13461);
xnor U13756 (N_13756,N_13402,N_13095);
and U13757 (N_13757,N_13459,N_13022);
and U13758 (N_13758,N_13451,N_13009);
nand U13759 (N_13759,N_13101,N_13391);
nand U13760 (N_13760,N_13298,N_13032);
or U13761 (N_13761,N_13445,N_13251);
nor U13762 (N_13762,N_13266,N_13453);
or U13763 (N_13763,N_13019,N_13120);
xnor U13764 (N_13764,N_13475,N_13168);
xnor U13765 (N_13765,N_13296,N_13390);
nor U13766 (N_13766,N_13276,N_13316);
nor U13767 (N_13767,N_13461,N_13251);
and U13768 (N_13768,N_13022,N_13423);
xor U13769 (N_13769,N_13177,N_13429);
nand U13770 (N_13770,N_13013,N_13090);
and U13771 (N_13771,N_13127,N_13492);
xnor U13772 (N_13772,N_13487,N_13093);
and U13773 (N_13773,N_13074,N_13002);
xnor U13774 (N_13774,N_13147,N_13042);
nor U13775 (N_13775,N_13277,N_13111);
nor U13776 (N_13776,N_13442,N_13000);
xnor U13777 (N_13777,N_13320,N_13221);
xor U13778 (N_13778,N_13312,N_13265);
nand U13779 (N_13779,N_13151,N_13482);
and U13780 (N_13780,N_13490,N_13376);
xor U13781 (N_13781,N_13233,N_13128);
or U13782 (N_13782,N_13304,N_13065);
xor U13783 (N_13783,N_13054,N_13334);
and U13784 (N_13784,N_13082,N_13172);
nand U13785 (N_13785,N_13322,N_13016);
nand U13786 (N_13786,N_13379,N_13188);
nand U13787 (N_13787,N_13245,N_13412);
xor U13788 (N_13788,N_13060,N_13456);
xnor U13789 (N_13789,N_13303,N_13141);
and U13790 (N_13790,N_13347,N_13395);
nand U13791 (N_13791,N_13119,N_13256);
nor U13792 (N_13792,N_13213,N_13174);
nor U13793 (N_13793,N_13060,N_13384);
or U13794 (N_13794,N_13129,N_13034);
nand U13795 (N_13795,N_13345,N_13166);
nand U13796 (N_13796,N_13274,N_13392);
or U13797 (N_13797,N_13226,N_13402);
nand U13798 (N_13798,N_13166,N_13379);
or U13799 (N_13799,N_13320,N_13026);
nand U13800 (N_13800,N_13473,N_13351);
and U13801 (N_13801,N_13170,N_13019);
and U13802 (N_13802,N_13495,N_13068);
nand U13803 (N_13803,N_13251,N_13415);
or U13804 (N_13804,N_13051,N_13373);
and U13805 (N_13805,N_13462,N_13063);
or U13806 (N_13806,N_13346,N_13165);
nand U13807 (N_13807,N_13286,N_13021);
nor U13808 (N_13808,N_13343,N_13441);
xnor U13809 (N_13809,N_13032,N_13039);
and U13810 (N_13810,N_13041,N_13067);
xnor U13811 (N_13811,N_13156,N_13210);
and U13812 (N_13812,N_13103,N_13375);
and U13813 (N_13813,N_13431,N_13401);
nand U13814 (N_13814,N_13417,N_13266);
nor U13815 (N_13815,N_13460,N_13474);
and U13816 (N_13816,N_13292,N_13447);
or U13817 (N_13817,N_13261,N_13224);
nor U13818 (N_13818,N_13448,N_13231);
nor U13819 (N_13819,N_13413,N_13379);
or U13820 (N_13820,N_13281,N_13230);
and U13821 (N_13821,N_13077,N_13292);
and U13822 (N_13822,N_13353,N_13169);
xor U13823 (N_13823,N_13388,N_13268);
and U13824 (N_13824,N_13486,N_13420);
xor U13825 (N_13825,N_13262,N_13401);
nor U13826 (N_13826,N_13459,N_13132);
nor U13827 (N_13827,N_13396,N_13116);
nand U13828 (N_13828,N_13010,N_13161);
nor U13829 (N_13829,N_13349,N_13178);
nor U13830 (N_13830,N_13276,N_13006);
xnor U13831 (N_13831,N_13271,N_13074);
nand U13832 (N_13832,N_13327,N_13341);
or U13833 (N_13833,N_13385,N_13454);
nor U13834 (N_13834,N_13050,N_13250);
and U13835 (N_13835,N_13340,N_13094);
nor U13836 (N_13836,N_13456,N_13437);
nand U13837 (N_13837,N_13371,N_13374);
and U13838 (N_13838,N_13233,N_13022);
or U13839 (N_13839,N_13192,N_13081);
nand U13840 (N_13840,N_13009,N_13452);
xnor U13841 (N_13841,N_13489,N_13130);
nand U13842 (N_13842,N_13106,N_13129);
nor U13843 (N_13843,N_13463,N_13075);
xor U13844 (N_13844,N_13075,N_13156);
nand U13845 (N_13845,N_13015,N_13088);
or U13846 (N_13846,N_13360,N_13373);
or U13847 (N_13847,N_13394,N_13363);
and U13848 (N_13848,N_13030,N_13279);
xor U13849 (N_13849,N_13458,N_13027);
and U13850 (N_13850,N_13433,N_13237);
xnor U13851 (N_13851,N_13034,N_13434);
xnor U13852 (N_13852,N_13349,N_13270);
and U13853 (N_13853,N_13233,N_13426);
xnor U13854 (N_13854,N_13104,N_13333);
or U13855 (N_13855,N_13195,N_13108);
nor U13856 (N_13856,N_13291,N_13413);
xnor U13857 (N_13857,N_13090,N_13318);
nand U13858 (N_13858,N_13244,N_13430);
or U13859 (N_13859,N_13070,N_13031);
and U13860 (N_13860,N_13054,N_13276);
nor U13861 (N_13861,N_13475,N_13025);
xnor U13862 (N_13862,N_13303,N_13384);
xnor U13863 (N_13863,N_13011,N_13196);
or U13864 (N_13864,N_13288,N_13274);
xnor U13865 (N_13865,N_13335,N_13310);
nand U13866 (N_13866,N_13002,N_13110);
nor U13867 (N_13867,N_13111,N_13137);
nor U13868 (N_13868,N_13134,N_13294);
and U13869 (N_13869,N_13329,N_13250);
nand U13870 (N_13870,N_13231,N_13167);
nand U13871 (N_13871,N_13366,N_13424);
xor U13872 (N_13872,N_13438,N_13136);
and U13873 (N_13873,N_13032,N_13313);
or U13874 (N_13874,N_13196,N_13309);
and U13875 (N_13875,N_13231,N_13198);
and U13876 (N_13876,N_13227,N_13461);
and U13877 (N_13877,N_13008,N_13236);
nor U13878 (N_13878,N_13226,N_13071);
nor U13879 (N_13879,N_13333,N_13344);
xnor U13880 (N_13880,N_13158,N_13477);
or U13881 (N_13881,N_13051,N_13131);
xnor U13882 (N_13882,N_13401,N_13441);
and U13883 (N_13883,N_13444,N_13091);
or U13884 (N_13884,N_13356,N_13318);
nor U13885 (N_13885,N_13243,N_13329);
or U13886 (N_13886,N_13094,N_13359);
nor U13887 (N_13887,N_13030,N_13477);
nor U13888 (N_13888,N_13373,N_13066);
and U13889 (N_13889,N_13093,N_13052);
nor U13890 (N_13890,N_13027,N_13381);
xnor U13891 (N_13891,N_13485,N_13214);
or U13892 (N_13892,N_13171,N_13069);
and U13893 (N_13893,N_13428,N_13002);
nand U13894 (N_13894,N_13456,N_13360);
nand U13895 (N_13895,N_13244,N_13424);
and U13896 (N_13896,N_13452,N_13208);
xnor U13897 (N_13897,N_13485,N_13179);
and U13898 (N_13898,N_13267,N_13271);
nand U13899 (N_13899,N_13315,N_13149);
or U13900 (N_13900,N_13431,N_13487);
xor U13901 (N_13901,N_13225,N_13378);
nor U13902 (N_13902,N_13197,N_13191);
xor U13903 (N_13903,N_13431,N_13002);
and U13904 (N_13904,N_13384,N_13029);
nand U13905 (N_13905,N_13304,N_13064);
nor U13906 (N_13906,N_13413,N_13041);
or U13907 (N_13907,N_13385,N_13498);
and U13908 (N_13908,N_13332,N_13448);
or U13909 (N_13909,N_13244,N_13440);
and U13910 (N_13910,N_13106,N_13285);
and U13911 (N_13911,N_13133,N_13173);
xor U13912 (N_13912,N_13187,N_13436);
nor U13913 (N_13913,N_13198,N_13460);
and U13914 (N_13914,N_13098,N_13078);
nand U13915 (N_13915,N_13065,N_13300);
xor U13916 (N_13916,N_13190,N_13170);
or U13917 (N_13917,N_13253,N_13440);
xnor U13918 (N_13918,N_13435,N_13208);
nand U13919 (N_13919,N_13090,N_13308);
nand U13920 (N_13920,N_13482,N_13086);
or U13921 (N_13921,N_13212,N_13220);
nor U13922 (N_13922,N_13103,N_13360);
xor U13923 (N_13923,N_13434,N_13252);
xnor U13924 (N_13924,N_13480,N_13046);
nand U13925 (N_13925,N_13180,N_13418);
nand U13926 (N_13926,N_13291,N_13077);
or U13927 (N_13927,N_13452,N_13475);
nand U13928 (N_13928,N_13218,N_13491);
nand U13929 (N_13929,N_13236,N_13186);
nand U13930 (N_13930,N_13282,N_13215);
nor U13931 (N_13931,N_13202,N_13369);
or U13932 (N_13932,N_13334,N_13381);
nand U13933 (N_13933,N_13358,N_13442);
or U13934 (N_13934,N_13017,N_13280);
nand U13935 (N_13935,N_13497,N_13455);
or U13936 (N_13936,N_13039,N_13167);
and U13937 (N_13937,N_13341,N_13071);
and U13938 (N_13938,N_13060,N_13161);
nor U13939 (N_13939,N_13465,N_13161);
or U13940 (N_13940,N_13209,N_13448);
xnor U13941 (N_13941,N_13378,N_13344);
xor U13942 (N_13942,N_13476,N_13283);
xnor U13943 (N_13943,N_13188,N_13172);
nand U13944 (N_13944,N_13177,N_13166);
nand U13945 (N_13945,N_13281,N_13185);
xor U13946 (N_13946,N_13330,N_13491);
and U13947 (N_13947,N_13460,N_13139);
xor U13948 (N_13948,N_13235,N_13077);
and U13949 (N_13949,N_13316,N_13416);
or U13950 (N_13950,N_13018,N_13073);
nor U13951 (N_13951,N_13255,N_13426);
nor U13952 (N_13952,N_13120,N_13090);
xnor U13953 (N_13953,N_13454,N_13163);
xor U13954 (N_13954,N_13169,N_13305);
or U13955 (N_13955,N_13042,N_13452);
nor U13956 (N_13956,N_13477,N_13492);
nor U13957 (N_13957,N_13060,N_13370);
or U13958 (N_13958,N_13101,N_13119);
xnor U13959 (N_13959,N_13272,N_13226);
xor U13960 (N_13960,N_13101,N_13489);
or U13961 (N_13961,N_13142,N_13011);
nand U13962 (N_13962,N_13021,N_13209);
nand U13963 (N_13963,N_13387,N_13146);
nor U13964 (N_13964,N_13042,N_13083);
or U13965 (N_13965,N_13268,N_13406);
xnor U13966 (N_13966,N_13246,N_13407);
and U13967 (N_13967,N_13008,N_13000);
and U13968 (N_13968,N_13142,N_13148);
nand U13969 (N_13969,N_13071,N_13027);
or U13970 (N_13970,N_13302,N_13325);
nor U13971 (N_13971,N_13115,N_13277);
xor U13972 (N_13972,N_13202,N_13494);
nand U13973 (N_13973,N_13099,N_13113);
nor U13974 (N_13974,N_13075,N_13178);
nor U13975 (N_13975,N_13107,N_13121);
nor U13976 (N_13976,N_13245,N_13367);
or U13977 (N_13977,N_13338,N_13326);
xor U13978 (N_13978,N_13498,N_13442);
and U13979 (N_13979,N_13096,N_13317);
nand U13980 (N_13980,N_13330,N_13376);
or U13981 (N_13981,N_13209,N_13199);
xnor U13982 (N_13982,N_13389,N_13006);
nand U13983 (N_13983,N_13326,N_13140);
or U13984 (N_13984,N_13052,N_13461);
or U13985 (N_13985,N_13003,N_13180);
xnor U13986 (N_13986,N_13240,N_13140);
and U13987 (N_13987,N_13057,N_13017);
nand U13988 (N_13988,N_13412,N_13329);
and U13989 (N_13989,N_13178,N_13214);
and U13990 (N_13990,N_13463,N_13023);
nand U13991 (N_13991,N_13037,N_13141);
and U13992 (N_13992,N_13287,N_13466);
nor U13993 (N_13993,N_13270,N_13028);
nor U13994 (N_13994,N_13221,N_13327);
nor U13995 (N_13995,N_13480,N_13396);
xor U13996 (N_13996,N_13243,N_13076);
and U13997 (N_13997,N_13096,N_13402);
and U13998 (N_13998,N_13066,N_13081);
nand U13999 (N_13999,N_13129,N_13132);
and U14000 (N_14000,N_13827,N_13526);
xnor U14001 (N_14001,N_13879,N_13966);
or U14002 (N_14002,N_13684,N_13780);
nand U14003 (N_14003,N_13979,N_13734);
nand U14004 (N_14004,N_13534,N_13824);
nor U14005 (N_14005,N_13978,N_13936);
nand U14006 (N_14006,N_13570,N_13582);
or U14007 (N_14007,N_13553,N_13653);
nand U14008 (N_14008,N_13655,N_13985);
and U14009 (N_14009,N_13941,N_13884);
and U14010 (N_14010,N_13916,N_13537);
and U14011 (N_14011,N_13829,N_13946);
nor U14012 (N_14012,N_13819,N_13642);
or U14013 (N_14013,N_13677,N_13831);
xor U14014 (N_14014,N_13701,N_13515);
nand U14015 (N_14015,N_13898,N_13588);
nand U14016 (N_14016,N_13787,N_13666);
and U14017 (N_14017,N_13718,N_13951);
and U14018 (N_14018,N_13735,N_13533);
or U14019 (N_14019,N_13933,N_13589);
xor U14020 (N_14020,N_13712,N_13602);
or U14021 (N_14021,N_13704,N_13867);
xnor U14022 (N_14022,N_13776,N_13806);
nand U14023 (N_14023,N_13516,N_13868);
nor U14024 (N_14024,N_13673,N_13648);
nand U14025 (N_14025,N_13762,N_13950);
and U14026 (N_14026,N_13889,N_13505);
or U14027 (N_14027,N_13927,N_13523);
nand U14028 (N_14028,N_13847,N_13721);
or U14029 (N_14029,N_13885,N_13859);
nor U14030 (N_14030,N_13938,N_13947);
or U14031 (N_14031,N_13805,N_13963);
or U14032 (N_14032,N_13679,N_13663);
xor U14033 (N_14033,N_13683,N_13973);
nand U14034 (N_14034,N_13914,N_13945);
xnor U14035 (N_14035,N_13940,N_13836);
nor U14036 (N_14036,N_13755,N_13915);
nor U14037 (N_14037,N_13576,N_13767);
or U14038 (N_14038,N_13658,N_13994);
xnor U14039 (N_14039,N_13906,N_13863);
and U14040 (N_14040,N_13844,N_13568);
nand U14041 (N_14041,N_13874,N_13580);
nand U14042 (N_14042,N_13625,N_13766);
and U14043 (N_14043,N_13764,N_13630);
and U14044 (N_14044,N_13561,N_13943);
nor U14045 (N_14045,N_13772,N_13886);
xnor U14046 (N_14046,N_13584,N_13837);
or U14047 (N_14047,N_13577,N_13817);
xnor U14048 (N_14048,N_13595,N_13619);
and U14049 (N_14049,N_13518,N_13904);
or U14050 (N_14050,N_13865,N_13717);
and U14051 (N_14051,N_13669,N_13761);
or U14052 (N_14052,N_13616,N_13590);
xnor U14053 (N_14053,N_13967,N_13850);
nor U14054 (N_14054,N_13681,N_13789);
and U14055 (N_14055,N_13647,N_13792);
or U14056 (N_14056,N_13809,N_13739);
nor U14057 (N_14057,N_13724,N_13990);
nor U14058 (N_14058,N_13769,N_13745);
and U14059 (N_14059,N_13935,N_13998);
and U14060 (N_14060,N_13543,N_13697);
or U14061 (N_14061,N_13921,N_13746);
xnor U14062 (N_14062,N_13965,N_13969);
or U14063 (N_14063,N_13797,N_13707);
and U14064 (N_14064,N_13615,N_13682);
nor U14065 (N_14065,N_13511,N_13928);
xnor U14066 (N_14066,N_13610,N_13917);
or U14067 (N_14067,N_13897,N_13725);
nor U14068 (N_14068,N_13854,N_13705);
xnor U14069 (N_14069,N_13905,N_13632);
nor U14070 (N_14070,N_13638,N_13680);
nand U14071 (N_14071,N_13864,N_13728);
nor U14072 (N_14072,N_13880,N_13617);
nor U14073 (N_14073,N_13782,N_13598);
nand U14074 (N_14074,N_13508,N_13506);
and U14075 (N_14075,N_13972,N_13895);
xor U14076 (N_14076,N_13975,N_13531);
nand U14077 (N_14077,N_13962,N_13667);
nor U14078 (N_14078,N_13609,N_13959);
and U14079 (N_14079,N_13737,N_13596);
or U14080 (N_14080,N_13779,N_13788);
nand U14081 (N_14081,N_13932,N_13507);
nand U14082 (N_14082,N_13845,N_13942);
xnor U14083 (N_14083,N_13643,N_13757);
nor U14084 (N_14084,N_13981,N_13876);
or U14085 (N_14085,N_13659,N_13800);
xor U14086 (N_14086,N_13548,N_13544);
or U14087 (N_14087,N_13887,N_13970);
or U14088 (N_14088,N_13798,N_13988);
or U14089 (N_14089,N_13821,N_13624);
nor U14090 (N_14090,N_13727,N_13991);
nor U14091 (N_14091,N_13605,N_13713);
nor U14092 (N_14092,N_13953,N_13563);
nand U14093 (N_14093,N_13695,N_13607);
or U14094 (N_14094,N_13784,N_13976);
or U14095 (N_14095,N_13670,N_13594);
nor U14096 (N_14096,N_13968,N_13881);
xnor U14097 (N_14097,N_13907,N_13900);
xor U14098 (N_14098,N_13752,N_13500);
nor U14099 (N_14099,N_13977,N_13891);
xnor U14100 (N_14100,N_13565,N_13536);
and U14101 (N_14101,N_13742,N_13649);
nor U14102 (N_14102,N_13944,N_13993);
nand U14103 (N_14103,N_13825,N_13586);
and U14104 (N_14104,N_13633,N_13983);
nand U14105 (N_14105,N_13542,N_13622);
or U14106 (N_14106,N_13753,N_13599);
nand U14107 (N_14107,N_13822,N_13640);
or U14108 (N_14108,N_13731,N_13853);
nand U14109 (N_14109,N_13730,N_13572);
xnor U14110 (N_14110,N_13860,N_13774);
nor U14111 (N_14111,N_13509,N_13939);
nor U14112 (N_14112,N_13581,N_13519);
nor U14113 (N_14113,N_13986,N_13587);
xor U14114 (N_14114,N_13634,N_13614);
nor U14115 (N_14115,N_13641,N_13971);
nor U14116 (N_14116,N_13583,N_13538);
and U14117 (N_14117,N_13956,N_13686);
nand U14118 (N_14118,N_13926,N_13901);
nand U14119 (N_14119,N_13654,N_13980);
xnor U14120 (N_14120,N_13961,N_13883);
nand U14121 (N_14121,N_13722,N_13660);
xor U14122 (N_14122,N_13613,N_13992);
xnor U14123 (N_14123,N_13744,N_13535);
xor U14124 (N_14124,N_13569,N_13620);
and U14125 (N_14125,N_13899,N_13996);
nor U14126 (N_14126,N_13549,N_13770);
or U14127 (N_14127,N_13575,N_13626);
nand U14128 (N_14128,N_13703,N_13521);
nor U14129 (N_14129,N_13591,N_13637);
and U14130 (N_14130,N_13893,N_13668);
and U14131 (N_14131,N_13842,N_13612);
and U14132 (N_14132,N_13715,N_13984);
nand U14133 (N_14133,N_13564,N_13960);
and U14134 (N_14134,N_13786,N_13803);
nor U14135 (N_14135,N_13987,N_13846);
nand U14136 (N_14136,N_13691,N_13794);
or U14137 (N_14137,N_13547,N_13878);
and U14138 (N_14138,N_13804,N_13711);
and U14139 (N_14139,N_13852,N_13541);
or U14140 (N_14140,N_13522,N_13818);
xnor U14141 (N_14141,N_13922,N_13957);
nor U14142 (N_14142,N_13514,N_13756);
nand U14143 (N_14143,N_13982,N_13559);
nand U14144 (N_14144,N_13801,N_13955);
nand U14145 (N_14145,N_13903,N_13925);
and U14146 (N_14146,N_13676,N_13750);
and U14147 (N_14147,N_13631,N_13934);
nand U14148 (N_14148,N_13823,N_13958);
nand U14149 (N_14149,N_13556,N_13820);
xnor U14150 (N_14150,N_13699,N_13608);
and U14151 (N_14151,N_13861,N_13989);
nor U14152 (N_14152,N_13738,N_13913);
xor U14153 (N_14153,N_13513,N_13775);
and U14154 (N_14154,N_13706,N_13758);
xnor U14155 (N_14155,N_13532,N_13740);
and U14156 (N_14156,N_13890,N_13689);
and U14157 (N_14157,N_13603,N_13768);
nand U14158 (N_14158,N_13636,N_13675);
and U14159 (N_14159,N_13645,N_13578);
xnor U14160 (N_14160,N_13835,N_13931);
or U14161 (N_14161,N_13554,N_13908);
nor U14162 (N_14162,N_13685,N_13520);
nand U14163 (N_14163,N_13719,N_13948);
nand U14164 (N_14164,N_13920,N_13688);
and U14165 (N_14165,N_13902,N_13802);
xor U14166 (N_14166,N_13919,N_13504);
or U14167 (N_14167,N_13964,N_13501);
nand U14168 (N_14168,N_13749,N_13952);
nand U14169 (N_14169,N_13664,N_13525);
and U14170 (N_14170,N_13585,N_13558);
nand U14171 (N_14171,N_13510,N_13692);
or U14172 (N_14172,N_13857,N_13754);
or U14173 (N_14173,N_13995,N_13657);
or U14174 (N_14174,N_13892,N_13644);
nor U14175 (N_14175,N_13877,N_13882);
nor U14176 (N_14176,N_13848,N_13579);
nand U14177 (N_14177,N_13635,N_13528);
and U14178 (N_14178,N_13833,N_13841);
nor U14179 (N_14179,N_13828,N_13791);
and U14180 (N_14180,N_13751,N_13714);
nor U14181 (N_14181,N_13838,N_13872);
or U14182 (N_14182,N_13816,N_13974);
or U14183 (N_14183,N_13709,N_13840);
nand U14184 (N_14184,N_13911,N_13650);
nor U14185 (N_14185,N_13623,N_13524);
nand U14186 (N_14186,N_13760,N_13812);
and U14187 (N_14187,N_13694,N_13503);
and U14188 (N_14188,N_13651,N_13672);
or U14189 (N_14189,N_13918,N_13855);
or U14190 (N_14190,N_13700,N_13869);
nor U14191 (N_14191,N_13807,N_13555);
xor U14192 (N_14192,N_13910,N_13567);
xnor U14193 (N_14193,N_13674,N_13796);
nor U14194 (N_14194,N_13593,N_13813);
nor U14195 (N_14195,N_13783,N_13997);
and U14196 (N_14196,N_13815,N_13870);
nand U14197 (N_14197,N_13562,N_13929);
nor U14198 (N_14198,N_13826,N_13873);
or U14199 (N_14199,N_13741,N_13811);
and U14200 (N_14200,N_13573,N_13832);
and U14201 (N_14201,N_13793,N_13646);
or U14202 (N_14202,N_13652,N_13571);
xor U14203 (N_14203,N_13665,N_13629);
nor U14204 (N_14204,N_13912,N_13875);
or U14205 (N_14205,N_13698,N_13759);
nor U14206 (N_14206,N_13687,N_13639);
and U14207 (N_14207,N_13763,N_13729);
nor U14208 (N_14208,N_13671,N_13512);
and U14209 (N_14209,N_13949,N_13662);
or U14210 (N_14210,N_13726,N_13628);
and U14211 (N_14211,N_13710,N_13527);
and U14212 (N_14212,N_13732,N_13856);
nor U14213 (N_14213,N_13690,N_13894);
nand U14214 (N_14214,N_13866,N_13723);
and U14215 (N_14215,N_13843,N_13862);
and U14216 (N_14216,N_13785,N_13849);
xor U14217 (N_14217,N_13773,N_13529);
nor U14218 (N_14218,N_13693,N_13778);
or U14219 (N_14219,N_13810,N_13808);
nand U14220 (N_14220,N_13871,N_13502);
nor U14221 (N_14221,N_13611,N_13574);
nor U14222 (N_14222,N_13799,N_13661);
or U14223 (N_14223,N_13597,N_13606);
and U14224 (N_14224,N_13736,N_13834);
nand U14225 (N_14225,N_13851,N_13777);
nand U14226 (N_14226,N_13546,N_13765);
and U14227 (N_14227,N_13696,N_13923);
or U14228 (N_14228,N_13937,N_13795);
or U14229 (N_14229,N_13708,N_13621);
nand U14230 (N_14230,N_13601,N_13743);
xnor U14231 (N_14231,N_13627,N_13771);
xnor U14232 (N_14232,N_13733,N_13814);
or U14233 (N_14233,N_13550,N_13566);
nand U14234 (N_14234,N_13517,N_13858);
xnor U14235 (N_14235,N_13552,N_13557);
or U14236 (N_14236,N_13560,N_13618);
nand U14237 (N_14237,N_13839,N_13781);
or U14238 (N_14238,N_13909,N_13702);
or U14239 (N_14239,N_13790,N_13600);
nor U14240 (N_14240,N_13592,N_13930);
and U14241 (N_14241,N_13830,N_13896);
or U14242 (N_14242,N_13545,N_13540);
or U14243 (N_14243,N_13530,N_13747);
and U14244 (N_14244,N_13604,N_13888);
or U14245 (N_14245,N_13748,N_13924);
and U14246 (N_14246,N_13656,N_13954);
and U14247 (N_14247,N_13678,N_13551);
and U14248 (N_14248,N_13539,N_13716);
and U14249 (N_14249,N_13999,N_13720);
nor U14250 (N_14250,N_13645,N_13835);
or U14251 (N_14251,N_13622,N_13907);
and U14252 (N_14252,N_13754,N_13502);
xor U14253 (N_14253,N_13908,N_13512);
xor U14254 (N_14254,N_13830,N_13626);
and U14255 (N_14255,N_13796,N_13824);
nand U14256 (N_14256,N_13564,N_13943);
xnor U14257 (N_14257,N_13979,N_13723);
nand U14258 (N_14258,N_13586,N_13870);
nor U14259 (N_14259,N_13563,N_13958);
or U14260 (N_14260,N_13673,N_13551);
or U14261 (N_14261,N_13968,N_13975);
and U14262 (N_14262,N_13979,N_13718);
nand U14263 (N_14263,N_13537,N_13726);
and U14264 (N_14264,N_13848,N_13911);
xnor U14265 (N_14265,N_13557,N_13986);
or U14266 (N_14266,N_13620,N_13994);
and U14267 (N_14267,N_13754,N_13635);
or U14268 (N_14268,N_13998,N_13563);
or U14269 (N_14269,N_13577,N_13744);
or U14270 (N_14270,N_13737,N_13858);
nor U14271 (N_14271,N_13818,N_13634);
and U14272 (N_14272,N_13761,N_13646);
nor U14273 (N_14273,N_13520,N_13690);
nor U14274 (N_14274,N_13517,N_13734);
nor U14275 (N_14275,N_13807,N_13567);
or U14276 (N_14276,N_13566,N_13719);
or U14277 (N_14277,N_13832,N_13908);
xor U14278 (N_14278,N_13953,N_13850);
or U14279 (N_14279,N_13842,N_13793);
nand U14280 (N_14280,N_13911,N_13571);
or U14281 (N_14281,N_13554,N_13695);
xor U14282 (N_14282,N_13588,N_13529);
xnor U14283 (N_14283,N_13851,N_13915);
nor U14284 (N_14284,N_13700,N_13791);
xor U14285 (N_14285,N_13933,N_13502);
or U14286 (N_14286,N_13565,N_13848);
nor U14287 (N_14287,N_13731,N_13888);
nand U14288 (N_14288,N_13800,N_13924);
xor U14289 (N_14289,N_13613,N_13637);
nand U14290 (N_14290,N_13685,N_13752);
nor U14291 (N_14291,N_13953,N_13786);
nand U14292 (N_14292,N_13859,N_13545);
nor U14293 (N_14293,N_13841,N_13509);
or U14294 (N_14294,N_13838,N_13660);
nor U14295 (N_14295,N_13741,N_13768);
xnor U14296 (N_14296,N_13615,N_13898);
nand U14297 (N_14297,N_13623,N_13548);
and U14298 (N_14298,N_13650,N_13967);
and U14299 (N_14299,N_13515,N_13980);
xor U14300 (N_14300,N_13858,N_13893);
and U14301 (N_14301,N_13609,N_13505);
xor U14302 (N_14302,N_13825,N_13520);
nand U14303 (N_14303,N_13861,N_13724);
nor U14304 (N_14304,N_13593,N_13726);
xnor U14305 (N_14305,N_13815,N_13647);
xor U14306 (N_14306,N_13849,N_13507);
and U14307 (N_14307,N_13945,N_13543);
xor U14308 (N_14308,N_13791,N_13891);
or U14309 (N_14309,N_13915,N_13507);
xor U14310 (N_14310,N_13695,N_13544);
nand U14311 (N_14311,N_13824,N_13773);
or U14312 (N_14312,N_13637,N_13846);
and U14313 (N_14313,N_13531,N_13558);
and U14314 (N_14314,N_13790,N_13933);
nor U14315 (N_14315,N_13734,N_13580);
or U14316 (N_14316,N_13890,N_13632);
nand U14317 (N_14317,N_13929,N_13784);
nor U14318 (N_14318,N_13669,N_13993);
nand U14319 (N_14319,N_13555,N_13970);
nand U14320 (N_14320,N_13619,N_13681);
or U14321 (N_14321,N_13653,N_13859);
and U14322 (N_14322,N_13733,N_13846);
nor U14323 (N_14323,N_13812,N_13992);
or U14324 (N_14324,N_13590,N_13646);
or U14325 (N_14325,N_13707,N_13595);
xor U14326 (N_14326,N_13506,N_13731);
xnor U14327 (N_14327,N_13650,N_13821);
nand U14328 (N_14328,N_13885,N_13770);
and U14329 (N_14329,N_13632,N_13602);
nor U14330 (N_14330,N_13932,N_13944);
and U14331 (N_14331,N_13918,N_13612);
and U14332 (N_14332,N_13888,N_13937);
and U14333 (N_14333,N_13513,N_13951);
nand U14334 (N_14334,N_13798,N_13790);
nor U14335 (N_14335,N_13938,N_13507);
or U14336 (N_14336,N_13604,N_13857);
or U14337 (N_14337,N_13524,N_13942);
nand U14338 (N_14338,N_13648,N_13549);
nor U14339 (N_14339,N_13842,N_13705);
or U14340 (N_14340,N_13612,N_13620);
nand U14341 (N_14341,N_13810,N_13629);
nor U14342 (N_14342,N_13543,N_13849);
and U14343 (N_14343,N_13527,N_13764);
nor U14344 (N_14344,N_13587,N_13639);
and U14345 (N_14345,N_13810,N_13833);
or U14346 (N_14346,N_13661,N_13979);
xnor U14347 (N_14347,N_13884,N_13771);
and U14348 (N_14348,N_13779,N_13831);
nand U14349 (N_14349,N_13537,N_13940);
nand U14350 (N_14350,N_13989,N_13511);
nor U14351 (N_14351,N_13960,N_13585);
xnor U14352 (N_14352,N_13561,N_13527);
xnor U14353 (N_14353,N_13691,N_13621);
nor U14354 (N_14354,N_13539,N_13681);
nand U14355 (N_14355,N_13567,N_13793);
or U14356 (N_14356,N_13648,N_13525);
nor U14357 (N_14357,N_13966,N_13955);
nand U14358 (N_14358,N_13782,N_13832);
nor U14359 (N_14359,N_13584,N_13535);
xnor U14360 (N_14360,N_13877,N_13694);
nand U14361 (N_14361,N_13706,N_13783);
and U14362 (N_14362,N_13773,N_13731);
nor U14363 (N_14363,N_13862,N_13975);
xor U14364 (N_14364,N_13705,N_13719);
nand U14365 (N_14365,N_13837,N_13663);
nor U14366 (N_14366,N_13982,N_13751);
nor U14367 (N_14367,N_13933,N_13539);
nand U14368 (N_14368,N_13529,N_13879);
xor U14369 (N_14369,N_13870,N_13544);
nand U14370 (N_14370,N_13998,N_13746);
nand U14371 (N_14371,N_13752,N_13507);
nand U14372 (N_14372,N_13568,N_13834);
nor U14373 (N_14373,N_13946,N_13967);
and U14374 (N_14374,N_13641,N_13586);
nor U14375 (N_14375,N_13576,N_13836);
nor U14376 (N_14376,N_13637,N_13765);
xor U14377 (N_14377,N_13631,N_13644);
and U14378 (N_14378,N_13733,N_13512);
or U14379 (N_14379,N_13939,N_13629);
and U14380 (N_14380,N_13500,N_13670);
nor U14381 (N_14381,N_13989,N_13909);
nand U14382 (N_14382,N_13655,N_13943);
or U14383 (N_14383,N_13727,N_13808);
nand U14384 (N_14384,N_13954,N_13591);
nor U14385 (N_14385,N_13777,N_13641);
nor U14386 (N_14386,N_13926,N_13989);
nand U14387 (N_14387,N_13985,N_13828);
and U14388 (N_14388,N_13916,N_13586);
nand U14389 (N_14389,N_13565,N_13852);
and U14390 (N_14390,N_13824,N_13799);
or U14391 (N_14391,N_13556,N_13834);
or U14392 (N_14392,N_13776,N_13795);
and U14393 (N_14393,N_13598,N_13956);
and U14394 (N_14394,N_13770,N_13950);
xnor U14395 (N_14395,N_13849,N_13667);
and U14396 (N_14396,N_13974,N_13817);
nand U14397 (N_14397,N_13895,N_13788);
nand U14398 (N_14398,N_13593,N_13603);
nand U14399 (N_14399,N_13702,N_13998);
and U14400 (N_14400,N_13672,N_13746);
nand U14401 (N_14401,N_13783,N_13816);
xnor U14402 (N_14402,N_13930,N_13816);
and U14403 (N_14403,N_13723,N_13831);
and U14404 (N_14404,N_13861,N_13870);
xnor U14405 (N_14405,N_13680,N_13961);
nand U14406 (N_14406,N_13739,N_13880);
nor U14407 (N_14407,N_13853,N_13970);
xnor U14408 (N_14408,N_13676,N_13580);
xor U14409 (N_14409,N_13513,N_13911);
nor U14410 (N_14410,N_13958,N_13751);
xor U14411 (N_14411,N_13748,N_13930);
or U14412 (N_14412,N_13558,N_13635);
or U14413 (N_14413,N_13991,N_13660);
and U14414 (N_14414,N_13815,N_13801);
nand U14415 (N_14415,N_13695,N_13998);
nor U14416 (N_14416,N_13929,N_13783);
nor U14417 (N_14417,N_13768,N_13542);
and U14418 (N_14418,N_13868,N_13751);
and U14419 (N_14419,N_13630,N_13821);
nand U14420 (N_14420,N_13821,N_13894);
and U14421 (N_14421,N_13980,N_13671);
or U14422 (N_14422,N_13980,N_13816);
xor U14423 (N_14423,N_13723,N_13581);
nand U14424 (N_14424,N_13790,N_13659);
xor U14425 (N_14425,N_13746,N_13704);
nor U14426 (N_14426,N_13944,N_13843);
or U14427 (N_14427,N_13717,N_13636);
or U14428 (N_14428,N_13807,N_13529);
nor U14429 (N_14429,N_13701,N_13853);
nand U14430 (N_14430,N_13539,N_13903);
xnor U14431 (N_14431,N_13643,N_13743);
xnor U14432 (N_14432,N_13544,N_13919);
nand U14433 (N_14433,N_13844,N_13755);
or U14434 (N_14434,N_13775,N_13539);
and U14435 (N_14435,N_13656,N_13613);
nand U14436 (N_14436,N_13919,N_13932);
nor U14437 (N_14437,N_13886,N_13915);
nand U14438 (N_14438,N_13758,N_13536);
nor U14439 (N_14439,N_13740,N_13512);
nor U14440 (N_14440,N_13628,N_13919);
or U14441 (N_14441,N_13529,N_13961);
nand U14442 (N_14442,N_13914,N_13607);
nor U14443 (N_14443,N_13510,N_13903);
nand U14444 (N_14444,N_13962,N_13748);
xor U14445 (N_14445,N_13918,N_13571);
nor U14446 (N_14446,N_13687,N_13704);
xnor U14447 (N_14447,N_13596,N_13934);
nand U14448 (N_14448,N_13713,N_13592);
xnor U14449 (N_14449,N_13736,N_13857);
xnor U14450 (N_14450,N_13762,N_13676);
or U14451 (N_14451,N_13875,N_13850);
or U14452 (N_14452,N_13814,N_13605);
nor U14453 (N_14453,N_13624,N_13731);
and U14454 (N_14454,N_13863,N_13840);
xor U14455 (N_14455,N_13807,N_13824);
nor U14456 (N_14456,N_13578,N_13758);
xnor U14457 (N_14457,N_13830,N_13878);
and U14458 (N_14458,N_13992,N_13869);
nand U14459 (N_14459,N_13729,N_13584);
nor U14460 (N_14460,N_13633,N_13713);
or U14461 (N_14461,N_13582,N_13816);
or U14462 (N_14462,N_13971,N_13615);
and U14463 (N_14463,N_13642,N_13529);
and U14464 (N_14464,N_13895,N_13628);
xnor U14465 (N_14465,N_13992,N_13967);
nor U14466 (N_14466,N_13729,N_13788);
and U14467 (N_14467,N_13893,N_13629);
or U14468 (N_14468,N_13822,N_13517);
nand U14469 (N_14469,N_13610,N_13794);
and U14470 (N_14470,N_13656,N_13896);
nand U14471 (N_14471,N_13902,N_13564);
or U14472 (N_14472,N_13827,N_13814);
nor U14473 (N_14473,N_13616,N_13906);
or U14474 (N_14474,N_13922,N_13658);
and U14475 (N_14475,N_13804,N_13698);
nand U14476 (N_14476,N_13853,N_13904);
nor U14477 (N_14477,N_13769,N_13853);
and U14478 (N_14478,N_13844,N_13959);
or U14479 (N_14479,N_13557,N_13651);
xnor U14480 (N_14480,N_13534,N_13917);
xnor U14481 (N_14481,N_13862,N_13695);
or U14482 (N_14482,N_13724,N_13899);
nor U14483 (N_14483,N_13896,N_13735);
or U14484 (N_14484,N_13906,N_13679);
nor U14485 (N_14485,N_13504,N_13838);
xnor U14486 (N_14486,N_13771,N_13780);
xnor U14487 (N_14487,N_13781,N_13673);
nor U14488 (N_14488,N_13857,N_13734);
nand U14489 (N_14489,N_13575,N_13679);
nand U14490 (N_14490,N_13770,N_13742);
or U14491 (N_14491,N_13549,N_13570);
or U14492 (N_14492,N_13964,N_13704);
xnor U14493 (N_14493,N_13769,N_13776);
nand U14494 (N_14494,N_13855,N_13507);
or U14495 (N_14495,N_13727,N_13629);
nor U14496 (N_14496,N_13759,N_13903);
and U14497 (N_14497,N_13841,N_13912);
and U14498 (N_14498,N_13999,N_13871);
xnor U14499 (N_14499,N_13574,N_13918);
nand U14500 (N_14500,N_14004,N_14390);
nor U14501 (N_14501,N_14361,N_14293);
or U14502 (N_14502,N_14074,N_14456);
nor U14503 (N_14503,N_14044,N_14119);
nor U14504 (N_14504,N_14473,N_14404);
xor U14505 (N_14505,N_14124,N_14481);
nand U14506 (N_14506,N_14024,N_14317);
nand U14507 (N_14507,N_14335,N_14178);
and U14508 (N_14508,N_14288,N_14498);
nand U14509 (N_14509,N_14331,N_14191);
and U14510 (N_14510,N_14077,N_14365);
xnor U14511 (N_14511,N_14064,N_14341);
nor U14512 (N_14512,N_14427,N_14165);
nor U14513 (N_14513,N_14027,N_14069);
xor U14514 (N_14514,N_14471,N_14387);
nand U14515 (N_14515,N_14136,N_14266);
nand U14516 (N_14516,N_14388,N_14426);
xor U14517 (N_14517,N_14056,N_14296);
nor U14518 (N_14518,N_14139,N_14182);
nand U14519 (N_14519,N_14096,N_14130);
xnor U14520 (N_14520,N_14194,N_14318);
nor U14521 (N_14521,N_14241,N_14003);
nand U14522 (N_14522,N_14314,N_14227);
or U14523 (N_14523,N_14445,N_14180);
or U14524 (N_14524,N_14402,N_14185);
nor U14525 (N_14525,N_14378,N_14416);
and U14526 (N_14526,N_14115,N_14057);
nand U14527 (N_14527,N_14391,N_14176);
and U14528 (N_14528,N_14034,N_14190);
xnor U14529 (N_14529,N_14030,N_14443);
xor U14530 (N_14530,N_14138,N_14422);
xnor U14531 (N_14531,N_14472,N_14411);
nor U14532 (N_14532,N_14497,N_14028);
xnor U14533 (N_14533,N_14073,N_14453);
and U14534 (N_14534,N_14281,N_14273);
xnor U14535 (N_14535,N_14109,N_14359);
and U14536 (N_14536,N_14389,N_14268);
nor U14537 (N_14537,N_14171,N_14491);
nor U14538 (N_14538,N_14320,N_14222);
nand U14539 (N_14539,N_14258,N_14032);
nor U14540 (N_14540,N_14282,N_14214);
nor U14541 (N_14541,N_14035,N_14110);
and U14542 (N_14542,N_14496,N_14257);
nand U14543 (N_14543,N_14099,N_14450);
or U14544 (N_14544,N_14249,N_14114);
and U14545 (N_14545,N_14458,N_14446);
nand U14546 (N_14546,N_14006,N_14184);
or U14547 (N_14547,N_14187,N_14368);
nand U14548 (N_14548,N_14019,N_14428);
and U14549 (N_14549,N_14488,N_14122);
xnor U14550 (N_14550,N_14403,N_14215);
and U14551 (N_14551,N_14183,N_14291);
nor U14552 (N_14552,N_14013,N_14094);
xor U14553 (N_14553,N_14287,N_14083);
nor U14554 (N_14554,N_14143,N_14343);
and U14555 (N_14555,N_14098,N_14058);
or U14556 (N_14556,N_14093,N_14052);
or U14557 (N_14557,N_14381,N_14080);
or U14558 (N_14558,N_14452,N_14434);
and U14559 (N_14559,N_14448,N_14468);
nor U14560 (N_14560,N_14285,N_14499);
xor U14561 (N_14561,N_14465,N_14418);
or U14562 (N_14562,N_14367,N_14276);
nand U14563 (N_14563,N_14256,N_14487);
xnor U14564 (N_14564,N_14095,N_14157);
or U14565 (N_14565,N_14239,N_14356);
or U14566 (N_14566,N_14442,N_14342);
xor U14567 (N_14567,N_14477,N_14147);
xor U14568 (N_14568,N_14436,N_14237);
xor U14569 (N_14569,N_14201,N_14437);
or U14570 (N_14570,N_14170,N_14104);
nand U14571 (N_14571,N_14090,N_14181);
xor U14572 (N_14572,N_14346,N_14449);
nor U14573 (N_14573,N_14008,N_14125);
xnor U14574 (N_14574,N_14290,N_14275);
nor U14575 (N_14575,N_14113,N_14020);
nand U14576 (N_14576,N_14200,N_14066);
and U14577 (N_14577,N_14357,N_14055);
nor U14578 (N_14578,N_14467,N_14349);
and U14579 (N_14579,N_14235,N_14304);
nor U14580 (N_14580,N_14204,N_14264);
nor U14581 (N_14581,N_14306,N_14313);
and U14582 (N_14582,N_14330,N_14039);
xor U14583 (N_14583,N_14021,N_14267);
nor U14584 (N_14584,N_14223,N_14360);
nor U14585 (N_14585,N_14482,N_14192);
xnor U14586 (N_14586,N_14326,N_14259);
xor U14587 (N_14587,N_14406,N_14302);
nand U14588 (N_14588,N_14203,N_14161);
and U14589 (N_14589,N_14144,N_14230);
nor U14590 (N_14590,N_14474,N_14175);
nor U14591 (N_14591,N_14242,N_14229);
nor U14592 (N_14592,N_14174,N_14251);
or U14593 (N_14593,N_14186,N_14345);
and U14594 (N_14594,N_14061,N_14071);
xor U14595 (N_14595,N_14451,N_14483);
and U14596 (N_14596,N_14172,N_14038);
nor U14597 (N_14597,N_14141,N_14211);
and U14598 (N_14598,N_14433,N_14134);
or U14599 (N_14599,N_14091,N_14219);
nor U14600 (N_14600,N_14475,N_14271);
and U14601 (N_14601,N_14196,N_14016);
or U14602 (N_14602,N_14392,N_14105);
nor U14603 (N_14603,N_14348,N_14375);
nor U14604 (N_14604,N_14148,N_14370);
nand U14605 (N_14605,N_14126,N_14455);
nor U14606 (N_14606,N_14207,N_14212);
and U14607 (N_14607,N_14396,N_14398);
nand U14608 (N_14608,N_14255,N_14407);
and U14609 (N_14609,N_14243,N_14344);
or U14610 (N_14610,N_14131,N_14492);
and U14611 (N_14611,N_14294,N_14250);
or U14612 (N_14612,N_14132,N_14233);
nor U14613 (N_14613,N_14197,N_14059);
xnor U14614 (N_14614,N_14202,N_14352);
nand U14615 (N_14615,N_14156,N_14060);
nand U14616 (N_14616,N_14459,N_14364);
and U14617 (N_14617,N_14167,N_14007);
nand U14618 (N_14618,N_14079,N_14189);
and U14619 (N_14619,N_14373,N_14009);
and U14620 (N_14620,N_14089,N_14305);
nor U14621 (N_14621,N_14307,N_14309);
nor U14622 (N_14622,N_14254,N_14031);
nand U14623 (N_14623,N_14046,N_14026);
xnor U14624 (N_14624,N_14253,N_14123);
nand U14625 (N_14625,N_14081,N_14311);
xor U14626 (N_14626,N_14133,N_14469);
or U14627 (N_14627,N_14193,N_14289);
nor U14628 (N_14628,N_14012,N_14308);
nor U14629 (N_14629,N_14128,N_14423);
nor U14630 (N_14630,N_14022,N_14333);
and U14631 (N_14631,N_14067,N_14414);
nor U14632 (N_14632,N_14100,N_14374);
or U14633 (N_14633,N_14236,N_14277);
xnor U14634 (N_14634,N_14260,N_14262);
nor U14635 (N_14635,N_14041,N_14279);
and U14636 (N_14636,N_14419,N_14023);
nand U14637 (N_14637,N_14085,N_14158);
xnor U14638 (N_14638,N_14142,N_14466);
or U14639 (N_14639,N_14232,N_14315);
and U14640 (N_14640,N_14199,N_14076);
nand U14641 (N_14641,N_14160,N_14429);
xor U14642 (N_14642,N_14238,N_14462);
nor U14643 (N_14643,N_14420,N_14018);
nand U14644 (N_14644,N_14447,N_14278);
nor U14645 (N_14645,N_14297,N_14301);
nor U14646 (N_14646,N_14351,N_14327);
nand U14647 (N_14647,N_14337,N_14412);
xnor U14648 (N_14648,N_14217,N_14065);
nand U14649 (N_14649,N_14086,N_14284);
and U14650 (N_14650,N_14213,N_14108);
xor U14651 (N_14651,N_14321,N_14051);
nand U14652 (N_14652,N_14169,N_14033);
xnor U14653 (N_14653,N_14394,N_14206);
xnor U14654 (N_14654,N_14386,N_14017);
nor U14655 (N_14655,N_14493,N_14188);
nor U14656 (N_14656,N_14303,N_14405);
nor U14657 (N_14657,N_14377,N_14036);
nand U14658 (N_14658,N_14154,N_14270);
nor U14659 (N_14659,N_14347,N_14298);
xor U14660 (N_14660,N_14216,N_14002);
and U14661 (N_14661,N_14140,N_14042);
and U14662 (N_14662,N_14478,N_14438);
and U14663 (N_14663,N_14400,N_14231);
or U14664 (N_14664,N_14265,N_14454);
nand U14665 (N_14665,N_14103,N_14162);
nor U14666 (N_14666,N_14116,N_14424);
and U14667 (N_14667,N_14362,N_14334);
nand U14668 (N_14668,N_14025,N_14261);
xnor U14669 (N_14669,N_14399,N_14484);
xor U14670 (N_14670,N_14149,N_14168);
nand U14671 (N_14671,N_14107,N_14226);
xnor U14672 (N_14672,N_14218,N_14379);
xnor U14673 (N_14673,N_14382,N_14111);
or U14674 (N_14674,N_14355,N_14470);
nor U14675 (N_14675,N_14152,N_14208);
xor U14676 (N_14676,N_14048,N_14247);
nor U14677 (N_14677,N_14040,N_14054);
xnor U14678 (N_14678,N_14118,N_14015);
nor U14679 (N_14679,N_14324,N_14310);
or U14680 (N_14680,N_14380,N_14353);
or U14681 (N_14681,N_14043,N_14408);
xnor U14682 (N_14682,N_14283,N_14430);
nor U14683 (N_14683,N_14363,N_14106);
nor U14684 (N_14684,N_14205,N_14441);
or U14685 (N_14685,N_14248,N_14316);
or U14686 (N_14686,N_14121,N_14485);
nand U14687 (N_14687,N_14486,N_14173);
or U14688 (N_14688,N_14409,N_14252);
or U14689 (N_14689,N_14244,N_14385);
xor U14690 (N_14690,N_14129,N_14120);
xor U14691 (N_14691,N_14461,N_14135);
nand U14692 (N_14692,N_14146,N_14371);
xnor U14693 (N_14693,N_14087,N_14166);
xnor U14694 (N_14694,N_14457,N_14228);
nor U14695 (N_14695,N_14300,N_14350);
or U14696 (N_14696,N_14417,N_14045);
xnor U14697 (N_14697,N_14401,N_14272);
xnor U14698 (N_14698,N_14490,N_14463);
nor U14699 (N_14699,N_14210,N_14274);
and U14700 (N_14700,N_14005,N_14383);
and U14701 (N_14701,N_14137,N_14101);
or U14702 (N_14702,N_14415,N_14397);
nand U14703 (N_14703,N_14286,N_14070);
xnor U14704 (N_14704,N_14435,N_14476);
nor U14705 (N_14705,N_14464,N_14332);
xor U14706 (N_14706,N_14376,N_14102);
xnor U14707 (N_14707,N_14280,N_14340);
or U14708 (N_14708,N_14323,N_14225);
nand U14709 (N_14709,N_14245,N_14092);
nor U14710 (N_14710,N_14037,N_14112);
xor U14711 (N_14711,N_14439,N_14117);
nor U14712 (N_14712,N_14068,N_14489);
nand U14713 (N_14713,N_14329,N_14495);
nor U14714 (N_14714,N_14440,N_14177);
nand U14715 (N_14715,N_14372,N_14047);
and U14716 (N_14716,N_14000,N_14049);
and U14717 (N_14717,N_14050,N_14369);
nand U14718 (N_14718,N_14011,N_14413);
or U14719 (N_14719,N_14336,N_14312);
nand U14720 (N_14720,N_14292,N_14153);
and U14721 (N_14721,N_14480,N_14322);
xnor U14722 (N_14722,N_14209,N_14339);
or U14723 (N_14723,N_14224,N_14240);
and U14724 (N_14724,N_14063,N_14150);
or U14725 (N_14725,N_14366,N_14159);
nor U14726 (N_14726,N_14421,N_14145);
and U14727 (N_14727,N_14299,N_14127);
or U14728 (N_14728,N_14384,N_14494);
or U14729 (N_14729,N_14395,N_14444);
or U14730 (N_14730,N_14269,N_14179);
or U14731 (N_14731,N_14460,N_14075);
and U14732 (N_14732,N_14151,N_14221);
nand U14733 (N_14733,N_14084,N_14164);
xnor U14734 (N_14734,N_14246,N_14078);
or U14735 (N_14735,N_14029,N_14014);
or U14736 (N_14736,N_14088,N_14234);
xnor U14737 (N_14737,N_14195,N_14053);
xor U14738 (N_14738,N_14001,N_14198);
and U14739 (N_14739,N_14295,N_14163);
xnor U14740 (N_14740,N_14425,N_14358);
xor U14741 (N_14741,N_14062,N_14082);
nand U14742 (N_14742,N_14010,N_14155);
xnor U14743 (N_14743,N_14325,N_14328);
and U14744 (N_14744,N_14097,N_14220);
nand U14745 (N_14745,N_14431,N_14263);
xor U14746 (N_14746,N_14393,N_14410);
or U14747 (N_14747,N_14354,N_14072);
nor U14748 (N_14748,N_14479,N_14338);
xor U14749 (N_14749,N_14432,N_14319);
and U14750 (N_14750,N_14218,N_14126);
nor U14751 (N_14751,N_14023,N_14204);
nand U14752 (N_14752,N_14066,N_14088);
xnor U14753 (N_14753,N_14122,N_14358);
and U14754 (N_14754,N_14401,N_14182);
xnor U14755 (N_14755,N_14073,N_14033);
nand U14756 (N_14756,N_14138,N_14482);
and U14757 (N_14757,N_14198,N_14069);
or U14758 (N_14758,N_14423,N_14232);
and U14759 (N_14759,N_14288,N_14467);
and U14760 (N_14760,N_14475,N_14297);
and U14761 (N_14761,N_14016,N_14164);
and U14762 (N_14762,N_14210,N_14080);
or U14763 (N_14763,N_14012,N_14406);
nor U14764 (N_14764,N_14081,N_14477);
and U14765 (N_14765,N_14437,N_14209);
nor U14766 (N_14766,N_14229,N_14160);
and U14767 (N_14767,N_14294,N_14184);
or U14768 (N_14768,N_14407,N_14280);
and U14769 (N_14769,N_14137,N_14390);
nor U14770 (N_14770,N_14043,N_14426);
xnor U14771 (N_14771,N_14468,N_14317);
or U14772 (N_14772,N_14172,N_14447);
nor U14773 (N_14773,N_14398,N_14203);
or U14774 (N_14774,N_14255,N_14473);
and U14775 (N_14775,N_14238,N_14176);
and U14776 (N_14776,N_14014,N_14172);
nor U14777 (N_14777,N_14442,N_14162);
and U14778 (N_14778,N_14164,N_14111);
xor U14779 (N_14779,N_14054,N_14201);
nand U14780 (N_14780,N_14187,N_14385);
xor U14781 (N_14781,N_14007,N_14420);
or U14782 (N_14782,N_14280,N_14366);
nor U14783 (N_14783,N_14166,N_14106);
nor U14784 (N_14784,N_14037,N_14110);
xor U14785 (N_14785,N_14156,N_14325);
xor U14786 (N_14786,N_14158,N_14494);
and U14787 (N_14787,N_14108,N_14066);
and U14788 (N_14788,N_14276,N_14112);
nand U14789 (N_14789,N_14307,N_14019);
xnor U14790 (N_14790,N_14131,N_14027);
nand U14791 (N_14791,N_14153,N_14120);
nor U14792 (N_14792,N_14083,N_14234);
nand U14793 (N_14793,N_14008,N_14013);
nor U14794 (N_14794,N_14274,N_14440);
or U14795 (N_14795,N_14195,N_14391);
nor U14796 (N_14796,N_14480,N_14469);
and U14797 (N_14797,N_14381,N_14373);
and U14798 (N_14798,N_14224,N_14270);
xnor U14799 (N_14799,N_14051,N_14139);
nand U14800 (N_14800,N_14028,N_14474);
nor U14801 (N_14801,N_14486,N_14109);
xor U14802 (N_14802,N_14106,N_14475);
and U14803 (N_14803,N_14072,N_14046);
nand U14804 (N_14804,N_14092,N_14141);
nor U14805 (N_14805,N_14488,N_14213);
nand U14806 (N_14806,N_14295,N_14106);
and U14807 (N_14807,N_14029,N_14260);
nand U14808 (N_14808,N_14095,N_14314);
and U14809 (N_14809,N_14377,N_14145);
nor U14810 (N_14810,N_14393,N_14040);
nor U14811 (N_14811,N_14217,N_14327);
xnor U14812 (N_14812,N_14127,N_14050);
nor U14813 (N_14813,N_14192,N_14494);
xnor U14814 (N_14814,N_14152,N_14047);
and U14815 (N_14815,N_14172,N_14027);
nand U14816 (N_14816,N_14162,N_14376);
and U14817 (N_14817,N_14439,N_14260);
or U14818 (N_14818,N_14227,N_14274);
nand U14819 (N_14819,N_14114,N_14380);
or U14820 (N_14820,N_14008,N_14379);
or U14821 (N_14821,N_14211,N_14156);
or U14822 (N_14822,N_14210,N_14132);
nand U14823 (N_14823,N_14403,N_14097);
or U14824 (N_14824,N_14449,N_14260);
nor U14825 (N_14825,N_14151,N_14405);
xnor U14826 (N_14826,N_14307,N_14097);
nand U14827 (N_14827,N_14457,N_14049);
nor U14828 (N_14828,N_14146,N_14123);
xnor U14829 (N_14829,N_14393,N_14250);
nand U14830 (N_14830,N_14034,N_14092);
nor U14831 (N_14831,N_14324,N_14315);
nand U14832 (N_14832,N_14082,N_14317);
nor U14833 (N_14833,N_14048,N_14000);
nor U14834 (N_14834,N_14148,N_14357);
or U14835 (N_14835,N_14345,N_14050);
or U14836 (N_14836,N_14388,N_14402);
xor U14837 (N_14837,N_14478,N_14331);
nand U14838 (N_14838,N_14078,N_14354);
nor U14839 (N_14839,N_14307,N_14258);
nor U14840 (N_14840,N_14437,N_14269);
nor U14841 (N_14841,N_14301,N_14232);
and U14842 (N_14842,N_14088,N_14002);
or U14843 (N_14843,N_14016,N_14305);
xnor U14844 (N_14844,N_14162,N_14022);
nor U14845 (N_14845,N_14009,N_14496);
nor U14846 (N_14846,N_14210,N_14314);
nor U14847 (N_14847,N_14099,N_14413);
or U14848 (N_14848,N_14483,N_14256);
nand U14849 (N_14849,N_14337,N_14354);
nand U14850 (N_14850,N_14368,N_14464);
nand U14851 (N_14851,N_14267,N_14371);
and U14852 (N_14852,N_14070,N_14209);
nand U14853 (N_14853,N_14363,N_14372);
nand U14854 (N_14854,N_14442,N_14291);
nor U14855 (N_14855,N_14311,N_14395);
or U14856 (N_14856,N_14487,N_14232);
and U14857 (N_14857,N_14269,N_14136);
xor U14858 (N_14858,N_14469,N_14401);
nand U14859 (N_14859,N_14114,N_14050);
xnor U14860 (N_14860,N_14450,N_14257);
xnor U14861 (N_14861,N_14311,N_14114);
nor U14862 (N_14862,N_14487,N_14455);
or U14863 (N_14863,N_14020,N_14491);
nand U14864 (N_14864,N_14333,N_14016);
and U14865 (N_14865,N_14130,N_14108);
xor U14866 (N_14866,N_14350,N_14307);
xor U14867 (N_14867,N_14367,N_14466);
and U14868 (N_14868,N_14275,N_14326);
or U14869 (N_14869,N_14069,N_14439);
nor U14870 (N_14870,N_14015,N_14022);
nor U14871 (N_14871,N_14110,N_14139);
nor U14872 (N_14872,N_14440,N_14402);
nor U14873 (N_14873,N_14066,N_14431);
nor U14874 (N_14874,N_14139,N_14042);
nor U14875 (N_14875,N_14278,N_14344);
nor U14876 (N_14876,N_14260,N_14074);
nor U14877 (N_14877,N_14434,N_14062);
nand U14878 (N_14878,N_14450,N_14034);
nor U14879 (N_14879,N_14132,N_14186);
nor U14880 (N_14880,N_14381,N_14487);
nor U14881 (N_14881,N_14294,N_14413);
and U14882 (N_14882,N_14239,N_14482);
nand U14883 (N_14883,N_14232,N_14432);
or U14884 (N_14884,N_14141,N_14239);
nor U14885 (N_14885,N_14188,N_14101);
or U14886 (N_14886,N_14162,N_14326);
nand U14887 (N_14887,N_14433,N_14231);
xnor U14888 (N_14888,N_14101,N_14403);
nor U14889 (N_14889,N_14443,N_14355);
and U14890 (N_14890,N_14401,N_14168);
or U14891 (N_14891,N_14193,N_14438);
xnor U14892 (N_14892,N_14321,N_14044);
nand U14893 (N_14893,N_14366,N_14419);
nand U14894 (N_14894,N_14118,N_14003);
nand U14895 (N_14895,N_14237,N_14462);
and U14896 (N_14896,N_14450,N_14202);
nor U14897 (N_14897,N_14420,N_14336);
nand U14898 (N_14898,N_14154,N_14007);
or U14899 (N_14899,N_14464,N_14013);
xor U14900 (N_14900,N_14054,N_14112);
nor U14901 (N_14901,N_14003,N_14306);
nor U14902 (N_14902,N_14462,N_14057);
nor U14903 (N_14903,N_14338,N_14298);
xor U14904 (N_14904,N_14489,N_14094);
or U14905 (N_14905,N_14230,N_14090);
or U14906 (N_14906,N_14364,N_14408);
xnor U14907 (N_14907,N_14388,N_14359);
nor U14908 (N_14908,N_14178,N_14341);
xor U14909 (N_14909,N_14358,N_14004);
and U14910 (N_14910,N_14120,N_14448);
and U14911 (N_14911,N_14357,N_14390);
and U14912 (N_14912,N_14012,N_14389);
or U14913 (N_14913,N_14254,N_14408);
xnor U14914 (N_14914,N_14382,N_14172);
or U14915 (N_14915,N_14225,N_14483);
xnor U14916 (N_14916,N_14074,N_14008);
or U14917 (N_14917,N_14081,N_14376);
and U14918 (N_14918,N_14115,N_14247);
nor U14919 (N_14919,N_14236,N_14405);
nor U14920 (N_14920,N_14246,N_14462);
nor U14921 (N_14921,N_14428,N_14287);
xor U14922 (N_14922,N_14393,N_14022);
and U14923 (N_14923,N_14292,N_14378);
nand U14924 (N_14924,N_14018,N_14010);
xor U14925 (N_14925,N_14018,N_14119);
or U14926 (N_14926,N_14473,N_14468);
nand U14927 (N_14927,N_14125,N_14342);
nand U14928 (N_14928,N_14428,N_14096);
or U14929 (N_14929,N_14285,N_14029);
and U14930 (N_14930,N_14021,N_14392);
or U14931 (N_14931,N_14038,N_14287);
and U14932 (N_14932,N_14022,N_14483);
nand U14933 (N_14933,N_14084,N_14243);
xor U14934 (N_14934,N_14410,N_14485);
and U14935 (N_14935,N_14099,N_14089);
nor U14936 (N_14936,N_14059,N_14445);
nand U14937 (N_14937,N_14026,N_14337);
nor U14938 (N_14938,N_14435,N_14176);
nor U14939 (N_14939,N_14303,N_14135);
nand U14940 (N_14940,N_14461,N_14499);
and U14941 (N_14941,N_14038,N_14191);
or U14942 (N_14942,N_14233,N_14089);
xnor U14943 (N_14943,N_14120,N_14481);
nor U14944 (N_14944,N_14185,N_14391);
and U14945 (N_14945,N_14162,N_14054);
nand U14946 (N_14946,N_14064,N_14018);
and U14947 (N_14947,N_14431,N_14474);
and U14948 (N_14948,N_14270,N_14327);
or U14949 (N_14949,N_14408,N_14206);
and U14950 (N_14950,N_14048,N_14361);
and U14951 (N_14951,N_14000,N_14478);
and U14952 (N_14952,N_14375,N_14153);
or U14953 (N_14953,N_14367,N_14362);
xnor U14954 (N_14954,N_14180,N_14487);
or U14955 (N_14955,N_14250,N_14412);
xor U14956 (N_14956,N_14068,N_14477);
or U14957 (N_14957,N_14299,N_14460);
xor U14958 (N_14958,N_14217,N_14117);
nor U14959 (N_14959,N_14395,N_14059);
or U14960 (N_14960,N_14148,N_14038);
xnor U14961 (N_14961,N_14373,N_14409);
and U14962 (N_14962,N_14165,N_14391);
xnor U14963 (N_14963,N_14294,N_14329);
and U14964 (N_14964,N_14323,N_14435);
or U14965 (N_14965,N_14042,N_14043);
or U14966 (N_14966,N_14037,N_14375);
and U14967 (N_14967,N_14115,N_14061);
nand U14968 (N_14968,N_14123,N_14159);
nand U14969 (N_14969,N_14367,N_14295);
and U14970 (N_14970,N_14138,N_14081);
or U14971 (N_14971,N_14496,N_14406);
xor U14972 (N_14972,N_14268,N_14197);
xnor U14973 (N_14973,N_14319,N_14368);
and U14974 (N_14974,N_14342,N_14224);
nand U14975 (N_14975,N_14329,N_14060);
and U14976 (N_14976,N_14335,N_14150);
nand U14977 (N_14977,N_14277,N_14497);
or U14978 (N_14978,N_14274,N_14347);
or U14979 (N_14979,N_14391,N_14038);
and U14980 (N_14980,N_14156,N_14250);
nand U14981 (N_14981,N_14068,N_14070);
and U14982 (N_14982,N_14069,N_14012);
nand U14983 (N_14983,N_14094,N_14252);
and U14984 (N_14984,N_14352,N_14296);
or U14985 (N_14985,N_14463,N_14233);
or U14986 (N_14986,N_14366,N_14188);
nor U14987 (N_14987,N_14014,N_14247);
xor U14988 (N_14988,N_14318,N_14423);
nand U14989 (N_14989,N_14283,N_14471);
or U14990 (N_14990,N_14157,N_14054);
and U14991 (N_14991,N_14388,N_14003);
and U14992 (N_14992,N_14281,N_14150);
xor U14993 (N_14993,N_14435,N_14395);
or U14994 (N_14994,N_14180,N_14221);
or U14995 (N_14995,N_14401,N_14416);
and U14996 (N_14996,N_14132,N_14301);
and U14997 (N_14997,N_14124,N_14008);
nor U14998 (N_14998,N_14487,N_14076);
or U14999 (N_14999,N_14265,N_14059);
or U15000 (N_15000,N_14921,N_14624);
nor U15001 (N_15001,N_14840,N_14774);
nand U15002 (N_15002,N_14877,N_14611);
nor U15003 (N_15003,N_14525,N_14502);
or U15004 (N_15004,N_14990,N_14958);
nor U15005 (N_15005,N_14541,N_14671);
and U15006 (N_15006,N_14759,N_14597);
nor U15007 (N_15007,N_14803,N_14581);
nor U15008 (N_15008,N_14507,N_14833);
nor U15009 (N_15009,N_14655,N_14792);
nor U15010 (N_15010,N_14549,N_14865);
nand U15011 (N_15011,N_14704,N_14646);
xor U15012 (N_15012,N_14657,N_14669);
nor U15013 (N_15013,N_14668,N_14588);
and U15014 (N_15014,N_14587,N_14500);
nand U15015 (N_15015,N_14640,N_14816);
and U15016 (N_15016,N_14690,N_14701);
and U15017 (N_15017,N_14828,N_14911);
nor U15018 (N_15018,N_14736,N_14749);
or U15019 (N_15019,N_14560,N_14880);
xor U15020 (N_15020,N_14805,N_14943);
and U15021 (N_15021,N_14707,N_14532);
nand U15022 (N_15022,N_14940,N_14686);
nor U15023 (N_15023,N_14658,N_14579);
and U15024 (N_15024,N_14798,N_14544);
nor U15025 (N_15025,N_14772,N_14815);
or U15026 (N_15026,N_14599,N_14741);
nor U15027 (N_15027,N_14819,N_14698);
or U15028 (N_15028,N_14562,N_14823);
nand U15029 (N_15029,N_14512,N_14786);
or U15030 (N_15030,N_14950,N_14710);
xor U15031 (N_15031,N_14547,N_14769);
xnor U15032 (N_15032,N_14553,N_14652);
xor U15033 (N_15033,N_14607,N_14945);
and U15034 (N_15034,N_14675,N_14585);
or U15035 (N_15035,N_14825,N_14610);
and U15036 (N_15036,N_14948,N_14648);
nor U15037 (N_15037,N_14746,N_14785);
or U15038 (N_15038,N_14586,N_14724);
nand U15039 (N_15039,N_14885,N_14670);
or U15040 (N_15040,N_14720,N_14901);
nand U15041 (N_15041,N_14931,N_14959);
xnor U15042 (N_15042,N_14888,N_14776);
or U15043 (N_15043,N_14723,N_14995);
or U15044 (N_15044,N_14807,N_14756);
and U15045 (N_15045,N_14519,N_14691);
and U15046 (N_15046,N_14784,N_14947);
nand U15047 (N_15047,N_14946,N_14837);
nand U15048 (N_15048,N_14557,N_14522);
nand U15049 (N_15049,N_14808,N_14893);
xor U15050 (N_15050,N_14683,N_14978);
nand U15051 (N_15051,N_14856,N_14956);
and U15052 (N_15052,N_14580,N_14713);
nand U15053 (N_15053,N_14732,N_14575);
xor U15054 (N_15054,N_14859,N_14853);
or U15055 (N_15055,N_14501,N_14666);
nand U15056 (N_15056,N_14700,N_14738);
nand U15057 (N_15057,N_14743,N_14902);
or U15058 (N_15058,N_14685,N_14899);
xnor U15059 (N_15059,N_14578,N_14509);
or U15060 (N_15060,N_14534,N_14747);
and U15061 (N_15061,N_14895,N_14603);
nor U15062 (N_15062,N_14829,N_14552);
xor U15063 (N_15063,N_14735,N_14886);
nor U15064 (N_15064,N_14768,N_14633);
xnor U15065 (N_15065,N_14625,N_14752);
or U15066 (N_15066,N_14684,N_14836);
and U15067 (N_15067,N_14653,N_14842);
and U15068 (N_15068,N_14524,N_14745);
nand U15069 (N_15069,N_14908,N_14674);
nand U15070 (N_15070,N_14764,N_14639);
nand U15071 (N_15071,N_14504,N_14518);
nor U15072 (N_15072,N_14744,N_14705);
nand U15073 (N_15073,N_14656,N_14935);
and U15074 (N_15074,N_14996,N_14844);
nor U15075 (N_15075,N_14926,N_14667);
nor U15076 (N_15076,N_14672,N_14876);
nand U15077 (N_15077,N_14916,N_14687);
and U15078 (N_15078,N_14697,N_14968);
nand U15079 (N_15079,N_14712,N_14716);
nand U15080 (N_15080,N_14878,N_14922);
and U15081 (N_15081,N_14788,N_14708);
nor U15082 (N_15082,N_14548,N_14917);
and U15083 (N_15083,N_14600,N_14527);
and U15084 (N_15084,N_14538,N_14702);
nor U15085 (N_15085,N_14944,N_14802);
xnor U15086 (N_15086,N_14626,N_14847);
or U15087 (N_15087,N_14750,N_14550);
and U15088 (N_15088,N_14602,N_14540);
nor U15089 (N_15089,N_14869,N_14554);
xnor U15090 (N_15090,N_14711,N_14559);
nor U15091 (N_15091,N_14595,N_14972);
and U15092 (N_15092,N_14883,N_14900);
xor U15093 (N_15093,N_14851,N_14887);
and U15094 (N_15094,N_14835,N_14634);
and U15095 (N_15095,N_14632,N_14766);
and U15096 (N_15096,N_14967,N_14546);
nor U15097 (N_15097,N_14521,N_14986);
nand U15098 (N_15098,N_14535,N_14635);
nand U15099 (N_15099,N_14574,N_14979);
or U15100 (N_15100,N_14678,N_14849);
and U15101 (N_15101,N_14755,N_14728);
or U15102 (N_15102,N_14934,N_14993);
or U15103 (N_15103,N_14629,N_14976);
or U15104 (N_15104,N_14693,N_14604);
or U15105 (N_15105,N_14841,N_14695);
nand U15106 (N_15106,N_14614,N_14918);
or U15107 (N_15107,N_14644,N_14962);
nor U15108 (N_15108,N_14520,N_14665);
and U15109 (N_15109,N_14928,N_14912);
xor U15110 (N_15110,N_14778,N_14866);
xor U15111 (N_15111,N_14981,N_14861);
nor U15112 (N_15112,N_14570,N_14742);
or U15113 (N_15113,N_14660,N_14894);
xor U15114 (N_15114,N_14858,N_14636);
and U15115 (N_15115,N_14622,N_14542);
and U15116 (N_15116,N_14960,N_14645);
nor U15117 (N_15117,N_14620,N_14564);
and U15118 (N_15118,N_14868,N_14761);
nor U15119 (N_15119,N_14970,N_14999);
xor U15120 (N_15120,N_14867,N_14654);
nor U15121 (N_15121,N_14925,N_14551);
xor U15122 (N_15122,N_14545,N_14757);
xor U15123 (N_15123,N_14814,N_14832);
nor U15124 (N_15124,N_14664,N_14923);
nand U15125 (N_15125,N_14590,N_14826);
nand U15126 (N_15126,N_14513,N_14619);
and U15127 (N_15127,N_14872,N_14838);
nand U15128 (N_15128,N_14642,N_14754);
or U15129 (N_15129,N_14677,N_14953);
nand U15130 (N_15130,N_14801,N_14572);
nor U15131 (N_15131,N_14992,N_14719);
and U15132 (N_15132,N_14966,N_14939);
and U15133 (N_15133,N_14909,N_14680);
xor U15134 (N_15134,N_14818,N_14884);
nand U15135 (N_15135,N_14739,N_14517);
nor U15136 (N_15136,N_14650,N_14827);
nor U15137 (N_15137,N_14523,N_14643);
and U15138 (N_15138,N_14563,N_14860);
nand U15139 (N_15139,N_14904,N_14806);
nand U15140 (N_15140,N_14810,N_14591);
and U15141 (N_15141,N_14601,N_14848);
or U15142 (N_15142,N_14651,N_14955);
xor U15143 (N_15143,N_14543,N_14906);
nand U15144 (N_15144,N_14773,N_14796);
or U15145 (N_15145,N_14717,N_14689);
nor U15146 (N_15146,N_14688,N_14714);
xor U15147 (N_15147,N_14526,N_14514);
nand U15148 (N_15148,N_14516,N_14852);
and U15149 (N_15149,N_14615,N_14982);
and U15150 (N_15150,N_14594,N_14973);
and U15151 (N_15151,N_14791,N_14751);
nor U15152 (N_15152,N_14977,N_14725);
xor U15153 (N_15153,N_14598,N_14617);
and U15154 (N_15154,N_14775,N_14910);
nand U15155 (N_15155,N_14539,N_14682);
xnor U15156 (N_15156,N_14567,N_14797);
xnor U15157 (N_15157,N_14609,N_14531);
or U15158 (N_15158,N_14936,N_14927);
and U15159 (N_15159,N_14941,N_14854);
xor U15160 (N_15160,N_14957,N_14506);
or U15161 (N_15161,N_14963,N_14627);
or U15162 (N_15162,N_14790,N_14729);
and U15163 (N_15163,N_14855,N_14718);
or U15164 (N_15164,N_14954,N_14997);
nand U15165 (N_15165,N_14882,N_14621);
nand U15166 (N_15166,N_14830,N_14932);
xor U15167 (N_15167,N_14795,N_14782);
or U15168 (N_15168,N_14577,N_14987);
nor U15169 (N_15169,N_14879,N_14951);
nor U15170 (N_15170,N_14613,N_14679);
nand U15171 (N_15171,N_14571,N_14845);
nand U15172 (N_15172,N_14793,N_14616);
xnor U15173 (N_15173,N_14813,N_14737);
or U15174 (N_15174,N_14989,N_14771);
nand U15175 (N_15175,N_14748,N_14920);
or U15176 (N_15176,N_14628,N_14804);
nor U15177 (N_15177,N_14789,N_14783);
and U15178 (N_15178,N_14794,N_14726);
nor U15179 (N_15179,N_14647,N_14905);
and U15180 (N_15180,N_14722,N_14938);
or U15181 (N_15181,N_14753,N_14965);
nand U15182 (N_15182,N_14529,N_14800);
nor U15183 (N_15183,N_14638,N_14846);
nor U15184 (N_15184,N_14843,N_14929);
xnor U15185 (N_15185,N_14873,N_14809);
xnor U15186 (N_15186,N_14781,N_14907);
or U15187 (N_15187,N_14662,N_14530);
nor U15188 (N_15188,N_14631,N_14508);
nand U15189 (N_15189,N_14582,N_14758);
nor U15190 (N_15190,N_14817,N_14555);
nor U15191 (N_15191,N_14676,N_14511);
nand U15192 (N_15192,N_14596,N_14949);
xnor U15193 (N_15193,N_14515,N_14974);
and U15194 (N_15194,N_14980,N_14566);
nand U15195 (N_15195,N_14891,N_14537);
xnor U15196 (N_15196,N_14780,N_14898);
or U15197 (N_15197,N_14767,N_14681);
and U15198 (N_15198,N_14975,N_14937);
xnor U15199 (N_15199,N_14952,N_14503);
and U15200 (N_15200,N_14994,N_14762);
nor U15201 (N_15201,N_14933,N_14623);
or U15202 (N_15202,N_14998,N_14839);
or U15203 (N_15203,N_14661,N_14770);
xnor U15204 (N_15204,N_14733,N_14914);
nand U15205 (N_15205,N_14734,N_14727);
or U15206 (N_15206,N_14881,N_14593);
nand U15207 (N_15207,N_14584,N_14897);
or U15208 (N_15208,N_14692,N_14696);
nor U15209 (N_15209,N_14663,N_14760);
nor U15210 (N_15210,N_14862,N_14558);
and U15211 (N_15211,N_14942,N_14533);
xor U15212 (N_15212,N_14569,N_14821);
nand U15213 (N_15213,N_14763,N_14592);
and U15214 (N_15214,N_14649,N_14820);
nor U15215 (N_15215,N_14694,N_14612);
nand U15216 (N_15216,N_14991,N_14703);
or U15217 (N_15217,N_14864,N_14988);
or U15218 (N_15218,N_14618,N_14870);
and U15219 (N_15219,N_14731,N_14874);
xor U15220 (N_15220,N_14984,N_14659);
nor U15221 (N_15221,N_14896,N_14699);
xor U15222 (N_15222,N_14871,N_14913);
nand U15223 (N_15223,N_14971,N_14779);
or U15224 (N_15224,N_14787,N_14589);
nor U15225 (N_15225,N_14857,N_14641);
nand U15226 (N_15226,N_14983,N_14583);
nand U15227 (N_15227,N_14969,N_14919);
xnor U15228 (N_15228,N_14824,N_14964);
or U15229 (N_15229,N_14889,N_14924);
xnor U15230 (N_15230,N_14930,N_14740);
or U15231 (N_15231,N_14721,N_14985);
or U15232 (N_15232,N_14961,N_14730);
xor U15233 (N_15233,N_14576,N_14765);
nor U15234 (N_15234,N_14556,N_14637);
or U15235 (N_15235,N_14811,N_14850);
nand U15236 (N_15236,N_14536,N_14715);
or U15237 (N_15237,N_14915,N_14510);
or U15238 (N_15238,N_14605,N_14777);
and U15239 (N_15239,N_14606,N_14528);
nand U15240 (N_15240,N_14863,N_14573);
nand U15241 (N_15241,N_14561,N_14831);
and U15242 (N_15242,N_14892,N_14568);
and U15243 (N_15243,N_14822,N_14706);
nor U15244 (N_15244,N_14890,N_14673);
and U15245 (N_15245,N_14812,N_14505);
or U15246 (N_15246,N_14834,N_14903);
or U15247 (N_15247,N_14630,N_14709);
nor U15248 (N_15248,N_14875,N_14565);
nor U15249 (N_15249,N_14608,N_14799);
nand U15250 (N_15250,N_14611,N_14908);
and U15251 (N_15251,N_14647,N_14653);
nand U15252 (N_15252,N_14871,N_14872);
xor U15253 (N_15253,N_14559,N_14585);
or U15254 (N_15254,N_14519,N_14949);
or U15255 (N_15255,N_14638,N_14777);
nand U15256 (N_15256,N_14688,N_14641);
and U15257 (N_15257,N_14779,N_14836);
nand U15258 (N_15258,N_14834,N_14805);
and U15259 (N_15259,N_14930,N_14965);
or U15260 (N_15260,N_14738,N_14504);
and U15261 (N_15261,N_14579,N_14927);
nor U15262 (N_15262,N_14772,N_14920);
or U15263 (N_15263,N_14793,N_14873);
nor U15264 (N_15264,N_14778,N_14555);
or U15265 (N_15265,N_14654,N_14730);
xor U15266 (N_15266,N_14596,N_14997);
or U15267 (N_15267,N_14983,N_14714);
nand U15268 (N_15268,N_14539,N_14992);
nor U15269 (N_15269,N_14687,N_14917);
xor U15270 (N_15270,N_14585,N_14792);
and U15271 (N_15271,N_14559,N_14766);
or U15272 (N_15272,N_14746,N_14892);
and U15273 (N_15273,N_14959,N_14755);
xnor U15274 (N_15274,N_14546,N_14788);
nor U15275 (N_15275,N_14958,N_14615);
and U15276 (N_15276,N_14555,N_14681);
and U15277 (N_15277,N_14649,N_14831);
or U15278 (N_15278,N_14741,N_14621);
or U15279 (N_15279,N_14555,N_14612);
nor U15280 (N_15280,N_14522,N_14694);
or U15281 (N_15281,N_14805,N_14810);
nor U15282 (N_15282,N_14969,N_14577);
nor U15283 (N_15283,N_14565,N_14891);
nor U15284 (N_15284,N_14818,N_14865);
xnor U15285 (N_15285,N_14577,N_14668);
xor U15286 (N_15286,N_14650,N_14704);
or U15287 (N_15287,N_14774,N_14682);
nor U15288 (N_15288,N_14781,N_14961);
or U15289 (N_15289,N_14974,N_14546);
nand U15290 (N_15290,N_14589,N_14971);
nor U15291 (N_15291,N_14825,N_14927);
xnor U15292 (N_15292,N_14674,N_14956);
or U15293 (N_15293,N_14968,N_14994);
or U15294 (N_15294,N_14749,N_14513);
xor U15295 (N_15295,N_14991,N_14510);
or U15296 (N_15296,N_14540,N_14988);
xor U15297 (N_15297,N_14828,N_14696);
nor U15298 (N_15298,N_14699,N_14860);
nor U15299 (N_15299,N_14576,N_14996);
and U15300 (N_15300,N_14770,N_14534);
and U15301 (N_15301,N_14554,N_14846);
xnor U15302 (N_15302,N_14973,N_14679);
xnor U15303 (N_15303,N_14679,N_14726);
or U15304 (N_15304,N_14777,N_14509);
nor U15305 (N_15305,N_14533,N_14895);
nand U15306 (N_15306,N_14598,N_14993);
xor U15307 (N_15307,N_14678,N_14838);
nor U15308 (N_15308,N_14803,N_14779);
xor U15309 (N_15309,N_14645,N_14700);
or U15310 (N_15310,N_14602,N_14876);
nor U15311 (N_15311,N_14979,N_14682);
nand U15312 (N_15312,N_14595,N_14636);
nor U15313 (N_15313,N_14527,N_14912);
nor U15314 (N_15314,N_14547,N_14647);
nand U15315 (N_15315,N_14855,N_14845);
nand U15316 (N_15316,N_14987,N_14894);
or U15317 (N_15317,N_14963,N_14796);
nor U15318 (N_15318,N_14609,N_14747);
and U15319 (N_15319,N_14756,N_14688);
xor U15320 (N_15320,N_14908,N_14632);
and U15321 (N_15321,N_14548,N_14945);
xnor U15322 (N_15322,N_14726,N_14627);
nand U15323 (N_15323,N_14859,N_14708);
nor U15324 (N_15324,N_14773,N_14575);
or U15325 (N_15325,N_14897,N_14874);
nand U15326 (N_15326,N_14879,N_14542);
or U15327 (N_15327,N_14500,N_14771);
and U15328 (N_15328,N_14942,N_14698);
xor U15329 (N_15329,N_14816,N_14949);
xor U15330 (N_15330,N_14829,N_14722);
or U15331 (N_15331,N_14972,N_14783);
nor U15332 (N_15332,N_14666,N_14838);
and U15333 (N_15333,N_14814,N_14684);
or U15334 (N_15334,N_14789,N_14987);
or U15335 (N_15335,N_14767,N_14869);
nand U15336 (N_15336,N_14727,N_14701);
or U15337 (N_15337,N_14607,N_14740);
nand U15338 (N_15338,N_14697,N_14772);
xor U15339 (N_15339,N_14785,N_14652);
and U15340 (N_15340,N_14883,N_14808);
or U15341 (N_15341,N_14667,N_14930);
nand U15342 (N_15342,N_14702,N_14700);
or U15343 (N_15343,N_14636,N_14535);
or U15344 (N_15344,N_14852,N_14602);
and U15345 (N_15345,N_14519,N_14927);
nor U15346 (N_15346,N_14561,N_14554);
nand U15347 (N_15347,N_14810,N_14709);
nand U15348 (N_15348,N_14655,N_14552);
nor U15349 (N_15349,N_14675,N_14895);
xor U15350 (N_15350,N_14628,N_14894);
and U15351 (N_15351,N_14930,N_14627);
or U15352 (N_15352,N_14850,N_14779);
or U15353 (N_15353,N_14710,N_14665);
nor U15354 (N_15354,N_14867,N_14656);
xnor U15355 (N_15355,N_14701,N_14910);
or U15356 (N_15356,N_14740,N_14757);
nand U15357 (N_15357,N_14921,N_14578);
and U15358 (N_15358,N_14945,N_14869);
nand U15359 (N_15359,N_14963,N_14508);
or U15360 (N_15360,N_14653,N_14905);
and U15361 (N_15361,N_14828,N_14603);
nand U15362 (N_15362,N_14659,N_14962);
xor U15363 (N_15363,N_14616,N_14973);
xnor U15364 (N_15364,N_14768,N_14716);
or U15365 (N_15365,N_14582,N_14983);
nand U15366 (N_15366,N_14893,N_14769);
or U15367 (N_15367,N_14614,N_14712);
and U15368 (N_15368,N_14943,N_14977);
or U15369 (N_15369,N_14988,N_14900);
or U15370 (N_15370,N_14627,N_14547);
or U15371 (N_15371,N_14889,N_14701);
or U15372 (N_15372,N_14701,N_14781);
xnor U15373 (N_15373,N_14780,N_14998);
nand U15374 (N_15374,N_14536,N_14709);
xnor U15375 (N_15375,N_14529,N_14790);
or U15376 (N_15376,N_14892,N_14785);
nor U15377 (N_15377,N_14727,N_14606);
nand U15378 (N_15378,N_14960,N_14713);
xor U15379 (N_15379,N_14861,N_14630);
and U15380 (N_15380,N_14942,N_14655);
nor U15381 (N_15381,N_14514,N_14737);
nand U15382 (N_15382,N_14823,N_14846);
or U15383 (N_15383,N_14863,N_14639);
nor U15384 (N_15384,N_14893,N_14792);
or U15385 (N_15385,N_14654,N_14638);
and U15386 (N_15386,N_14944,N_14528);
or U15387 (N_15387,N_14637,N_14566);
nor U15388 (N_15388,N_14906,N_14823);
and U15389 (N_15389,N_14670,N_14792);
or U15390 (N_15390,N_14936,N_14839);
nand U15391 (N_15391,N_14943,N_14742);
and U15392 (N_15392,N_14720,N_14827);
and U15393 (N_15393,N_14897,N_14671);
or U15394 (N_15394,N_14983,N_14708);
and U15395 (N_15395,N_14775,N_14980);
or U15396 (N_15396,N_14655,N_14866);
nor U15397 (N_15397,N_14791,N_14833);
or U15398 (N_15398,N_14970,N_14733);
xor U15399 (N_15399,N_14717,N_14550);
nor U15400 (N_15400,N_14904,N_14950);
nand U15401 (N_15401,N_14548,N_14905);
nand U15402 (N_15402,N_14843,N_14681);
nor U15403 (N_15403,N_14601,N_14916);
and U15404 (N_15404,N_14745,N_14612);
or U15405 (N_15405,N_14651,N_14839);
nand U15406 (N_15406,N_14804,N_14836);
nand U15407 (N_15407,N_14980,N_14655);
nand U15408 (N_15408,N_14929,N_14985);
nand U15409 (N_15409,N_14667,N_14697);
nand U15410 (N_15410,N_14532,N_14576);
nor U15411 (N_15411,N_14625,N_14868);
or U15412 (N_15412,N_14798,N_14846);
and U15413 (N_15413,N_14703,N_14661);
or U15414 (N_15414,N_14647,N_14669);
nand U15415 (N_15415,N_14527,N_14898);
or U15416 (N_15416,N_14984,N_14687);
xnor U15417 (N_15417,N_14638,N_14954);
and U15418 (N_15418,N_14611,N_14982);
xor U15419 (N_15419,N_14862,N_14903);
and U15420 (N_15420,N_14728,N_14698);
nand U15421 (N_15421,N_14586,N_14547);
xor U15422 (N_15422,N_14646,N_14898);
or U15423 (N_15423,N_14997,N_14996);
or U15424 (N_15424,N_14867,N_14942);
or U15425 (N_15425,N_14742,N_14759);
nor U15426 (N_15426,N_14890,N_14967);
and U15427 (N_15427,N_14736,N_14554);
nand U15428 (N_15428,N_14593,N_14545);
xnor U15429 (N_15429,N_14827,N_14627);
or U15430 (N_15430,N_14736,N_14763);
or U15431 (N_15431,N_14685,N_14596);
nand U15432 (N_15432,N_14858,N_14691);
nor U15433 (N_15433,N_14861,N_14770);
xnor U15434 (N_15434,N_14839,N_14899);
and U15435 (N_15435,N_14943,N_14715);
or U15436 (N_15436,N_14812,N_14632);
xor U15437 (N_15437,N_14598,N_14533);
or U15438 (N_15438,N_14797,N_14886);
nor U15439 (N_15439,N_14804,N_14898);
nand U15440 (N_15440,N_14956,N_14575);
or U15441 (N_15441,N_14816,N_14558);
and U15442 (N_15442,N_14791,N_14610);
nand U15443 (N_15443,N_14991,N_14997);
nand U15444 (N_15444,N_14593,N_14737);
and U15445 (N_15445,N_14500,N_14795);
or U15446 (N_15446,N_14982,N_14547);
or U15447 (N_15447,N_14967,N_14574);
xor U15448 (N_15448,N_14571,N_14797);
nor U15449 (N_15449,N_14856,N_14790);
and U15450 (N_15450,N_14858,N_14913);
nand U15451 (N_15451,N_14993,N_14763);
xor U15452 (N_15452,N_14833,N_14859);
nand U15453 (N_15453,N_14735,N_14926);
and U15454 (N_15454,N_14719,N_14780);
and U15455 (N_15455,N_14788,N_14654);
nand U15456 (N_15456,N_14724,N_14520);
nand U15457 (N_15457,N_14877,N_14508);
xnor U15458 (N_15458,N_14512,N_14770);
xnor U15459 (N_15459,N_14681,N_14805);
nand U15460 (N_15460,N_14510,N_14501);
xor U15461 (N_15461,N_14602,N_14806);
or U15462 (N_15462,N_14948,N_14996);
nand U15463 (N_15463,N_14794,N_14981);
xnor U15464 (N_15464,N_14790,N_14660);
nor U15465 (N_15465,N_14781,N_14733);
and U15466 (N_15466,N_14612,N_14906);
xnor U15467 (N_15467,N_14661,N_14584);
or U15468 (N_15468,N_14725,N_14628);
nor U15469 (N_15469,N_14807,N_14906);
xor U15470 (N_15470,N_14683,N_14810);
nor U15471 (N_15471,N_14882,N_14765);
nand U15472 (N_15472,N_14855,N_14959);
nand U15473 (N_15473,N_14870,N_14513);
or U15474 (N_15474,N_14801,N_14799);
nand U15475 (N_15475,N_14804,N_14687);
nor U15476 (N_15476,N_14746,N_14719);
and U15477 (N_15477,N_14932,N_14834);
nand U15478 (N_15478,N_14890,N_14992);
and U15479 (N_15479,N_14985,N_14760);
nand U15480 (N_15480,N_14967,N_14640);
xor U15481 (N_15481,N_14672,N_14788);
and U15482 (N_15482,N_14911,N_14891);
xor U15483 (N_15483,N_14686,N_14954);
nand U15484 (N_15484,N_14853,N_14722);
or U15485 (N_15485,N_14895,N_14758);
nand U15486 (N_15486,N_14568,N_14961);
xor U15487 (N_15487,N_14943,N_14914);
nand U15488 (N_15488,N_14942,N_14713);
nand U15489 (N_15489,N_14588,N_14517);
xnor U15490 (N_15490,N_14978,N_14720);
or U15491 (N_15491,N_14523,N_14729);
nor U15492 (N_15492,N_14646,N_14937);
or U15493 (N_15493,N_14937,N_14844);
nand U15494 (N_15494,N_14670,N_14982);
and U15495 (N_15495,N_14800,N_14759);
nor U15496 (N_15496,N_14699,N_14621);
xnor U15497 (N_15497,N_14856,N_14680);
and U15498 (N_15498,N_14743,N_14573);
or U15499 (N_15499,N_14832,N_14855);
or U15500 (N_15500,N_15130,N_15424);
nand U15501 (N_15501,N_15292,N_15320);
nand U15502 (N_15502,N_15276,N_15112);
xor U15503 (N_15503,N_15416,N_15012);
or U15504 (N_15504,N_15370,N_15286);
xnor U15505 (N_15505,N_15306,N_15022);
or U15506 (N_15506,N_15060,N_15102);
or U15507 (N_15507,N_15021,N_15158);
xor U15508 (N_15508,N_15036,N_15188);
xnor U15509 (N_15509,N_15434,N_15323);
xnor U15510 (N_15510,N_15109,N_15342);
xnor U15511 (N_15511,N_15468,N_15146);
or U15512 (N_15512,N_15097,N_15033);
and U15513 (N_15513,N_15088,N_15346);
nor U15514 (N_15514,N_15423,N_15023);
nor U15515 (N_15515,N_15390,N_15402);
and U15516 (N_15516,N_15181,N_15343);
or U15517 (N_15517,N_15160,N_15428);
nor U15518 (N_15518,N_15357,N_15392);
and U15519 (N_15519,N_15307,N_15330);
or U15520 (N_15520,N_15144,N_15284);
xor U15521 (N_15521,N_15381,N_15134);
nor U15522 (N_15522,N_15004,N_15103);
or U15523 (N_15523,N_15426,N_15249);
or U15524 (N_15524,N_15304,N_15059);
or U15525 (N_15525,N_15162,N_15173);
nor U15526 (N_15526,N_15192,N_15274);
xor U15527 (N_15527,N_15216,N_15484);
and U15528 (N_15528,N_15049,N_15353);
and U15529 (N_15529,N_15115,N_15187);
nor U15530 (N_15530,N_15007,N_15106);
or U15531 (N_15531,N_15120,N_15350);
nor U15532 (N_15532,N_15020,N_15494);
and U15533 (N_15533,N_15364,N_15064);
or U15534 (N_15534,N_15324,N_15356);
nand U15535 (N_15535,N_15482,N_15457);
and U15536 (N_15536,N_15190,N_15301);
and U15537 (N_15537,N_15326,N_15451);
nor U15538 (N_15538,N_15002,N_15231);
and U15539 (N_15539,N_15200,N_15001);
nand U15540 (N_15540,N_15465,N_15375);
and U15541 (N_15541,N_15252,N_15498);
xor U15542 (N_15542,N_15495,N_15168);
nand U15543 (N_15543,N_15308,N_15491);
xor U15544 (N_15544,N_15054,N_15362);
or U15545 (N_15545,N_15037,N_15430);
and U15546 (N_15546,N_15179,N_15417);
xor U15547 (N_15547,N_15221,N_15340);
nor U15548 (N_15548,N_15358,N_15116);
nor U15549 (N_15549,N_15113,N_15199);
or U15550 (N_15550,N_15311,N_15366);
nor U15551 (N_15551,N_15272,N_15337);
or U15552 (N_15552,N_15039,N_15185);
or U15553 (N_15553,N_15486,N_15177);
and U15554 (N_15554,N_15458,N_15204);
or U15555 (N_15555,N_15136,N_15352);
and U15556 (N_15556,N_15461,N_15123);
and U15557 (N_15557,N_15280,N_15262);
xor U15558 (N_15558,N_15497,N_15046);
and U15559 (N_15559,N_15018,N_15069);
or U15560 (N_15560,N_15260,N_15379);
nand U15561 (N_15561,N_15309,N_15041);
xnor U15562 (N_15562,N_15319,N_15124);
xnor U15563 (N_15563,N_15202,N_15266);
nor U15564 (N_15564,N_15030,N_15407);
and U15565 (N_15565,N_15325,N_15025);
and U15566 (N_15566,N_15251,N_15044);
nor U15567 (N_15567,N_15338,N_15183);
nand U15568 (N_15568,N_15403,N_15386);
or U15569 (N_15569,N_15446,N_15072);
or U15570 (N_15570,N_15290,N_15108);
nor U15571 (N_15571,N_15282,N_15387);
xor U15572 (N_15572,N_15076,N_15091);
nand U15573 (N_15573,N_15253,N_15332);
xnor U15574 (N_15574,N_15475,N_15126);
nand U15575 (N_15575,N_15299,N_15289);
nand U15576 (N_15576,N_15125,N_15087);
nand U15577 (N_15577,N_15198,N_15207);
or U15578 (N_15578,N_15077,N_15015);
nand U15579 (N_15579,N_15333,N_15441);
nor U15580 (N_15580,N_15217,N_15034);
or U15581 (N_15581,N_15003,N_15454);
xor U15582 (N_15582,N_15053,N_15111);
or U15583 (N_15583,N_15361,N_15396);
or U15584 (N_15584,N_15226,N_15328);
xor U15585 (N_15585,N_15354,N_15388);
or U15586 (N_15586,N_15070,N_15157);
xnor U15587 (N_15587,N_15310,N_15418);
or U15588 (N_15588,N_15377,N_15421);
nor U15589 (N_15589,N_15476,N_15344);
and U15590 (N_15590,N_15410,N_15211);
or U15591 (N_15591,N_15232,N_15149);
xnor U15592 (N_15592,N_15271,N_15100);
or U15593 (N_15593,N_15071,N_15479);
nor U15594 (N_15594,N_15477,N_15161);
xor U15595 (N_15595,N_15398,N_15051);
and U15596 (N_15596,N_15341,N_15006);
nand U15597 (N_15597,N_15425,N_15128);
nand U15598 (N_15598,N_15055,N_15209);
or U15599 (N_15599,N_15101,N_15027);
xor U15600 (N_15600,N_15096,N_15219);
xor U15601 (N_15601,N_15118,N_15114);
xor U15602 (N_15602,N_15212,N_15224);
nand U15603 (N_15603,N_15011,N_15061);
and U15604 (N_15604,N_15026,N_15277);
nand U15605 (N_15605,N_15449,N_15078);
nor U15606 (N_15606,N_15184,N_15073);
nand U15607 (N_15607,N_15234,N_15327);
nor U15608 (N_15608,N_15110,N_15315);
and U15609 (N_15609,N_15401,N_15245);
xor U15610 (N_15610,N_15294,N_15107);
nor U15611 (N_15611,N_15139,N_15239);
xnor U15612 (N_15612,N_15483,N_15229);
nor U15613 (N_15613,N_15029,N_15269);
nand U15614 (N_15614,N_15360,N_15452);
and U15615 (N_15615,N_15005,N_15348);
xor U15616 (N_15616,N_15191,N_15223);
xor U15617 (N_15617,N_15296,N_15135);
xnor U15618 (N_15618,N_15246,N_15099);
and U15619 (N_15619,N_15121,N_15043);
or U15620 (N_15620,N_15368,N_15405);
or U15621 (N_15621,N_15305,N_15156);
or U15622 (N_15622,N_15176,N_15470);
xor U15623 (N_15623,N_15165,N_15167);
nor U15624 (N_15624,N_15056,N_15445);
xnor U15625 (N_15625,N_15389,N_15197);
xor U15626 (N_15626,N_15238,N_15195);
xnor U15627 (N_15627,N_15429,N_15303);
nand U15628 (N_15628,N_15263,N_15242);
or U15629 (N_15629,N_15066,N_15329);
nor U15630 (N_15630,N_15488,N_15086);
or U15631 (N_15631,N_15464,N_15119);
nor U15632 (N_15632,N_15275,N_15467);
nand U15633 (N_15633,N_15435,N_15104);
nand U15634 (N_15634,N_15152,N_15383);
or U15635 (N_15635,N_15351,N_15267);
nand U15636 (N_15636,N_15017,N_15492);
nand U15637 (N_15637,N_15058,N_15084);
nor U15638 (N_15638,N_15098,N_15016);
nand U15639 (N_15639,N_15178,N_15230);
nand U15640 (N_15640,N_15057,N_15240);
nand U15641 (N_15641,N_15474,N_15092);
nand U15642 (N_15642,N_15228,N_15137);
nand U15643 (N_15643,N_15283,N_15172);
or U15644 (N_15644,N_15414,N_15322);
or U15645 (N_15645,N_15335,N_15359);
and U15646 (N_15646,N_15153,N_15369);
xnor U15647 (N_15647,N_15075,N_15175);
nand U15648 (N_15648,N_15438,N_15481);
nor U15649 (N_15649,N_15024,N_15145);
xor U15650 (N_15650,N_15433,N_15317);
nand U15651 (N_15651,N_15105,N_15141);
nor U15652 (N_15652,N_15093,N_15159);
nand U15653 (N_15653,N_15117,N_15273);
nor U15654 (N_15654,N_15081,N_15248);
or U15655 (N_15655,N_15288,N_15493);
nand U15656 (N_15656,N_15496,N_15347);
and U15657 (N_15657,N_15122,N_15456);
and U15658 (N_15658,N_15000,N_15450);
nor U15659 (N_15659,N_15473,N_15278);
xnor U15660 (N_15660,N_15063,N_15244);
or U15661 (N_15661,N_15259,N_15371);
or U15662 (N_15662,N_15432,N_15062);
and U15663 (N_15663,N_15411,N_15180);
nand U15664 (N_15664,N_15400,N_15265);
xnor U15665 (N_15665,N_15469,N_15455);
and U15666 (N_15666,N_15170,N_15067);
or U15667 (N_15667,N_15095,N_15336);
and U15668 (N_15668,N_15166,N_15163);
xnor U15669 (N_15669,N_15205,N_15487);
nand U15670 (N_15670,N_15302,N_15052);
or U15671 (N_15671,N_15279,N_15236);
or U15672 (N_15672,N_15079,N_15408);
or U15673 (N_15673,N_15264,N_15300);
nor U15674 (N_15674,N_15250,N_15437);
nand U15675 (N_15675,N_15089,N_15142);
nor U15676 (N_15676,N_15147,N_15349);
xor U15677 (N_15677,N_15148,N_15384);
and U15678 (N_15678,N_15345,N_15222);
nand U15679 (N_15679,N_15009,N_15313);
and U15680 (N_15680,N_15422,N_15440);
and U15681 (N_15681,N_15443,N_15237);
nand U15682 (N_15682,N_15065,N_15132);
nor U15683 (N_15683,N_15466,N_15164);
nand U15684 (N_15684,N_15406,N_15255);
xnor U15685 (N_15685,N_15420,N_15032);
and U15686 (N_15686,N_15127,N_15131);
or U15687 (N_15687,N_15129,N_15367);
xor U15688 (N_15688,N_15047,N_15213);
or U15689 (N_15689,N_15042,N_15462);
nand U15690 (N_15690,N_15080,N_15436);
and U15691 (N_15691,N_15485,N_15448);
and U15692 (N_15692,N_15243,N_15028);
and U15693 (N_15693,N_15241,N_15459);
nand U15694 (N_15694,N_15404,N_15365);
nand U15695 (N_15695,N_15094,N_15155);
nand U15696 (N_15696,N_15298,N_15254);
xnor U15697 (N_15697,N_15385,N_15394);
nor U15698 (N_15698,N_15220,N_15439);
xor U15699 (N_15699,N_15151,N_15334);
nor U15700 (N_15700,N_15233,N_15373);
nor U15701 (N_15701,N_15419,N_15363);
xnor U15702 (N_15702,N_15499,N_15268);
or U15703 (N_15703,N_15035,N_15186);
and U15704 (N_15704,N_15196,N_15409);
or U15705 (N_15705,N_15208,N_15090);
nand U15706 (N_15706,N_15182,N_15447);
xor U15707 (N_15707,N_15321,N_15395);
or U15708 (N_15708,N_15193,N_15463);
nand U15709 (N_15709,N_15478,N_15019);
nor U15710 (N_15710,N_15083,N_15214);
nor U15711 (N_15711,N_15285,N_15235);
or U15712 (N_15712,N_15203,N_15314);
or U15713 (N_15713,N_15374,N_15189);
or U15714 (N_15714,N_15480,N_15206);
nor U15715 (N_15715,N_15143,N_15415);
and U15716 (N_15716,N_15171,N_15225);
and U15717 (N_15717,N_15201,N_15442);
nor U15718 (N_15718,N_15331,N_15460);
or U15719 (N_15719,N_15397,N_15378);
or U15720 (N_15720,N_15045,N_15297);
nand U15721 (N_15721,N_15391,N_15074);
and U15722 (N_15722,N_15372,N_15194);
or U15723 (N_15723,N_15287,N_15247);
or U15724 (N_15724,N_15169,N_15472);
or U15725 (N_15725,N_15210,N_15444);
nor U15726 (N_15726,N_15393,N_15085);
and U15727 (N_15727,N_15316,N_15010);
and U15728 (N_15728,N_15355,N_15014);
nand U15729 (N_15729,N_15453,N_15312);
and U15730 (N_15730,N_15227,N_15293);
nand U15731 (N_15731,N_15382,N_15008);
nor U15732 (N_15732,N_15174,N_15218);
or U15733 (N_15733,N_15261,N_15013);
and U15734 (N_15734,N_15281,N_15427);
and U15735 (N_15735,N_15270,N_15138);
xnor U15736 (N_15736,N_15031,N_15471);
nor U15737 (N_15737,N_15215,N_15490);
or U15738 (N_15738,N_15339,N_15154);
and U15739 (N_15739,N_15489,N_15150);
and U15740 (N_15740,N_15050,N_15258);
nand U15741 (N_15741,N_15040,N_15295);
xor U15742 (N_15742,N_15399,N_15133);
nor U15743 (N_15743,N_15413,N_15380);
xor U15744 (N_15744,N_15318,N_15431);
and U15745 (N_15745,N_15376,N_15140);
or U15746 (N_15746,N_15412,N_15068);
xnor U15747 (N_15747,N_15038,N_15291);
nor U15748 (N_15748,N_15256,N_15082);
nand U15749 (N_15749,N_15257,N_15048);
xnor U15750 (N_15750,N_15033,N_15022);
and U15751 (N_15751,N_15322,N_15160);
and U15752 (N_15752,N_15290,N_15105);
or U15753 (N_15753,N_15192,N_15366);
xor U15754 (N_15754,N_15396,N_15123);
or U15755 (N_15755,N_15360,N_15161);
and U15756 (N_15756,N_15183,N_15002);
nor U15757 (N_15757,N_15278,N_15443);
and U15758 (N_15758,N_15416,N_15210);
nand U15759 (N_15759,N_15015,N_15433);
or U15760 (N_15760,N_15068,N_15299);
and U15761 (N_15761,N_15368,N_15138);
and U15762 (N_15762,N_15448,N_15307);
xor U15763 (N_15763,N_15098,N_15126);
or U15764 (N_15764,N_15223,N_15071);
and U15765 (N_15765,N_15497,N_15317);
nand U15766 (N_15766,N_15114,N_15098);
and U15767 (N_15767,N_15120,N_15344);
or U15768 (N_15768,N_15221,N_15344);
nand U15769 (N_15769,N_15045,N_15277);
and U15770 (N_15770,N_15243,N_15306);
and U15771 (N_15771,N_15382,N_15453);
and U15772 (N_15772,N_15021,N_15356);
xor U15773 (N_15773,N_15496,N_15112);
and U15774 (N_15774,N_15452,N_15051);
nand U15775 (N_15775,N_15491,N_15257);
and U15776 (N_15776,N_15285,N_15392);
and U15777 (N_15777,N_15314,N_15212);
or U15778 (N_15778,N_15104,N_15310);
or U15779 (N_15779,N_15125,N_15048);
xnor U15780 (N_15780,N_15352,N_15082);
or U15781 (N_15781,N_15241,N_15389);
nand U15782 (N_15782,N_15354,N_15233);
nor U15783 (N_15783,N_15134,N_15435);
and U15784 (N_15784,N_15374,N_15405);
nor U15785 (N_15785,N_15248,N_15241);
xnor U15786 (N_15786,N_15305,N_15060);
and U15787 (N_15787,N_15298,N_15325);
and U15788 (N_15788,N_15499,N_15029);
nor U15789 (N_15789,N_15233,N_15036);
nor U15790 (N_15790,N_15196,N_15352);
nor U15791 (N_15791,N_15367,N_15151);
and U15792 (N_15792,N_15069,N_15474);
nand U15793 (N_15793,N_15401,N_15396);
xor U15794 (N_15794,N_15217,N_15015);
xnor U15795 (N_15795,N_15250,N_15092);
xnor U15796 (N_15796,N_15086,N_15354);
and U15797 (N_15797,N_15052,N_15309);
nand U15798 (N_15798,N_15252,N_15096);
or U15799 (N_15799,N_15478,N_15091);
and U15800 (N_15800,N_15139,N_15101);
nor U15801 (N_15801,N_15085,N_15301);
nand U15802 (N_15802,N_15431,N_15294);
nand U15803 (N_15803,N_15157,N_15334);
and U15804 (N_15804,N_15182,N_15243);
and U15805 (N_15805,N_15097,N_15493);
xnor U15806 (N_15806,N_15170,N_15075);
nor U15807 (N_15807,N_15229,N_15398);
and U15808 (N_15808,N_15036,N_15062);
or U15809 (N_15809,N_15190,N_15423);
xor U15810 (N_15810,N_15499,N_15043);
nand U15811 (N_15811,N_15442,N_15325);
nand U15812 (N_15812,N_15422,N_15184);
or U15813 (N_15813,N_15356,N_15499);
or U15814 (N_15814,N_15318,N_15329);
nor U15815 (N_15815,N_15095,N_15142);
or U15816 (N_15816,N_15220,N_15139);
or U15817 (N_15817,N_15451,N_15178);
xor U15818 (N_15818,N_15424,N_15417);
xor U15819 (N_15819,N_15294,N_15083);
and U15820 (N_15820,N_15359,N_15138);
xnor U15821 (N_15821,N_15166,N_15175);
xor U15822 (N_15822,N_15495,N_15100);
nor U15823 (N_15823,N_15091,N_15203);
xor U15824 (N_15824,N_15060,N_15062);
or U15825 (N_15825,N_15081,N_15445);
nor U15826 (N_15826,N_15184,N_15249);
nor U15827 (N_15827,N_15153,N_15193);
nand U15828 (N_15828,N_15151,N_15383);
and U15829 (N_15829,N_15488,N_15402);
xor U15830 (N_15830,N_15318,N_15326);
nor U15831 (N_15831,N_15291,N_15476);
or U15832 (N_15832,N_15283,N_15350);
nor U15833 (N_15833,N_15361,N_15353);
or U15834 (N_15834,N_15440,N_15465);
or U15835 (N_15835,N_15179,N_15260);
xor U15836 (N_15836,N_15259,N_15325);
nand U15837 (N_15837,N_15092,N_15395);
xor U15838 (N_15838,N_15036,N_15250);
nor U15839 (N_15839,N_15318,N_15188);
nand U15840 (N_15840,N_15161,N_15499);
nor U15841 (N_15841,N_15050,N_15107);
or U15842 (N_15842,N_15148,N_15301);
nor U15843 (N_15843,N_15013,N_15050);
xnor U15844 (N_15844,N_15326,N_15202);
nand U15845 (N_15845,N_15257,N_15438);
nor U15846 (N_15846,N_15444,N_15142);
nor U15847 (N_15847,N_15088,N_15151);
or U15848 (N_15848,N_15351,N_15019);
and U15849 (N_15849,N_15420,N_15449);
or U15850 (N_15850,N_15080,N_15173);
xnor U15851 (N_15851,N_15012,N_15068);
and U15852 (N_15852,N_15013,N_15127);
nand U15853 (N_15853,N_15263,N_15338);
and U15854 (N_15854,N_15455,N_15418);
nor U15855 (N_15855,N_15466,N_15187);
nor U15856 (N_15856,N_15454,N_15483);
xor U15857 (N_15857,N_15233,N_15186);
and U15858 (N_15858,N_15217,N_15412);
and U15859 (N_15859,N_15018,N_15453);
or U15860 (N_15860,N_15311,N_15449);
nand U15861 (N_15861,N_15151,N_15023);
and U15862 (N_15862,N_15067,N_15043);
and U15863 (N_15863,N_15287,N_15074);
xnor U15864 (N_15864,N_15005,N_15116);
and U15865 (N_15865,N_15413,N_15374);
nand U15866 (N_15866,N_15046,N_15456);
nor U15867 (N_15867,N_15455,N_15012);
nor U15868 (N_15868,N_15055,N_15486);
or U15869 (N_15869,N_15430,N_15198);
nand U15870 (N_15870,N_15206,N_15299);
nor U15871 (N_15871,N_15265,N_15416);
xnor U15872 (N_15872,N_15276,N_15243);
nand U15873 (N_15873,N_15350,N_15007);
xnor U15874 (N_15874,N_15344,N_15152);
xor U15875 (N_15875,N_15386,N_15245);
or U15876 (N_15876,N_15458,N_15026);
or U15877 (N_15877,N_15052,N_15313);
nand U15878 (N_15878,N_15012,N_15073);
xnor U15879 (N_15879,N_15158,N_15319);
xor U15880 (N_15880,N_15253,N_15145);
or U15881 (N_15881,N_15199,N_15235);
nor U15882 (N_15882,N_15176,N_15003);
and U15883 (N_15883,N_15245,N_15286);
xnor U15884 (N_15884,N_15122,N_15347);
nor U15885 (N_15885,N_15237,N_15283);
nand U15886 (N_15886,N_15429,N_15033);
or U15887 (N_15887,N_15046,N_15005);
nor U15888 (N_15888,N_15393,N_15081);
nor U15889 (N_15889,N_15286,N_15405);
xnor U15890 (N_15890,N_15198,N_15439);
nor U15891 (N_15891,N_15081,N_15185);
nand U15892 (N_15892,N_15027,N_15166);
or U15893 (N_15893,N_15188,N_15203);
or U15894 (N_15894,N_15151,N_15045);
nand U15895 (N_15895,N_15167,N_15308);
and U15896 (N_15896,N_15419,N_15160);
and U15897 (N_15897,N_15402,N_15406);
nand U15898 (N_15898,N_15241,N_15072);
nand U15899 (N_15899,N_15324,N_15389);
nor U15900 (N_15900,N_15402,N_15487);
nor U15901 (N_15901,N_15250,N_15055);
nor U15902 (N_15902,N_15303,N_15461);
nor U15903 (N_15903,N_15336,N_15335);
xnor U15904 (N_15904,N_15494,N_15212);
or U15905 (N_15905,N_15111,N_15181);
and U15906 (N_15906,N_15304,N_15495);
xor U15907 (N_15907,N_15025,N_15462);
nand U15908 (N_15908,N_15414,N_15206);
and U15909 (N_15909,N_15436,N_15194);
xnor U15910 (N_15910,N_15186,N_15196);
nor U15911 (N_15911,N_15368,N_15203);
nand U15912 (N_15912,N_15109,N_15200);
nand U15913 (N_15913,N_15161,N_15335);
nor U15914 (N_15914,N_15499,N_15069);
nor U15915 (N_15915,N_15421,N_15485);
and U15916 (N_15916,N_15002,N_15353);
or U15917 (N_15917,N_15265,N_15195);
nand U15918 (N_15918,N_15191,N_15128);
and U15919 (N_15919,N_15423,N_15445);
nor U15920 (N_15920,N_15386,N_15330);
nor U15921 (N_15921,N_15046,N_15219);
or U15922 (N_15922,N_15174,N_15323);
and U15923 (N_15923,N_15229,N_15211);
and U15924 (N_15924,N_15464,N_15242);
xor U15925 (N_15925,N_15139,N_15282);
xnor U15926 (N_15926,N_15429,N_15280);
nand U15927 (N_15927,N_15022,N_15352);
and U15928 (N_15928,N_15247,N_15348);
and U15929 (N_15929,N_15316,N_15458);
or U15930 (N_15930,N_15325,N_15167);
xnor U15931 (N_15931,N_15245,N_15256);
xor U15932 (N_15932,N_15256,N_15357);
or U15933 (N_15933,N_15086,N_15238);
nor U15934 (N_15934,N_15108,N_15226);
xnor U15935 (N_15935,N_15122,N_15043);
xor U15936 (N_15936,N_15067,N_15235);
and U15937 (N_15937,N_15301,N_15110);
or U15938 (N_15938,N_15309,N_15100);
and U15939 (N_15939,N_15206,N_15266);
xnor U15940 (N_15940,N_15038,N_15394);
nand U15941 (N_15941,N_15346,N_15451);
nor U15942 (N_15942,N_15282,N_15114);
xor U15943 (N_15943,N_15021,N_15029);
nand U15944 (N_15944,N_15356,N_15059);
nor U15945 (N_15945,N_15256,N_15350);
nand U15946 (N_15946,N_15467,N_15133);
nand U15947 (N_15947,N_15046,N_15165);
xor U15948 (N_15948,N_15247,N_15081);
nand U15949 (N_15949,N_15025,N_15039);
nand U15950 (N_15950,N_15174,N_15192);
nand U15951 (N_15951,N_15247,N_15359);
nand U15952 (N_15952,N_15335,N_15370);
and U15953 (N_15953,N_15149,N_15021);
nor U15954 (N_15954,N_15025,N_15215);
or U15955 (N_15955,N_15079,N_15406);
or U15956 (N_15956,N_15337,N_15404);
or U15957 (N_15957,N_15055,N_15270);
xnor U15958 (N_15958,N_15282,N_15322);
nand U15959 (N_15959,N_15145,N_15436);
nand U15960 (N_15960,N_15343,N_15037);
xnor U15961 (N_15961,N_15135,N_15060);
nand U15962 (N_15962,N_15371,N_15083);
and U15963 (N_15963,N_15498,N_15469);
or U15964 (N_15964,N_15212,N_15149);
nand U15965 (N_15965,N_15336,N_15049);
nand U15966 (N_15966,N_15117,N_15376);
nand U15967 (N_15967,N_15287,N_15012);
xnor U15968 (N_15968,N_15235,N_15382);
nand U15969 (N_15969,N_15057,N_15450);
nor U15970 (N_15970,N_15032,N_15242);
xor U15971 (N_15971,N_15461,N_15409);
and U15972 (N_15972,N_15193,N_15201);
nor U15973 (N_15973,N_15330,N_15069);
nor U15974 (N_15974,N_15427,N_15313);
nor U15975 (N_15975,N_15477,N_15358);
nor U15976 (N_15976,N_15261,N_15413);
xnor U15977 (N_15977,N_15186,N_15092);
nand U15978 (N_15978,N_15095,N_15418);
nand U15979 (N_15979,N_15187,N_15373);
and U15980 (N_15980,N_15289,N_15469);
and U15981 (N_15981,N_15060,N_15379);
nor U15982 (N_15982,N_15409,N_15167);
or U15983 (N_15983,N_15255,N_15164);
nor U15984 (N_15984,N_15493,N_15498);
nor U15985 (N_15985,N_15227,N_15145);
or U15986 (N_15986,N_15486,N_15331);
or U15987 (N_15987,N_15363,N_15301);
or U15988 (N_15988,N_15209,N_15121);
xor U15989 (N_15989,N_15257,N_15184);
nand U15990 (N_15990,N_15101,N_15458);
xor U15991 (N_15991,N_15205,N_15405);
nand U15992 (N_15992,N_15394,N_15460);
nor U15993 (N_15993,N_15047,N_15371);
nor U15994 (N_15994,N_15173,N_15042);
and U15995 (N_15995,N_15230,N_15419);
or U15996 (N_15996,N_15386,N_15014);
or U15997 (N_15997,N_15153,N_15144);
nand U15998 (N_15998,N_15272,N_15325);
or U15999 (N_15999,N_15215,N_15133);
and U16000 (N_16000,N_15597,N_15637);
or U16001 (N_16001,N_15559,N_15959);
or U16002 (N_16002,N_15754,N_15605);
nor U16003 (N_16003,N_15638,N_15592);
and U16004 (N_16004,N_15750,N_15766);
nand U16005 (N_16005,N_15629,N_15529);
xnor U16006 (N_16006,N_15916,N_15833);
and U16007 (N_16007,N_15543,N_15552);
and U16008 (N_16008,N_15712,N_15650);
xor U16009 (N_16009,N_15512,N_15777);
nor U16010 (N_16010,N_15781,N_15539);
nor U16011 (N_16011,N_15955,N_15632);
and U16012 (N_16012,N_15644,N_15794);
and U16013 (N_16013,N_15940,N_15731);
and U16014 (N_16014,N_15818,N_15627);
or U16015 (N_16015,N_15937,N_15520);
nor U16016 (N_16016,N_15949,N_15697);
nand U16017 (N_16017,N_15655,N_15802);
or U16018 (N_16018,N_15545,N_15670);
nand U16019 (N_16019,N_15922,N_15981);
and U16020 (N_16020,N_15945,N_15809);
xor U16021 (N_16021,N_15847,N_15960);
nand U16022 (N_16022,N_15679,N_15946);
nor U16023 (N_16023,N_15815,N_15792);
nor U16024 (N_16024,N_15852,N_15640);
xnor U16025 (N_16025,N_15894,N_15993);
xnor U16026 (N_16026,N_15983,N_15669);
xnor U16027 (N_16027,N_15694,N_15649);
or U16028 (N_16028,N_15865,N_15851);
xor U16029 (N_16029,N_15727,N_15749);
and U16030 (N_16030,N_15821,N_15598);
nand U16031 (N_16031,N_15584,N_15528);
and U16032 (N_16032,N_15660,N_15561);
and U16033 (N_16033,N_15630,N_15868);
xor U16034 (N_16034,N_15728,N_15775);
nand U16035 (N_16035,N_15530,N_15501);
nor U16036 (N_16036,N_15635,N_15932);
and U16037 (N_16037,N_15850,N_15500);
and U16038 (N_16038,N_15641,N_15832);
nor U16039 (N_16039,N_15891,N_15623);
nor U16040 (N_16040,N_15909,N_15579);
nand U16041 (N_16041,N_15594,N_15606);
nor U16042 (N_16042,N_15857,N_15678);
nand U16043 (N_16043,N_15789,N_15692);
and U16044 (N_16044,N_15763,N_15642);
nand U16045 (N_16045,N_15682,N_15843);
or U16046 (N_16046,N_15668,N_15665);
and U16047 (N_16047,N_15869,N_15967);
nand U16048 (N_16048,N_15717,N_15703);
xor U16049 (N_16049,N_15908,N_15854);
nor U16050 (N_16050,N_15544,N_15782);
or U16051 (N_16051,N_15830,N_15713);
xor U16052 (N_16052,N_15951,N_15824);
or U16053 (N_16053,N_15730,N_15663);
nor U16054 (N_16054,N_15760,N_15620);
nor U16055 (N_16055,N_15624,N_15872);
nand U16056 (N_16056,N_15705,N_15819);
xor U16057 (N_16057,N_15564,N_15925);
nor U16058 (N_16058,N_15643,N_15701);
nor U16059 (N_16059,N_15577,N_15688);
nand U16060 (N_16060,N_15842,N_15513);
xor U16061 (N_16061,N_15877,N_15799);
or U16062 (N_16062,N_15591,N_15783);
or U16063 (N_16063,N_15774,N_15652);
nor U16064 (N_16064,N_15785,N_15651);
or U16065 (N_16065,N_15999,N_15700);
nand U16066 (N_16066,N_15662,N_15575);
nor U16067 (N_16067,N_15826,N_15803);
and U16068 (N_16068,N_15913,N_15621);
nand U16069 (N_16069,N_15910,N_15957);
nand U16070 (N_16070,N_15812,N_15690);
and U16071 (N_16071,N_15714,N_15979);
xnor U16072 (N_16072,N_15975,N_15954);
xnor U16073 (N_16073,N_15840,N_15965);
nand U16074 (N_16074,N_15570,N_15657);
xnor U16075 (N_16075,N_15767,N_15617);
nand U16076 (N_16076,N_15733,N_15732);
nor U16077 (N_16077,N_15648,N_15875);
nand U16078 (N_16078,N_15631,N_15709);
or U16079 (N_16079,N_15654,N_15893);
and U16080 (N_16080,N_15645,N_15969);
and U16081 (N_16081,N_15685,N_15736);
nand U16082 (N_16082,N_15737,N_15885);
or U16083 (N_16083,N_15985,N_15686);
or U16084 (N_16084,N_15827,N_15795);
xnor U16085 (N_16085,N_15920,N_15542);
nand U16086 (N_16086,N_15698,N_15687);
nor U16087 (N_16087,N_15810,N_15836);
or U16088 (N_16088,N_15518,N_15771);
xnor U16089 (N_16089,N_15786,N_15888);
and U16090 (N_16090,N_15950,N_15906);
nand U16091 (N_16091,N_15556,N_15515);
nand U16092 (N_16092,N_15667,N_15917);
nor U16093 (N_16093,N_15859,N_15574);
xor U16094 (N_16094,N_15876,N_15846);
nor U16095 (N_16095,N_15525,N_15791);
nand U16096 (N_16096,N_15800,N_15510);
nor U16097 (N_16097,N_15647,N_15941);
xor U16098 (N_16098,N_15784,N_15633);
xnor U16099 (N_16099,N_15793,N_15862);
xor U16100 (N_16100,N_15693,N_15744);
and U16101 (N_16101,N_15604,N_15984);
or U16102 (N_16102,N_15961,N_15905);
nand U16103 (N_16103,N_15933,N_15820);
or U16104 (N_16104,N_15535,N_15702);
nor U16105 (N_16105,N_15808,N_15549);
xnor U16106 (N_16106,N_15557,N_15589);
or U16107 (N_16107,N_15540,N_15801);
nor U16108 (N_16108,N_15867,N_15751);
nor U16109 (N_16109,N_15676,N_15882);
or U16110 (N_16110,N_15672,N_15581);
xnor U16111 (N_16111,N_15968,N_15938);
nor U16112 (N_16112,N_15666,N_15722);
nand U16113 (N_16113,N_15926,N_15616);
or U16114 (N_16114,N_15822,N_15806);
xnor U16115 (N_16115,N_15560,N_15998);
and U16116 (N_16116,N_15580,N_15860);
nand U16117 (N_16117,N_15707,N_15919);
nand U16118 (N_16118,N_15886,N_15978);
nor U16119 (N_16119,N_15571,N_15729);
xor U16120 (N_16120,N_15986,N_15680);
xnor U16121 (N_16121,N_15989,N_15546);
nor U16122 (N_16122,N_15918,N_15689);
nor U16123 (N_16123,N_15547,N_15684);
nand U16124 (N_16124,N_15970,N_15823);
xor U16125 (N_16125,N_15898,N_15849);
or U16126 (N_16126,N_15817,N_15996);
xnor U16127 (N_16127,N_15704,N_15895);
xnor U16128 (N_16128,N_15952,N_15582);
xnor U16129 (N_16129,N_15613,N_15814);
nand U16130 (N_16130,N_15927,N_15864);
nor U16131 (N_16131,N_15677,N_15602);
or U16132 (N_16132,N_15588,N_15856);
nor U16133 (N_16133,N_15931,N_15761);
and U16134 (N_16134,N_15790,N_15639);
and U16135 (N_16135,N_15711,N_15966);
and U16136 (N_16136,N_15871,N_15673);
nand U16137 (N_16137,N_15896,N_15508);
nor U16138 (N_16138,N_15534,N_15912);
and U16139 (N_16139,N_15719,N_15994);
nand U16140 (N_16140,N_15524,N_15841);
nor U16141 (N_16141,N_15742,N_15900);
nor U16142 (N_16142,N_15930,N_15537);
and U16143 (N_16143,N_15990,N_15626);
nor U16144 (N_16144,N_15921,N_15765);
nand U16145 (N_16145,N_15747,N_15567);
xor U16146 (N_16146,N_15987,N_15887);
nor U16147 (N_16147,N_15725,N_15904);
xor U16148 (N_16148,N_15554,N_15992);
xnor U16149 (N_16149,N_15972,N_15797);
nor U16150 (N_16150,N_15958,N_15615);
xor U16151 (N_16151,N_15805,N_15929);
or U16152 (N_16152,N_15699,N_15756);
nor U16153 (N_16153,N_15691,N_15748);
and U16154 (N_16154,N_15618,N_15716);
xor U16155 (N_16155,N_15759,N_15787);
xor U16156 (N_16156,N_15504,N_15681);
nand U16157 (N_16157,N_15956,N_15531);
xor U16158 (N_16158,N_15599,N_15746);
nor U16159 (N_16159,N_15724,N_15590);
nand U16160 (N_16160,N_15770,N_15915);
or U16161 (N_16161,N_15595,N_15671);
xnor U16162 (N_16162,N_15745,N_15514);
nand U16163 (N_16163,N_15884,N_15656);
and U16164 (N_16164,N_15923,N_15548);
xor U16165 (N_16165,N_15664,N_15942);
or U16166 (N_16166,N_15991,N_15934);
xor U16167 (N_16167,N_15735,N_15828);
or U16168 (N_16168,N_15502,N_15988);
and U16169 (N_16169,N_15683,N_15511);
nand U16170 (N_16170,N_15612,N_15878);
and U16171 (N_16171,N_15708,N_15522);
nand U16172 (N_16172,N_15553,N_15939);
nor U16173 (N_16173,N_15734,N_15541);
nor U16174 (N_16174,N_15562,N_15558);
nand U16175 (N_16175,N_15715,N_15569);
and U16176 (N_16176,N_15611,N_15710);
or U16177 (N_16177,N_15899,N_15723);
and U16178 (N_16178,N_15813,N_15902);
and U16179 (N_16179,N_15924,N_15720);
nand U16180 (N_16180,N_15995,N_15769);
and U16181 (N_16181,N_15890,N_15622);
nand U16182 (N_16182,N_15536,N_15578);
or U16183 (N_16183,N_15976,N_15757);
or U16184 (N_16184,N_15675,N_15527);
xor U16185 (N_16185,N_15646,N_15576);
and U16186 (N_16186,N_15943,N_15870);
or U16187 (N_16187,N_15773,N_15634);
and U16188 (N_16188,N_15653,N_15838);
xor U16189 (N_16189,N_15658,N_15533);
or U16190 (N_16190,N_15889,N_15780);
nand U16191 (N_16191,N_15980,N_15948);
and U16192 (N_16192,N_15523,N_15892);
and U16193 (N_16193,N_15739,N_15517);
nor U16194 (N_16194,N_15831,N_15914);
xnor U16195 (N_16195,N_15901,N_15526);
nor U16196 (N_16196,N_15565,N_15811);
xnor U16197 (N_16197,N_15964,N_15897);
and U16198 (N_16198,N_15762,N_15855);
or U16199 (N_16199,N_15977,N_15962);
xnor U16200 (N_16200,N_15509,N_15609);
and U16201 (N_16201,N_15778,N_15614);
nor U16202 (N_16202,N_15997,N_15971);
or U16203 (N_16203,N_15873,N_15726);
or U16204 (N_16204,N_15573,N_15858);
nand U16205 (N_16205,N_15911,N_15953);
or U16206 (N_16206,N_15768,N_15844);
and U16207 (N_16207,N_15555,N_15519);
xor U16208 (N_16208,N_15973,N_15874);
nor U16209 (N_16209,N_15974,N_15796);
nor U16210 (N_16210,N_15752,N_15879);
nor U16211 (N_16211,N_15861,N_15798);
and U16212 (N_16212,N_15607,N_15585);
and U16213 (N_16213,N_15863,N_15521);
and U16214 (N_16214,N_15721,N_15600);
or U16215 (N_16215,N_15566,N_15807);
nor U16216 (N_16216,N_15866,N_15848);
nand U16217 (N_16217,N_15776,N_15880);
xor U16218 (N_16218,N_15881,N_15853);
and U16219 (N_16219,N_15718,N_15608);
or U16220 (N_16220,N_15772,N_15695);
nand U16221 (N_16221,N_15740,N_15839);
and U16222 (N_16222,N_15593,N_15568);
or U16223 (N_16223,N_15935,N_15659);
or U16224 (N_16224,N_15503,N_15741);
nor U16225 (N_16225,N_15758,N_15661);
nand U16226 (N_16226,N_15804,N_15596);
nor U16227 (N_16227,N_15636,N_15944);
nor U16228 (N_16228,N_15696,N_15829);
xor U16229 (N_16229,N_15538,N_15507);
xnor U16230 (N_16230,N_15816,N_15845);
nand U16231 (N_16231,N_15505,N_15837);
nor U16232 (N_16232,N_15583,N_15610);
nor U16233 (N_16233,N_15788,N_15825);
nand U16234 (N_16234,N_15563,N_15764);
nor U16235 (N_16235,N_15834,N_15936);
nor U16236 (N_16236,N_15628,N_15947);
and U16237 (N_16237,N_15551,N_15753);
xor U16238 (N_16238,N_15603,N_15779);
nand U16239 (N_16239,N_15755,N_15550);
nor U16240 (N_16240,N_15674,N_15619);
nor U16241 (N_16241,N_15706,N_15738);
xnor U16242 (N_16242,N_15963,N_15532);
and U16243 (N_16243,N_15625,N_15572);
and U16244 (N_16244,N_15743,N_15516);
nand U16245 (N_16245,N_15586,N_15835);
nand U16246 (N_16246,N_15982,N_15928);
nor U16247 (N_16247,N_15506,N_15907);
or U16248 (N_16248,N_15587,N_15903);
or U16249 (N_16249,N_15601,N_15883);
and U16250 (N_16250,N_15741,N_15806);
xor U16251 (N_16251,N_15933,N_15894);
nand U16252 (N_16252,N_15886,N_15644);
nor U16253 (N_16253,N_15854,N_15888);
or U16254 (N_16254,N_15708,N_15958);
and U16255 (N_16255,N_15739,N_15650);
and U16256 (N_16256,N_15847,N_15569);
or U16257 (N_16257,N_15662,N_15854);
xnor U16258 (N_16258,N_15843,N_15780);
and U16259 (N_16259,N_15797,N_15664);
nor U16260 (N_16260,N_15635,N_15564);
nor U16261 (N_16261,N_15628,N_15584);
nand U16262 (N_16262,N_15602,N_15848);
nand U16263 (N_16263,N_15534,N_15755);
nor U16264 (N_16264,N_15657,N_15660);
xor U16265 (N_16265,N_15838,N_15700);
nor U16266 (N_16266,N_15736,N_15676);
or U16267 (N_16267,N_15967,N_15660);
and U16268 (N_16268,N_15789,N_15877);
nand U16269 (N_16269,N_15856,N_15685);
and U16270 (N_16270,N_15763,N_15727);
xor U16271 (N_16271,N_15611,N_15502);
xnor U16272 (N_16272,N_15547,N_15638);
xnor U16273 (N_16273,N_15708,N_15562);
xnor U16274 (N_16274,N_15877,N_15719);
or U16275 (N_16275,N_15912,N_15670);
or U16276 (N_16276,N_15776,N_15509);
xnor U16277 (N_16277,N_15642,N_15858);
or U16278 (N_16278,N_15573,N_15770);
nor U16279 (N_16279,N_15611,N_15510);
nand U16280 (N_16280,N_15995,N_15722);
and U16281 (N_16281,N_15792,N_15515);
or U16282 (N_16282,N_15525,N_15607);
and U16283 (N_16283,N_15773,N_15930);
or U16284 (N_16284,N_15641,N_15629);
nand U16285 (N_16285,N_15864,N_15597);
nand U16286 (N_16286,N_15533,N_15815);
nor U16287 (N_16287,N_15731,N_15760);
xnor U16288 (N_16288,N_15908,N_15570);
or U16289 (N_16289,N_15504,N_15600);
nand U16290 (N_16290,N_15596,N_15995);
xor U16291 (N_16291,N_15851,N_15809);
xor U16292 (N_16292,N_15831,N_15507);
nand U16293 (N_16293,N_15812,N_15867);
and U16294 (N_16294,N_15535,N_15947);
and U16295 (N_16295,N_15625,N_15864);
nor U16296 (N_16296,N_15975,N_15608);
nand U16297 (N_16297,N_15503,N_15763);
nand U16298 (N_16298,N_15916,N_15927);
nor U16299 (N_16299,N_15591,N_15697);
and U16300 (N_16300,N_15597,N_15639);
or U16301 (N_16301,N_15807,N_15948);
or U16302 (N_16302,N_15696,N_15593);
xor U16303 (N_16303,N_15512,N_15868);
and U16304 (N_16304,N_15622,N_15661);
nor U16305 (N_16305,N_15942,N_15910);
nor U16306 (N_16306,N_15581,N_15732);
nor U16307 (N_16307,N_15753,N_15692);
nor U16308 (N_16308,N_15576,N_15882);
xnor U16309 (N_16309,N_15673,N_15885);
nand U16310 (N_16310,N_15754,N_15531);
nand U16311 (N_16311,N_15996,N_15820);
and U16312 (N_16312,N_15574,N_15534);
and U16313 (N_16313,N_15708,N_15748);
and U16314 (N_16314,N_15987,N_15778);
and U16315 (N_16315,N_15539,N_15537);
nand U16316 (N_16316,N_15672,N_15567);
nand U16317 (N_16317,N_15552,N_15844);
nor U16318 (N_16318,N_15980,N_15705);
xor U16319 (N_16319,N_15626,N_15659);
nor U16320 (N_16320,N_15589,N_15780);
and U16321 (N_16321,N_15823,N_15835);
and U16322 (N_16322,N_15898,N_15515);
nand U16323 (N_16323,N_15834,N_15856);
nor U16324 (N_16324,N_15826,N_15754);
xnor U16325 (N_16325,N_15800,N_15767);
or U16326 (N_16326,N_15816,N_15761);
and U16327 (N_16327,N_15992,N_15605);
xnor U16328 (N_16328,N_15935,N_15795);
nor U16329 (N_16329,N_15547,N_15812);
and U16330 (N_16330,N_15988,N_15970);
nor U16331 (N_16331,N_15861,N_15817);
nand U16332 (N_16332,N_15956,N_15789);
nand U16333 (N_16333,N_15885,N_15650);
and U16334 (N_16334,N_15943,N_15710);
xnor U16335 (N_16335,N_15817,N_15864);
xnor U16336 (N_16336,N_15752,N_15945);
nand U16337 (N_16337,N_15998,N_15733);
nor U16338 (N_16338,N_15638,N_15883);
nand U16339 (N_16339,N_15667,N_15776);
xnor U16340 (N_16340,N_15569,N_15818);
nand U16341 (N_16341,N_15640,N_15694);
xor U16342 (N_16342,N_15889,N_15716);
or U16343 (N_16343,N_15837,N_15754);
nor U16344 (N_16344,N_15649,N_15511);
nand U16345 (N_16345,N_15562,N_15771);
xnor U16346 (N_16346,N_15911,N_15619);
and U16347 (N_16347,N_15738,N_15763);
xnor U16348 (N_16348,N_15835,N_15589);
nand U16349 (N_16349,N_15505,N_15530);
nand U16350 (N_16350,N_15934,N_15658);
and U16351 (N_16351,N_15651,N_15847);
and U16352 (N_16352,N_15907,N_15693);
or U16353 (N_16353,N_15925,N_15979);
xor U16354 (N_16354,N_15836,N_15853);
nor U16355 (N_16355,N_15929,N_15755);
nand U16356 (N_16356,N_15862,N_15564);
nand U16357 (N_16357,N_15590,N_15750);
nor U16358 (N_16358,N_15744,N_15649);
xnor U16359 (N_16359,N_15590,N_15730);
and U16360 (N_16360,N_15662,N_15880);
nand U16361 (N_16361,N_15912,N_15509);
xor U16362 (N_16362,N_15773,N_15954);
or U16363 (N_16363,N_15791,N_15766);
and U16364 (N_16364,N_15957,N_15628);
nand U16365 (N_16365,N_15989,N_15966);
or U16366 (N_16366,N_15777,N_15714);
nand U16367 (N_16367,N_15725,N_15827);
or U16368 (N_16368,N_15772,N_15941);
nand U16369 (N_16369,N_15785,N_15963);
nand U16370 (N_16370,N_15627,N_15605);
or U16371 (N_16371,N_15720,N_15528);
xnor U16372 (N_16372,N_15807,N_15977);
xor U16373 (N_16373,N_15617,N_15516);
or U16374 (N_16374,N_15810,N_15625);
nor U16375 (N_16375,N_15711,N_15881);
nand U16376 (N_16376,N_15637,N_15744);
or U16377 (N_16377,N_15610,N_15661);
xnor U16378 (N_16378,N_15563,N_15534);
nor U16379 (N_16379,N_15946,N_15727);
or U16380 (N_16380,N_15775,N_15582);
and U16381 (N_16381,N_15640,N_15915);
nor U16382 (N_16382,N_15941,N_15867);
nor U16383 (N_16383,N_15791,N_15663);
nand U16384 (N_16384,N_15586,N_15883);
nor U16385 (N_16385,N_15837,N_15742);
and U16386 (N_16386,N_15767,N_15643);
nor U16387 (N_16387,N_15701,N_15602);
or U16388 (N_16388,N_15793,N_15620);
xor U16389 (N_16389,N_15542,N_15591);
nand U16390 (N_16390,N_15813,N_15807);
or U16391 (N_16391,N_15867,N_15613);
nor U16392 (N_16392,N_15987,N_15561);
or U16393 (N_16393,N_15648,N_15696);
nor U16394 (N_16394,N_15562,N_15931);
xor U16395 (N_16395,N_15555,N_15918);
or U16396 (N_16396,N_15851,N_15957);
nor U16397 (N_16397,N_15956,N_15995);
xor U16398 (N_16398,N_15518,N_15948);
nor U16399 (N_16399,N_15596,N_15926);
xor U16400 (N_16400,N_15968,N_15807);
nand U16401 (N_16401,N_15699,N_15738);
xnor U16402 (N_16402,N_15693,N_15769);
nand U16403 (N_16403,N_15789,N_15859);
and U16404 (N_16404,N_15796,N_15601);
and U16405 (N_16405,N_15613,N_15788);
or U16406 (N_16406,N_15972,N_15859);
nor U16407 (N_16407,N_15567,N_15877);
and U16408 (N_16408,N_15533,N_15941);
xnor U16409 (N_16409,N_15610,N_15733);
or U16410 (N_16410,N_15685,N_15588);
nand U16411 (N_16411,N_15601,N_15963);
nand U16412 (N_16412,N_15526,N_15565);
nor U16413 (N_16413,N_15504,N_15912);
or U16414 (N_16414,N_15710,N_15949);
nand U16415 (N_16415,N_15931,N_15977);
xnor U16416 (N_16416,N_15763,N_15606);
and U16417 (N_16417,N_15636,N_15876);
nor U16418 (N_16418,N_15717,N_15504);
xnor U16419 (N_16419,N_15845,N_15679);
and U16420 (N_16420,N_15646,N_15720);
and U16421 (N_16421,N_15764,N_15998);
xor U16422 (N_16422,N_15675,N_15821);
nor U16423 (N_16423,N_15791,N_15917);
or U16424 (N_16424,N_15974,N_15634);
nand U16425 (N_16425,N_15529,N_15783);
or U16426 (N_16426,N_15552,N_15611);
nand U16427 (N_16427,N_15976,N_15855);
and U16428 (N_16428,N_15838,N_15903);
xnor U16429 (N_16429,N_15670,N_15639);
or U16430 (N_16430,N_15626,N_15696);
xor U16431 (N_16431,N_15673,N_15870);
and U16432 (N_16432,N_15753,N_15966);
and U16433 (N_16433,N_15544,N_15676);
xor U16434 (N_16434,N_15525,N_15747);
xor U16435 (N_16435,N_15723,N_15947);
nor U16436 (N_16436,N_15842,N_15613);
nand U16437 (N_16437,N_15622,N_15550);
or U16438 (N_16438,N_15747,N_15988);
and U16439 (N_16439,N_15739,N_15778);
nand U16440 (N_16440,N_15769,N_15512);
and U16441 (N_16441,N_15824,N_15859);
nand U16442 (N_16442,N_15643,N_15980);
or U16443 (N_16443,N_15968,N_15995);
or U16444 (N_16444,N_15638,N_15822);
xor U16445 (N_16445,N_15720,N_15584);
or U16446 (N_16446,N_15778,N_15699);
or U16447 (N_16447,N_15559,N_15901);
xnor U16448 (N_16448,N_15984,N_15869);
or U16449 (N_16449,N_15624,N_15599);
nand U16450 (N_16450,N_15707,N_15603);
and U16451 (N_16451,N_15981,N_15781);
and U16452 (N_16452,N_15645,N_15600);
nor U16453 (N_16453,N_15806,N_15999);
and U16454 (N_16454,N_15515,N_15995);
and U16455 (N_16455,N_15620,N_15530);
nor U16456 (N_16456,N_15998,N_15567);
xnor U16457 (N_16457,N_15729,N_15667);
and U16458 (N_16458,N_15955,N_15579);
nor U16459 (N_16459,N_15517,N_15729);
nor U16460 (N_16460,N_15637,N_15526);
nand U16461 (N_16461,N_15767,N_15798);
or U16462 (N_16462,N_15672,N_15753);
nand U16463 (N_16463,N_15605,N_15577);
or U16464 (N_16464,N_15812,N_15843);
and U16465 (N_16465,N_15963,N_15625);
nand U16466 (N_16466,N_15630,N_15886);
nand U16467 (N_16467,N_15945,N_15773);
xnor U16468 (N_16468,N_15833,N_15677);
nor U16469 (N_16469,N_15675,N_15826);
nor U16470 (N_16470,N_15552,N_15784);
nor U16471 (N_16471,N_15969,N_15770);
or U16472 (N_16472,N_15792,N_15835);
and U16473 (N_16473,N_15594,N_15727);
xnor U16474 (N_16474,N_15961,N_15505);
and U16475 (N_16475,N_15501,N_15970);
nand U16476 (N_16476,N_15545,N_15503);
nand U16477 (N_16477,N_15922,N_15835);
xnor U16478 (N_16478,N_15549,N_15921);
xor U16479 (N_16479,N_15837,N_15889);
xor U16480 (N_16480,N_15555,N_15890);
and U16481 (N_16481,N_15529,N_15804);
and U16482 (N_16482,N_15867,N_15551);
or U16483 (N_16483,N_15888,N_15581);
or U16484 (N_16484,N_15898,N_15984);
or U16485 (N_16485,N_15859,N_15539);
or U16486 (N_16486,N_15570,N_15790);
nand U16487 (N_16487,N_15967,N_15573);
nand U16488 (N_16488,N_15647,N_15572);
xnor U16489 (N_16489,N_15518,N_15659);
nor U16490 (N_16490,N_15579,N_15616);
xor U16491 (N_16491,N_15931,N_15715);
nand U16492 (N_16492,N_15929,N_15886);
nor U16493 (N_16493,N_15787,N_15598);
nand U16494 (N_16494,N_15636,N_15754);
or U16495 (N_16495,N_15779,N_15911);
xor U16496 (N_16496,N_15643,N_15907);
nor U16497 (N_16497,N_15551,N_15652);
nand U16498 (N_16498,N_15735,N_15620);
and U16499 (N_16499,N_15685,N_15557);
xnor U16500 (N_16500,N_16135,N_16022);
nor U16501 (N_16501,N_16004,N_16292);
nor U16502 (N_16502,N_16437,N_16358);
nand U16503 (N_16503,N_16368,N_16092);
nand U16504 (N_16504,N_16265,N_16290);
and U16505 (N_16505,N_16408,N_16277);
xnor U16506 (N_16506,N_16248,N_16212);
nand U16507 (N_16507,N_16220,N_16475);
nand U16508 (N_16508,N_16268,N_16060);
nor U16509 (N_16509,N_16132,N_16012);
xnor U16510 (N_16510,N_16481,N_16474);
nor U16511 (N_16511,N_16080,N_16199);
nor U16512 (N_16512,N_16215,N_16353);
nand U16513 (N_16513,N_16233,N_16315);
nor U16514 (N_16514,N_16355,N_16445);
nand U16515 (N_16515,N_16056,N_16057);
nor U16516 (N_16516,N_16103,N_16007);
nand U16517 (N_16517,N_16403,N_16304);
nand U16518 (N_16518,N_16381,N_16407);
or U16519 (N_16519,N_16446,N_16145);
or U16520 (N_16520,N_16066,N_16010);
nor U16521 (N_16521,N_16061,N_16226);
xor U16522 (N_16522,N_16418,N_16089);
and U16523 (N_16523,N_16404,N_16105);
nand U16524 (N_16524,N_16297,N_16399);
xnor U16525 (N_16525,N_16114,N_16318);
nor U16526 (N_16526,N_16207,N_16347);
nor U16527 (N_16527,N_16062,N_16458);
nor U16528 (N_16528,N_16093,N_16067);
or U16529 (N_16529,N_16468,N_16161);
nor U16530 (N_16530,N_16043,N_16371);
xnor U16531 (N_16531,N_16213,N_16117);
nand U16532 (N_16532,N_16175,N_16072);
nand U16533 (N_16533,N_16470,N_16225);
nor U16534 (N_16534,N_16227,N_16050);
and U16535 (N_16535,N_16413,N_16183);
nor U16536 (N_16536,N_16477,N_16473);
or U16537 (N_16537,N_16307,N_16359);
nor U16538 (N_16538,N_16234,N_16037);
nand U16539 (N_16539,N_16003,N_16260);
or U16540 (N_16540,N_16375,N_16008);
xnor U16541 (N_16541,N_16452,N_16025);
xnor U16542 (N_16542,N_16148,N_16074);
xnor U16543 (N_16543,N_16224,N_16163);
nor U16544 (N_16544,N_16389,N_16172);
xor U16545 (N_16545,N_16366,N_16186);
nand U16546 (N_16546,N_16208,N_16121);
or U16547 (N_16547,N_16480,N_16002);
or U16548 (N_16548,N_16270,N_16082);
xnor U16549 (N_16549,N_16306,N_16115);
xnor U16550 (N_16550,N_16461,N_16137);
nor U16551 (N_16551,N_16210,N_16152);
or U16552 (N_16552,N_16125,N_16372);
or U16553 (N_16553,N_16143,N_16344);
nand U16554 (N_16554,N_16127,N_16239);
or U16555 (N_16555,N_16426,N_16046);
and U16556 (N_16556,N_16419,N_16450);
and U16557 (N_16557,N_16476,N_16054);
nand U16558 (N_16558,N_16332,N_16222);
and U16559 (N_16559,N_16424,N_16126);
xor U16560 (N_16560,N_16243,N_16442);
and U16561 (N_16561,N_16231,N_16241);
nor U16562 (N_16562,N_16487,N_16354);
nor U16563 (N_16563,N_16469,N_16052);
xor U16564 (N_16564,N_16406,N_16328);
nor U16565 (N_16565,N_16288,N_16324);
and U16566 (N_16566,N_16451,N_16484);
xor U16567 (N_16567,N_16258,N_16174);
and U16568 (N_16568,N_16298,N_16109);
and U16569 (N_16569,N_16144,N_16496);
nor U16570 (N_16570,N_16078,N_16216);
xnor U16571 (N_16571,N_16077,N_16108);
nand U16572 (N_16572,N_16266,N_16032);
and U16573 (N_16573,N_16123,N_16369);
nand U16574 (N_16574,N_16017,N_16176);
and U16575 (N_16575,N_16420,N_16486);
and U16576 (N_16576,N_16257,N_16203);
nand U16577 (N_16577,N_16036,N_16141);
nor U16578 (N_16578,N_16015,N_16088);
and U16579 (N_16579,N_16201,N_16422);
nor U16580 (N_16580,N_16416,N_16149);
or U16581 (N_16581,N_16086,N_16223);
xor U16582 (N_16582,N_16081,N_16031);
and U16583 (N_16583,N_16417,N_16357);
or U16584 (N_16584,N_16342,N_16168);
or U16585 (N_16585,N_16471,N_16099);
and U16586 (N_16586,N_16439,N_16205);
and U16587 (N_16587,N_16073,N_16443);
xnor U16588 (N_16588,N_16158,N_16444);
nor U16589 (N_16589,N_16494,N_16423);
xor U16590 (N_16590,N_16402,N_16398);
and U16591 (N_16591,N_16206,N_16460);
nand U16592 (N_16592,N_16281,N_16181);
nor U16593 (N_16593,N_16409,N_16323);
nor U16594 (N_16594,N_16156,N_16498);
or U16595 (N_16595,N_16334,N_16346);
or U16596 (N_16596,N_16111,N_16244);
nand U16597 (N_16597,N_16440,N_16090);
xnor U16598 (N_16598,N_16285,N_16302);
and U16599 (N_16599,N_16236,N_16000);
nor U16600 (N_16600,N_16335,N_16329);
nand U16601 (N_16601,N_16033,N_16263);
or U16602 (N_16602,N_16142,N_16383);
nand U16603 (N_16603,N_16068,N_16278);
nor U16604 (N_16604,N_16179,N_16316);
xnor U16605 (N_16605,N_16110,N_16364);
and U16606 (N_16606,N_16493,N_16049);
nand U16607 (N_16607,N_16096,N_16211);
and U16608 (N_16608,N_16479,N_16178);
xnor U16609 (N_16609,N_16262,N_16330);
xnor U16610 (N_16610,N_16360,N_16427);
nor U16611 (N_16611,N_16284,N_16345);
nand U16612 (N_16612,N_16151,N_16162);
xor U16613 (N_16613,N_16497,N_16245);
nand U16614 (N_16614,N_16412,N_16275);
nor U16615 (N_16615,N_16251,N_16140);
xor U16616 (N_16616,N_16113,N_16386);
and U16617 (N_16617,N_16079,N_16261);
nor U16618 (N_16618,N_16028,N_16130);
or U16619 (N_16619,N_16349,N_16352);
or U16620 (N_16620,N_16177,N_16035);
nand U16621 (N_16621,N_16048,N_16188);
or U16622 (N_16622,N_16184,N_16038);
xnor U16623 (N_16623,N_16485,N_16146);
nand U16624 (N_16624,N_16454,N_16271);
nor U16625 (N_16625,N_16456,N_16308);
or U16626 (N_16626,N_16235,N_16467);
nand U16627 (N_16627,N_16014,N_16134);
nor U16628 (N_16628,N_16321,N_16378);
and U16629 (N_16629,N_16387,N_16361);
and U16630 (N_16630,N_16438,N_16120);
nand U16631 (N_16631,N_16400,N_16018);
nor U16632 (N_16632,N_16465,N_16291);
and U16633 (N_16633,N_16180,N_16217);
or U16634 (N_16634,N_16129,N_16436);
nand U16635 (N_16635,N_16097,N_16299);
nor U16636 (N_16636,N_16122,N_16191);
and U16637 (N_16637,N_16295,N_16457);
and U16638 (N_16638,N_16491,N_16382);
or U16639 (N_16639,N_16350,N_16197);
or U16640 (N_16640,N_16071,N_16273);
nand U16641 (N_16641,N_16160,N_16166);
and U16642 (N_16642,N_16429,N_16193);
xnor U16643 (N_16643,N_16076,N_16139);
or U16644 (N_16644,N_16393,N_16055);
xor U16645 (N_16645,N_16376,N_16356);
nand U16646 (N_16646,N_16392,N_16098);
nor U16647 (N_16647,N_16325,N_16362);
xor U16648 (N_16648,N_16252,N_16200);
xor U16649 (N_16649,N_16319,N_16034);
nand U16650 (N_16650,N_16185,N_16026);
and U16651 (N_16651,N_16101,N_16276);
nand U16652 (N_16652,N_16187,N_16322);
and U16653 (N_16653,N_16247,N_16040);
nor U16654 (N_16654,N_16274,N_16489);
nor U16655 (N_16655,N_16434,N_16464);
and U16656 (N_16656,N_16320,N_16459);
and U16657 (N_16657,N_16296,N_16059);
and U16658 (N_16658,N_16410,N_16432);
nor U16659 (N_16659,N_16029,N_16374);
nor U16660 (N_16660,N_16448,N_16384);
or U16661 (N_16661,N_16391,N_16138);
or U16662 (N_16662,N_16041,N_16006);
xor U16663 (N_16663,N_16255,N_16395);
nor U16664 (N_16664,N_16100,N_16287);
nor U16665 (N_16665,N_16147,N_16001);
nand U16666 (N_16666,N_16131,N_16337);
or U16667 (N_16667,N_16058,N_16069);
nor U16668 (N_16668,N_16280,N_16343);
or U16669 (N_16669,N_16300,N_16085);
or U16670 (N_16670,N_16020,N_16202);
or U16671 (N_16671,N_16194,N_16164);
xor U16672 (N_16672,N_16351,N_16240);
nor U16673 (N_16673,N_16190,N_16312);
xnor U16674 (N_16674,N_16167,N_16023);
and U16675 (N_16675,N_16198,N_16310);
nand U16676 (N_16676,N_16107,N_16195);
nor U16677 (N_16677,N_16118,N_16254);
nand U16678 (N_16678,N_16431,N_16153);
nor U16679 (N_16679,N_16363,N_16326);
nor U16680 (N_16680,N_16030,N_16094);
nand U16681 (N_16681,N_16182,N_16380);
or U16682 (N_16682,N_16449,N_16064);
or U16683 (N_16683,N_16331,N_16169);
or U16684 (N_16684,N_16051,N_16045);
nor U16685 (N_16685,N_16411,N_16478);
xnor U16686 (N_16686,N_16013,N_16367);
xnor U16687 (N_16687,N_16259,N_16070);
xor U16688 (N_16688,N_16441,N_16294);
nand U16689 (N_16689,N_16242,N_16425);
nand U16690 (N_16690,N_16430,N_16472);
nand U16691 (N_16691,N_16124,N_16104);
nand U16692 (N_16692,N_16133,N_16087);
nor U16693 (N_16693,N_16253,N_16112);
xor U16694 (N_16694,N_16196,N_16024);
xnor U16695 (N_16695,N_16394,N_16170);
and U16696 (N_16696,N_16229,N_16221);
or U16697 (N_16697,N_16490,N_16075);
and U16698 (N_16698,N_16483,N_16218);
nor U16699 (N_16699,N_16303,N_16039);
and U16700 (N_16700,N_16401,N_16173);
nor U16701 (N_16701,N_16269,N_16267);
or U16702 (N_16702,N_16305,N_16165);
or U16703 (N_16703,N_16171,N_16341);
and U16704 (N_16704,N_16495,N_16027);
and U16705 (N_16705,N_16447,N_16011);
nand U16706 (N_16706,N_16421,N_16116);
nand U16707 (N_16707,N_16053,N_16047);
or U16708 (N_16708,N_16150,N_16466);
nand U16709 (N_16709,N_16232,N_16327);
or U16710 (N_16710,N_16189,N_16388);
and U16711 (N_16711,N_16293,N_16377);
or U16712 (N_16712,N_16102,N_16311);
xor U16713 (N_16713,N_16462,N_16415);
or U16714 (N_16714,N_16065,N_16044);
and U16715 (N_16715,N_16042,N_16095);
xor U16716 (N_16716,N_16209,N_16228);
nand U16717 (N_16717,N_16286,N_16021);
xnor U16718 (N_16718,N_16317,N_16264);
nand U16719 (N_16719,N_16405,N_16414);
xnor U16720 (N_16720,N_16279,N_16385);
xnor U16721 (N_16721,N_16009,N_16390);
or U16722 (N_16722,N_16428,N_16063);
nor U16723 (N_16723,N_16301,N_16091);
nor U16724 (N_16724,N_16433,N_16453);
and U16725 (N_16725,N_16339,N_16373);
nand U16726 (N_16726,N_16237,N_16155);
or U16727 (N_16727,N_16005,N_16219);
xnor U16728 (N_16728,N_16492,N_16499);
nand U16729 (N_16729,N_16333,N_16379);
nor U16730 (N_16730,N_16282,N_16313);
nor U16731 (N_16731,N_16340,N_16157);
xor U16732 (N_16732,N_16246,N_16230);
or U16733 (N_16733,N_16019,N_16136);
nand U16734 (N_16734,N_16159,N_16314);
xor U16735 (N_16735,N_16397,N_16192);
nor U16736 (N_16736,N_16482,N_16083);
xor U16737 (N_16737,N_16365,N_16435);
nand U16738 (N_16738,N_16128,N_16283);
nand U16739 (N_16739,N_16154,N_16106);
nand U16740 (N_16740,N_16348,N_16272);
and U16741 (N_16741,N_16119,N_16309);
and U16742 (N_16742,N_16249,N_16338);
or U16743 (N_16743,N_16016,N_16289);
nand U16744 (N_16744,N_16336,N_16370);
nand U16745 (N_16745,N_16084,N_16396);
nor U16746 (N_16746,N_16256,N_16455);
and U16747 (N_16747,N_16204,N_16488);
or U16748 (N_16748,N_16250,N_16463);
or U16749 (N_16749,N_16214,N_16238);
xor U16750 (N_16750,N_16116,N_16342);
nand U16751 (N_16751,N_16328,N_16226);
and U16752 (N_16752,N_16398,N_16134);
xnor U16753 (N_16753,N_16172,N_16179);
nor U16754 (N_16754,N_16354,N_16360);
nand U16755 (N_16755,N_16362,N_16072);
or U16756 (N_16756,N_16363,N_16134);
and U16757 (N_16757,N_16367,N_16394);
nor U16758 (N_16758,N_16050,N_16058);
nor U16759 (N_16759,N_16238,N_16162);
and U16760 (N_16760,N_16395,N_16289);
nor U16761 (N_16761,N_16314,N_16418);
and U16762 (N_16762,N_16148,N_16016);
xnor U16763 (N_16763,N_16427,N_16225);
nand U16764 (N_16764,N_16449,N_16017);
nand U16765 (N_16765,N_16317,N_16193);
and U16766 (N_16766,N_16030,N_16132);
or U16767 (N_16767,N_16429,N_16186);
nor U16768 (N_16768,N_16449,N_16167);
and U16769 (N_16769,N_16218,N_16470);
nand U16770 (N_16770,N_16442,N_16194);
or U16771 (N_16771,N_16198,N_16073);
and U16772 (N_16772,N_16431,N_16103);
xnor U16773 (N_16773,N_16288,N_16088);
and U16774 (N_16774,N_16152,N_16063);
nor U16775 (N_16775,N_16283,N_16184);
or U16776 (N_16776,N_16405,N_16136);
xor U16777 (N_16777,N_16007,N_16379);
xnor U16778 (N_16778,N_16226,N_16107);
nand U16779 (N_16779,N_16154,N_16287);
nand U16780 (N_16780,N_16028,N_16179);
or U16781 (N_16781,N_16009,N_16487);
or U16782 (N_16782,N_16405,N_16478);
nor U16783 (N_16783,N_16012,N_16097);
or U16784 (N_16784,N_16318,N_16413);
nor U16785 (N_16785,N_16269,N_16490);
nand U16786 (N_16786,N_16351,N_16329);
or U16787 (N_16787,N_16286,N_16491);
nor U16788 (N_16788,N_16410,N_16115);
xnor U16789 (N_16789,N_16433,N_16249);
or U16790 (N_16790,N_16379,N_16370);
xor U16791 (N_16791,N_16350,N_16285);
or U16792 (N_16792,N_16465,N_16273);
nand U16793 (N_16793,N_16338,N_16074);
or U16794 (N_16794,N_16132,N_16383);
xnor U16795 (N_16795,N_16407,N_16023);
nor U16796 (N_16796,N_16218,N_16115);
xor U16797 (N_16797,N_16029,N_16455);
nand U16798 (N_16798,N_16295,N_16463);
and U16799 (N_16799,N_16492,N_16460);
or U16800 (N_16800,N_16046,N_16160);
nor U16801 (N_16801,N_16289,N_16384);
nor U16802 (N_16802,N_16398,N_16336);
or U16803 (N_16803,N_16434,N_16033);
nand U16804 (N_16804,N_16056,N_16002);
and U16805 (N_16805,N_16170,N_16132);
xnor U16806 (N_16806,N_16440,N_16281);
nand U16807 (N_16807,N_16461,N_16132);
and U16808 (N_16808,N_16043,N_16022);
nor U16809 (N_16809,N_16046,N_16247);
xor U16810 (N_16810,N_16242,N_16498);
xor U16811 (N_16811,N_16106,N_16067);
nor U16812 (N_16812,N_16391,N_16283);
nand U16813 (N_16813,N_16462,N_16242);
nand U16814 (N_16814,N_16382,N_16337);
or U16815 (N_16815,N_16288,N_16356);
xnor U16816 (N_16816,N_16052,N_16132);
nor U16817 (N_16817,N_16485,N_16140);
nand U16818 (N_16818,N_16298,N_16033);
xnor U16819 (N_16819,N_16232,N_16337);
nand U16820 (N_16820,N_16400,N_16392);
nor U16821 (N_16821,N_16061,N_16222);
nor U16822 (N_16822,N_16464,N_16123);
or U16823 (N_16823,N_16352,N_16001);
or U16824 (N_16824,N_16371,N_16088);
xnor U16825 (N_16825,N_16190,N_16493);
nand U16826 (N_16826,N_16468,N_16363);
xor U16827 (N_16827,N_16325,N_16176);
or U16828 (N_16828,N_16298,N_16059);
and U16829 (N_16829,N_16025,N_16078);
nand U16830 (N_16830,N_16282,N_16469);
and U16831 (N_16831,N_16222,N_16201);
or U16832 (N_16832,N_16278,N_16423);
and U16833 (N_16833,N_16040,N_16499);
xor U16834 (N_16834,N_16174,N_16039);
xor U16835 (N_16835,N_16243,N_16076);
and U16836 (N_16836,N_16122,N_16235);
nor U16837 (N_16837,N_16496,N_16299);
and U16838 (N_16838,N_16204,N_16450);
or U16839 (N_16839,N_16103,N_16167);
or U16840 (N_16840,N_16399,N_16374);
nand U16841 (N_16841,N_16118,N_16320);
or U16842 (N_16842,N_16035,N_16301);
nor U16843 (N_16843,N_16243,N_16310);
nand U16844 (N_16844,N_16102,N_16424);
and U16845 (N_16845,N_16170,N_16077);
nand U16846 (N_16846,N_16218,N_16414);
or U16847 (N_16847,N_16080,N_16191);
nor U16848 (N_16848,N_16497,N_16336);
nor U16849 (N_16849,N_16085,N_16124);
nor U16850 (N_16850,N_16015,N_16005);
and U16851 (N_16851,N_16408,N_16475);
xnor U16852 (N_16852,N_16180,N_16190);
and U16853 (N_16853,N_16380,N_16156);
xor U16854 (N_16854,N_16429,N_16357);
and U16855 (N_16855,N_16263,N_16425);
xnor U16856 (N_16856,N_16292,N_16105);
or U16857 (N_16857,N_16137,N_16373);
xnor U16858 (N_16858,N_16382,N_16219);
and U16859 (N_16859,N_16222,N_16497);
nor U16860 (N_16860,N_16025,N_16077);
xnor U16861 (N_16861,N_16353,N_16144);
nor U16862 (N_16862,N_16031,N_16295);
xnor U16863 (N_16863,N_16300,N_16093);
and U16864 (N_16864,N_16145,N_16310);
and U16865 (N_16865,N_16161,N_16475);
and U16866 (N_16866,N_16261,N_16185);
and U16867 (N_16867,N_16144,N_16430);
and U16868 (N_16868,N_16493,N_16172);
nand U16869 (N_16869,N_16302,N_16033);
nor U16870 (N_16870,N_16346,N_16305);
nand U16871 (N_16871,N_16056,N_16102);
or U16872 (N_16872,N_16282,N_16306);
xnor U16873 (N_16873,N_16134,N_16264);
nor U16874 (N_16874,N_16496,N_16244);
or U16875 (N_16875,N_16283,N_16393);
xor U16876 (N_16876,N_16086,N_16458);
nor U16877 (N_16877,N_16465,N_16164);
and U16878 (N_16878,N_16499,N_16482);
xor U16879 (N_16879,N_16225,N_16312);
or U16880 (N_16880,N_16053,N_16044);
xor U16881 (N_16881,N_16284,N_16250);
nand U16882 (N_16882,N_16294,N_16351);
xor U16883 (N_16883,N_16034,N_16214);
nor U16884 (N_16884,N_16457,N_16458);
or U16885 (N_16885,N_16348,N_16394);
nor U16886 (N_16886,N_16430,N_16075);
xnor U16887 (N_16887,N_16086,N_16300);
nand U16888 (N_16888,N_16419,N_16260);
xor U16889 (N_16889,N_16135,N_16404);
or U16890 (N_16890,N_16325,N_16470);
and U16891 (N_16891,N_16286,N_16219);
xor U16892 (N_16892,N_16239,N_16265);
or U16893 (N_16893,N_16207,N_16316);
nor U16894 (N_16894,N_16080,N_16124);
or U16895 (N_16895,N_16183,N_16089);
nor U16896 (N_16896,N_16049,N_16223);
nand U16897 (N_16897,N_16114,N_16049);
xor U16898 (N_16898,N_16266,N_16093);
nor U16899 (N_16899,N_16081,N_16159);
and U16900 (N_16900,N_16182,N_16047);
nor U16901 (N_16901,N_16487,N_16159);
nand U16902 (N_16902,N_16052,N_16041);
nand U16903 (N_16903,N_16309,N_16450);
or U16904 (N_16904,N_16074,N_16005);
nand U16905 (N_16905,N_16307,N_16329);
nor U16906 (N_16906,N_16143,N_16092);
or U16907 (N_16907,N_16389,N_16055);
nand U16908 (N_16908,N_16016,N_16031);
nand U16909 (N_16909,N_16424,N_16053);
and U16910 (N_16910,N_16128,N_16231);
nor U16911 (N_16911,N_16092,N_16390);
and U16912 (N_16912,N_16116,N_16013);
nor U16913 (N_16913,N_16149,N_16469);
nor U16914 (N_16914,N_16289,N_16326);
nor U16915 (N_16915,N_16175,N_16292);
nand U16916 (N_16916,N_16010,N_16347);
and U16917 (N_16917,N_16081,N_16251);
and U16918 (N_16918,N_16325,N_16255);
nand U16919 (N_16919,N_16103,N_16397);
or U16920 (N_16920,N_16144,N_16349);
and U16921 (N_16921,N_16428,N_16202);
xnor U16922 (N_16922,N_16073,N_16310);
or U16923 (N_16923,N_16019,N_16110);
xnor U16924 (N_16924,N_16167,N_16212);
and U16925 (N_16925,N_16385,N_16337);
xor U16926 (N_16926,N_16113,N_16189);
nand U16927 (N_16927,N_16359,N_16054);
nor U16928 (N_16928,N_16335,N_16181);
and U16929 (N_16929,N_16431,N_16470);
nand U16930 (N_16930,N_16104,N_16487);
nor U16931 (N_16931,N_16048,N_16077);
nand U16932 (N_16932,N_16028,N_16277);
xnor U16933 (N_16933,N_16421,N_16104);
or U16934 (N_16934,N_16446,N_16373);
or U16935 (N_16935,N_16044,N_16274);
xor U16936 (N_16936,N_16101,N_16286);
nand U16937 (N_16937,N_16387,N_16213);
and U16938 (N_16938,N_16229,N_16172);
nor U16939 (N_16939,N_16129,N_16474);
nand U16940 (N_16940,N_16096,N_16274);
xnor U16941 (N_16941,N_16300,N_16114);
or U16942 (N_16942,N_16220,N_16348);
xor U16943 (N_16943,N_16057,N_16213);
nand U16944 (N_16944,N_16112,N_16106);
and U16945 (N_16945,N_16033,N_16212);
nor U16946 (N_16946,N_16120,N_16461);
and U16947 (N_16947,N_16012,N_16249);
nand U16948 (N_16948,N_16395,N_16336);
xnor U16949 (N_16949,N_16385,N_16165);
or U16950 (N_16950,N_16381,N_16383);
xor U16951 (N_16951,N_16057,N_16113);
nand U16952 (N_16952,N_16331,N_16258);
xnor U16953 (N_16953,N_16237,N_16273);
and U16954 (N_16954,N_16407,N_16322);
nor U16955 (N_16955,N_16405,N_16357);
nand U16956 (N_16956,N_16230,N_16153);
and U16957 (N_16957,N_16342,N_16343);
xnor U16958 (N_16958,N_16091,N_16444);
or U16959 (N_16959,N_16406,N_16421);
nand U16960 (N_16960,N_16153,N_16231);
xnor U16961 (N_16961,N_16499,N_16065);
xor U16962 (N_16962,N_16073,N_16215);
nor U16963 (N_16963,N_16132,N_16066);
nand U16964 (N_16964,N_16427,N_16413);
and U16965 (N_16965,N_16355,N_16028);
or U16966 (N_16966,N_16399,N_16038);
or U16967 (N_16967,N_16174,N_16150);
nor U16968 (N_16968,N_16382,N_16147);
nand U16969 (N_16969,N_16164,N_16371);
nand U16970 (N_16970,N_16398,N_16073);
xnor U16971 (N_16971,N_16408,N_16462);
xnor U16972 (N_16972,N_16393,N_16392);
or U16973 (N_16973,N_16195,N_16379);
and U16974 (N_16974,N_16321,N_16392);
nand U16975 (N_16975,N_16241,N_16256);
and U16976 (N_16976,N_16286,N_16079);
xor U16977 (N_16977,N_16487,N_16380);
nor U16978 (N_16978,N_16258,N_16466);
or U16979 (N_16979,N_16050,N_16392);
xnor U16980 (N_16980,N_16127,N_16073);
or U16981 (N_16981,N_16015,N_16033);
nand U16982 (N_16982,N_16335,N_16427);
and U16983 (N_16983,N_16400,N_16194);
and U16984 (N_16984,N_16427,N_16399);
nor U16985 (N_16985,N_16237,N_16217);
nand U16986 (N_16986,N_16084,N_16373);
and U16987 (N_16987,N_16306,N_16090);
and U16988 (N_16988,N_16370,N_16243);
nand U16989 (N_16989,N_16163,N_16410);
and U16990 (N_16990,N_16030,N_16462);
nor U16991 (N_16991,N_16014,N_16196);
and U16992 (N_16992,N_16003,N_16074);
and U16993 (N_16993,N_16254,N_16185);
nor U16994 (N_16994,N_16084,N_16270);
or U16995 (N_16995,N_16289,N_16373);
or U16996 (N_16996,N_16468,N_16489);
or U16997 (N_16997,N_16006,N_16160);
xor U16998 (N_16998,N_16100,N_16088);
xor U16999 (N_16999,N_16040,N_16426);
or U17000 (N_17000,N_16537,N_16971);
xnor U17001 (N_17001,N_16792,N_16618);
or U17002 (N_17002,N_16521,N_16536);
xor U17003 (N_17003,N_16833,N_16579);
and U17004 (N_17004,N_16892,N_16730);
nor U17005 (N_17005,N_16816,N_16791);
nor U17006 (N_17006,N_16852,N_16704);
and U17007 (N_17007,N_16800,N_16986);
nand U17008 (N_17008,N_16864,N_16566);
or U17009 (N_17009,N_16809,N_16847);
or U17010 (N_17010,N_16534,N_16661);
and U17011 (N_17011,N_16738,N_16538);
and U17012 (N_17012,N_16645,N_16637);
or U17013 (N_17013,N_16855,N_16894);
or U17014 (N_17014,N_16502,N_16983);
xnor U17015 (N_17015,N_16587,N_16743);
xor U17016 (N_17016,N_16844,N_16780);
nand U17017 (N_17017,N_16557,N_16575);
xor U17018 (N_17018,N_16735,N_16762);
or U17019 (N_17019,N_16509,N_16741);
and U17020 (N_17020,N_16520,N_16649);
or U17021 (N_17021,N_16760,N_16937);
nor U17022 (N_17022,N_16736,N_16962);
and U17023 (N_17023,N_16872,N_16769);
and U17024 (N_17024,N_16943,N_16912);
nor U17025 (N_17025,N_16646,N_16705);
or U17026 (N_17026,N_16569,N_16626);
or U17027 (N_17027,N_16694,N_16977);
and U17028 (N_17028,N_16878,N_16553);
and U17029 (N_17029,N_16643,N_16710);
xor U17030 (N_17030,N_16856,N_16776);
xor U17031 (N_17031,N_16834,N_16673);
and U17032 (N_17032,N_16934,N_16529);
xnor U17033 (N_17033,N_16748,N_16805);
xor U17034 (N_17034,N_16850,N_16863);
or U17035 (N_17035,N_16562,N_16770);
nand U17036 (N_17036,N_16953,N_16758);
or U17037 (N_17037,N_16820,N_16518);
nor U17038 (N_17038,N_16706,N_16714);
nor U17039 (N_17039,N_16788,N_16727);
and U17040 (N_17040,N_16884,N_16978);
xor U17041 (N_17041,N_16530,N_16604);
nor U17042 (N_17042,N_16556,N_16775);
or U17043 (N_17043,N_16558,N_16565);
and U17044 (N_17044,N_16582,N_16806);
or U17045 (N_17045,N_16860,N_16511);
and U17046 (N_17046,N_16592,N_16890);
nor U17047 (N_17047,N_16628,N_16919);
nor U17048 (N_17048,N_16550,N_16989);
nor U17049 (N_17049,N_16915,N_16612);
nor U17050 (N_17050,N_16940,N_16923);
and U17051 (N_17051,N_16564,N_16808);
xor U17052 (N_17052,N_16602,N_16638);
xor U17053 (N_17053,N_16795,N_16754);
nand U17054 (N_17054,N_16528,N_16688);
nand U17055 (N_17055,N_16990,N_16681);
nand U17056 (N_17056,N_16910,N_16984);
xnor U17057 (N_17057,N_16596,N_16887);
nand U17058 (N_17058,N_16512,N_16655);
and U17059 (N_17059,N_16695,N_16902);
or U17060 (N_17060,N_16929,N_16563);
nand U17061 (N_17061,N_16689,N_16682);
or U17062 (N_17062,N_16680,N_16924);
nand U17063 (N_17063,N_16866,N_16697);
nand U17064 (N_17064,N_16969,N_16621);
and U17065 (N_17065,N_16801,N_16551);
nor U17066 (N_17066,N_16731,N_16876);
and U17067 (N_17067,N_16614,N_16519);
or U17068 (N_17068,N_16939,N_16664);
and U17069 (N_17069,N_16747,N_16718);
nand U17070 (N_17070,N_16812,N_16843);
and U17071 (N_17071,N_16609,N_16574);
and U17072 (N_17072,N_16669,N_16639);
and U17073 (N_17073,N_16584,N_16685);
and U17074 (N_17074,N_16968,N_16693);
or U17075 (N_17075,N_16822,N_16837);
nand U17076 (N_17076,N_16959,N_16598);
nand U17077 (N_17077,N_16981,N_16901);
xor U17078 (N_17078,N_16601,N_16828);
or U17079 (N_17079,N_16572,N_16514);
or U17080 (N_17080,N_16963,N_16524);
and U17081 (N_17081,N_16737,N_16966);
and U17082 (N_17082,N_16607,N_16961);
xor U17083 (N_17083,N_16802,N_16883);
nand U17084 (N_17084,N_16672,N_16952);
nand U17085 (N_17085,N_16796,N_16829);
xnor U17086 (N_17086,N_16996,N_16577);
nand U17087 (N_17087,N_16980,N_16641);
xnor U17088 (N_17088,N_16836,N_16650);
nor U17089 (N_17089,N_16542,N_16555);
nor U17090 (N_17090,N_16900,N_16867);
nand U17091 (N_17091,N_16955,N_16616);
nand U17092 (N_17092,N_16576,N_16667);
or U17093 (N_17093,N_16956,N_16723);
nand U17094 (N_17094,N_16753,N_16819);
xor U17095 (N_17095,N_16677,N_16831);
and U17096 (N_17096,N_16648,N_16993);
nor U17097 (N_17097,N_16913,N_16657);
nor U17098 (N_17098,N_16728,N_16504);
xnor U17099 (N_17099,N_16505,N_16586);
nor U17100 (N_17100,N_16666,N_16580);
and U17101 (N_17101,N_16513,N_16713);
xnor U17102 (N_17102,N_16692,N_16789);
and U17103 (N_17103,N_16948,N_16578);
or U17104 (N_17104,N_16599,N_16739);
xor U17105 (N_17105,N_16658,N_16818);
xnor U17106 (N_17106,N_16740,N_16585);
xnor U17107 (N_17107,N_16691,N_16659);
nor U17108 (N_17108,N_16597,N_16708);
or U17109 (N_17109,N_16916,N_16671);
and U17110 (N_17110,N_16782,N_16832);
nor U17111 (N_17111,N_16633,N_16627);
nand U17112 (N_17112,N_16868,N_16749);
and U17113 (N_17113,N_16531,N_16732);
or U17114 (N_17114,N_16768,N_16701);
or U17115 (N_17115,N_16991,N_16975);
nand U17116 (N_17116,N_16532,N_16539);
xnor U17117 (N_17117,N_16613,N_16676);
and U17118 (N_17118,N_16783,N_16931);
nand U17119 (N_17119,N_16651,N_16547);
and U17120 (N_17120,N_16759,N_16696);
xor U17121 (N_17121,N_16640,N_16811);
nor U17122 (N_17122,N_16567,N_16583);
and U17123 (N_17123,N_16814,N_16798);
or U17124 (N_17124,N_16620,N_16665);
or U17125 (N_17125,N_16914,N_16548);
or U17126 (N_17126,N_16570,N_16979);
nand U17127 (N_17127,N_16930,N_16686);
nor U17128 (N_17128,N_16862,N_16830);
nand U17129 (N_17129,N_16715,N_16810);
or U17130 (N_17130,N_16687,N_16938);
xor U17131 (N_17131,N_16644,N_16871);
xor U17132 (N_17132,N_16772,N_16908);
nor U17133 (N_17133,N_16857,N_16917);
nor U17134 (N_17134,N_16985,N_16660);
or U17135 (N_17135,N_16560,N_16543);
nand U17136 (N_17136,N_16624,N_16561);
xnor U17137 (N_17137,N_16763,N_16522);
or U17138 (N_17138,N_16733,N_16779);
and U17139 (N_17139,N_16711,N_16839);
xor U17140 (N_17140,N_16652,N_16925);
nand U17141 (N_17141,N_16717,N_16859);
nor U17142 (N_17142,N_16703,N_16675);
or U17143 (N_17143,N_16552,N_16720);
nand U17144 (N_17144,N_16778,N_16851);
xnor U17145 (N_17145,N_16882,N_16593);
or U17146 (N_17146,N_16588,N_16960);
or U17147 (N_17147,N_16840,N_16623);
nand U17148 (N_17148,N_16813,N_16881);
or U17149 (N_17149,N_16744,N_16619);
nand U17150 (N_17150,N_16764,N_16610);
xnor U17151 (N_17151,N_16794,N_16972);
nor U17152 (N_17152,N_16950,N_16865);
nand U17153 (N_17153,N_16909,N_16899);
nor U17154 (N_17154,N_16523,N_16995);
xnor U17155 (N_17155,N_16501,N_16507);
or U17156 (N_17156,N_16726,N_16880);
and U17157 (N_17157,N_16589,N_16988);
nor U17158 (N_17158,N_16936,N_16678);
xor U17159 (N_17159,N_16510,N_16886);
nor U17160 (N_17160,N_16911,N_16891);
xnor U17161 (N_17161,N_16729,N_16841);
or U17162 (N_17162,N_16721,N_16949);
xnor U17163 (N_17163,N_16750,N_16893);
or U17164 (N_17164,N_16635,N_16757);
nor U17165 (N_17165,N_16875,N_16670);
nor U17166 (N_17166,N_16874,N_16947);
or U17167 (N_17167,N_16853,N_16964);
xor U17168 (N_17168,N_16656,N_16973);
and U17169 (N_17169,N_16581,N_16611);
xnor U17170 (N_17170,N_16545,N_16752);
nand U17171 (N_17171,N_16516,N_16642);
nor U17172 (N_17172,N_16858,N_16674);
nand U17173 (N_17173,N_16998,N_16889);
or U17174 (N_17174,N_16719,N_16571);
nor U17175 (N_17175,N_16906,N_16987);
or U17176 (N_17176,N_16515,N_16605);
and U17177 (N_17177,N_16815,N_16756);
and U17178 (N_17178,N_16927,N_16594);
xnor U17179 (N_17179,N_16653,N_16544);
or U17180 (N_17180,N_16785,N_16921);
nor U17181 (N_17181,N_16821,N_16781);
nor U17182 (N_17182,N_16679,N_16974);
nor U17183 (N_17183,N_16625,N_16848);
or U17184 (N_17184,N_16767,N_16707);
nand U17185 (N_17185,N_16541,N_16928);
xor U17186 (N_17186,N_16970,N_16994);
xor U17187 (N_17187,N_16699,N_16745);
xnor U17188 (N_17188,N_16765,N_16976);
or U17189 (N_17189,N_16634,N_16944);
or U17190 (N_17190,N_16957,N_16500);
nor U17191 (N_17191,N_16662,N_16700);
nor U17192 (N_17192,N_16709,N_16842);
nand U17193 (N_17193,N_16722,N_16845);
or U17194 (N_17194,N_16824,N_16907);
or U17195 (N_17195,N_16941,N_16965);
nand U17196 (N_17196,N_16517,N_16797);
nor U17197 (N_17197,N_16873,N_16967);
nand U17198 (N_17198,N_16904,N_16590);
and U17199 (N_17199,N_16896,N_16793);
nand U17200 (N_17200,N_16631,N_16647);
and U17201 (N_17201,N_16942,N_16849);
nor U17202 (N_17202,N_16826,N_16698);
and U17203 (N_17203,N_16905,N_16958);
and U17204 (N_17204,N_16807,N_16506);
xor U17205 (N_17205,N_16982,N_16823);
and U17206 (N_17206,N_16997,N_16766);
nor U17207 (N_17207,N_16526,N_16636);
nand U17208 (N_17208,N_16918,N_16835);
xor U17209 (N_17209,N_16746,N_16885);
xnor U17210 (N_17210,N_16724,N_16725);
nor U17211 (N_17211,N_16773,N_16926);
nor U17212 (N_17212,N_16922,N_16568);
and U17213 (N_17213,N_16603,N_16898);
and U17214 (N_17214,N_16559,N_16771);
or U17215 (N_17215,N_16615,N_16549);
nand U17216 (N_17216,N_16663,N_16895);
xnor U17217 (N_17217,N_16654,N_16879);
nand U17218 (N_17218,N_16702,N_16854);
xor U17219 (N_17219,N_16533,N_16712);
and U17220 (N_17220,N_16827,N_16825);
nor U17221 (N_17221,N_16755,N_16784);
and U17222 (N_17222,N_16668,N_16888);
xnor U17223 (N_17223,N_16992,N_16690);
xor U17224 (N_17224,N_16932,N_16527);
and U17225 (N_17225,N_16632,N_16608);
xor U17226 (N_17226,N_16799,N_16573);
xnor U17227 (N_17227,N_16846,N_16946);
nor U17228 (N_17228,N_16540,N_16503);
and U17229 (N_17229,N_16751,N_16999);
nand U17230 (N_17230,N_16804,N_16617);
or U17231 (N_17231,N_16683,N_16595);
nor U17232 (N_17232,N_16803,N_16933);
nor U17233 (N_17233,N_16525,N_16838);
xor U17234 (N_17234,N_16546,N_16629);
nor U17235 (N_17235,N_16869,N_16777);
or U17236 (N_17236,N_16897,N_16954);
xnor U17237 (N_17237,N_16817,N_16945);
nor U17238 (N_17238,N_16554,N_16508);
nor U17239 (N_17239,N_16684,N_16734);
and U17240 (N_17240,N_16790,N_16716);
and U17241 (N_17241,N_16951,N_16861);
nor U17242 (N_17242,N_16591,N_16903);
nor U17243 (N_17243,N_16786,N_16535);
nor U17244 (N_17244,N_16774,N_16787);
or U17245 (N_17245,N_16630,N_16742);
or U17246 (N_17246,N_16935,N_16600);
nor U17247 (N_17247,N_16622,N_16877);
and U17248 (N_17248,N_16761,N_16606);
nand U17249 (N_17249,N_16870,N_16920);
and U17250 (N_17250,N_16769,N_16563);
nor U17251 (N_17251,N_16546,N_16990);
xor U17252 (N_17252,N_16663,N_16633);
nand U17253 (N_17253,N_16510,N_16744);
and U17254 (N_17254,N_16958,N_16909);
or U17255 (N_17255,N_16848,N_16884);
nand U17256 (N_17256,N_16732,N_16919);
nand U17257 (N_17257,N_16996,N_16505);
nor U17258 (N_17258,N_16733,N_16560);
or U17259 (N_17259,N_16548,N_16653);
xnor U17260 (N_17260,N_16944,N_16773);
nor U17261 (N_17261,N_16976,N_16747);
nand U17262 (N_17262,N_16703,N_16839);
or U17263 (N_17263,N_16962,N_16661);
or U17264 (N_17264,N_16623,N_16755);
nand U17265 (N_17265,N_16842,N_16927);
nand U17266 (N_17266,N_16823,N_16837);
and U17267 (N_17267,N_16527,N_16976);
or U17268 (N_17268,N_16774,N_16875);
and U17269 (N_17269,N_16524,N_16754);
or U17270 (N_17270,N_16570,N_16642);
nand U17271 (N_17271,N_16573,N_16644);
and U17272 (N_17272,N_16675,N_16939);
nor U17273 (N_17273,N_16907,N_16993);
and U17274 (N_17274,N_16634,N_16533);
and U17275 (N_17275,N_16593,N_16627);
nand U17276 (N_17276,N_16809,N_16990);
or U17277 (N_17277,N_16852,N_16761);
or U17278 (N_17278,N_16768,N_16724);
and U17279 (N_17279,N_16789,N_16516);
nand U17280 (N_17280,N_16696,N_16698);
nand U17281 (N_17281,N_16708,N_16693);
nor U17282 (N_17282,N_16924,N_16709);
nand U17283 (N_17283,N_16889,N_16999);
nand U17284 (N_17284,N_16632,N_16593);
or U17285 (N_17285,N_16979,N_16865);
nor U17286 (N_17286,N_16718,N_16716);
xnor U17287 (N_17287,N_16597,N_16726);
xor U17288 (N_17288,N_16732,N_16687);
nor U17289 (N_17289,N_16910,N_16821);
and U17290 (N_17290,N_16947,N_16645);
nand U17291 (N_17291,N_16746,N_16685);
nor U17292 (N_17292,N_16704,N_16876);
and U17293 (N_17293,N_16608,N_16934);
nor U17294 (N_17294,N_16805,N_16791);
and U17295 (N_17295,N_16983,N_16882);
nor U17296 (N_17296,N_16631,N_16593);
nor U17297 (N_17297,N_16560,N_16511);
nand U17298 (N_17298,N_16682,N_16822);
or U17299 (N_17299,N_16645,N_16769);
nand U17300 (N_17300,N_16594,N_16508);
nand U17301 (N_17301,N_16670,N_16944);
nor U17302 (N_17302,N_16703,N_16930);
nor U17303 (N_17303,N_16555,N_16863);
or U17304 (N_17304,N_16811,N_16759);
and U17305 (N_17305,N_16958,N_16850);
and U17306 (N_17306,N_16524,N_16544);
and U17307 (N_17307,N_16956,N_16538);
nand U17308 (N_17308,N_16806,N_16947);
or U17309 (N_17309,N_16546,N_16684);
nand U17310 (N_17310,N_16670,N_16785);
xor U17311 (N_17311,N_16610,N_16622);
or U17312 (N_17312,N_16841,N_16860);
or U17313 (N_17313,N_16661,N_16586);
or U17314 (N_17314,N_16766,N_16873);
and U17315 (N_17315,N_16562,N_16635);
nor U17316 (N_17316,N_16718,N_16974);
and U17317 (N_17317,N_16719,N_16760);
and U17318 (N_17318,N_16685,N_16981);
or U17319 (N_17319,N_16858,N_16731);
or U17320 (N_17320,N_16995,N_16862);
nand U17321 (N_17321,N_16692,N_16505);
and U17322 (N_17322,N_16591,N_16815);
or U17323 (N_17323,N_16862,N_16971);
and U17324 (N_17324,N_16814,N_16809);
and U17325 (N_17325,N_16629,N_16685);
xor U17326 (N_17326,N_16682,N_16677);
nand U17327 (N_17327,N_16775,N_16914);
nor U17328 (N_17328,N_16840,N_16564);
and U17329 (N_17329,N_16849,N_16714);
nand U17330 (N_17330,N_16907,N_16509);
nand U17331 (N_17331,N_16948,N_16931);
or U17332 (N_17332,N_16793,N_16741);
xor U17333 (N_17333,N_16903,N_16899);
or U17334 (N_17334,N_16877,N_16589);
nor U17335 (N_17335,N_16849,N_16872);
nand U17336 (N_17336,N_16835,N_16603);
and U17337 (N_17337,N_16767,N_16579);
xnor U17338 (N_17338,N_16862,N_16575);
xor U17339 (N_17339,N_16507,N_16635);
nand U17340 (N_17340,N_16803,N_16619);
or U17341 (N_17341,N_16612,N_16895);
nor U17342 (N_17342,N_16875,N_16504);
or U17343 (N_17343,N_16572,N_16552);
nand U17344 (N_17344,N_16571,N_16698);
nor U17345 (N_17345,N_16777,N_16593);
nand U17346 (N_17346,N_16548,N_16987);
nand U17347 (N_17347,N_16939,N_16737);
xor U17348 (N_17348,N_16660,N_16871);
and U17349 (N_17349,N_16977,N_16810);
or U17350 (N_17350,N_16685,N_16787);
nor U17351 (N_17351,N_16556,N_16510);
nor U17352 (N_17352,N_16970,N_16794);
or U17353 (N_17353,N_16601,N_16679);
and U17354 (N_17354,N_16911,N_16598);
nand U17355 (N_17355,N_16686,N_16794);
nor U17356 (N_17356,N_16703,N_16516);
nor U17357 (N_17357,N_16959,N_16743);
and U17358 (N_17358,N_16610,N_16665);
and U17359 (N_17359,N_16547,N_16918);
and U17360 (N_17360,N_16862,N_16756);
nand U17361 (N_17361,N_16918,N_16914);
or U17362 (N_17362,N_16575,N_16656);
xnor U17363 (N_17363,N_16698,N_16798);
or U17364 (N_17364,N_16708,N_16805);
nor U17365 (N_17365,N_16952,N_16567);
nand U17366 (N_17366,N_16917,N_16978);
xor U17367 (N_17367,N_16734,N_16686);
and U17368 (N_17368,N_16725,N_16972);
xor U17369 (N_17369,N_16951,N_16735);
nand U17370 (N_17370,N_16687,N_16637);
or U17371 (N_17371,N_16656,N_16953);
and U17372 (N_17372,N_16605,N_16936);
nand U17373 (N_17373,N_16646,N_16892);
and U17374 (N_17374,N_16838,N_16683);
nor U17375 (N_17375,N_16954,N_16961);
and U17376 (N_17376,N_16771,N_16598);
nor U17377 (N_17377,N_16753,N_16588);
or U17378 (N_17378,N_16909,N_16598);
nand U17379 (N_17379,N_16845,N_16718);
and U17380 (N_17380,N_16607,N_16724);
xnor U17381 (N_17381,N_16597,N_16951);
xnor U17382 (N_17382,N_16998,N_16938);
nand U17383 (N_17383,N_16717,N_16514);
or U17384 (N_17384,N_16674,N_16744);
or U17385 (N_17385,N_16667,N_16510);
or U17386 (N_17386,N_16569,N_16856);
nand U17387 (N_17387,N_16695,N_16866);
xor U17388 (N_17388,N_16823,N_16578);
nor U17389 (N_17389,N_16982,N_16731);
nand U17390 (N_17390,N_16822,N_16713);
or U17391 (N_17391,N_16995,N_16704);
xnor U17392 (N_17392,N_16717,N_16587);
nor U17393 (N_17393,N_16971,N_16749);
nor U17394 (N_17394,N_16955,N_16756);
or U17395 (N_17395,N_16770,N_16785);
nor U17396 (N_17396,N_16654,N_16849);
nand U17397 (N_17397,N_16854,N_16977);
or U17398 (N_17398,N_16680,N_16697);
or U17399 (N_17399,N_16861,N_16664);
nor U17400 (N_17400,N_16646,N_16998);
xor U17401 (N_17401,N_16755,N_16896);
xnor U17402 (N_17402,N_16792,N_16642);
or U17403 (N_17403,N_16865,N_16524);
nand U17404 (N_17404,N_16535,N_16870);
nor U17405 (N_17405,N_16734,N_16509);
nor U17406 (N_17406,N_16853,N_16818);
and U17407 (N_17407,N_16878,N_16519);
xor U17408 (N_17408,N_16600,N_16876);
and U17409 (N_17409,N_16591,N_16987);
or U17410 (N_17410,N_16947,N_16636);
nand U17411 (N_17411,N_16561,N_16942);
nand U17412 (N_17412,N_16543,N_16715);
xnor U17413 (N_17413,N_16758,N_16971);
nor U17414 (N_17414,N_16990,N_16913);
or U17415 (N_17415,N_16905,N_16916);
xor U17416 (N_17416,N_16996,N_16581);
xor U17417 (N_17417,N_16545,N_16601);
xnor U17418 (N_17418,N_16725,N_16932);
xnor U17419 (N_17419,N_16790,N_16767);
nor U17420 (N_17420,N_16560,N_16547);
xor U17421 (N_17421,N_16885,N_16859);
nand U17422 (N_17422,N_16951,N_16619);
and U17423 (N_17423,N_16525,N_16821);
nand U17424 (N_17424,N_16511,N_16825);
and U17425 (N_17425,N_16543,N_16654);
nor U17426 (N_17426,N_16624,N_16633);
nor U17427 (N_17427,N_16552,N_16837);
nand U17428 (N_17428,N_16936,N_16639);
xnor U17429 (N_17429,N_16568,N_16713);
or U17430 (N_17430,N_16627,N_16737);
nand U17431 (N_17431,N_16691,N_16935);
or U17432 (N_17432,N_16550,N_16903);
nand U17433 (N_17433,N_16610,N_16612);
nor U17434 (N_17434,N_16550,N_16540);
and U17435 (N_17435,N_16888,N_16615);
nor U17436 (N_17436,N_16596,N_16601);
nand U17437 (N_17437,N_16577,N_16997);
or U17438 (N_17438,N_16979,N_16715);
nand U17439 (N_17439,N_16524,N_16961);
or U17440 (N_17440,N_16848,N_16569);
xnor U17441 (N_17441,N_16749,N_16578);
xor U17442 (N_17442,N_16778,N_16991);
or U17443 (N_17443,N_16610,N_16683);
nand U17444 (N_17444,N_16789,N_16577);
nor U17445 (N_17445,N_16677,N_16704);
xor U17446 (N_17446,N_16826,N_16906);
nor U17447 (N_17447,N_16604,N_16675);
nand U17448 (N_17448,N_16655,N_16618);
nand U17449 (N_17449,N_16989,N_16887);
nand U17450 (N_17450,N_16893,N_16724);
nor U17451 (N_17451,N_16820,N_16903);
xor U17452 (N_17452,N_16774,N_16604);
nor U17453 (N_17453,N_16983,N_16716);
and U17454 (N_17454,N_16786,N_16929);
or U17455 (N_17455,N_16543,N_16699);
and U17456 (N_17456,N_16506,N_16707);
xnor U17457 (N_17457,N_16727,N_16598);
or U17458 (N_17458,N_16524,N_16912);
xnor U17459 (N_17459,N_16981,N_16522);
nor U17460 (N_17460,N_16915,N_16968);
and U17461 (N_17461,N_16938,N_16812);
and U17462 (N_17462,N_16697,N_16985);
nand U17463 (N_17463,N_16717,N_16808);
or U17464 (N_17464,N_16652,N_16836);
and U17465 (N_17465,N_16893,N_16744);
or U17466 (N_17466,N_16655,N_16647);
and U17467 (N_17467,N_16701,N_16609);
nor U17468 (N_17468,N_16683,N_16705);
xnor U17469 (N_17469,N_16986,N_16526);
or U17470 (N_17470,N_16816,N_16763);
nand U17471 (N_17471,N_16885,N_16635);
or U17472 (N_17472,N_16980,N_16753);
nand U17473 (N_17473,N_16662,N_16678);
or U17474 (N_17474,N_16727,N_16871);
and U17475 (N_17475,N_16943,N_16853);
nand U17476 (N_17476,N_16609,N_16729);
nand U17477 (N_17477,N_16991,N_16881);
xor U17478 (N_17478,N_16717,N_16555);
and U17479 (N_17479,N_16694,N_16741);
or U17480 (N_17480,N_16853,N_16874);
xor U17481 (N_17481,N_16960,N_16514);
nand U17482 (N_17482,N_16806,N_16521);
or U17483 (N_17483,N_16693,N_16856);
or U17484 (N_17484,N_16997,N_16519);
or U17485 (N_17485,N_16951,N_16668);
or U17486 (N_17486,N_16963,N_16853);
or U17487 (N_17487,N_16633,N_16887);
nand U17488 (N_17488,N_16758,N_16760);
and U17489 (N_17489,N_16873,N_16623);
nand U17490 (N_17490,N_16993,N_16780);
or U17491 (N_17491,N_16643,N_16602);
xnor U17492 (N_17492,N_16918,N_16825);
nand U17493 (N_17493,N_16948,N_16537);
nand U17494 (N_17494,N_16691,N_16840);
nor U17495 (N_17495,N_16799,N_16701);
and U17496 (N_17496,N_16749,N_16664);
or U17497 (N_17497,N_16909,N_16544);
nor U17498 (N_17498,N_16945,N_16950);
and U17499 (N_17499,N_16532,N_16502);
or U17500 (N_17500,N_17078,N_17269);
nor U17501 (N_17501,N_17168,N_17325);
or U17502 (N_17502,N_17285,N_17034);
xor U17503 (N_17503,N_17341,N_17134);
and U17504 (N_17504,N_17301,N_17310);
and U17505 (N_17505,N_17473,N_17090);
or U17506 (N_17506,N_17165,N_17164);
or U17507 (N_17507,N_17131,N_17471);
nand U17508 (N_17508,N_17496,N_17457);
or U17509 (N_17509,N_17385,N_17076);
or U17510 (N_17510,N_17304,N_17235);
or U17511 (N_17511,N_17350,N_17336);
and U17512 (N_17512,N_17431,N_17262);
nor U17513 (N_17513,N_17247,N_17191);
and U17514 (N_17514,N_17458,N_17037);
xnor U17515 (N_17515,N_17383,N_17278);
xor U17516 (N_17516,N_17241,N_17053);
or U17517 (N_17517,N_17029,N_17010);
xor U17518 (N_17518,N_17342,N_17483);
and U17519 (N_17519,N_17218,N_17254);
and U17520 (N_17520,N_17358,N_17049);
nor U17521 (N_17521,N_17230,N_17048);
xnor U17522 (N_17522,N_17129,N_17020);
or U17523 (N_17523,N_17347,N_17410);
or U17524 (N_17524,N_17246,N_17427);
nor U17525 (N_17525,N_17374,N_17356);
xor U17526 (N_17526,N_17038,N_17467);
nor U17527 (N_17527,N_17245,N_17368);
nor U17528 (N_17528,N_17450,N_17058);
nor U17529 (N_17529,N_17415,N_17080);
and U17530 (N_17530,N_17276,N_17443);
nand U17531 (N_17531,N_17302,N_17295);
or U17532 (N_17532,N_17171,N_17217);
and U17533 (N_17533,N_17343,N_17184);
nand U17534 (N_17534,N_17127,N_17194);
or U17535 (N_17535,N_17101,N_17202);
and U17536 (N_17536,N_17114,N_17242);
xnor U17537 (N_17537,N_17142,N_17210);
or U17538 (N_17538,N_17287,N_17154);
nor U17539 (N_17539,N_17438,N_17461);
xor U17540 (N_17540,N_17050,N_17331);
nand U17541 (N_17541,N_17187,N_17209);
xnor U17542 (N_17542,N_17139,N_17157);
nor U17543 (N_17543,N_17416,N_17082);
or U17544 (N_17544,N_17063,N_17019);
and U17545 (N_17545,N_17222,N_17452);
and U17546 (N_17546,N_17201,N_17231);
xnor U17547 (N_17547,N_17261,N_17051);
xnor U17548 (N_17548,N_17266,N_17440);
and U17549 (N_17549,N_17337,N_17401);
or U17550 (N_17550,N_17024,N_17221);
nand U17551 (N_17551,N_17313,N_17229);
and U17552 (N_17552,N_17225,N_17004);
and U17553 (N_17553,N_17213,N_17015);
and U17554 (N_17554,N_17257,N_17444);
xnor U17555 (N_17555,N_17064,N_17196);
nor U17556 (N_17556,N_17095,N_17062);
xor U17557 (N_17557,N_17224,N_17378);
xnor U17558 (N_17558,N_17094,N_17039);
nand U17559 (N_17559,N_17459,N_17115);
nor U17560 (N_17560,N_17043,N_17429);
xor U17561 (N_17561,N_17435,N_17002);
or U17562 (N_17562,N_17130,N_17354);
and U17563 (N_17563,N_17409,N_17366);
nor U17564 (N_17564,N_17016,N_17248);
nor U17565 (N_17565,N_17298,N_17071);
or U17566 (N_17566,N_17036,N_17012);
xnor U17567 (N_17567,N_17267,N_17315);
or U17568 (N_17568,N_17380,N_17283);
xnor U17569 (N_17569,N_17092,N_17156);
or U17570 (N_17570,N_17441,N_17422);
and U17571 (N_17571,N_17372,N_17151);
and U17572 (N_17572,N_17279,N_17484);
and U17573 (N_17573,N_17057,N_17469);
or U17574 (N_17574,N_17203,N_17322);
or U17575 (N_17575,N_17137,N_17204);
or U17576 (N_17576,N_17085,N_17143);
or U17577 (N_17577,N_17338,N_17111);
nand U17578 (N_17578,N_17121,N_17237);
xnor U17579 (N_17579,N_17112,N_17390);
nand U17580 (N_17580,N_17316,N_17386);
or U17581 (N_17581,N_17398,N_17491);
or U17582 (N_17582,N_17182,N_17146);
and U17583 (N_17583,N_17373,N_17494);
and U17584 (N_17584,N_17055,N_17328);
nand U17585 (N_17585,N_17286,N_17096);
xor U17586 (N_17586,N_17432,N_17250);
nor U17587 (N_17587,N_17120,N_17075);
or U17588 (N_17588,N_17158,N_17258);
nand U17589 (N_17589,N_17056,N_17077);
nand U17590 (N_17590,N_17207,N_17308);
nor U17591 (N_17591,N_17288,N_17417);
and U17592 (N_17592,N_17255,N_17447);
and U17593 (N_17593,N_17348,N_17284);
nand U17594 (N_17594,N_17205,N_17044);
and U17595 (N_17595,N_17349,N_17307);
and U17596 (N_17596,N_17355,N_17321);
nand U17597 (N_17597,N_17070,N_17200);
nor U17598 (N_17598,N_17406,N_17472);
xnor U17599 (N_17599,N_17361,N_17352);
or U17600 (N_17600,N_17376,N_17296);
xnor U17601 (N_17601,N_17489,N_17499);
and U17602 (N_17602,N_17495,N_17268);
xor U17603 (N_17603,N_17228,N_17454);
and U17604 (N_17604,N_17052,N_17482);
nor U17605 (N_17605,N_17149,N_17370);
and U17606 (N_17606,N_17125,N_17180);
nand U17607 (N_17607,N_17176,N_17192);
xor U17608 (N_17608,N_17041,N_17161);
xor U17609 (N_17609,N_17403,N_17317);
nor U17610 (N_17610,N_17000,N_17303);
nor U17611 (N_17611,N_17346,N_17379);
and U17612 (N_17612,N_17323,N_17189);
and U17613 (N_17613,N_17446,N_17185);
nor U17614 (N_17614,N_17453,N_17277);
or U17615 (N_17615,N_17104,N_17018);
or U17616 (N_17616,N_17497,N_17170);
and U17617 (N_17617,N_17026,N_17272);
or U17618 (N_17618,N_17397,N_17420);
nor U17619 (N_17619,N_17419,N_17297);
nand U17620 (N_17620,N_17309,N_17177);
nor U17621 (N_17621,N_17226,N_17208);
xor U17622 (N_17622,N_17344,N_17421);
nor U17623 (N_17623,N_17271,N_17061);
and U17624 (N_17624,N_17334,N_17167);
nor U17625 (N_17625,N_17214,N_17294);
xnor U17626 (N_17626,N_17387,N_17032);
nand U17627 (N_17627,N_17381,N_17488);
nor U17628 (N_17628,N_17211,N_17088);
and U17629 (N_17629,N_17363,N_17470);
and U17630 (N_17630,N_17172,N_17033);
xnor U17631 (N_17631,N_17195,N_17364);
and U17632 (N_17632,N_17093,N_17478);
and U17633 (N_17633,N_17490,N_17147);
nor U17634 (N_17634,N_17493,N_17007);
or U17635 (N_17635,N_17253,N_17117);
and U17636 (N_17636,N_17320,N_17199);
and U17637 (N_17637,N_17227,N_17216);
or U17638 (N_17638,N_17008,N_17067);
nor U17639 (N_17639,N_17232,N_17181);
and U17640 (N_17640,N_17163,N_17155);
xnor U17641 (N_17641,N_17135,N_17219);
and U17642 (N_17642,N_17079,N_17263);
or U17643 (N_17643,N_17106,N_17109);
xor U17644 (N_17644,N_17116,N_17188);
and U17645 (N_17645,N_17332,N_17264);
nand U17646 (N_17646,N_17448,N_17396);
or U17647 (N_17647,N_17474,N_17175);
and U17648 (N_17648,N_17119,N_17353);
and U17649 (N_17649,N_17339,N_17006);
nor U17650 (N_17650,N_17244,N_17265);
nor U17651 (N_17651,N_17252,N_17141);
xnor U17652 (N_17652,N_17169,N_17423);
nand U17653 (N_17653,N_17392,N_17463);
nand U17654 (N_17654,N_17282,N_17426);
nand U17655 (N_17655,N_17148,N_17027);
nor U17656 (N_17656,N_17005,N_17351);
or U17657 (N_17657,N_17395,N_17060);
xnor U17658 (N_17658,N_17300,N_17414);
nor U17659 (N_17659,N_17233,N_17025);
xor U17660 (N_17660,N_17333,N_17260);
nand U17661 (N_17661,N_17314,N_17404);
xnor U17662 (N_17662,N_17412,N_17462);
nand U17663 (N_17663,N_17306,N_17400);
or U17664 (N_17664,N_17011,N_17305);
and U17665 (N_17665,N_17434,N_17485);
and U17666 (N_17666,N_17240,N_17273);
nand U17667 (N_17667,N_17186,N_17281);
or U17668 (N_17668,N_17152,N_17487);
or U17669 (N_17669,N_17413,N_17001);
or U17670 (N_17670,N_17212,N_17108);
or U17671 (N_17671,N_17105,N_17291);
nor U17672 (N_17672,N_17357,N_17091);
xor U17673 (N_17673,N_17206,N_17407);
and U17674 (N_17674,N_17198,N_17133);
nand U17675 (N_17675,N_17371,N_17428);
or U17676 (N_17676,N_17046,N_17031);
or U17677 (N_17677,N_17072,N_17464);
nor U17678 (N_17678,N_17477,N_17123);
nor U17679 (N_17679,N_17173,N_17359);
nand U17680 (N_17680,N_17293,N_17099);
nand U17681 (N_17681,N_17220,N_17100);
nand U17682 (N_17682,N_17292,N_17047);
or U17683 (N_17683,N_17113,N_17086);
and U17684 (N_17684,N_17081,N_17476);
xnor U17685 (N_17685,N_17022,N_17311);
nor U17686 (N_17686,N_17174,N_17160);
nand U17687 (N_17687,N_17451,N_17003);
and U17688 (N_17688,N_17367,N_17084);
and U17689 (N_17689,N_17340,N_17492);
xor U17690 (N_17690,N_17107,N_17437);
nand U17691 (N_17691,N_17394,N_17425);
or U17692 (N_17692,N_17445,N_17236);
and U17693 (N_17693,N_17399,N_17498);
xnor U17694 (N_17694,N_17249,N_17068);
or U17695 (N_17695,N_17098,N_17162);
xor U17696 (N_17696,N_17197,N_17193);
xnor U17697 (N_17697,N_17030,N_17393);
or U17698 (N_17698,N_17468,N_17330);
nor U17699 (N_17699,N_17140,N_17159);
and U17700 (N_17700,N_17382,N_17365);
and U17701 (N_17701,N_17017,N_17375);
nor U17702 (N_17702,N_17456,N_17251);
and U17703 (N_17703,N_17065,N_17054);
or U17704 (N_17704,N_17436,N_17234);
nor U17705 (N_17705,N_17256,N_17035);
or U17706 (N_17706,N_17045,N_17405);
nand U17707 (N_17707,N_17318,N_17223);
nor U17708 (N_17708,N_17360,N_17183);
or U17709 (N_17709,N_17083,N_17418);
and U17710 (N_17710,N_17299,N_17118);
nand U17711 (N_17711,N_17424,N_17097);
or U17712 (N_17712,N_17465,N_17275);
xor U17713 (N_17713,N_17132,N_17126);
or U17714 (N_17714,N_17238,N_17259);
nand U17715 (N_17715,N_17377,N_17089);
or U17716 (N_17716,N_17144,N_17215);
or U17717 (N_17717,N_17466,N_17329);
and U17718 (N_17718,N_17442,N_17369);
and U17719 (N_17719,N_17280,N_17486);
or U17720 (N_17720,N_17239,N_17074);
and U17721 (N_17721,N_17391,N_17040);
and U17722 (N_17722,N_17327,N_17480);
and U17723 (N_17723,N_17274,N_17475);
and U17724 (N_17724,N_17124,N_17319);
and U17725 (N_17725,N_17021,N_17178);
xor U17726 (N_17726,N_17430,N_17122);
or U17727 (N_17727,N_17110,N_17312);
xor U17728 (N_17728,N_17014,N_17153);
xor U17729 (N_17729,N_17166,N_17028);
nor U17730 (N_17730,N_17059,N_17479);
and U17731 (N_17731,N_17066,N_17324);
or U17732 (N_17732,N_17013,N_17270);
nand U17733 (N_17733,N_17384,N_17150);
xor U17734 (N_17734,N_17460,N_17335);
xnor U17735 (N_17735,N_17402,N_17023);
nor U17736 (N_17736,N_17073,N_17102);
nor U17737 (N_17737,N_17362,N_17009);
or U17738 (N_17738,N_17439,N_17326);
nand U17739 (N_17739,N_17449,N_17136);
nor U17740 (N_17740,N_17243,N_17138);
nor U17741 (N_17741,N_17103,N_17408);
and U17742 (N_17742,N_17455,N_17388);
or U17743 (N_17743,N_17481,N_17069);
xnor U17744 (N_17744,N_17145,N_17433);
nand U17745 (N_17745,N_17128,N_17389);
nor U17746 (N_17746,N_17190,N_17411);
or U17747 (N_17747,N_17087,N_17042);
xnor U17748 (N_17748,N_17290,N_17179);
and U17749 (N_17749,N_17345,N_17289);
nor U17750 (N_17750,N_17311,N_17471);
and U17751 (N_17751,N_17202,N_17469);
xnor U17752 (N_17752,N_17282,N_17035);
nand U17753 (N_17753,N_17499,N_17117);
nand U17754 (N_17754,N_17370,N_17277);
nand U17755 (N_17755,N_17277,N_17142);
nor U17756 (N_17756,N_17150,N_17155);
nand U17757 (N_17757,N_17073,N_17004);
xnor U17758 (N_17758,N_17188,N_17318);
and U17759 (N_17759,N_17349,N_17364);
or U17760 (N_17760,N_17456,N_17064);
and U17761 (N_17761,N_17280,N_17192);
and U17762 (N_17762,N_17052,N_17409);
nand U17763 (N_17763,N_17104,N_17026);
xnor U17764 (N_17764,N_17381,N_17258);
and U17765 (N_17765,N_17352,N_17062);
xor U17766 (N_17766,N_17449,N_17386);
and U17767 (N_17767,N_17499,N_17355);
or U17768 (N_17768,N_17353,N_17341);
nor U17769 (N_17769,N_17459,N_17181);
xor U17770 (N_17770,N_17041,N_17065);
nand U17771 (N_17771,N_17366,N_17096);
and U17772 (N_17772,N_17140,N_17102);
or U17773 (N_17773,N_17326,N_17070);
nor U17774 (N_17774,N_17115,N_17371);
nand U17775 (N_17775,N_17224,N_17314);
and U17776 (N_17776,N_17381,N_17442);
and U17777 (N_17777,N_17235,N_17379);
nor U17778 (N_17778,N_17449,N_17457);
or U17779 (N_17779,N_17357,N_17077);
and U17780 (N_17780,N_17042,N_17298);
nor U17781 (N_17781,N_17401,N_17190);
or U17782 (N_17782,N_17458,N_17372);
or U17783 (N_17783,N_17468,N_17245);
nor U17784 (N_17784,N_17208,N_17189);
and U17785 (N_17785,N_17492,N_17199);
xor U17786 (N_17786,N_17209,N_17303);
nor U17787 (N_17787,N_17211,N_17058);
xor U17788 (N_17788,N_17253,N_17027);
or U17789 (N_17789,N_17463,N_17107);
or U17790 (N_17790,N_17356,N_17133);
nand U17791 (N_17791,N_17147,N_17387);
or U17792 (N_17792,N_17007,N_17306);
or U17793 (N_17793,N_17498,N_17077);
or U17794 (N_17794,N_17152,N_17408);
nor U17795 (N_17795,N_17381,N_17387);
nor U17796 (N_17796,N_17181,N_17122);
or U17797 (N_17797,N_17002,N_17282);
xor U17798 (N_17798,N_17137,N_17277);
and U17799 (N_17799,N_17203,N_17227);
nand U17800 (N_17800,N_17432,N_17330);
nor U17801 (N_17801,N_17107,N_17223);
nor U17802 (N_17802,N_17048,N_17161);
or U17803 (N_17803,N_17248,N_17074);
and U17804 (N_17804,N_17221,N_17017);
or U17805 (N_17805,N_17216,N_17005);
xnor U17806 (N_17806,N_17355,N_17439);
or U17807 (N_17807,N_17083,N_17228);
xor U17808 (N_17808,N_17081,N_17352);
or U17809 (N_17809,N_17246,N_17419);
nor U17810 (N_17810,N_17317,N_17015);
nand U17811 (N_17811,N_17266,N_17441);
nor U17812 (N_17812,N_17315,N_17302);
and U17813 (N_17813,N_17367,N_17011);
xnor U17814 (N_17814,N_17392,N_17219);
xor U17815 (N_17815,N_17225,N_17241);
nor U17816 (N_17816,N_17292,N_17460);
or U17817 (N_17817,N_17338,N_17017);
xor U17818 (N_17818,N_17070,N_17348);
or U17819 (N_17819,N_17379,N_17369);
xnor U17820 (N_17820,N_17430,N_17109);
nor U17821 (N_17821,N_17030,N_17159);
nand U17822 (N_17822,N_17410,N_17452);
nand U17823 (N_17823,N_17360,N_17071);
nand U17824 (N_17824,N_17338,N_17136);
and U17825 (N_17825,N_17241,N_17486);
or U17826 (N_17826,N_17431,N_17141);
nor U17827 (N_17827,N_17002,N_17353);
or U17828 (N_17828,N_17013,N_17048);
or U17829 (N_17829,N_17293,N_17351);
nor U17830 (N_17830,N_17468,N_17424);
nand U17831 (N_17831,N_17300,N_17012);
or U17832 (N_17832,N_17274,N_17495);
and U17833 (N_17833,N_17215,N_17387);
xor U17834 (N_17834,N_17302,N_17084);
and U17835 (N_17835,N_17451,N_17301);
and U17836 (N_17836,N_17372,N_17351);
or U17837 (N_17837,N_17121,N_17014);
xnor U17838 (N_17838,N_17151,N_17271);
and U17839 (N_17839,N_17099,N_17025);
nor U17840 (N_17840,N_17355,N_17081);
or U17841 (N_17841,N_17388,N_17461);
or U17842 (N_17842,N_17227,N_17010);
or U17843 (N_17843,N_17084,N_17154);
nand U17844 (N_17844,N_17496,N_17448);
nand U17845 (N_17845,N_17006,N_17086);
nand U17846 (N_17846,N_17461,N_17292);
nand U17847 (N_17847,N_17133,N_17451);
and U17848 (N_17848,N_17010,N_17197);
nor U17849 (N_17849,N_17410,N_17225);
or U17850 (N_17850,N_17082,N_17361);
nor U17851 (N_17851,N_17133,N_17077);
nand U17852 (N_17852,N_17415,N_17248);
and U17853 (N_17853,N_17155,N_17362);
nand U17854 (N_17854,N_17317,N_17213);
or U17855 (N_17855,N_17163,N_17150);
nand U17856 (N_17856,N_17103,N_17039);
or U17857 (N_17857,N_17005,N_17184);
nand U17858 (N_17858,N_17435,N_17333);
nand U17859 (N_17859,N_17431,N_17307);
xor U17860 (N_17860,N_17143,N_17485);
xor U17861 (N_17861,N_17084,N_17201);
nand U17862 (N_17862,N_17421,N_17181);
and U17863 (N_17863,N_17451,N_17096);
or U17864 (N_17864,N_17290,N_17095);
nand U17865 (N_17865,N_17277,N_17340);
nand U17866 (N_17866,N_17344,N_17227);
xnor U17867 (N_17867,N_17371,N_17268);
nand U17868 (N_17868,N_17036,N_17167);
and U17869 (N_17869,N_17184,N_17118);
or U17870 (N_17870,N_17168,N_17210);
xor U17871 (N_17871,N_17041,N_17072);
nand U17872 (N_17872,N_17083,N_17239);
nor U17873 (N_17873,N_17494,N_17471);
xor U17874 (N_17874,N_17422,N_17443);
or U17875 (N_17875,N_17232,N_17498);
and U17876 (N_17876,N_17238,N_17367);
and U17877 (N_17877,N_17203,N_17014);
xor U17878 (N_17878,N_17072,N_17431);
or U17879 (N_17879,N_17208,N_17095);
nor U17880 (N_17880,N_17145,N_17321);
and U17881 (N_17881,N_17245,N_17028);
xnor U17882 (N_17882,N_17332,N_17287);
or U17883 (N_17883,N_17245,N_17403);
and U17884 (N_17884,N_17134,N_17211);
nand U17885 (N_17885,N_17215,N_17362);
and U17886 (N_17886,N_17240,N_17154);
and U17887 (N_17887,N_17474,N_17326);
xnor U17888 (N_17888,N_17150,N_17437);
and U17889 (N_17889,N_17066,N_17096);
and U17890 (N_17890,N_17478,N_17274);
xnor U17891 (N_17891,N_17088,N_17294);
nor U17892 (N_17892,N_17210,N_17469);
and U17893 (N_17893,N_17129,N_17011);
nor U17894 (N_17894,N_17377,N_17366);
nand U17895 (N_17895,N_17023,N_17297);
and U17896 (N_17896,N_17030,N_17002);
and U17897 (N_17897,N_17382,N_17127);
nand U17898 (N_17898,N_17077,N_17111);
xor U17899 (N_17899,N_17292,N_17425);
xnor U17900 (N_17900,N_17489,N_17065);
and U17901 (N_17901,N_17387,N_17466);
and U17902 (N_17902,N_17171,N_17235);
nor U17903 (N_17903,N_17097,N_17316);
and U17904 (N_17904,N_17250,N_17235);
nor U17905 (N_17905,N_17180,N_17474);
and U17906 (N_17906,N_17352,N_17426);
xor U17907 (N_17907,N_17364,N_17274);
nor U17908 (N_17908,N_17154,N_17490);
or U17909 (N_17909,N_17491,N_17114);
nor U17910 (N_17910,N_17393,N_17151);
xor U17911 (N_17911,N_17303,N_17399);
xor U17912 (N_17912,N_17037,N_17485);
or U17913 (N_17913,N_17273,N_17328);
nor U17914 (N_17914,N_17487,N_17249);
or U17915 (N_17915,N_17219,N_17149);
or U17916 (N_17916,N_17388,N_17219);
xor U17917 (N_17917,N_17074,N_17108);
xnor U17918 (N_17918,N_17192,N_17120);
or U17919 (N_17919,N_17150,N_17300);
nand U17920 (N_17920,N_17055,N_17131);
xor U17921 (N_17921,N_17273,N_17163);
xnor U17922 (N_17922,N_17183,N_17189);
nand U17923 (N_17923,N_17182,N_17030);
xnor U17924 (N_17924,N_17250,N_17089);
and U17925 (N_17925,N_17171,N_17233);
xnor U17926 (N_17926,N_17045,N_17435);
xor U17927 (N_17927,N_17253,N_17064);
xor U17928 (N_17928,N_17149,N_17244);
xnor U17929 (N_17929,N_17037,N_17117);
or U17930 (N_17930,N_17491,N_17374);
nor U17931 (N_17931,N_17254,N_17302);
nand U17932 (N_17932,N_17198,N_17038);
and U17933 (N_17933,N_17331,N_17413);
nand U17934 (N_17934,N_17227,N_17484);
xnor U17935 (N_17935,N_17369,N_17348);
nand U17936 (N_17936,N_17472,N_17010);
nor U17937 (N_17937,N_17271,N_17166);
xnor U17938 (N_17938,N_17408,N_17238);
nor U17939 (N_17939,N_17056,N_17298);
nand U17940 (N_17940,N_17453,N_17309);
and U17941 (N_17941,N_17065,N_17051);
nand U17942 (N_17942,N_17449,N_17064);
xnor U17943 (N_17943,N_17463,N_17050);
and U17944 (N_17944,N_17444,N_17322);
nor U17945 (N_17945,N_17049,N_17219);
and U17946 (N_17946,N_17094,N_17018);
xnor U17947 (N_17947,N_17116,N_17187);
nand U17948 (N_17948,N_17009,N_17294);
and U17949 (N_17949,N_17057,N_17025);
xor U17950 (N_17950,N_17278,N_17055);
nand U17951 (N_17951,N_17293,N_17483);
nor U17952 (N_17952,N_17446,N_17463);
and U17953 (N_17953,N_17251,N_17043);
and U17954 (N_17954,N_17252,N_17454);
xor U17955 (N_17955,N_17113,N_17229);
or U17956 (N_17956,N_17058,N_17011);
xnor U17957 (N_17957,N_17325,N_17285);
or U17958 (N_17958,N_17227,N_17006);
or U17959 (N_17959,N_17346,N_17099);
xnor U17960 (N_17960,N_17339,N_17440);
nor U17961 (N_17961,N_17358,N_17332);
xnor U17962 (N_17962,N_17451,N_17170);
xor U17963 (N_17963,N_17330,N_17376);
xor U17964 (N_17964,N_17320,N_17398);
or U17965 (N_17965,N_17322,N_17328);
nor U17966 (N_17966,N_17245,N_17094);
nand U17967 (N_17967,N_17290,N_17489);
or U17968 (N_17968,N_17134,N_17082);
nand U17969 (N_17969,N_17131,N_17272);
or U17970 (N_17970,N_17011,N_17479);
nor U17971 (N_17971,N_17263,N_17035);
xnor U17972 (N_17972,N_17143,N_17013);
nor U17973 (N_17973,N_17133,N_17095);
nand U17974 (N_17974,N_17255,N_17337);
nor U17975 (N_17975,N_17114,N_17289);
nand U17976 (N_17976,N_17183,N_17382);
or U17977 (N_17977,N_17002,N_17268);
nor U17978 (N_17978,N_17408,N_17042);
and U17979 (N_17979,N_17367,N_17096);
or U17980 (N_17980,N_17332,N_17457);
nor U17981 (N_17981,N_17449,N_17334);
nor U17982 (N_17982,N_17026,N_17212);
and U17983 (N_17983,N_17423,N_17226);
nand U17984 (N_17984,N_17083,N_17229);
xnor U17985 (N_17985,N_17324,N_17141);
or U17986 (N_17986,N_17262,N_17498);
or U17987 (N_17987,N_17159,N_17142);
or U17988 (N_17988,N_17370,N_17342);
nand U17989 (N_17989,N_17031,N_17155);
nand U17990 (N_17990,N_17019,N_17485);
nor U17991 (N_17991,N_17093,N_17337);
nand U17992 (N_17992,N_17093,N_17210);
nor U17993 (N_17993,N_17361,N_17395);
or U17994 (N_17994,N_17084,N_17412);
nand U17995 (N_17995,N_17119,N_17498);
nor U17996 (N_17996,N_17291,N_17464);
nand U17997 (N_17997,N_17490,N_17108);
or U17998 (N_17998,N_17081,N_17479);
xnor U17999 (N_17999,N_17354,N_17260);
nor U18000 (N_18000,N_17854,N_17579);
or U18001 (N_18001,N_17869,N_17931);
and U18002 (N_18002,N_17681,N_17734);
and U18003 (N_18003,N_17574,N_17862);
nand U18004 (N_18004,N_17843,N_17639);
or U18005 (N_18005,N_17771,N_17563);
and U18006 (N_18006,N_17654,N_17740);
nor U18007 (N_18007,N_17608,N_17956);
or U18008 (N_18008,N_17819,N_17599);
and U18009 (N_18009,N_17852,N_17850);
nand U18010 (N_18010,N_17834,N_17913);
or U18011 (N_18011,N_17925,N_17641);
nor U18012 (N_18012,N_17992,N_17618);
or U18013 (N_18013,N_17543,N_17676);
and U18014 (N_18014,N_17761,N_17742);
and U18015 (N_18015,N_17706,N_17929);
and U18016 (N_18016,N_17737,N_17841);
nand U18017 (N_18017,N_17633,N_17508);
and U18018 (N_18018,N_17610,N_17947);
or U18019 (N_18019,N_17952,N_17770);
or U18020 (N_18020,N_17711,N_17533);
nor U18021 (N_18021,N_17939,N_17612);
or U18022 (N_18022,N_17875,N_17899);
or U18023 (N_18023,N_17860,N_17648);
xor U18024 (N_18024,N_17564,N_17851);
nor U18025 (N_18025,N_17921,N_17928);
and U18026 (N_18026,N_17999,N_17754);
and U18027 (N_18027,N_17751,N_17691);
or U18028 (N_18028,N_17795,N_17876);
nand U18029 (N_18029,N_17807,N_17859);
nand U18030 (N_18030,N_17664,N_17853);
nor U18031 (N_18031,N_17526,N_17988);
nor U18032 (N_18032,N_17932,N_17958);
nor U18033 (N_18033,N_17720,N_17614);
nand U18034 (N_18034,N_17799,N_17512);
xnor U18035 (N_18035,N_17796,N_17979);
nand U18036 (N_18036,N_17987,N_17870);
or U18037 (N_18037,N_17885,N_17678);
nor U18038 (N_18038,N_17683,N_17700);
nand U18039 (N_18039,N_17809,N_17946);
or U18040 (N_18040,N_17652,N_17872);
nand U18041 (N_18041,N_17686,N_17601);
or U18042 (N_18042,N_17624,N_17553);
xnor U18043 (N_18043,N_17889,N_17840);
or U18044 (N_18044,N_17516,N_17719);
nor U18045 (N_18045,N_17730,N_17837);
or U18046 (N_18046,N_17699,N_17513);
nand U18047 (N_18047,N_17983,N_17835);
nand U18048 (N_18048,N_17715,N_17726);
nor U18049 (N_18049,N_17621,N_17708);
nand U18050 (N_18050,N_17907,N_17558);
nand U18051 (N_18051,N_17709,N_17606);
nor U18052 (N_18052,N_17504,N_17970);
or U18053 (N_18053,N_17521,N_17896);
or U18054 (N_18054,N_17758,N_17724);
nor U18055 (N_18055,N_17961,N_17856);
xor U18056 (N_18056,N_17694,N_17634);
and U18057 (N_18057,N_17857,N_17908);
and U18058 (N_18058,N_17944,N_17650);
xnor U18059 (N_18059,N_17735,N_17756);
or U18060 (N_18060,N_17917,N_17984);
nand U18061 (N_18061,N_17714,N_17600);
xnor U18062 (N_18062,N_17670,N_17888);
and U18063 (N_18063,N_17651,N_17914);
nand U18064 (N_18064,N_17747,N_17598);
or U18065 (N_18065,N_17990,N_17653);
or U18066 (N_18066,N_17702,N_17590);
and U18067 (N_18067,N_17994,N_17657);
or U18068 (N_18068,N_17717,N_17895);
nand U18069 (N_18069,N_17525,N_17948);
or U18070 (N_18070,N_17636,N_17713);
xor U18071 (N_18071,N_17530,N_17855);
nor U18072 (N_18072,N_17559,N_17844);
nor U18073 (N_18073,N_17682,N_17592);
nand U18074 (N_18074,N_17980,N_17968);
or U18075 (N_18075,N_17849,N_17620);
and U18076 (N_18076,N_17845,N_17551);
and U18077 (N_18077,N_17630,N_17707);
and U18078 (N_18078,N_17868,N_17831);
or U18079 (N_18079,N_17692,N_17560);
nand U18080 (N_18080,N_17838,N_17976);
xnor U18081 (N_18081,N_17775,N_17631);
nor U18082 (N_18082,N_17922,N_17773);
and U18083 (N_18083,N_17673,N_17514);
and U18084 (N_18084,N_17776,N_17864);
or U18085 (N_18085,N_17718,N_17605);
xnor U18086 (N_18086,N_17552,N_17915);
and U18087 (N_18087,N_17566,N_17750);
nor U18088 (N_18088,N_17873,N_17957);
nor U18089 (N_18089,N_17832,N_17541);
nand U18090 (N_18090,N_17562,N_17800);
xnor U18091 (N_18091,N_17905,N_17585);
nand U18092 (N_18092,N_17950,N_17522);
or U18093 (N_18093,N_17741,N_17898);
and U18094 (N_18094,N_17936,N_17866);
and U18095 (N_18095,N_17762,N_17536);
and U18096 (N_18096,N_17926,N_17623);
nand U18097 (N_18097,N_17812,N_17828);
nand U18098 (N_18098,N_17960,N_17632);
nand U18099 (N_18099,N_17759,N_17797);
nor U18100 (N_18100,N_17660,N_17910);
and U18101 (N_18101,N_17671,N_17723);
nand U18102 (N_18102,N_17666,N_17540);
and U18103 (N_18103,N_17802,N_17625);
and U18104 (N_18104,N_17943,N_17519);
xnor U18105 (N_18105,N_17847,N_17836);
or U18106 (N_18106,N_17535,N_17745);
nand U18107 (N_18107,N_17688,N_17981);
nor U18108 (N_18108,N_17906,N_17748);
or U18109 (N_18109,N_17953,N_17749);
xor U18110 (N_18110,N_17712,N_17767);
xor U18111 (N_18111,N_17586,N_17545);
nor U18112 (N_18112,N_17507,N_17962);
nand U18113 (N_18113,N_17959,N_17877);
and U18114 (N_18114,N_17615,N_17902);
and U18115 (N_18115,N_17509,N_17788);
nor U18116 (N_18116,N_17659,N_17611);
nor U18117 (N_18117,N_17995,N_17934);
nand U18118 (N_18118,N_17817,N_17668);
and U18119 (N_18119,N_17532,N_17774);
nand U18120 (N_18120,N_17777,N_17500);
or U18121 (N_18121,N_17893,N_17806);
and U18122 (N_18122,N_17753,N_17594);
xnor U18123 (N_18123,N_17863,N_17803);
and U18124 (N_18124,N_17768,N_17697);
or U18125 (N_18125,N_17695,N_17782);
nand U18126 (N_18126,N_17627,N_17675);
xor U18127 (N_18127,N_17635,N_17982);
or U18128 (N_18128,N_17501,N_17881);
nor U18129 (N_18129,N_17555,N_17798);
xor U18130 (N_18130,N_17821,N_17649);
and U18131 (N_18131,N_17661,N_17813);
or U18132 (N_18132,N_17705,N_17880);
nor U18133 (N_18133,N_17871,N_17546);
or U18134 (N_18134,N_17972,N_17757);
xnor U18135 (N_18135,N_17569,N_17567);
nor U18136 (N_18136,N_17531,N_17572);
and U18137 (N_18137,N_17710,N_17544);
nand U18138 (N_18138,N_17576,N_17942);
xnor U18139 (N_18139,N_17517,N_17538);
and U18140 (N_18140,N_17858,N_17728);
and U18141 (N_18141,N_17825,N_17933);
xor U18142 (N_18142,N_17698,N_17548);
and U18143 (N_18143,N_17901,N_17772);
or U18144 (N_18144,N_17674,N_17897);
and U18145 (N_18145,N_17642,N_17924);
nand U18146 (N_18146,N_17690,N_17738);
nor U18147 (N_18147,N_17619,N_17583);
and U18148 (N_18148,N_17549,N_17998);
xnor U18149 (N_18149,N_17573,N_17963);
and U18150 (N_18150,N_17556,N_17954);
nand U18151 (N_18151,N_17785,N_17892);
or U18152 (N_18152,N_17511,N_17584);
nor U18153 (N_18153,N_17811,N_17765);
and U18154 (N_18154,N_17510,N_17593);
and U18155 (N_18155,N_17539,N_17964);
or U18156 (N_18156,N_17582,N_17565);
nand U18157 (N_18157,N_17701,N_17833);
or U18158 (N_18158,N_17966,N_17945);
or U18159 (N_18159,N_17923,N_17663);
and U18160 (N_18160,N_17528,N_17989);
or U18161 (N_18161,N_17769,N_17729);
nor U18162 (N_18162,N_17703,N_17515);
and U18163 (N_18163,N_17965,N_17940);
nor U18164 (N_18164,N_17882,N_17679);
and U18165 (N_18165,N_17804,N_17829);
nor U18166 (N_18166,N_17716,N_17523);
nor U18167 (N_18167,N_17602,N_17909);
nor U18168 (N_18168,N_17746,N_17846);
or U18169 (N_18169,N_17808,N_17577);
and U18170 (N_18170,N_17779,N_17919);
and U18171 (N_18171,N_17725,N_17597);
or U18172 (N_18172,N_17554,N_17763);
or U18173 (N_18173,N_17561,N_17626);
and U18174 (N_18174,N_17722,N_17935);
nor U18175 (N_18175,N_17778,N_17638);
nand U18176 (N_18176,N_17542,N_17662);
nand U18177 (N_18177,N_17878,N_17974);
nand U18178 (N_18178,N_17822,N_17865);
and U18179 (N_18179,N_17781,N_17971);
and U18180 (N_18180,N_17684,N_17520);
and U18181 (N_18181,N_17644,N_17916);
nor U18182 (N_18182,N_17704,N_17529);
nand U18183 (N_18183,N_17884,N_17890);
nor U18184 (N_18184,N_17912,N_17733);
or U18185 (N_18185,N_17911,N_17685);
nor U18186 (N_18186,N_17793,N_17839);
xor U18187 (N_18187,N_17524,N_17887);
and U18188 (N_18188,N_17930,N_17607);
or U18189 (N_18189,N_17827,N_17830);
or U18190 (N_18190,N_17629,N_17587);
nand U18191 (N_18191,N_17588,N_17687);
and U18192 (N_18192,N_17672,N_17604);
nor U18193 (N_18193,N_17580,N_17978);
nand U18194 (N_18194,N_17640,N_17732);
nor U18195 (N_18195,N_17789,N_17680);
and U18196 (N_18196,N_17689,N_17570);
nor U18197 (N_18197,N_17886,N_17760);
xnor U18198 (N_18198,N_17903,N_17609);
xor U18199 (N_18199,N_17628,N_17967);
or U18200 (N_18200,N_17727,N_17616);
xnor U18201 (N_18201,N_17527,N_17975);
xor U18202 (N_18202,N_17792,N_17646);
and U18203 (N_18203,N_17973,N_17900);
nand U18204 (N_18204,N_17596,N_17891);
nand U18205 (N_18205,N_17883,N_17617);
and U18206 (N_18206,N_17842,N_17810);
or U18207 (N_18207,N_17787,N_17997);
nor U18208 (N_18208,N_17874,N_17815);
xor U18209 (N_18209,N_17665,N_17669);
nand U18210 (N_18210,N_17791,N_17731);
and U18211 (N_18211,N_17918,N_17667);
or U18212 (N_18212,N_17647,N_17790);
xor U18213 (N_18213,N_17996,N_17784);
xnor U18214 (N_18214,N_17658,N_17955);
xnor U18215 (N_18215,N_17693,N_17949);
and U18216 (N_18216,N_17645,N_17986);
or U18217 (N_18217,N_17991,N_17937);
xor U18218 (N_18218,N_17755,N_17938);
nor U18219 (N_18219,N_17894,N_17879);
xor U18220 (N_18220,N_17622,N_17603);
nand U18221 (N_18221,N_17656,N_17993);
nor U18222 (N_18222,N_17861,N_17848);
and U18223 (N_18223,N_17518,N_17571);
xnor U18224 (N_18224,N_17613,N_17502);
nand U18225 (N_18225,N_17820,N_17537);
nor U18226 (N_18226,N_17826,N_17786);
or U18227 (N_18227,N_17801,N_17783);
and U18228 (N_18228,N_17655,N_17739);
xnor U18229 (N_18229,N_17503,N_17818);
or U18230 (N_18230,N_17589,N_17985);
or U18231 (N_18231,N_17534,N_17547);
nand U18232 (N_18232,N_17744,N_17505);
xnor U18233 (N_18233,N_17581,N_17927);
nand U18234 (N_18234,N_17766,N_17920);
xnor U18235 (N_18235,N_17752,N_17568);
and U18236 (N_18236,N_17764,N_17696);
nand U18237 (N_18237,N_17550,N_17794);
and U18238 (N_18238,N_17867,N_17951);
nor U18239 (N_18239,N_17977,N_17969);
or U18240 (N_18240,N_17578,N_17941);
or U18241 (N_18241,N_17904,N_17677);
nand U18242 (N_18242,N_17575,N_17824);
xor U18243 (N_18243,N_17591,N_17557);
nor U18244 (N_18244,N_17721,N_17816);
or U18245 (N_18245,N_17823,N_17805);
and U18246 (N_18246,N_17595,N_17637);
and U18247 (N_18247,N_17743,N_17814);
and U18248 (N_18248,N_17506,N_17780);
or U18249 (N_18249,N_17643,N_17736);
or U18250 (N_18250,N_17948,N_17871);
nand U18251 (N_18251,N_17999,N_17785);
nand U18252 (N_18252,N_17878,N_17655);
or U18253 (N_18253,N_17731,N_17879);
or U18254 (N_18254,N_17960,N_17883);
nor U18255 (N_18255,N_17511,N_17722);
and U18256 (N_18256,N_17754,N_17751);
or U18257 (N_18257,N_17526,N_17590);
or U18258 (N_18258,N_17617,N_17582);
and U18259 (N_18259,N_17821,N_17566);
and U18260 (N_18260,N_17743,N_17847);
nor U18261 (N_18261,N_17759,N_17882);
nor U18262 (N_18262,N_17541,N_17762);
and U18263 (N_18263,N_17506,N_17816);
nand U18264 (N_18264,N_17770,N_17898);
xor U18265 (N_18265,N_17624,N_17926);
nor U18266 (N_18266,N_17612,N_17926);
or U18267 (N_18267,N_17532,N_17554);
or U18268 (N_18268,N_17708,N_17950);
and U18269 (N_18269,N_17644,N_17582);
nor U18270 (N_18270,N_17867,N_17941);
nor U18271 (N_18271,N_17576,N_17586);
or U18272 (N_18272,N_17883,N_17591);
and U18273 (N_18273,N_17600,N_17605);
or U18274 (N_18274,N_17543,N_17900);
xor U18275 (N_18275,N_17847,N_17612);
nor U18276 (N_18276,N_17840,N_17800);
or U18277 (N_18277,N_17698,N_17618);
and U18278 (N_18278,N_17623,N_17809);
and U18279 (N_18279,N_17876,N_17625);
or U18280 (N_18280,N_17607,N_17546);
xnor U18281 (N_18281,N_17815,N_17723);
or U18282 (N_18282,N_17810,N_17688);
or U18283 (N_18283,N_17659,N_17540);
and U18284 (N_18284,N_17883,N_17551);
nand U18285 (N_18285,N_17884,N_17811);
xor U18286 (N_18286,N_17666,N_17957);
nand U18287 (N_18287,N_17796,N_17593);
and U18288 (N_18288,N_17515,N_17985);
and U18289 (N_18289,N_17721,N_17672);
and U18290 (N_18290,N_17738,N_17603);
xnor U18291 (N_18291,N_17952,N_17756);
and U18292 (N_18292,N_17931,N_17944);
or U18293 (N_18293,N_17855,N_17993);
and U18294 (N_18294,N_17841,N_17782);
and U18295 (N_18295,N_17629,N_17789);
nand U18296 (N_18296,N_17916,N_17555);
and U18297 (N_18297,N_17851,N_17820);
or U18298 (N_18298,N_17796,N_17580);
nor U18299 (N_18299,N_17716,N_17652);
xnor U18300 (N_18300,N_17706,N_17590);
or U18301 (N_18301,N_17557,N_17756);
or U18302 (N_18302,N_17968,N_17666);
xor U18303 (N_18303,N_17602,N_17738);
nand U18304 (N_18304,N_17663,N_17711);
nand U18305 (N_18305,N_17998,N_17609);
xnor U18306 (N_18306,N_17989,N_17613);
and U18307 (N_18307,N_17985,N_17689);
xor U18308 (N_18308,N_17848,N_17611);
and U18309 (N_18309,N_17875,N_17792);
and U18310 (N_18310,N_17751,N_17822);
and U18311 (N_18311,N_17903,N_17737);
xor U18312 (N_18312,N_17775,N_17677);
or U18313 (N_18313,N_17530,N_17940);
xnor U18314 (N_18314,N_17614,N_17842);
nor U18315 (N_18315,N_17780,N_17508);
xnor U18316 (N_18316,N_17839,N_17996);
and U18317 (N_18317,N_17574,N_17950);
or U18318 (N_18318,N_17922,N_17735);
xor U18319 (N_18319,N_17951,N_17550);
nand U18320 (N_18320,N_17990,N_17806);
nor U18321 (N_18321,N_17932,N_17944);
nor U18322 (N_18322,N_17885,N_17854);
xnor U18323 (N_18323,N_17930,N_17551);
nand U18324 (N_18324,N_17900,N_17983);
nor U18325 (N_18325,N_17703,N_17760);
or U18326 (N_18326,N_17625,N_17905);
and U18327 (N_18327,N_17946,N_17821);
nand U18328 (N_18328,N_17545,N_17504);
and U18329 (N_18329,N_17760,N_17850);
nor U18330 (N_18330,N_17756,N_17572);
nand U18331 (N_18331,N_17898,N_17647);
nor U18332 (N_18332,N_17750,N_17556);
or U18333 (N_18333,N_17951,N_17786);
nand U18334 (N_18334,N_17898,N_17539);
and U18335 (N_18335,N_17548,N_17674);
nor U18336 (N_18336,N_17819,N_17918);
nor U18337 (N_18337,N_17610,N_17728);
nand U18338 (N_18338,N_17768,N_17614);
nor U18339 (N_18339,N_17891,N_17514);
xor U18340 (N_18340,N_17776,N_17660);
nor U18341 (N_18341,N_17690,N_17857);
or U18342 (N_18342,N_17820,N_17863);
and U18343 (N_18343,N_17916,N_17514);
or U18344 (N_18344,N_17947,N_17730);
nor U18345 (N_18345,N_17758,N_17829);
or U18346 (N_18346,N_17588,N_17711);
nor U18347 (N_18347,N_17595,N_17923);
and U18348 (N_18348,N_17665,N_17709);
nand U18349 (N_18349,N_17586,N_17989);
nor U18350 (N_18350,N_17642,N_17652);
and U18351 (N_18351,N_17992,N_17604);
or U18352 (N_18352,N_17836,N_17931);
xor U18353 (N_18353,N_17511,N_17620);
nand U18354 (N_18354,N_17924,N_17633);
nor U18355 (N_18355,N_17898,N_17849);
or U18356 (N_18356,N_17635,N_17680);
nor U18357 (N_18357,N_17507,N_17737);
nor U18358 (N_18358,N_17822,N_17544);
nor U18359 (N_18359,N_17900,N_17704);
xor U18360 (N_18360,N_17617,N_17802);
nor U18361 (N_18361,N_17977,N_17725);
nand U18362 (N_18362,N_17975,N_17596);
nor U18363 (N_18363,N_17841,N_17632);
nor U18364 (N_18364,N_17742,N_17960);
or U18365 (N_18365,N_17964,N_17721);
xnor U18366 (N_18366,N_17917,N_17961);
or U18367 (N_18367,N_17575,N_17984);
and U18368 (N_18368,N_17867,N_17943);
or U18369 (N_18369,N_17622,N_17785);
or U18370 (N_18370,N_17581,N_17671);
or U18371 (N_18371,N_17831,N_17990);
and U18372 (N_18372,N_17827,N_17584);
and U18373 (N_18373,N_17606,N_17509);
nand U18374 (N_18374,N_17653,N_17934);
and U18375 (N_18375,N_17593,N_17771);
and U18376 (N_18376,N_17653,N_17591);
or U18377 (N_18377,N_17842,N_17686);
and U18378 (N_18378,N_17653,N_17984);
or U18379 (N_18379,N_17652,N_17670);
nand U18380 (N_18380,N_17631,N_17598);
nand U18381 (N_18381,N_17953,N_17832);
nand U18382 (N_18382,N_17740,N_17595);
xnor U18383 (N_18383,N_17583,N_17865);
xnor U18384 (N_18384,N_17927,N_17651);
nor U18385 (N_18385,N_17788,N_17567);
xor U18386 (N_18386,N_17738,N_17626);
nor U18387 (N_18387,N_17833,N_17869);
nand U18388 (N_18388,N_17758,N_17764);
or U18389 (N_18389,N_17889,N_17825);
or U18390 (N_18390,N_17766,N_17690);
or U18391 (N_18391,N_17601,N_17943);
or U18392 (N_18392,N_17763,N_17759);
nor U18393 (N_18393,N_17961,N_17700);
xor U18394 (N_18394,N_17932,N_17689);
or U18395 (N_18395,N_17739,N_17972);
and U18396 (N_18396,N_17638,N_17575);
and U18397 (N_18397,N_17559,N_17940);
or U18398 (N_18398,N_17676,N_17533);
and U18399 (N_18399,N_17538,N_17530);
or U18400 (N_18400,N_17835,N_17853);
xnor U18401 (N_18401,N_17715,N_17662);
nor U18402 (N_18402,N_17897,N_17603);
or U18403 (N_18403,N_17611,N_17700);
nand U18404 (N_18404,N_17886,N_17812);
and U18405 (N_18405,N_17823,N_17758);
xor U18406 (N_18406,N_17853,N_17647);
and U18407 (N_18407,N_17902,N_17939);
xnor U18408 (N_18408,N_17554,N_17559);
or U18409 (N_18409,N_17677,N_17551);
nand U18410 (N_18410,N_17519,N_17958);
nand U18411 (N_18411,N_17836,N_17964);
and U18412 (N_18412,N_17853,N_17791);
nor U18413 (N_18413,N_17671,N_17953);
and U18414 (N_18414,N_17924,N_17623);
or U18415 (N_18415,N_17558,N_17992);
nand U18416 (N_18416,N_17785,N_17988);
nand U18417 (N_18417,N_17744,N_17995);
or U18418 (N_18418,N_17569,N_17622);
nand U18419 (N_18419,N_17996,N_17556);
xnor U18420 (N_18420,N_17985,N_17685);
nor U18421 (N_18421,N_17532,N_17612);
nand U18422 (N_18422,N_17546,N_17550);
xnor U18423 (N_18423,N_17532,N_17732);
nand U18424 (N_18424,N_17904,N_17963);
and U18425 (N_18425,N_17910,N_17677);
and U18426 (N_18426,N_17521,N_17939);
nor U18427 (N_18427,N_17791,N_17662);
xor U18428 (N_18428,N_17833,N_17664);
or U18429 (N_18429,N_17843,N_17808);
and U18430 (N_18430,N_17521,N_17536);
nand U18431 (N_18431,N_17743,N_17736);
nand U18432 (N_18432,N_17879,N_17821);
xor U18433 (N_18433,N_17663,N_17772);
or U18434 (N_18434,N_17648,N_17652);
and U18435 (N_18435,N_17542,N_17594);
or U18436 (N_18436,N_17663,N_17554);
or U18437 (N_18437,N_17837,N_17948);
nor U18438 (N_18438,N_17512,N_17962);
and U18439 (N_18439,N_17551,N_17890);
nor U18440 (N_18440,N_17769,N_17652);
xor U18441 (N_18441,N_17933,N_17712);
or U18442 (N_18442,N_17770,N_17625);
and U18443 (N_18443,N_17692,N_17844);
or U18444 (N_18444,N_17900,N_17507);
xnor U18445 (N_18445,N_17516,N_17979);
or U18446 (N_18446,N_17669,N_17809);
nand U18447 (N_18447,N_17666,N_17896);
and U18448 (N_18448,N_17806,N_17846);
xnor U18449 (N_18449,N_17852,N_17848);
nand U18450 (N_18450,N_17958,N_17594);
or U18451 (N_18451,N_17734,N_17861);
nor U18452 (N_18452,N_17679,N_17599);
or U18453 (N_18453,N_17883,N_17943);
and U18454 (N_18454,N_17826,N_17851);
and U18455 (N_18455,N_17575,N_17662);
xnor U18456 (N_18456,N_17778,N_17510);
xnor U18457 (N_18457,N_17932,N_17741);
or U18458 (N_18458,N_17922,N_17991);
or U18459 (N_18459,N_17975,N_17809);
xnor U18460 (N_18460,N_17950,N_17943);
nand U18461 (N_18461,N_17752,N_17876);
nand U18462 (N_18462,N_17604,N_17800);
or U18463 (N_18463,N_17675,N_17506);
nand U18464 (N_18464,N_17999,N_17540);
nand U18465 (N_18465,N_17944,N_17556);
or U18466 (N_18466,N_17817,N_17581);
nor U18467 (N_18467,N_17787,N_17990);
and U18468 (N_18468,N_17793,N_17936);
and U18469 (N_18469,N_17731,N_17993);
nor U18470 (N_18470,N_17986,N_17980);
nand U18471 (N_18471,N_17546,N_17503);
nand U18472 (N_18472,N_17914,N_17563);
nor U18473 (N_18473,N_17553,N_17563);
xnor U18474 (N_18474,N_17866,N_17609);
and U18475 (N_18475,N_17958,N_17866);
nor U18476 (N_18476,N_17932,N_17904);
nor U18477 (N_18477,N_17523,N_17631);
xor U18478 (N_18478,N_17619,N_17541);
xor U18479 (N_18479,N_17825,N_17537);
and U18480 (N_18480,N_17536,N_17588);
nor U18481 (N_18481,N_17699,N_17729);
and U18482 (N_18482,N_17506,N_17708);
nand U18483 (N_18483,N_17791,N_17759);
and U18484 (N_18484,N_17762,N_17654);
nor U18485 (N_18485,N_17559,N_17539);
xnor U18486 (N_18486,N_17972,N_17667);
or U18487 (N_18487,N_17530,N_17874);
or U18488 (N_18488,N_17658,N_17568);
or U18489 (N_18489,N_17696,N_17823);
and U18490 (N_18490,N_17568,N_17992);
xnor U18491 (N_18491,N_17921,N_17555);
xor U18492 (N_18492,N_17638,N_17648);
nand U18493 (N_18493,N_17797,N_17601);
nor U18494 (N_18494,N_17594,N_17814);
xor U18495 (N_18495,N_17996,N_17774);
or U18496 (N_18496,N_17675,N_17757);
nand U18497 (N_18497,N_17823,N_17522);
and U18498 (N_18498,N_17544,N_17612);
or U18499 (N_18499,N_17572,N_17838);
and U18500 (N_18500,N_18359,N_18421);
nand U18501 (N_18501,N_18459,N_18230);
nor U18502 (N_18502,N_18193,N_18494);
or U18503 (N_18503,N_18398,N_18465);
and U18504 (N_18504,N_18012,N_18029);
and U18505 (N_18505,N_18276,N_18483);
or U18506 (N_18506,N_18122,N_18091);
nor U18507 (N_18507,N_18070,N_18259);
or U18508 (N_18508,N_18019,N_18165);
nor U18509 (N_18509,N_18034,N_18128);
or U18510 (N_18510,N_18110,N_18151);
xnor U18511 (N_18511,N_18144,N_18011);
xor U18512 (N_18512,N_18094,N_18160);
and U18513 (N_18513,N_18123,N_18079);
nand U18514 (N_18514,N_18106,N_18025);
xor U18515 (N_18515,N_18493,N_18124);
or U18516 (N_18516,N_18308,N_18114);
nand U18517 (N_18517,N_18197,N_18142);
or U18518 (N_18518,N_18480,N_18407);
nand U18519 (N_18519,N_18309,N_18060);
or U18520 (N_18520,N_18280,N_18246);
and U18521 (N_18521,N_18120,N_18245);
xor U18522 (N_18522,N_18209,N_18496);
nor U18523 (N_18523,N_18254,N_18208);
nand U18524 (N_18524,N_18098,N_18044);
or U18525 (N_18525,N_18210,N_18361);
and U18526 (N_18526,N_18453,N_18214);
nor U18527 (N_18527,N_18075,N_18300);
or U18528 (N_18528,N_18267,N_18164);
or U18529 (N_18529,N_18184,N_18024);
xor U18530 (N_18530,N_18458,N_18474);
xor U18531 (N_18531,N_18454,N_18009);
and U18532 (N_18532,N_18443,N_18037);
nand U18533 (N_18533,N_18258,N_18022);
nor U18534 (N_18534,N_18190,N_18358);
nor U18535 (N_18535,N_18482,N_18220);
nor U18536 (N_18536,N_18261,N_18176);
xor U18537 (N_18537,N_18240,N_18416);
and U18538 (N_18538,N_18340,N_18158);
nand U18539 (N_18539,N_18227,N_18335);
and U18540 (N_18540,N_18048,N_18112);
nor U18541 (N_18541,N_18129,N_18385);
xor U18542 (N_18542,N_18036,N_18351);
and U18543 (N_18543,N_18005,N_18362);
xnor U18544 (N_18544,N_18279,N_18413);
nor U18545 (N_18545,N_18440,N_18139);
nor U18546 (N_18546,N_18052,N_18076);
and U18547 (N_18547,N_18017,N_18107);
nand U18548 (N_18548,N_18399,N_18326);
nand U18549 (N_18549,N_18140,N_18430);
xor U18550 (N_18550,N_18004,N_18175);
nand U18551 (N_18551,N_18379,N_18368);
nand U18552 (N_18552,N_18477,N_18093);
nand U18553 (N_18553,N_18232,N_18381);
or U18554 (N_18554,N_18272,N_18397);
nand U18555 (N_18555,N_18087,N_18305);
or U18556 (N_18556,N_18307,N_18287);
nand U18557 (N_18557,N_18263,N_18321);
xor U18558 (N_18558,N_18071,N_18242);
nand U18559 (N_18559,N_18143,N_18218);
xor U18560 (N_18560,N_18095,N_18035);
nor U18561 (N_18561,N_18334,N_18337);
nand U18562 (N_18562,N_18181,N_18378);
nor U18563 (N_18563,N_18319,N_18330);
nand U18564 (N_18564,N_18270,N_18360);
nand U18565 (N_18565,N_18391,N_18324);
xor U18566 (N_18566,N_18409,N_18366);
and U18567 (N_18567,N_18150,N_18341);
xnor U18568 (N_18568,N_18414,N_18467);
xnor U18569 (N_18569,N_18251,N_18295);
nor U18570 (N_18570,N_18006,N_18344);
nor U18571 (N_18571,N_18301,N_18406);
nand U18572 (N_18572,N_18473,N_18350);
and U18573 (N_18573,N_18073,N_18269);
and U18574 (N_18574,N_18081,N_18404);
nand U18575 (N_18575,N_18135,N_18316);
nor U18576 (N_18576,N_18283,N_18431);
xnor U18577 (N_18577,N_18105,N_18375);
and U18578 (N_18578,N_18348,N_18429);
nand U18579 (N_18579,N_18274,N_18086);
xnor U18580 (N_18580,N_18053,N_18304);
and U18581 (N_18581,N_18395,N_18322);
xor U18582 (N_18582,N_18312,N_18464);
or U18583 (N_18583,N_18339,N_18302);
and U18584 (N_18584,N_18161,N_18441);
nor U18585 (N_18585,N_18016,N_18002);
or U18586 (N_18586,N_18067,N_18329);
or U18587 (N_18587,N_18174,N_18255);
xnor U18588 (N_18588,N_18222,N_18457);
xor U18589 (N_18589,N_18207,N_18491);
nand U18590 (N_18590,N_18401,N_18061);
xnor U18591 (N_18591,N_18294,N_18394);
nor U18592 (N_18592,N_18213,N_18043);
xor U18593 (N_18593,N_18266,N_18066);
nand U18594 (N_18594,N_18058,N_18239);
nand U18595 (N_18595,N_18127,N_18231);
xor U18596 (N_18596,N_18059,N_18342);
and U18597 (N_18597,N_18063,N_18159);
nor U18598 (N_18598,N_18096,N_18487);
xnor U18599 (N_18599,N_18115,N_18108);
nand U18600 (N_18600,N_18383,N_18403);
and U18601 (N_18601,N_18198,N_18126);
or U18602 (N_18602,N_18498,N_18288);
nand U18603 (N_18603,N_18206,N_18082);
and U18604 (N_18604,N_18026,N_18187);
xor U18605 (N_18605,N_18476,N_18444);
or U18606 (N_18606,N_18237,N_18328);
nor U18607 (N_18607,N_18363,N_18196);
xnor U18608 (N_18608,N_18172,N_18439);
nor U18609 (N_18609,N_18428,N_18460);
and U18610 (N_18610,N_18417,N_18078);
nor U18611 (N_18611,N_18433,N_18296);
nor U18612 (N_18612,N_18233,N_18281);
nand U18613 (N_18613,N_18103,N_18148);
or U18614 (N_18614,N_18130,N_18185);
and U18615 (N_18615,N_18250,N_18147);
and U18616 (N_18616,N_18177,N_18492);
nor U18617 (N_18617,N_18099,N_18286);
nand U18618 (N_18618,N_18212,N_18471);
xor U18619 (N_18619,N_18027,N_18345);
nor U18620 (N_18620,N_18021,N_18040);
nor U18621 (N_18621,N_18092,N_18215);
xor U18622 (N_18622,N_18370,N_18065);
nor U18623 (N_18623,N_18020,N_18434);
xnor U18624 (N_18624,N_18396,N_18199);
nand U18625 (N_18625,N_18072,N_18303);
and U18626 (N_18626,N_18365,N_18264);
nor U18627 (N_18627,N_18064,N_18111);
nand U18628 (N_18628,N_18117,N_18014);
or U18629 (N_18629,N_18317,N_18331);
or U18630 (N_18630,N_18438,N_18008);
xor U18631 (N_18631,N_18163,N_18424);
or U18632 (N_18632,N_18188,N_18173);
nor U18633 (N_18633,N_18315,N_18380);
and U18634 (N_18634,N_18134,N_18118);
or U18635 (N_18635,N_18113,N_18262);
nand U18636 (N_18636,N_18427,N_18167);
nand U18637 (N_18637,N_18353,N_18432);
nand U18638 (N_18638,N_18412,N_18488);
xnor U18639 (N_18639,N_18179,N_18311);
or U18640 (N_18640,N_18372,N_18131);
and U18641 (N_18641,N_18408,N_18442);
xnor U18642 (N_18642,N_18224,N_18382);
xor U18643 (N_18643,N_18384,N_18320);
xor U18644 (N_18644,N_18205,N_18201);
nand U18645 (N_18645,N_18191,N_18486);
or U18646 (N_18646,N_18141,N_18074);
nand U18647 (N_18647,N_18448,N_18050);
or U18648 (N_18648,N_18223,N_18297);
xnor U18649 (N_18649,N_18485,N_18449);
xor U18650 (N_18650,N_18364,N_18244);
xnor U18651 (N_18651,N_18478,N_18354);
nand U18652 (N_18652,N_18186,N_18418);
xor U18653 (N_18653,N_18282,N_18102);
nor U18654 (N_18654,N_18475,N_18219);
and U18655 (N_18655,N_18293,N_18371);
or U18656 (N_18656,N_18265,N_18042);
xor U18657 (N_18657,N_18194,N_18292);
xnor U18658 (N_18658,N_18247,N_18195);
and U18659 (N_18659,N_18435,N_18100);
xor U18660 (N_18660,N_18470,N_18390);
nor U18661 (N_18661,N_18310,N_18425);
xor U18662 (N_18662,N_18387,N_18437);
nor U18663 (N_18663,N_18484,N_18133);
nor U18664 (N_18664,N_18277,N_18033);
nor U18665 (N_18665,N_18489,N_18271);
nand U18666 (N_18666,N_18080,N_18462);
nor U18667 (N_18667,N_18055,N_18374);
nand U18668 (N_18668,N_18388,N_18152);
xnor U18669 (N_18669,N_18400,N_18039);
and U18670 (N_18670,N_18211,N_18355);
xor U18671 (N_18671,N_18204,N_18101);
xor U18672 (N_18672,N_18285,N_18289);
nor U18673 (N_18673,N_18411,N_18146);
nor U18674 (N_18674,N_18273,N_18069);
nor U18675 (N_18675,N_18490,N_18192);
or U18676 (N_18676,N_18062,N_18162);
nor U18677 (N_18677,N_18238,N_18221);
and U18678 (N_18678,N_18253,N_18038);
xnor U18679 (N_18679,N_18479,N_18155);
or U18680 (N_18680,N_18156,N_18234);
or U18681 (N_18681,N_18137,N_18090);
xor U18682 (N_18682,N_18356,N_18125);
and U18683 (N_18683,N_18313,N_18089);
nand U18684 (N_18684,N_18386,N_18229);
xor U18685 (N_18685,N_18169,N_18119);
nor U18686 (N_18686,N_18138,N_18419);
and U18687 (N_18687,N_18000,N_18182);
xor U18688 (N_18688,N_18171,N_18389);
xor U18689 (N_18689,N_18447,N_18347);
nor U18690 (N_18690,N_18007,N_18183);
nor U18691 (N_18691,N_18466,N_18290);
xnor U18692 (N_18692,N_18249,N_18499);
and U18693 (N_18693,N_18333,N_18023);
or U18694 (N_18694,N_18497,N_18367);
and U18695 (N_18695,N_18116,N_18085);
nor U18696 (N_18696,N_18452,N_18268);
nor U18697 (N_18697,N_18084,N_18415);
and U18698 (N_18698,N_18083,N_18260);
and U18699 (N_18699,N_18015,N_18045);
xor U18700 (N_18700,N_18109,N_18291);
and U18701 (N_18701,N_18077,N_18469);
and U18702 (N_18702,N_18088,N_18166);
and U18703 (N_18703,N_18041,N_18031);
nor U18704 (N_18704,N_18001,N_18472);
nand U18705 (N_18705,N_18357,N_18299);
and U18706 (N_18706,N_18420,N_18068);
nor U18707 (N_18707,N_18243,N_18018);
nand U18708 (N_18708,N_18495,N_18189);
and U18709 (N_18709,N_18104,N_18010);
nand U18710 (N_18710,N_18323,N_18170);
and U18711 (N_18711,N_18200,N_18252);
or U18712 (N_18712,N_18047,N_18393);
xor U18713 (N_18713,N_18168,N_18373);
and U18714 (N_18714,N_18468,N_18256);
and U18715 (N_18715,N_18402,N_18450);
and U18716 (N_18716,N_18216,N_18275);
or U18717 (N_18717,N_18056,N_18013);
nor U18718 (N_18718,N_18376,N_18003);
and U18719 (N_18719,N_18180,N_18145);
or U18720 (N_18720,N_18057,N_18455);
xor U18721 (N_18721,N_18225,N_18318);
nand U18722 (N_18722,N_18257,N_18392);
xor U18723 (N_18723,N_18423,N_18306);
nor U18724 (N_18724,N_18054,N_18157);
nand U18725 (N_18725,N_18284,N_18456);
nor U18726 (N_18726,N_18178,N_18332);
or U18727 (N_18727,N_18369,N_18132);
nand U18728 (N_18728,N_18248,N_18451);
or U18729 (N_18729,N_18422,N_18236);
nor U18730 (N_18730,N_18445,N_18121);
or U18731 (N_18731,N_18377,N_18327);
and U18732 (N_18732,N_18346,N_18336);
nor U18733 (N_18733,N_18149,N_18032);
nand U18734 (N_18734,N_18049,N_18325);
or U18735 (N_18735,N_18046,N_18481);
xor U18736 (N_18736,N_18426,N_18352);
and U18737 (N_18737,N_18338,N_18410);
or U18738 (N_18738,N_18028,N_18463);
or U18739 (N_18739,N_18136,N_18051);
xor U18740 (N_18740,N_18235,N_18349);
and U18741 (N_18741,N_18153,N_18228);
nor U18742 (N_18742,N_18217,N_18154);
nor U18743 (N_18743,N_18030,N_18097);
xor U18744 (N_18744,N_18314,N_18446);
nor U18745 (N_18745,N_18436,N_18203);
and U18746 (N_18746,N_18241,N_18405);
xor U18747 (N_18747,N_18278,N_18461);
xor U18748 (N_18748,N_18298,N_18226);
xor U18749 (N_18749,N_18202,N_18343);
and U18750 (N_18750,N_18085,N_18036);
nor U18751 (N_18751,N_18386,N_18433);
nor U18752 (N_18752,N_18470,N_18173);
xor U18753 (N_18753,N_18438,N_18449);
nand U18754 (N_18754,N_18032,N_18154);
nor U18755 (N_18755,N_18266,N_18471);
xnor U18756 (N_18756,N_18247,N_18124);
nand U18757 (N_18757,N_18348,N_18162);
nor U18758 (N_18758,N_18182,N_18266);
or U18759 (N_18759,N_18304,N_18407);
or U18760 (N_18760,N_18363,N_18472);
nor U18761 (N_18761,N_18138,N_18297);
or U18762 (N_18762,N_18071,N_18328);
xor U18763 (N_18763,N_18185,N_18451);
nand U18764 (N_18764,N_18047,N_18069);
and U18765 (N_18765,N_18247,N_18291);
nor U18766 (N_18766,N_18115,N_18117);
or U18767 (N_18767,N_18412,N_18465);
and U18768 (N_18768,N_18445,N_18097);
xor U18769 (N_18769,N_18267,N_18403);
nor U18770 (N_18770,N_18307,N_18401);
nor U18771 (N_18771,N_18231,N_18495);
xnor U18772 (N_18772,N_18111,N_18079);
nor U18773 (N_18773,N_18469,N_18109);
or U18774 (N_18774,N_18079,N_18479);
xor U18775 (N_18775,N_18178,N_18453);
nor U18776 (N_18776,N_18382,N_18180);
nand U18777 (N_18777,N_18079,N_18399);
nor U18778 (N_18778,N_18353,N_18325);
and U18779 (N_18779,N_18145,N_18018);
xnor U18780 (N_18780,N_18375,N_18152);
xor U18781 (N_18781,N_18030,N_18331);
or U18782 (N_18782,N_18314,N_18454);
xnor U18783 (N_18783,N_18499,N_18430);
xor U18784 (N_18784,N_18026,N_18313);
xnor U18785 (N_18785,N_18337,N_18433);
nand U18786 (N_18786,N_18115,N_18112);
nand U18787 (N_18787,N_18223,N_18225);
nand U18788 (N_18788,N_18275,N_18295);
xor U18789 (N_18789,N_18355,N_18210);
nand U18790 (N_18790,N_18006,N_18254);
or U18791 (N_18791,N_18406,N_18434);
nand U18792 (N_18792,N_18325,N_18244);
nor U18793 (N_18793,N_18151,N_18387);
nor U18794 (N_18794,N_18171,N_18045);
and U18795 (N_18795,N_18467,N_18181);
nand U18796 (N_18796,N_18384,N_18452);
nand U18797 (N_18797,N_18280,N_18249);
nand U18798 (N_18798,N_18463,N_18002);
nor U18799 (N_18799,N_18376,N_18091);
nor U18800 (N_18800,N_18443,N_18253);
xor U18801 (N_18801,N_18010,N_18336);
xor U18802 (N_18802,N_18071,N_18380);
nor U18803 (N_18803,N_18404,N_18312);
xor U18804 (N_18804,N_18402,N_18132);
xor U18805 (N_18805,N_18338,N_18024);
xor U18806 (N_18806,N_18469,N_18475);
or U18807 (N_18807,N_18159,N_18275);
and U18808 (N_18808,N_18220,N_18185);
or U18809 (N_18809,N_18432,N_18480);
nand U18810 (N_18810,N_18116,N_18349);
xor U18811 (N_18811,N_18194,N_18025);
nand U18812 (N_18812,N_18085,N_18004);
xnor U18813 (N_18813,N_18460,N_18192);
or U18814 (N_18814,N_18298,N_18255);
nor U18815 (N_18815,N_18157,N_18300);
or U18816 (N_18816,N_18425,N_18188);
nor U18817 (N_18817,N_18491,N_18271);
nor U18818 (N_18818,N_18053,N_18381);
and U18819 (N_18819,N_18118,N_18188);
nand U18820 (N_18820,N_18093,N_18157);
xor U18821 (N_18821,N_18307,N_18452);
and U18822 (N_18822,N_18364,N_18012);
or U18823 (N_18823,N_18250,N_18299);
xnor U18824 (N_18824,N_18245,N_18032);
nor U18825 (N_18825,N_18302,N_18263);
and U18826 (N_18826,N_18366,N_18133);
nand U18827 (N_18827,N_18462,N_18124);
or U18828 (N_18828,N_18345,N_18334);
xnor U18829 (N_18829,N_18286,N_18167);
and U18830 (N_18830,N_18239,N_18145);
nor U18831 (N_18831,N_18135,N_18453);
nor U18832 (N_18832,N_18196,N_18323);
xnor U18833 (N_18833,N_18239,N_18401);
and U18834 (N_18834,N_18278,N_18172);
nor U18835 (N_18835,N_18010,N_18369);
nand U18836 (N_18836,N_18261,N_18498);
and U18837 (N_18837,N_18077,N_18132);
nor U18838 (N_18838,N_18047,N_18401);
nor U18839 (N_18839,N_18379,N_18100);
nor U18840 (N_18840,N_18466,N_18334);
nand U18841 (N_18841,N_18060,N_18155);
nand U18842 (N_18842,N_18192,N_18429);
nand U18843 (N_18843,N_18186,N_18244);
xor U18844 (N_18844,N_18432,N_18049);
xnor U18845 (N_18845,N_18146,N_18275);
xor U18846 (N_18846,N_18145,N_18088);
nand U18847 (N_18847,N_18342,N_18474);
or U18848 (N_18848,N_18098,N_18170);
or U18849 (N_18849,N_18009,N_18119);
nand U18850 (N_18850,N_18133,N_18453);
nor U18851 (N_18851,N_18056,N_18261);
or U18852 (N_18852,N_18163,N_18131);
xor U18853 (N_18853,N_18019,N_18492);
and U18854 (N_18854,N_18147,N_18071);
or U18855 (N_18855,N_18327,N_18076);
nor U18856 (N_18856,N_18413,N_18304);
nor U18857 (N_18857,N_18434,N_18129);
and U18858 (N_18858,N_18146,N_18165);
and U18859 (N_18859,N_18101,N_18231);
xor U18860 (N_18860,N_18117,N_18159);
and U18861 (N_18861,N_18424,N_18056);
nand U18862 (N_18862,N_18330,N_18458);
nand U18863 (N_18863,N_18010,N_18330);
nand U18864 (N_18864,N_18474,N_18293);
nor U18865 (N_18865,N_18255,N_18087);
nor U18866 (N_18866,N_18237,N_18404);
nand U18867 (N_18867,N_18358,N_18357);
or U18868 (N_18868,N_18180,N_18363);
xor U18869 (N_18869,N_18425,N_18348);
xnor U18870 (N_18870,N_18252,N_18324);
xor U18871 (N_18871,N_18123,N_18294);
and U18872 (N_18872,N_18282,N_18476);
or U18873 (N_18873,N_18177,N_18055);
and U18874 (N_18874,N_18384,N_18376);
nand U18875 (N_18875,N_18397,N_18317);
xor U18876 (N_18876,N_18232,N_18050);
and U18877 (N_18877,N_18071,N_18236);
nor U18878 (N_18878,N_18132,N_18485);
nor U18879 (N_18879,N_18409,N_18150);
or U18880 (N_18880,N_18016,N_18127);
or U18881 (N_18881,N_18191,N_18079);
and U18882 (N_18882,N_18197,N_18298);
or U18883 (N_18883,N_18222,N_18039);
or U18884 (N_18884,N_18449,N_18092);
or U18885 (N_18885,N_18329,N_18081);
and U18886 (N_18886,N_18140,N_18319);
nand U18887 (N_18887,N_18348,N_18439);
nor U18888 (N_18888,N_18025,N_18138);
nand U18889 (N_18889,N_18482,N_18030);
xor U18890 (N_18890,N_18131,N_18239);
xor U18891 (N_18891,N_18148,N_18461);
nand U18892 (N_18892,N_18187,N_18307);
xnor U18893 (N_18893,N_18223,N_18074);
or U18894 (N_18894,N_18094,N_18045);
nor U18895 (N_18895,N_18142,N_18003);
or U18896 (N_18896,N_18427,N_18110);
xor U18897 (N_18897,N_18315,N_18283);
nand U18898 (N_18898,N_18474,N_18251);
and U18899 (N_18899,N_18466,N_18159);
xor U18900 (N_18900,N_18471,N_18216);
nand U18901 (N_18901,N_18377,N_18245);
nand U18902 (N_18902,N_18198,N_18350);
or U18903 (N_18903,N_18124,N_18080);
nor U18904 (N_18904,N_18046,N_18065);
xnor U18905 (N_18905,N_18199,N_18494);
nor U18906 (N_18906,N_18357,N_18138);
xnor U18907 (N_18907,N_18365,N_18383);
and U18908 (N_18908,N_18142,N_18039);
nor U18909 (N_18909,N_18035,N_18279);
nor U18910 (N_18910,N_18078,N_18180);
nand U18911 (N_18911,N_18073,N_18356);
and U18912 (N_18912,N_18038,N_18310);
and U18913 (N_18913,N_18029,N_18225);
xor U18914 (N_18914,N_18179,N_18116);
nand U18915 (N_18915,N_18324,N_18216);
nand U18916 (N_18916,N_18422,N_18169);
and U18917 (N_18917,N_18389,N_18073);
and U18918 (N_18918,N_18354,N_18028);
and U18919 (N_18919,N_18285,N_18151);
xor U18920 (N_18920,N_18402,N_18272);
or U18921 (N_18921,N_18333,N_18051);
and U18922 (N_18922,N_18185,N_18318);
nor U18923 (N_18923,N_18475,N_18419);
nand U18924 (N_18924,N_18298,N_18081);
and U18925 (N_18925,N_18092,N_18083);
and U18926 (N_18926,N_18457,N_18006);
or U18927 (N_18927,N_18316,N_18172);
nor U18928 (N_18928,N_18376,N_18067);
and U18929 (N_18929,N_18147,N_18127);
xnor U18930 (N_18930,N_18157,N_18166);
or U18931 (N_18931,N_18213,N_18064);
nor U18932 (N_18932,N_18177,N_18451);
nor U18933 (N_18933,N_18362,N_18422);
nand U18934 (N_18934,N_18490,N_18005);
xor U18935 (N_18935,N_18162,N_18285);
nand U18936 (N_18936,N_18448,N_18386);
or U18937 (N_18937,N_18263,N_18129);
nor U18938 (N_18938,N_18321,N_18431);
or U18939 (N_18939,N_18413,N_18442);
nor U18940 (N_18940,N_18113,N_18188);
xor U18941 (N_18941,N_18127,N_18124);
xnor U18942 (N_18942,N_18151,N_18235);
or U18943 (N_18943,N_18192,N_18098);
nand U18944 (N_18944,N_18076,N_18244);
or U18945 (N_18945,N_18295,N_18148);
nor U18946 (N_18946,N_18128,N_18495);
and U18947 (N_18947,N_18309,N_18038);
xor U18948 (N_18948,N_18016,N_18241);
nor U18949 (N_18949,N_18453,N_18340);
nor U18950 (N_18950,N_18308,N_18280);
nand U18951 (N_18951,N_18008,N_18387);
nand U18952 (N_18952,N_18022,N_18372);
nor U18953 (N_18953,N_18055,N_18101);
nand U18954 (N_18954,N_18405,N_18114);
or U18955 (N_18955,N_18224,N_18026);
or U18956 (N_18956,N_18051,N_18340);
xnor U18957 (N_18957,N_18421,N_18031);
and U18958 (N_18958,N_18003,N_18073);
and U18959 (N_18959,N_18347,N_18062);
xnor U18960 (N_18960,N_18103,N_18318);
or U18961 (N_18961,N_18179,N_18412);
or U18962 (N_18962,N_18435,N_18091);
xor U18963 (N_18963,N_18203,N_18111);
nand U18964 (N_18964,N_18302,N_18066);
nor U18965 (N_18965,N_18490,N_18336);
xor U18966 (N_18966,N_18422,N_18125);
or U18967 (N_18967,N_18142,N_18005);
nand U18968 (N_18968,N_18363,N_18177);
nand U18969 (N_18969,N_18329,N_18147);
xnor U18970 (N_18970,N_18497,N_18203);
and U18971 (N_18971,N_18089,N_18197);
and U18972 (N_18972,N_18262,N_18425);
nand U18973 (N_18973,N_18340,N_18037);
or U18974 (N_18974,N_18214,N_18038);
or U18975 (N_18975,N_18094,N_18210);
nand U18976 (N_18976,N_18118,N_18408);
nor U18977 (N_18977,N_18453,N_18099);
nor U18978 (N_18978,N_18194,N_18080);
nor U18979 (N_18979,N_18431,N_18113);
nand U18980 (N_18980,N_18104,N_18065);
or U18981 (N_18981,N_18431,N_18377);
nand U18982 (N_18982,N_18405,N_18079);
xor U18983 (N_18983,N_18279,N_18088);
and U18984 (N_18984,N_18142,N_18420);
nor U18985 (N_18985,N_18403,N_18415);
nand U18986 (N_18986,N_18017,N_18019);
and U18987 (N_18987,N_18017,N_18247);
xnor U18988 (N_18988,N_18380,N_18393);
xnor U18989 (N_18989,N_18186,N_18068);
nor U18990 (N_18990,N_18015,N_18200);
nand U18991 (N_18991,N_18234,N_18159);
and U18992 (N_18992,N_18381,N_18451);
xnor U18993 (N_18993,N_18266,N_18092);
and U18994 (N_18994,N_18392,N_18023);
or U18995 (N_18995,N_18337,N_18116);
nor U18996 (N_18996,N_18239,N_18263);
or U18997 (N_18997,N_18352,N_18129);
or U18998 (N_18998,N_18393,N_18196);
nand U18999 (N_18999,N_18461,N_18421);
or U19000 (N_19000,N_18956,N_18938);
or U19001 (N_19001,N_18958,N_18627);
nand U19002 (N_19002,N_18661,N_18903);
or U19003 (N_19003,N_18794,N_18869);
or U19004 (N_19004,N_18749,N_18633);
or U19005 (N_19005,N_18930,N_18970);
xor U19006 (N_19006,N_18675,N_18734);
and U19007 (N_19007,N_18888,N_18584);
and U19008 (N_19008,N_18978,N_18530);
nand U19009 (N_19009,N_18981,N_18542);
xor U19010 (N_19010,N_18748,N_18580);
nand U19011 (N_19011,N_18630,N_18901);
or U19012 (N_19012,N_18613,N_18925);
or U19013 (N_19013,N_18685,N_18744);
nand U19014 (N_19014,N_18880,N_18800);
or U19015 (N_19015,N_18691,N_18550);
nor U19016 (N_19016,N_18861,N_18926);
xor U19017 (N_19017,N_18902,N_18558);
nor U19018 (N_19018,N_18750,N_18563);
nand U19019 (N_19019,N_18738,N_18731);
or U19020 (N_19020,N_18673,N_18910);
nor U19021 (N_19021,N_18585,N_18789);
nor U19022 (N_19022,N_18747,N_18737);
nor U19023 (N_19023,N_18727,N_18988);
xor U19024 (N_19024,N_18877,N_18569);
and U19025 (N_19025,N_18672,N_18856);
xor U19026 (N_19026,N_18649,N_18959);
or U19027 (N_19027,N_18500,N_18610);
and U19028 (N_19028,N_18532,N_18946);
xnor U19029 (N_19029,N_18803,N_18527);
or U19030 (N_19030,N_18729,N_18684);
xnor U19031 (N_19031,N_18928,N_18617);
and U19032 (N_19032,N_18984,N_18881);
xnor U19033 (N_19033,N_18813,N_18689);
nor U19034 (N_19034,N_18581,N_18574);
and U19035 (N_19035,N_18885,N_18510);
nand U19036 (N_19036,N_18785,N_18908);
or U19037 (N_19037,N_18882,N_18784);
xnor U19038 (N_19038,N_18577,N_18915);
nor U19039 (N_19039,N_18918,N_18892);
and U19040 (N_19040,N_18551,N_18890);
or U19041 (N_19041,N_18690,N_18507);
nor U19042 (N_19042,N_18629,N_18643);
nor U19043 (N_19043,N_18963,N_18600);
xor U19044 (N_19044,N_18625,N_18674);
and U19045 (N_19045,N_18611,N_18695);
or U19046 (N_19046,N_18536,N_18945);
and U19047 (N_19047,N_18982,N_18607);
xor U19048 (N_19048,N_18855,N_18572);
nor U19049 (N_19049,N_18835,N_18664);
nor U19050 (N_19050,N_18904,N_18503);
nand U19051 (N_19051,N_18848,N_18917);
or U19052 (N_19052,N_18752,N_18667);
and U19053 (N_19053,N_18557,N_18893);
nor U19054 (N_19054,N_18829,N_18628);
nand U19055 (N_19055,N_18966,N_18823);
or U19056 (N_19056,N_18780,N_18875);
or U19057 (N_19057,N_18548,N_18941);
xor U19058 (N_19058,N_18758,N_18878);
and U19059 (N_19059,N_18570,N_18701);
or U19060 (N_19060,N_18555,N_18773);
or U19061 (N_19061,N_18631,N_18936);
nor U19062 (N_19062,N_18740,N_18726);
xnor U19063 (N_19063,N_18797,N_18920);
nor U19064 (N_19064,N_18509,N_18900);
xnor U19065 (N_19065,N_18652,N_18775);
or U19066 (N_19066,N_18967,N_18522);
xnor U19067 (N_19067,N_18772,N_18670);
xnor U19068 (N_19068,N_18896,N_18801);
and U19069 (N_19069,N_18683,N_18994);
xor U19070 (N_19070,N_18924,N_18779);
and U19071 (N_19071,N_18699,N_18634);
nor U19072 (N_19072,N_18663,N_18646);
or U19073 (N_19073,N_18912,N_18921);
and U19074 (N_19074,N_18537,N_18682);
nand U19075 (N_19075,N_18874,N_18680);
nor U19076 (N_19076,N_18565,N_18761);
nor U19077 (N_19077,N_18931,N_18608);
and U19078 (N_19078,N_18647,N_18521);
and U19079 (N_19079,N_18913,N_18907);
nand U19080 (N_19080,N_18582,N_18826);
nor U19081 (N_19081,N_18753,N_18567);
and U19082 (N_19082,N_18944,N_18774);
nor U19083 (N_19083,N_18865,N_18899);
and U19084 (N_19084,N_18711,N_18622);
xnor U19085 (N_19085,N_18820,N_18626);
and U19086 (N_19086,N_18762,N_18668);
nand U19087 (N_19087,N_18817,N_18722);
and U19088 (N_19088,N_18725,N_18976);
xnor U19089 (N_19089,N_18755,N_18515);
nor U19090 (N_19090,N_18937,N_18854);
or U19091 (N_19091,N_18995,N_18886);
and U19092 (N_19092,N_18942,N_18528);
nor U19093 (N_19093,N_18905,N_18706);
xor U19094 (N_19094,N_18589,N_18703);
xnor U19095 (N_19095,N_18843,N_18642);
nor U19096 (N_19096,N_18853,N_18822);
nor U19097 (N_19097,N_18952,N_18524);
xnor U19098 (N_19098,N_18810,N_18662);
xnor U19099 (N_19099,N_18992,N_18681);
nand U19100 (N_19100,N_18836,N_18825);
and U19101 (N_19101,N_18506,N_18766);
nor U19102 (N_19102,N_18788,N_18897);
xnor U19103 (N_19103,N_18732,N_18957);
nand U19104 (N_19104,N_18980,N_18929);
nor U19105 (N_19105,N_18940,N_18791);
xor U19106 (N_19106,N_18720,N_18769);
nand U19107 (N_19107,N_18669,N_18623);
xor U19108 (N_19108,N_18827,N_18741);
nor U19109 (N_19109,N_18594,N_18559);
or U19110 (N_19110,N_18989,N_18760);
nand U19111 (N_19111,N_18841,N_18786);
nor U19112 (N_19112,N_18949,N_18964);
nor U19113 (N_19113,N_18847,N_18534);
nand U19114 (N_19114,N_18891,N_18838);
nand U19115 (N_19115,N_18651,N_18955);
xor U19116 (N_19116,N_18696,N_18612);
or U19117 (N_19117,N_18714,N_18776);
nand U19118 (N_19118,N_18806,N_18543);
xor U19119 (N_19119,N_18873,N_18832);
or U19120 (N_19120,N_18606,N_18638);
or U19121 (N_19121,N_18974,N_18533);
nor U19122 (N_19122,N_18933,N_18860);
or U19123 (N_19123,N_18849,N_18516);
or U19124 (N_19124,N_18615,N_18590);
nand U19125 (N_19125,N_18636,N_18824);
and U19126 (N_19126,N_18644,N_18923);
nor U19127 (N_19127,N_18592,N_18561);
xor U19128 (N_19128,N_18987,N_18520);
xnor U19129 (N_19129,N_18764,N_18721);
xor U19130 (N_19130,N_18811,N_18887);
nor U19131 (N_19131,N_18588,N_18807);
xor U19132 (N_19132,N_18906,N_18951);
or U19133 (N_19133,N_18916,N_18990);
and U19134 (N_19134,N_18517,N_18919);
xnor U19135 (N_19135,N_18717,N_18932);
nand U19136 (N_19136,N_18724,N_18778);
nor U19137 (N_19137,N_18637,N_18743);
xnor U19138 (N_19138,N_18914,N_18553);
and U19139 (N_19139,N_18809,N_18851);
nor U19140 (N_19140,N_18660,N_18770);
xor U19141 (N_19141,N_18983,N_18993);
nor U19142 (N_19142,N_18739,N_18834);
or U19143 (N_19143,N_18546,N_18979);
nor U19144 (N_19144,N_18697,N_18519);
nand U19145 (N_19145,N_18889,N_18692);
nor U19146 (N_19146,N_18895,N_18568);
xnor U19147 (N_19147,N_18996,N_18560);
nor U19148 (N_19148,N_18969,N_18604);
nor U19149 (N_19149,N_18547,N_18705);
and U19150 (N_19150,N_18704,N_18716);
or U19151 (N_19151,N_18531,N_18818);
and U19152 (N_19152,N_18525,N_18977);
or U19153 (N_19153,N_18894,N_18972);
nand U19154 (N_19154,N_18975,N_18635);
nand U19155 (N_19155,N_18523,N_18845);
and U19156 (N_19156,N_18998,N_18573);
xnor U19157 (N_19157,N_18624,N_18783);
and U19158 (N_19158,N_18922,N_18709);
and U19159 (N_19159,N_18618,N_18583);
or U19160 (N_19160,N_18549,N_18767);
nor U19161 (N_19161,N_18540,N_18757);
or U19162 (N_19162,N_18700,N_18962);
xnor U19163 (N_19163,N_18787,N_18965);
or U19164 (N_19164,N_18603,N_18986);
xnor U19165 (N_19165,N_18535,N_18564);
nor U19166 (N_19166,N_18934,N_18708);
and U19167 (N_19167,N_18614,N_18686);
nand U19168 (N_19168,N_18508,N_18842);
xnor U19169 (N_19169,N_18514,N_18587);
nor U19170 (N_19170,N_18768,N_18719);
or U19171 (N_19171,N_18973,N_18545);
and U19172 (N_19172,N_18609,N_18812);
nand U19173 (N_19173,N_18620,N_18883);
or U19174 (N_19174,N_18805,N_18850);
nor U19175 (N_19175,N_18911,N_18593);
or U19176 (N_19176,N_18596,N_18728);
nor U19177 (N_19177,N_18833,N_18529);
or U19178 (N_19178,N_18718,N_18698);
xor U19179 (N_19179,N_18763,N_18948);
and U19180 (N_19180,N_18552,N_18968);
and U19181 (N_19181,N_18526,N_18745);
and U19182 (N_19182,N_18601,N_18960);
nor U19183 (N_19183,N_18586,N_18971);
or U19184 (N_19184,N_18579,N_18597);
or U19185 (N_19185,N_18616,N_18777);
xnor U19186 (N_19186,N_18591,N_18950);
xnor U19187 (N_19187,N_18985,N_18864);
or U19188 (N_19188,N_18804,N_18665);
nand U19189 (N_19189,N_18713,N_18802);
nor U19190 (N_19190,N_18679,N_18751);
nor U19191 (N_19191,N_18688,N_18798);
nor U19192 (N_19192,N_18702,N_18939);
or U19193 (N_19193,N_18815,N_18867);
nor U19194 (N_19194,N_18641,N_18733);
nand U19195 (N_19195,N_18909,N_18655);
nand U19196 (N_19196,N_18640,N_18676);
or U19197 (N_19197,N_18666,N_18659);
nand U19198 (N_19198,N_18539,N_18723);
nor U19199 (N_19199,N_18879,N_18504);
or U19200 (N_19200,N_18961,N_18678);
and U19201 (N_19201,N_18793,N_18839);
xor U19202 (N_19202,N_18884,N_18671);
nor U19203 (N_19203,N_18715,N_18857);
nand U19204 (N_19204,N_18754,N_18656);
nor U19205 (N_19205,N_18599,N_18538);
and U19206 (N_19206,N_18602,N_18648);
xnor U19207 (N_19207,N_18759,N_18710);
and U19208 (N_19208,N_18677,N_18650);
nor U19209 (N_19209,N_18571,N_18866);
xor U19210 (N_19210,N_18796,N_18876);
nor U19211 (N_19211,N_18619,N_18837);
xor U19212 (N_19212,N_18771,N_18566);
nor U19213 (N_19213,N_18872,N_18870);
nand U19214 (N_19214,N_18575,N_18846);
nand U19215 (N_19215,N_18512,N_18578);
and U19216 (N_19216,N_18694,N_18999);
nor U19217 (N_19217,N_18862,N_18859);
and U19218 (N_19218,N_18595,N_18947);
and U19219 (N_19219,N_18657,N_18863);
and U19220 (N_19220,N_18799,N_18605);
nor U19221 (N_19221,N_18513,N_18953);
xnor U19222 (N_19222,N_18935,N_18621);
nand U19223 (N_19223,N_18576,N_18518);
and U19224 (N_19224,N_18782,N_18840);
nor U19225 (N_19225,N_18639,N_18556);
and U19226 (N_19226,N_18868,N_18831);
nor U19227 (N_19227,N_18654,N_18735);
or U19228 (N_19228,N_18632,N_18790);
or U19229 (N_19229,N_18687,N_18991);
and U19230 (N_19230,N_18554,N_18927);
xnor U19231 (N_19231,N_18653,N_18852);
or U19232 (N_19232,N_18746,N_18795);
and U19233 (N_19233,N_18830,N_18598);
nor U19234 (N_19234,N_18712,N_18541);
nor U19235 (N_19235,N_18693,N_18781);
nand U19236 (N_19236,N_18544,N_18943);
xor U19237 (N_19237,N_18645,N_18502);
or U19238 (N_19238,N_18819,N_18814);
or U19239 (N_19239,N_18898,N_18730);
nor U19240 (N_19240,N_18954,N_18765);
and U19241 (N_19241,N_18858,N_18511);
xnor U19242 (N_19242,N_18828,N_18844);
nor U19243 (N_19243,N_18736,N_18821);
and U19244 (N_19244,N_18816,N_18501);
nand U19245 (N_19245,N_18742,N_18756);
xor U19246 (N_19246,N_18505,N_18808);
nand U19247 (N_19247,N_18871,N_18562);
and U19248 (N_19248,N_18792,N_18707);
nand U19249 (N_19249,N_18997,N_18658);
xor U19250 (N_19250,N_18805,N_18566);
nor U19251 (N_19251,N_18611,N_18768);
xor U19252 (N_19252,N_18547,N_18986);
and U19253 (N_19253,N_18564,N_18543);
or U19254 (N_19254,N_18800,N_18599);
nor U19255 (N_19255,N_18872,N_18606);
xor U19256 (N_19256,N_18672,N_18989);
xor U19257 (N_19257,N_18935,N_18692);
or U19258 (N_19258,N_18698,N_18657);
nor U19259 (N_19259,N_18783,N_18535);
nand U19260 (N_19260,N_18799,N_18899);
xor U19261 (N_19261,N_18545,N_18585);
nor U19262 (N_19262,N_18561,N_18583);
xor U19263 (N_19263,N_18666,N_18538);
or U19264 (N_19264,N_18669,N_18725);
nor U19265 (N_19265,N_18927,N_18895);
nor U19266 (N_19266,N_18612,N_18736);
nor U19267 (N_19267,N_18919,N_18984);
or U19268 (N_19268,N_18876,N_18771);
and U19269 (N_19269,N_18532,N_18748);
xnor U19270 (N_19270,N_18830,N_18885);
or U19271 (N_19271,N_18856,N_18568);
or U19272 (N_19272,N_18616,N_18533);
nand U19273 (N_19273,N_18878,N_18914);
xor U19274 (N_19274,N_18702,N_18928);
xor U19275 (N_19275,N_18727,N_18545);
or U19276 (N_19276,N_18627,N_18916);
xnor U19277 (N_19277,N_18518,N_18624);
nor U19278 (N_19278,N_18607,N_18734);
and U19279 (N_19279,N_18836,N_18863);
and U19280 (N_19280,N_18969,N_18572);
or U19281 (N_19281,N_18902,N_18675);
and U19282 (N_19282,N_18911,N_18769);
and U19283 (N_19283,N_18625,N_18546);
and U19284 (N_19284,N_18620,N_18581);
or U19285 (N_19285,N_18839,N_18790);
nand U19286 (N_19286,N_18556,N_18946);
or U19287 (N_19287,N_18990,N_18782);
and U19288 (N_19288,N_18952,N_18608);
nor U19289 (N_19289,N_18858,N_18983);
nand U19290 (N_19290,N_18912,N_18757);
nor U19291 (N_19291,N_18724,N_18738);
nand U19292 (N_19292,N_18580,N_18860);
or U19293 (N_19293,N_18869,N_18717);
or U19294 (N_19294,N_18899,N_18617);
nor U19295 (N_19295,N_18970,N_18738);
nand U19296 (N_19296,N_18893,N_18905);
nand U19297 (N_19297,N_18822,N_18988);
nand U19298 (N_19298,N_18524,N_18622);
or U19299 (N_19299,N_18512,N_18630);
nand U19300 (N_19300,N_18611,N_18820);
xor U19301 (N_19301,N_18913,N_18884);
or U19302 (N_19302,N_18568,N_18517);
xor U19303 (N_19303,N_18849,N_18583);
and U19304 (N_19304,N_18524,N_18506);
or U19305 (N_19305,N_18857,N_18733);
nor U19306 (N_19306,N_18990,N_18840);
and U19307 (N_19307,N_18917,N_18538);
or U19308 (N_19308,N_18819,N_18541);
nor U19309 (N_19309,N_18763,N_18593);
or U19310 (N_19310,N_18699,N_18592);
nor U19311 (N_19311,N_18598,N_18612);
or U19312 (N_19312,N_18653,N_18562);
and U19313 (N_19313,N_18979,N_18720);
nand U19314 (N_19314,N_18873,N_18772);
xnor U19315 (N_19315,N_18516,N_18688);
or U19316 (N_19316,N_18773,N_18865);
xnor U19317 (N_19317,N_18933,N_18833);
nand U19318 (N_19318,N_18546,N_18629);
xor U19319 (N_19319,N_18639,N_18792);
nor U19320 (N_19320,N_18653,N_18750);
nor U19321 (N_19321,N_18781,N_18811);
or U19322 (N_19322,N_18981,N_18694);
nand U19323 (N_19323,N_18626,N_18760);
and U19324 (N_19324,N_18826,N_18778);
xnor U19325 (N_19325,N_18998,N_18798);
xor U19326 (N_19326,N_18869,N_18501);
nor U19327 (N_19327,N_18908,N_18521);
nor U19328 (N_19328,N_18681,N_18684);
and U19329 (N_19329,N_18524,N_18557);
nor U19330 (N_19330,N_18629,N_18709);
and U19331 (N_19331,N_18880,N_18515);
nor U19332 (N_19332,N_18708,N_18909);
and U19333 (N_19333,N_18716,N_18573);
or U19334 (N_19334,N_18608,N_18896);
xnor U19335 (N_19335,N_18805,N_18705);
nor U19336 (N_19336,N_18772,N_18717);
nand U19337 (N_19337,N_18939,N_18844);
xor U19338 (N_19338,N_18951,N_18910);
xnor U19339 (N_19339,N_18646,N_18860);
nand U19340 (N_19340,N_18835,N_18520);
xor U19341 (N_19341,N_18745,N_18984);
and U19342 (N_19342,N_18840,N_18741);
or U19343 (N_19343,N_18864,N_18920);
and U19344 (N_19344,N_18621,N_18879);
or U19345 (N_19345,N_18584,N_18718);
and U19346 (N_19346,N_18602,N_18502);
or U19347 (N_19347,N_18639,N_18893);
xor U19348 (N_19348,N_18508,N_18560);
nand U19349 (N_19349,N_18831,N_18788);
xor U19350 (N_19350,N_18747,N_18814);
xor U19351 (N_19351,N_18594,N_18843);
xnor U19352 (N_19352,N_18880,N_18731);
nand U19353 (N_19353,N_18613,N_18697);
nor U19354 (N_19354,N_18987,N_18939);
nand U19355 (N_19355,N_18905,N_18599);
and U19356 (N_19356,N_18585,N_18561);
nand U19357 (N_19357,N_18930,N_18858);
nor U19358 (N_19358,N_18945,N_18676);
and U19359 (N_19359,N_18516,N_18812);
nor U19360 (N_19360,N_18797,N_18953);
and U19361 (N_19361,N_18858,N_18746);
nor U19362 (N_19362,N_18867,N_18786);
nor U19363 (N_19363,N_18913,N_18516);
xor U19364 (N_19364,N_18862,N_18544);
or U19365 (N_19365,N_18735,N_18653);
and U19366 (N_19366,N_18504,N_18567);
xnor U19367 (N_19367,N_18616,N_18764);
or U19368 (N_19368,N_18962,N_18819);
and U19369 (N_19369,N_18664,N_18799);
xnor U19370 (N_19370,N_18768,N_18635);
xnor U19371 (N_19371,N_18913,N_18773);
nor U19372 (N_19372,N_18664,N_18880);
or U19373 (N_19373,N_18876,N_18648);
nor U19374 (N_19374,N_18594,N_18905);
nand U19375 (N_19375,N_18589,N_18777);
nand U19376 (N_19376,N_18716,N_18571);
xnor U19377 (N_19377,N_18882,N_18621);
nor U19378 (N_19378,N_18701,N_18962);
xnor U19379 (N_19379,N_18508,N_18628);
nand U19380 (N_19380,N_18756,N_18839);
nand U19381 (N_19381,N_18904,N_18944);
or U19382 (N_19382,N_18943,N_18815);
xnor U19383 (N_19383,N_18609,N_18830);
or U19384 (N_19384,N_18694,N_18937);
or U19385 (N_19385,N_18531,N_18897);
nor U19386 (N_19386,N_18623,N_18570);
nand U19387 (N_19387,N_18933,N_18920);
and U19388 (N_19388,N_18537,N_18582);
xnor U19389 (N_19389,N_18807,N_18960);
or U19390 (N_19390,N_18985,N_18953);
and U19391 (N_19391,N_18759,N_18711);
or U19392 (N_19392,N_18955,N_18831);
and U19393 (N_19393,N_18866,N_18850);
xnor U19394 (N_19394,N_18672,N_18653);
nor U19395 (N_19395,N_18507,N_18817);
xor U19396 (N_19396,N_18907,N_18953);
nor U19397 (N_19397,N_18887,N_18951);
or U19398 (N_19398,N_18938,N_18631);
nor U19399 (N_19399,N_18639,N_18803);
nor U19400 (N_19400,N_18731,N_18584);
nor U19401 (N_19401,N_18702,N_18539);
or U19402 (N_19402,N_18789,N_18516);
nand U19403 (N_19403,N_18549,N_18564);
and U19404 (N_19404,N_18679,N_18674);
xnor U19405 (N_19405,N_18752,N_18978);
xnor U19406 (N_19406,N_18569,N_18857);
and U19407 (N_19407,N_18743,N_18663);
nor U19408 (N_19408,N_18896,N_18506);
nand U19409 (N_19409,N_18620,N_18724);
or U19410 (N_19410,N_18558,N_18671);
and U19411 (N_19411,N_18818,N_18601);
nand U19412 (N_19412,N_18973,N_18924);
nand U19413 (N_19413,N_18993,N_18663);
nand U19414 (N_19414,N_18580,N_18979);
nor U19415 (N_19415,N_18591,N_18988);
xnor U19416 (N_19416,N_18742,N_18908);
nand U19417 (N_19417,N_18738,N_18614);
and U19418 (N_19418,N_18747,N_18569);
or U19419 (N_19419,N_18545,N_18618);
nand U19420 (N_19420,N_18655,N_18931);
and U19421 (N_19421,N_18625,N_18680);
nor U19422 (N_19422,N_18731,N_18744);
nor U19423 (N_19423,N_18614,N_18587);
or U19424 (N_19424,N_18756,N_18829);
and U19425 (N_19425,N_18932,N_18706);
nor U19426 (N_19426,N_18877,N_18940);
and U19427 (N_19427,N_18649,N_18749);
xnor U19428 (N_19428,N_18970,N_18647);
xor U19429 (N_19429,N_18768,N_18625);
nor U19430 (N_19430,N_18751,N_18547);
or U19431 (N_19431,N_18668,N_18916);
or U19432 (N_19432,N_18684,N_18664);
and U19433 (N_19433,N_18924,N_18939);
nand U19434 (N_19434,N_18806,N_18890);
and U19435 (N_19435,N_18523,N_18869);
or U19436 (N_19436,N_18867,N_18720);
or U19437 (N_19437,N_18800,N_18520);
xnor U19438 (N_19438,N_18876,N_18906);
nor U19439 (N_19439,N_18935,N_18786);
xor U19440 (N_19440,N_18567,N_18871);
or U19441 (N_19441,N_18931,N_18967);
nand U19442 (N_19442,N_18640,N_18721);
xor U19443 (N_19443,N_18561,N_18551);
and U19444 (N_19444,N_18757,N_18684);
or U19445 (N_19445,N_18642,N_18998);
nand U19446 (N_19446,N_18654,N_18685);
xor U19447 (N_19447,N_18589,N_18732);
nand U19448 (N_19448,N_18531,N_18750);
nand U19449 (N_19449,N_18583,N_18902);
nand U19450 (N_19450,N_18980,N_18727);
and U19451 (N_19451,N_18825,N_18896);
and U19452 (N_19452,N_18684,N_18979);
nor U19453 (N_19453,N_18649,N_18914);
and U19454 (N_19454,N_18994,N_18945);
and U19455 (N_19455,N_18948,N_18683);
nor U19456 (N_19456,N_18882,N_18542);
nand U19457 (N_19457,N_18845,N_18723);
xnor U19458 (N_19458,N_18859,N_18991);
xnor U19459 (N_19459,N_18654,N_18728);
and U19460 (N_19460,N_18585,N_18912);
or U19461 (N_19461,N_18818,N_18931);
nand U19462 (N_19462,N_18706,N_18748);
or U19463 (N_19463,N_18735,N_18815);
nor U19464 (N_19464,N_18503,N_18854);
nor U19465 (N_19465,N_18686,N_18823);
xor U19466 (N_19466,N_18626,N_18694);
xor U19467 (N_19467,N_18970,N_18702);
nand U19468 (N_19468,N_18971,N_18604);
nand U19469 (N_19469,N_18810,N_18536);
xnor U19470 (N_19470,N_18899,N_18876);
nor U19471 (N_19471,N_18771,N_18971);
and U19472 (N_19472,N_18985,N_18944);
and U19473 (N_19473,N_18867,N_18882);
xor U19474 (N_19474,N_18763,N_18701);
and U19475 (N_19475,N_18865,N_18513);
nand U19476 (N_19476,N_18508,N_18911);
and U19477 (N_19477,N_18986,N_18725);
xor U19478 (N_19478,N_18545,N_18795);
xor U19479 (N_19479,N_18513,N_18715);
and U19480 (N_19480,N_18915,N_18679);
nand U19481 (N_19481,N_18591,N_18616);
nor U19482 (N_19482,N_18919,N_18862);
or U19483 (N_19483,N_18832,N_18631);
or U19484 (N_19484,N_18989,N_18695);
xnor U19485 (N_19485,N_18675,N_18663);
nor U19486 (N_19486,N_18726,N_18948);
nand U19487 (N_19487,N_18754,N_18581);
nand U19488 (N_19488,N_18904,N_18902);
and U19489 (N_19489,N_18940,N_18833);
or U19490 (N_19490,N_18571,N_18925);
nand U19491 (N_19491,N_18654,N_18964);
and U19492 (N_19492,N_18788,N_18860);
and U19493 (N_19493,N_18870,N_18605);
xnor U19494 (N_19494,N_18679,N_18932);
nor U19495 (N_19495,N_18911,N_18546);
or U19496 (N_19496,N_18621,N_18573);
nand U19497 (N_19497,N_18525,N_18846);
nand U19498 (N_19498,N_18984,N_18702);
xor U19499 (N_19499,N_18790,N_18989);
or U19500 (N_19500,N_19313,N_19338);
nor U19501 (N_19501,N_19054,N_19112);
or U19502 (N_19502,N_19439,N_19470);
xnor U19503 (N_19503,N_19438,N_19312);
nor U19504 (N_19504,N_19225,N_19076);
nand U19505 (N_19505,N_19375,N_19094);
or U19506 (N_19506,N_19431,N_19302);
nand U19507 (N_19507,N_19473,N_19210);
or U19508 (N_19508,N_19046,N_19056);
nand U19509 (N_19509,N_19357,N_19218);
xor U19510 (N_19510,N_19186,N_19150);
nand U19511 (N_19511,N_19477,N_19257);
xor U19512 (N_19512,N_19039,N_19194);
and U19513 (N_19513,N_19295,N_19195);
xnor U19514 (N_19514,N_19367,N_19396);
and U19515 (N_19515,N_19403,N_19486);
nand U19516 (N_19516,N_19081,N_19024);
and U19517 (N_19517,N_19131,N_19065);
nor U19518 (N_19518,N_19219,N_19404);
xor U19519 (N_19519,N_19304,N_19258);
nor U19520 (N_19520,N_19422,N_19037);
and U19521 (N_19521,N_19060,N_19467);
nand U19522 (N_19522,N_19482,N_19251);
nor U19523 (N_19523,N_19173,N_19216);
nor U19524 (N_19524,N_19018,N_19346);
xnor U19525 (N_19525,N_19306,N_19266);
or U19526 (N_19526,N_19455,N_19461);
or U19527 (N_19527,N_19248,N_19017);
nor U19528 (N_19528,N_19072,N_19007);
nand U19529 (N_19529,N_19337,N_19031);
nand U19530 (N_19530,N_19256,N_19016);
xor U19531 (N_19531,N_19179,N_19328);
nor U19532 (N_19532,N_19409,N_19005);
and U19533 (N_19533,N_19330,N_19185);
nand U19534 (N_19534,N_19062,N_19296);
and U19535 (N_19535,N_19270,N_19188);
nand U19536 (N_19536,N_19155,N_19309);
and U19537 (N_19537,N_19288,N_19325);
and U19538 (N_19538,N_19026,N_19428);
and U19539 (N_19539,N_19141,N_19310);
nor U19540 (N_19540,N_19265,N_19269);
and U19541 (N_19541,N_19279,N_19245);
and U19542 (N_19542,N_19293,N_19456);
or U19543 (N_19543,N_19014,N_19427);
xnor U19544 (N_19544,N_19490,N_19029);
xnor U19545 (N_19545,N_19169,N_19458);
and U19546 (N_19546,N_19499,N_19451);
xnor U19547 (N_19547,N_19174,N_19144);
nand U19548 (N_19548,N_19246,N_19061);
nor U19549 (N_19549,N_19154,N_19344);
nor U19550 (N_19550,N_19317,N_19229);
or U19551 (N_19551,N_19095,N_19276);
xor U19552 (N_19552,N_19290,N_19423);
xor U19553 (N_19553,N_19078,N_19469);
nor U19554 (N_19554,N_19006,N_19388);
xnor U19555 (N_19555,N_19285,N_19274);
nand U19556 (N_19556,N_19096,N_19215);
xnor U19557 (N_19557,N_19410,N_19432);
xor U19558 (N_19558,N_19091,N_19119);
or U19559 (N_19559,N_19320,N_19101);
or U19560 (N_19560,N_19275,N_19394);
xor U19561 (N_19561,N_19373,N_19097);
nand U19562 (N_19562,N_19098,N_19314);
nor U19563 (N_19563,N_19299,N_19308);
nor U19564 (N_19564,N_19377,N_19329);
xnor U19565 (N_19565,N_19381,N_19231);
xor U19566 (N_19566,N_19012,N_19408);
and U19567 (N_19567,N_19494,N_19075);
nand U19568 (N_19568,N_19391,N_19462);
nand U19569 (N_19569,N_19064,N_19379);
and U19570 (N_19570,N_19468,N_19291);
xnor U19571 (N_19571,N_19238,N_19208);
nand U19572 (N_19572,N_19497,N_19389);
xor U19573 (N_19573,N_19335,N_19387);
and U19574 (N_19574,N_19230,N_19484);
and U19575 (N_19575,N_19315,N_19492);
nor U19576 (N_19576,N_19452,N_19003);
nand U19577 (N_19577,N_19079,N_19444);
nor U19578 (N_19578,N_19134,N_19085);
and U19579 (N_19579,N_19434,N_19033);
xor U19580 (N_19580,N_19465,N_19192);
and U19581 (N_19581,N_19104,N_19298);
nor U19582 (N_19582,N_19178,N_19340);
or U19583 (N_19583,N_19413,N_19025);
xnor U19584 (N_19584,N_19415,N_19398);
nand U19585 (N_19585,N_19022,N_19083);
nor U19586 (N_19586,N_19476,N_19435);
xor U19587 (N_19587,N_19167,N_19372);
and U19588 (N_19588,N_19148,N_19264);
nand U19589 (N_19589,N_19009,N_19425);
nand U19590 (N_19590,N_19013,N_19294);
nand U19591 (N_19591,N_19202,N_19472);
and U19592 (N_19592,N_19390,N_19496);
and U19593 (N_19593,N_19201,N_19114);
nor U19594 (N_19594,N_19153,N_19177);
and U19595 (N_19595,N_19158,N_19129);
nand U19596 (N_19596,N_19287,N_19030);
nand U19597 (N_19597,N_19015,N_19135);
and U19598 (N_19598,N_19019,N_19371);
or U19599 (N_19599,N_19399,N_19401);
xor U19600 (N_19600,N_19149,N_19397);
xor U19601 (N_19601,N_19261,N_19147);
xnor U19602 (N_19602,N_19226,N_19426);
nor U19603 (N_19603,N_19175,N_19115);
or U19604 (N_19604,N_19326,N_19350);
nand U19605 (N_19605,N_19412,N_19355);
nor U19606 (N_19606,N_19368,N_19464);
and U19607 (N_19607,N_19199,N_19223);
or U19608 (N_19608,N_19289,N_19164);
nand U19609 (N_19609,N_19093,N_19204);
nor U19610 (N_19610,N_19400,N_19262);
and U19611 (N_19611,N_19385,N_19239);
nand U19612 (N_19612,N_19419,N_19190);
or U19613 (N_19613,N_19240,N_19362);
nor U19614 (N_19614,N_19145,N_19117);
xnor U19615 (N_19615,N_19331,N_19143);
nand U19616 (N_19616,N_19442,N_19366);
and U19617 (N_19617,N_19086,N_19234);
or U19618 (N_19618,N_19020,N_19139);
nand U19619 (N_19619,N_19034,N_19040);
nand U19620 (N_19620,N_19142,N_19152);
nor U19621 (N_19621,N_19004,N_19102);
nor U19622 (N_19622,N_19200,N_19235);
nand U19623 (N_19623,N_19196,N_19336);
or U19624 (N_19624,N_19332,N_19100);
nor U19625 (N_19625,N_19084,N_19352);
and U19626 (N_19626,N_19043,N_19354);
nand U19627 (N_19627,N_19303,N_19123);
and U19628 (N_19628,N_19126,N_19137);
xor U19629 (N_19629,N_19322,N_19217);
nor U19630 (N_19630,N_19417,N_19487);
or U19631 (N_19631,N_19050,N_19203);
and U19632 (N_19632,N_19171,N_19181);
or U19633 (N_19633,N_19059,N_19443);
and U19634 (N_19634,N_19446,N_19207);
or U19635 (N_19635,N_19485,N_19250);
and U19636 (N_19636,N_19369,N_19454);
nor U19637 (N_19637,N_19108,N_19133);
xnor U19638 (N_19638,N_19405,N_19478);
or U19639 (N_19639,N_19067,N_19267);
or U19640 (N_19640,N_19105,N_19323);
or U19641 (N_19641,N_19392,N_19474);
nand U19642 (N_19642,N_19182,N_19305);
and U19643 (N_19643,N_19277,N_19437);
xnor U19644 (N_19644,N_19068,N_19424);
nor U19645 (N_19645,N_19090,N_19286);
nand U19646 (N_19646,N_19316,N_19071);
nand U19647 (N_19647,N_19436,N_19023);
or U19648 (N_19648,N_19051,N_19138);
nor U19649 (N_19649,N_19271,N_19198);
xnor U19650 (N_19650,N_19342,N_19224);
nor U19651 (N_19651,N_19383,N_19341);
xor U19652 (N_19652,N_19088,N_19162);
and U19653 (N_19653,N_19421,N_19483);
and U19654 (N_19654,N_19430,N_19418);
nand U19655 (N_19655,N_19197,N_19159);
or U19656 (N_19656,N_19236,N_19318);
nand U19657 (N_19657,N_19106,N_19363);
and U19658 (N_19658,N_19211,N_19471);
xnor U19659 (N_19659,N_19376,N_19121);
nor U19660 (N_19660,N_19146,N_19089);
nand U19661 (N_19661,N_19327,N_19498);
or U19662 (N_19662,N_19120,N_19480);
and U19663 (N_19663,N_19082,N_19395);
and U19664 (N_19664,N_19053,N_19130);
or U19665 (N_19665,N_19283,N_19360);
nand U19666 (N_19666,N_19457,N_19221);
nor U19667 (N_19667,N_19281,N_19349);
and U19668 (N_19668,N_19166,N_19386);
nor U19669 (N_19669,N_19345,N_19252);
and U19670 (N_19670,N_19347,N_19011);
nor U19671 (N_19671,N_19193,N_19339);
xnor U19672 (N_19672,N_19364,N_19184);
or U19673 (N_19673,N_19021,N_19254);
or U19674 (N_19674,N_19172,N_19348);
nor U19675 (N_19675,N_19242,N_19282);
nor U19676 (N_19676,N_19365,N_19220);
xor U19677 (N_19677,N_19124,N_19228);
xnor U19678 (N_19678,N_19116,N_19370);
and U19679 (N_19679,N_19010,N_19466);
xnor U19680 (N_19680,N_19479,N_19263);
and U19681 (N_19681,N_19132,N_19488);
nor U19682 (N_19682,N_19351,N_19069);
and U19683 (N_19683,N_19393,N_19212);
nand U19684 (N_19684,N_19187,N_19002);
and U19685 (N_19685,N_19092,N_19284);
or U19686 (N_19686,N_19047,N_19247);
and U19687 (N_19687,N_19253,N_19000);
nand U19688 (N_19688,N_19268,N_19384);
nor U19689 (N_19689,N_19232,N_19045);
or U19690 (N_19690,N_19361,N_19463);
nor U19691 (N_19691,N_19440,N_19353);
nand U19692 (N_19692,N_19297,N_19300);
and U19693 (N_19693,N_19140,N_19118);
nor U19694 (N_19694,N_19481,N_19380);
xnor U19695 (N_19695,N_19170,N_19099);
and U19696 (N_19696,N_19445,N_19001);
nor U19697 (N_19697,N_19008,N_19416);
xnor U19698 (N_19698,N_19449,N_19278);
nand U19699 (N_19699,N_19382,N_19151);
nand U19700 (N_19700,N_19205,N_19087);
or U19701 (N_19701,N_19109,N_19324);
nand U19702 (N_19702,N_19049,N_19074);
nor U19703 (N_19703,N_19333,N_19191);
xnor U19704 (N_19704,N_19209,N_19110);
xnor U19705 (N_19705,N_19107,N_19493);
and U19706 (N_19706,N_19402,N_19113);
xnor U19707 (N_19707,N_19334,N_19292);
nor U19708 (N_19708,N_19259,N_19041);
xor U19709 (N_19709,N_19272,N_19168);
nor U19710 (N_19710,N_19244,N_19032);
nor U19711 (N_19711,N_19378,N_19111);
xor U19712 (N_19712,N_19280,N_19180);
xnor U19713 (N_19713,N_19495,N_19206);
or U19714 (N_19714,N_19447,N_19359);
or U19715 (N_19715,N_19183,N_19237);
or U19716 (N_19716,N_19163,N_19077);
or U19717 (N_19717,N_19358,N_19165);
xnor U19718 (N_19718,N_19214,N_19311);
xor U19719 (N_19719,N_19055,N_19255);
nand U19720 (N_19720,N_19073,N_19066);
nor U19721 (N_19721,N_19319,N_19489);
nand U19722 (N_19722,N_19420,N_19241);
nor U19723 (N_19723,N_19450,N_19156);
and U19724 (N_19724,N_19433,N_19070);
or U19725 (N_19725,N_19028,N_19122);
nor U19726 (N_19726,N_19103,N_19160);
nor U19727 (N_19727,N_19044,N_19189);
nand U19728 (N_19728,N_19035,N_19036);
xnor U19729 (N_19729,N_19057,N_19052);
and U19730 (N_19730,N_19260,N_19301);
nand U19731 (N_19731,N_19128,N_19321);
xnor U19732 (N_19732,N_19407,N_19356);
nor U19733 (N_19733,N_19406,N_19249);
nand U19734 (N_19734,N_19491,N_19161);
and U19735 (N_19735,N_19411,N_19227);
xor U19736 (N_19736,N_19374,N_19058);
nand U19737 (N_19737,N_19048,N_19063);
xnor U19738 (N_19738,N_19127,N_19222);
nand U19739 (N_19739,N_19459,N_19136);
nand U19740 (N_19740,N_19176,N_19460);
nand U19741 (N_19741,N_19080,N_19213);
nand U19742 (N_19742,N_19233,N_19448);
xor U19743 (N_19743,N_19429,N_19243);
or U19744 (N_19744,N_19273,N_19453);
nor U19745 (N_19745,N_19307,N_19475);
and U19746 (N_19746,N_19414,N_19157);
xor U19747 (N_19747,N_19441,N_19038);
xnor U19748 (N_19748,N_19027,N_19042);
and U19749 (N_19749,N_19125,N_19343);
and U19750 (N_19750,N_19285,N_19341);
xor U19751 (N_19751,N_19160,N_19282);
nor U19752 (N_19752,N_19179,N_19068);
or U19753 (N_19753,N_19125,N_19378);
or U19754 (N_19754,N_19158,N_19160);
nand U19755 (N_19755,N_19220,N_19409);
or U19756 (N_19756,N_19351,N_19342);
xnor U19757 (N_19757,N_19209,N_19350);
or U19758 (N_19758,N_19074,N_19423);
nand U19759 (N_19759,N_19434,N_19121);
xor U19760 (N_19760,N_19291,N_19202);
or U19761 (N_19761,N_19031,N_19307);
nor U19762 (N_19762,N_19151,N_19289);
and U19763 (N_19763,N_19360,N_19130);
nor U19764 (N_19764,N_19159,N_19074);
xor U19765 (N_19765,N_19469,N_19015);
nor U19766 (N_19766,N_19188,N_19444);
nand U19767 (N_19767,N_19361,N_19471);
nor U19768 (N_19768,N_19480,N_19007);
xnor U19769 (N_19769,N_19072,N_19350);
nand U19770 (N_19770,N_19155,N_19024);
or U19771 (N_19771,N_19289,N_19036);
or U19772 (N_19772,N_19398,N_19362);
nand U19773 (N_19773,N_19092,N_19479);
and U19774 (N_19774,N_19262,N_19497);
or U19775 (N_19775,N_19449,N_19419);
or U19776 (N_19776,N_19108,N_19173);
xnor U19777 (N_19777,N_19485,N_19449);
and U19778 (N_19778,N_19186,N_19246);
nor U19779 (N_19779,N_19250,N_19449);
xor U19780 (N_19780,N_19479,N_19166);
nand U19781 (N_19781,N_19138,N_19062);
or U19782 (N_19782,N_19481,N_19047);
or U19783 (N_19783,N_19279,N_19150);
xnor U19784 (N_19784,N_19336,N_19402);
nand U19785 (N_19785,N_19152,N_19375);
nand U19786 (N_19786,N_19114,N_19064);
xor U19787 (N_19787,N_19203,N_19375);
or U19788 (N_19788,N_19022,N_19173);
nand U19789 (N_19789,N_19341,N_19273);
xnor U19790 (N_19790,N_19058,N_19338);
nor U19791 (N_19791,N_19033,N_19020);
or U19792 (N_19792,N_19325,N_19084);
and U19793 (N_19793,N_19444,N_19143);
xnor U19794 (N_19794,N_19229,N_19451);
xnor U19795 (N_19795,N_19370,N_19094);
xor U19796 (N_19796,N_19298,N_19172);
and U19797 (N_19797,N_19034,N_19184);
nand U19798 (N_19798,N_19021,N_19237);
or U19799 (N_19799,N_19476,N_19032);
nor U19800 (N_19800,N_19011,N_19245);
nor U19801 (N_19801,N_19136,N_19267);
nor U19802 (N_19802,N_19273,N_19461);
or U19803 (N_19803,N_19028,N_19170);
xnor U19804 (N_19804,N_19418,N_19410);
and U19805 (N_19805,N_19291,N_19209);
or U19806 (N_19806,N_19242,N_19491);
nand U19807 (N_19807,N_19453,N_19421);
xnor U19808 (N_19808,N_19065,N_19076);
or U19809 (N_19809,N_19135,N_19157);
nor U19810 (N_19810,N_19442,N_19198);
and U19811 (N_19811,N_19176,N_19214);
nand U19812 (N_19812,N_19100,N_19417);
nand U19813 (N_19813,N_19044,N_19009);
xor U19814 (N_19814,N_19355,N_19090);
nor U19815 (N_19815,N_19466,N_19096);
and U19816 (N_19816,N_19183,N_19243);
nor U19817 (N_19817,N_19082,N_19229);
and U19818 (N_19818,N_19189,N_19343);
and U19819 (N_19819,N_19127,N_19141);
xor U19820 (N_19820,N_19332,N_19423);
nand U19821 (N_19821,N_19300,N_19070);
nand U19822 (N_19822,N_19074,N_19487);
and U19823 (N_19823,N_19183,N_19066);
nor U19824 (N_19824,N_19215,N_19451);
nor U19825 (N_19825,N_19295,N_19311);
nand U19826 (N_19826,N_19218,N_19041);
and U19827 (N_19827,N_19108,N_19459);
xor U19828 (N_19828,N_19463,N_19478);
xnor U19829 (N_19829,N_19121,N_19410);
or U19830 (N_19830,N_19004,N_19284);
xnor U19831 (N_19831,N_19107,N_19185);
nor U19832 (N_19832,N_19399,N_19258);
xor U19833 (N_19833,N_19401,N_19371);
xnor U19834 (N_19834,N_19194,N_19489);
nor U19835 (N_19835,N_19427,N_19280);
xnor U19836 (N_19836,N_19474,N_19466);
nand U19837 (N_19837,N_19055,N_19438);
nor U19838 (N_19838,N_19134,N_19122);
xor U19839 (N_19839,N_19394,N_19254);
xnor U19840 (N_19840,N_19097,N_19462);
nor U19841 (N_19841,N_19008,N_19314);
or U19842 (N_19842,N_19372,N_19323);
and U19843 (N_19843,N_19149,N_19151);
nand U19844 (N_19844,N_19288,N_19392);
and U19845 (N_19845,N_19023,N_19348);
or U19846 (N_19846,N_19432,N_19055);
or U19847 (N_19847,N_19012,N_19185);
nor U19848 (N_19848,N_19389,N_19476);
nor U19849 (N_19849,N_19340,N_19225);
or U19850 (N_19850,N_19206,N_19310);
and U19851 (N_19851,N_19235,N_19000);
xor U19852 (N_19852,N_19438,N_19066);
nand U19853 (N_19853,N_19071,N_19439);
nor U19854 (N_19854,N_19468,N_19026);
nand U19855 (N_19855,N_19081,N_19357);
and U19856 (N_19856,N_19332,N_19402);
nand U19857 (N_19857,N_19168,N_19452);
and U19858 (N_19858,N_19088,N_19042);
nor U19859 (N_19859,N_19302,N_19007);
nand U19860 (N_19860,N_19156,N_19124);
or U19861 (N_19861,N_19485,N_19096);
or U19862 (N_19862,N_19299,N_19398);
and U19863 (N_19863,N_19477,N_19321);
xor U19864 (N_19864,N_19072,N_19390);
nand U19865 (N_19865,N_19325,N_19315);
nand U19866 (N_19866,N_19428,N_19377);
nor U19867 (N_19867,N_19351,N_19381);
nor U19868 (N_19868,N_19240,N_19024);
and U19869 (N_19869,N_19060,N_19442);
xor U19870 (N_19870,N_19299,N_19269);
and U19871 (N_19871,N_19166,N_19134);
xor U19872 (N_19872,N_19130,N_19221);
and U19873 (N_19873,N_19199,N_19312);
nor U19874 (N_19874,N_19430,N_19199);
or U19875 (N_19875,N_19235,N_19240);
nand U19876 (N_19876,N_19013,N_19202);
nand U19877 (N_19877,N_19336,N_19407);
nor U19878 (N_19878,N_19460,N_19140);
nor U19879 (N_19879,N_19350,N_19048);
or U19880 (N_19880,N_19251,N_19355);
or U19881 (N_19881,N_19201,N_19486);
nand U19882 (N_19882,N_19268,N_19261);
xnor U19883 (N_19883,N_19297,N_19282);
or U19884 (N_19884,N_19099,N_19385);
and U19885 (N_19885,N_19411,N_19478);
and U19886 (N_19886,N_19452,N_19259);
nor U19887 (N_19887,N_19434,N_19399);
nand U19888 (N_19888,N_19132,N_19189);
nor U19889 (N_19889,N_19226,N_19046);
and U19890 (N_19890,N_19443,N_19211);
nand U19891 (N_19891,N_19114,N_19128);
or U19892 (N_19892,N_19408,N_19042);
or U19893 (N_19893,N_19451,N_19331);
xor U19894 (N_19894,N_19416,N_19381);
nand U19895 (N_19895,N_19319,N_19377);
nor U19896 (N_19896,N_19358,N_19359);
xnor U19897 (N_19897,N_19203,N_19112);
xor U19898 (N_19898,N_19055,N_19189);
nor U19899 (N_19899,N_19067,N_19096);
nor U19900 (N_19900,N_19201,N_19043);
and U19901 (N_19901,N_19268,N_19463);
nand U19902 (N_19902,N_19353,N_19191);
xnor U19903 (N_19903,N_19328,N_19476);
nand U19904 (N_19904,N_19323,N_19227);
and U19905 (N_19905,N_19101,N_19137);
nor U19906 (N_19906,N_19319,N_19253);
and U19907 (N_19907,N_19034,N_19148);
and U19908 (N_19908,N_19234,N_19449);
nand U19909 (N_19909,N_19232,N_19087);
nor U19910 (N_19910,N_19179,N_19143);
nand U19911 (N_19911,N_19275,N_19145);
and U19912 (N_19912,N_19043,N_19117);
or U19913 (N_19913,N_19381,N_19236);
and U19914 (N_19914,N_19331,N_19110);
nand U19915 (N_19915,N_19494,N_19275);
and U19916 (N_19916,N_19080,N_19382);
and U19917 (N_19917,N_19491,N_19021);
or U19918 (N_19918,N_19396,N_19123);
and U19919 (N_19919,N_19407,N_19062);
nand U19920 (N_19920,N_19356,N_19395);
xor U19921 (N_19921,N_19319,N_19408);
nand U19922 (N_19922,N_19322,N_19382);
xnor U19923 (N_19923,N_19189,N_19052);
nand U19924 (N_19924,N_19444,N_19283);
nand U19925 (N_19925,N_19037,N_19257);
nand U19926 (N_19926,N_19419,N_19126);
nor U19927 (N_19927,N_19478,N_19169);
nand U19928 (N_19928,N_19161,N_19167);
xor U19929 (N_19929,N_19237,N_19311);
or U19930 (N_19930,N_19476,N_19188);
nand U19931 (N_19931,N_19137,N_19458);
xnor U19932 (N_19932,N_19431,N_19352);
or U19933 (N_19933,N_19219,N_19352);
xnor U19934 (N_19934,N_19126,N_19138);
and U19935 (N_19935,N_19421,N_19048);
nor U19936 (N_19936,N_19122,N_19294);
xor U19937 (N_19937,N_19394,N_19055);
xnor U19938 (N_19938,N_19404,N_19104);
and U19939 (N_19939,N_19167,N_19406);
or U19940 (N_19940,N_19154,N_19317);
nor U19941 (N_19941,N_19138,N_19183);
nand U19942 (N_19942,N_19417,N_19471);
nand U19943 (N_19943,N_19297,N_19167);
or U19944 (N_19944,N_19358,N_19009);
and U19945 (N_19945,N_19095,N_19323);
nor U19946 (N_19946,N_19243,N_19069);
and U19947 (N_19947,N_19218,N_19309);
and U19948 (N_19948,N_19422,N_19284);
or U19949 (N_19949,N_19020,N_19332);
xnor U19950 (N_19950,N_19022,N_19286);
or U19951 (N_19951,N_19134,N_19146);
nor U19952 (N_19952,N_19120,N_19324);
xnor U19953 (N_19953,N_19255,N_19492);
nand U19954 (N_19954,N_19358,N_19385);
nand U19955 (N_19955,N_19017,N_19296);
nand U19956 (N_19956,N_19057,N_19114);
nand U19957 (N_19957,N_19426,N_19020);
nor U19958 (N_19958,N_19471,N_19488);
nand U19959 (N_19959,N_19104,N_19182);
and U19960 (N_19960,N_19395,N_19367);
and U19961 (N_19961,N_19101,N_19427);
or U19962 (N_19962,N_19440,N_19315);
xnor U19963 (N_19963,N_19494,N_19215);
xor U19964 (N_19964,N_19321,N_19352);
and U19965 (N_19965,N_19218,N_19362);
and U19966 (N_19966,N_19251,N_19483);
nand U19967 (N_19967,N_19393,N_19258);
nor U19968 (N_19968,N_19043,N_19108);
nor U19969 (N_19969,N_19097,N_19105);
and U19970 (N_19970,N_19002,N_19018);
xor U19971 (N_19971,N_19368,N_19004);
and U19972 (N_19972,N_19296,N_19431);
xor U19973 (N_19973,N_19134,N_19260);
or U19974 (N_19974,N_19491,N_19499);
nand U19975 (N_19975,N_19117,N_19324);
xor U19976 (N_19976,N_19386,N_19366);
and U19977 (N_19977,N_19212,N_19010);
or U19978 (N_19978,N_19301,N_19175);
xor U19979 (N_19979,N_19274,N_19021);
nor U19980 (N_19980,N_19276,N_19192);
nor U19981 (N_19981,N_19468,N_19330);
nand U19982 (N_19982,N_19403,N_19475);
nand U19983 (N_19983,N_19102,N_19125);
nor U19984 (N_19984,N_19498,N_19320);
or U19985 (N_19985,N_19467,N_19093);
nor U19986 (N_19986,N_19365,N_19054);
nor U19987 (N_19987,N_19029,N_19152);
and U19988 (N_19988,N_19262,N_19369);
nor U19989 (N_19989,N_19217,N_19358);
and U19990 (N_19990,N_19444,N_19198);
or U19991 (N_19991,N_19047,N_19410);
nor U19992 (N_19992,N_19378,N_19308);
xor U19993 (N_19993,N_19058,N_19437);
nor U19994 (N_19994,N_19465,N_19401);
and U19995 (N_19995,N_19154,N_19167);
or U19996 (N_19996,N_19219,N_19376);
nand U19997 (N_19997,N_19133,N_19250);
or U19998 (N_19998,N_19437,N_19413);
nor U19999 (N_19999,N_19390,N_19415);
nor U20000 (N_20000,N_19840,N_19787);
nand U20001 (N_20001,N_19667,N_19841);
or U20002 (N_20002,N_19554,N_19936);
xor U20003 (N_20003,N_19806,N_19907);
nand U20004 (N_20004,N_19716,N_19924);
nand U20005 (N_20005,N_19659,N_19705);
nand U20006 (N_20006,N_19995,N_19950);
or U20007 (N_20007,N_19576,N_19635);
and U20008 (N_20008,N_19676,N_19827);
or U20009 (N_20009,N_19690,N_19550);
nor U20010 (N_20010,N_19894,N_19958);
nor U20011 (N_20011,N_19551,N_19509);
or U20012 (N_20012,N_19504,N_19696);
nand U20013 (N_20013,N_19570,N_19955);
nor U20014 (N_20014,N_19636,N_19988);
nand U20015 (N_20015,N_19784,N_19712);
nor U20016 (N_20016,N_19915,N_19796);
xnor U20017 (N_20017,N_19653,N_19852);
nand U20018 (N_20018,N_19885,N_19822);
nor U20019 (N_20019,N_19641,N_19855);
xor U20020 (N_20020,N_19600,N_19561);
nand U20021 (N_20021,N_19780,N_19668);
and U20022 (N_20022,N_19908,N_19802);
and U20023 (N_20023,N_19591,N_19864);
xnor U20024 (N_20024,N_19813,N_19596);
nor U20025 (N_20025,N_19726,N_19850);
and U20026 (N_20026,N_19881,N_19771);
nor U20027 (N_20027,N_19516,N_19730);
and U20028 (N_20028,N_19700,N_19633);
nand U20029 (N_20029,N_19931,N_19986);
nand U20030 (N_20030,N_19876,N_19692);
and U20031 (N_20031,N_19835,N_19513);
xnor U20032 (N_20032,N_19875,N_19662);
and U20033 (N_20033,N_19526,N_19845);
nor U20034 (N_20034,N_19744,N_19597);
nand U20035 (N_20035,N_19706,N_19899);
and U20036 (N_20036,N_19863,N_19564);
xor U20037 (N_20037,N_19521,N_19539);
nor U20038 (N_20038,N_19929,N_19742);
or U20039 (N_20039,N_19632,N_19946);
nor U20040 (N_20040,N_19650,N_19556);
nor U20041 (N_20041,N_19501,N_19804);
nand U20042 (N_20042,N_19949,N_19951);
nor U20043 (N_20043,N_19703,N_19790);
nor U20044 (N_20044,N_19954,N_19938);
xnor U20045 (N_20045,N_19540,N_19699);
xnor U20046 (N_20046,N_19525,N_19506);
nor U20047 (N_20047,N_19584,N_19971);
nor U20048 (N_20048,N_19595,N_19891);
nand U20049 (N_20049,N_19625,N_19531);
xnor U20050 (N_20050,N_19638,N_19725);
or U20051 (N_20051,N_19837,N_19945);
nor U20052 (N_20052,N_19957,N_19555);
nand U20053 (N_20053,N_19631,N_19895);
and U20054 (N_20054,N_19919,N_19882);
nand U20055 (N_20055,N_19970,N_19524);
and U20056 (N_20056,N_19634,N_19964);
nor U20057 (N_20057,N_19642,N_19861);
xnor U20058 (N_20058,N_19752,N_19508);
and U20059 (N_20059,N_19962,N_19602);
xnor U20060 (N_20060,N_19646,N_19824);
nor U20061 (N_20061,N_19708,N_19905);
or U20062 (N_20062,N_19767,N_19893);
nor U20063 (N_20063,N_19888,N_19750);
or U20064 (N_20064,N_19967,N_19663);
xor U20065 (N_20065,N_19758,N_19562);
and U20066 (N_20066,N_19735,N_19694);
nor U20067 (N_20067,N_19917,N_19973);
nor U20068 (N_20068,N_19503,N_19765);
nand U20069 (N_20069,N_19665,N_19715);
xnor U20070 (N_20070,N_19768,N_19808);
and U20071 (N_20071,N_19598,N_19603);
and U20072 (N_20072,N_19916,N_19713);
xor U20073 (N_20073,N_19507,N_19728);
nor U20074 (N_20074,N_19857,N_19607);
nand U20075 (N_20075,N_19710,N_19543);
nor U20076 (N_20076,N_19831,N_19669);
and U20077 (N_20077,N_19582,N_19877);
nor U20078 (N_20078,N_19989,N_19909);
nand U20079 (N_20079,N_19658,N_19781);
and U20080 (N_20080,N_19686,N_19736);
and U20081 (N_20081,N_19817,N_19886);
or U20082 (N_20082,N_19872,N_19546);
nand U20083 (N_20083,N_19741,N_19997);
xnor U20084 (N_20084,N_19772,N_19969);
xnor U20085 (N_20085,N_19568,N_19579);
and U20086 (N_20086,N_19604,N_19552);
nor U20087 (N_20087,N_19775,N_19626);
nor U20088 (N_20088,N_19542,N_19810);
xnor U20089 (N_20089,N_19627,N_19677);
nor U20090 (N_20090,N_19902,N_19981);
or U20091 (N_20091,N_19614,N_19874);
xor U20092 (N_20092,N_19776,N_19510);
or U20093 (N_20093,N_19849,N_19559);
or U20094 (N_20094,N_19724,N_19578);
xor U20095 (N_20095,N_19980,N_19976);
and U20096 (N_20096,N_19618,N_19900);
nand U20097 (N_20097,N_19953,N_19571);
nand U20098 (N_20098,N_19826,N_19994);
and U20099 (N_20099,N_19865,N_19847);
xnor U20100 (N_20100,N_19737,N_19975);
xnor U20101 (N_20101,N_19657,N_19610);
xor U20102 (N_20102,N_19577,N_19580);
and U20103 (N_20103,N_19698,N_19755);
nand U20104 (N_20104,N_19572,N_19718);
nor U20105 (N_20105,N_19536,N_19856);
or U20106 (N_20106,N_19911,N_19651);
xnor U20107 (N_20107,N_19647,N_19733);
nand U20108 (N_20108,N_19854,N_19910);
xnor U20109 (N_20109,N_19760,N_19678);
or U20110 (N_20110,N_19585,N_19639);
xor U20111 (N_20111,N_19828,N_19789);
nand U20112 (N_20112,N_19652,N_19544);
xor U20113 (N_20113,N_19688,N_19518);
or U20114 (N_20114,N_19927,N_19519);
nor U20115 (N_20115,N_19846,N_19811);
nand U20116 (N_20116,N_19966,N_19628);
nand U20117 (N_20117,N_19999,N_19948);
xor U20118 (N_20118,N_19795,N_19693);
xnor U20119 (N_20119,N_19901,N_19500);
nor U20120 (N_20120,N_19574,N_19939);
and U20121 (N_20121,N_19853,N_19581);
nand U20122 (N_20122,N_19926,N_19921);
nand U20123 (N_20123,N_19793,N_19606);
xor U20124 (N_20124,N_19943,N_19517);
xor U20125 (N_20125,N_19714,N_19723);
or U20126 (N_20126,N_19720,N_19739);
nand U20127 (N_20127,N_19512,N_19821);
or U20128 (N_20128,N_19890,N_19673);
nand U20129 (N_20129,N_19529,N_19851);
nand U20130 (N_20130,N_19738,N_19541);
and U20131 (N_20131,N_19952,N_19812);
nand U20132 (N_20132,N_19680,N_19611);
nand U20133 (N_20133,N_19629,N_19879);
nor U20134 (N_20134,N_19779,N_19920);
nor U20135 (N_20135,N_19898,N_19537);
and U20136 (N_20136,N_19871,N_19757);
and U20137 (N_20137,N_19887,N_19523);
and U20138 (N_20138,N_19640,N_19753);
nor U20139 (N_20139,N_19833,N_19731);
nor U20140 (N_20140,N_19996,N_19684);
xnor U20141 (N_20141,N_19515,N_19534);
nand U20142 (N_20142,N_19834,N_19560);
and U20143 (N_20143,N_19985,N_19773);
and U20144 (N_20144,N_19704,N_19990);
or U20145 (N_20145,N_19977,N_19545);
nand U20146 (N_20146,N_19982,N_19589);
or U20147 (N_20147,N_19538,N_19583);
or U20148 (N_20148,N_19791,N_19956);
nand U20149 (N_20149,N_19533,N_19830);
and U20150 (N_20150,N_19889,N_19514);
or U20151 (N_20151,N_19532,N_19896);
xnor U20152 (N_20152,N_19528,N_19649);
xor U20153 (N_20153,N_19594,N_19617);
and U20154 (N_20154,N_19880,N_19884);
nand U20155 (N_20155,N_19527,N_19944);
nand U20156 (N_20156,N_19838,N_19588);
nand U20157 (N_20157,N_19599,N_19839);
and U20158 (N_20158,N_19749,N_19930);
or U20159 (N_20159,N_19695,N_19801);
nor U20160 (N_20160,N_19520,N_19843);
and U20161 (N_20161,N_19923,N_19707);
xor U20162 (N_20162,N_19530,N_19732);
or U20163 (N_20163,N_19683,N_19759);
and U20164 (N_20164,N_19859,N_19820);
xnor U20165 (N_20165,N_19987,N_19809);
nand U20166 (N_20166,N_19660,N_19866);
or U20167 (N_20167,N_19609,N_19687);
or U20168 (N_20168,N_19858,N_19746);
xnor U20169 (N_20169,N_19800,N_19783);
and U20170 (N_20170,N_19797,N_19832);
nor U20171 (N_20171,N_19643,N_19645);
xnor U20172 (N_20172,N_19942,N_19756);
xor U20173 (N_20173,N_19937,N_19816);
xnor U20174 (N_20174,N_19786,N_19666);
nor U20175 (N_20175,N_19778,N_19807);
nand U20176 (N_20176,N_19814,N_19553);
nor U20177 (N_20177,N_19549,N_19522);
xnor U20178 (N_20178,N_19612,N_19547);
or U20179 (N_20179,N_19815,N_19794);
xor U20180 (N_20180,N_19656,N_19675);
and U20181 (N_20181,N_19892,N_19566);
nand U20182 (N_20182,N_19615,N_19965);
or U20183 (N_20183,N_19903,N_19819);
and U20184 (N_20184,N_19648,N_19593);
nand U20185 (N_20185,N_19557,N_19586);
nand U20186 (N_20186,N_19761,N_19993);
and U20187 (N_20187,N_19674,N_19829);
and U20188 (N_20188,N_19587,N_19747);
xor U20189 (N_20189,N_19621,N_19869);
nor U20190 (N_20190,N_19630,N_19721);
and U20191 (N_20191,N_19748,N_19672);
nor U20192 (N_20192,N_19719,N_19754);
or U20193 (N_20193,N_19912,N_19722);
xor U20194 (N_20194,N_19535,N_19984);
or U20195 (N_20195,N_19671,N_19868);
nand U20196 (N_20196,N_19883,N_19601);
or U20197 (N_20197,N_19928,N_19569);
nor U20198 (N_20198,N_19782,N_19682);
and U20199 (N_20199,N_19691,N_19979);
and U20200 (N_20200,N_19613,N_19842);
xor U20201 (N_20201,N_19679,N_19836);
nand U20202 (N_20202,N_19961,N_19959);
nand U20203 (N_20203,N_19978,N_19803);
xor U20204 (N_20204,N_19914,N_19573);
xor U20205 (N_20205,N_19654,N_19644);
nand U20206 (N_20206,N_19727,N_19637);
xnor U20207 (N_20207,N_19922,N_19992);
xor U20208 (N_20208,N_19897,N_19825);
and U20209 (N_20209,N_19785,N_19717);
and U20210 (N_20210,N_19935,N_19991);
xnor U20211 (N_20211,N_19616,N_19702);
or U20212 (N_20212,N_19511,N_19619);
nand U20213 (N_20213,N_19940,N_19563);
xor U20214 (N_20214,N_19777,N_19867);
and U20215 (N_20215,N_19711,N_19968);
nor U20216 (N_20216,N_19548,N_19623);
nand U20217 (N_20217,N_19823,N_19941);
nor U20218 (N_20218,N_19934,N_19998);
nor U20219 (N_20219,N_19862,N_19873);
nand U20220 (N_20220,N_19655,N_19701);
or U20221 (N_20221,N_19743,N_19913);
and U20222 (N_20222,N_19918,N_19947);
nor U20223 (N_20223,N_19764,N_19974);
and U20224 (N_20224,N_19792,N_19818);
nand U20225 (N_20225,N_19925,N_19670);
or U20226 (N_20226,N_19624,N_19799);
and U20227 (N_20227,N_19729,N_19661);
and U20228 (N_20228,N_19762,N_19870);
nand U20229 (N_20229,N_19960,N_19685);
xor U20230 (N_20230,N_19567,N_19608);
and U20231 (N_20231,N_19565,N_19734);
or U20232 (N_20232,N_19664,N_19605);
or U20233 (N_20233,N_19774,N_19590);
and U20234 (N_20234,N_19740,N_19620);
or U20235 (N_20235,N_19681,N_19709);
and U20236 (N_20236,N_19860,N_19769);
xor U20237 (N_20237,N_19788,N_19622);
xnor U20238 (N_20238,N_19805,N_19763);
nor U20239 (N_20239,N_19505,N_19798);
or U20240 (N_20240,N_19904,N_19575);
xnor U20241 (N_20241,N_19592,N_19558);
nor U20242 (N_20242,N_19697,N_19770);
xnor U20243 (N_20243,N_19963,N_19878);
nor U20244 (N_20244,N_19766,N_19933);
nand U20245 (N_20245,N_19848,N_19502);
xor U20246 (N_20246,N_19745,N_19751);
nand U20247 (N_20247,N_19983,N_19972);
and U20248 (N_20248,N_19906,N_19689);
or U20249 (N_20249,N_19932,N_19844);
nor U20250 (N_20250,N_19966,N_19597);
xnor U20251 (N_20251,N_19703,N_19692);
and U20252 (N_20252,N_19660,N_19778);
nand U20253 (N_20253,N_19707,N_19789);
nand U20254 (N_20254,N_19950,N_19731);
xnor U20255 (N_20255,N_19709,N_19738);
nor U20256 (N_20256,N_19798,N_19719);
and U20257 (N_20257,N_19610,N_19574);
nand U20258 (N_20258,N_19885,N_19710);
xor U20259 (N_20259,N_19769,N_19944);
nand U20260 (N_20260,N_19594,N_19692);
nor U20261 (N_20261,N_19578,N_19902);
and U20262 (N_20262,N_19852,N_19968);
or U20263 (N_20263,N_19907,N_19830);
nor U20264 (N_20264,N_19978,N_19507);
nand U20265 (N_20265,N_19807,N_19789);
xor U20266 (N_20266,N_19614,N_19643);
or U20267 (N_20267,N_19865,N_19961);
xor U20268 (N_20268,N_19987,N_19878);
or U20269 (N_20269,N_19939,N_19507);
and U20270 (N_20270,N_19741,N_19809);
and U20271 (N_20271,N_19999,N_19604);
nor U20272 (N_20272,N_19681,N_19581);
nand U20273 (N_20273,N_19925,N_19912);
xnor U20274 (N_20274,N_19554,N_19715);
nand U20275 (N_20275,N_19819,N_19949);
nand U20276 (N_20276,N_19929,N_19755);
or U20277 (N_20277,N_19999,N_19554);
and U20278 (N_20278,N_19608,N_19580);
xnor U20279 (N_20279,N_19848,N_19570);
and U20280 (N_20280,N_19961,N_19954);
and U20281 (N_20281,N_19552,N_19565);
nand U20282 (N_20282,N_19936,N_19969);
nand U20283 (N_20283,N_19895,N_19782);
nor U20284 (N_20284,N_19912,N_19518);
or U20285 (N_20285,N_19639,N_19864);
xor U20286 (N_20286,N_19842,N_19629);
nor U20287 (N_20287,N_19743,N_19742);
or U20288 (N_20288,N_19536,N_19849);
and U20289 (N_20289,N_19775,N_19695);
xnor U20290 (N_20290,N_19979,N_19592);
and U20291 (N_20291,N_19838,N_19983);
nor U20292 (N_20292,N_19953,N_19868);
and U20293 (N_20293,N_19970,N_19659);
nand U20294 (N_20294,N_19620,N_19833);
nand U20295 (N_20295,N_19701,N_19629);
and U20296 (N_20296,N_19527,N_19511);
or U20297 (N_20297,N_19715,N_19596);
nor U20298 (N_20298,N_19834,N_19544);
and U20299 (N_20299,N_19673,N_19559);
xnor U20300 (N_20300,N_19855,N_19867);
or U20301 (N_20301,N_19767,N_19827);
nand U20302 (N_20302,N_19908,N_19621);
nor U20303 (N_20303,N_19744,N_19603);
nand U20304 (N_20304,N_19658,N_19748);
nand U20305 (N_20305,N_19788,N_19794);
nand U20306 (N_20306,N_19798,N_19891);
or U20307 (N_20307,N_19545,N_19853);
nor U20308 (N_20308,N_19905,N_19917);
xor U20309 (N_20309,N_19622,N_19654);
or U20310 (N_20310,N_19517,N_19712);
and U20311 (N_20311,N_19593,N_19965);
nor U20312 (N_20312,N_19513,N_19590);
or U20313 (N_20313,N_19743,N_19737);
nand U20314 (N_20314,N_19605,N_19706);
or U20315 (N_20315,N_19945,N_19886);
nand U20316 (N_20316,N_19519,N_19714);
nand U20317 (N_20317,N_19687,N_19726);
nor U20318 (N_20318,N_19744,N_19626);
nand U20319 (N_20319,N_19979,N_19955);
xnor U20320 (N_20320,N_19889,N_19986);
nor U20321 (N_20321,N_19882,N_19848);
nor U20322 (N_20322,N_19802,N_19642);
nor U20323 (N_20323,N_19638,N_19681);
nand U20324 (N_20324,N_19631,N_19579);
or U20325 (N_20325,N_19906,N_19630);
nand U20326 (N_20326,N_19641,N_19602);
nand U20327 (N_20327,N_19778,N_19815);
nand U20328 (N_20328,N_19963,N_19577);
and U20329 (N_20329,N_19570,N_19884);
or U20330 (N_20330,N_19774,N_19859);
nand U20331 (N_20331,N_19661,N_19505);
nor U20332 (N_20332,N_19583,N_19727);
nor U20333 (N_20333,N_19755,N_19786);
or U20334 (N_20334,N_19920,N_19788);
nor U20335 (N_20335,N_19719,N_19833);
or U20336 (N_20336,N_19832,N_19890);
and U20337 (N_20337,N_19583,N_19656);
nand U20338 (N_20338,N_19655,N_19503);
or U20339 (N_20339,N_19957,N_19886);
nor U20340 (N_20340,N_19935,N_19988);
nand U20341 (N_20341,N_19871,N_19949);
and U20342 (N_20342,N_19633,N_19692);
xnor U20343 (N_20343,N_19544,N_19533);
or U20344 (N_20344,N_19766,N_19686);
xnor U20345 (N_20345,N_19726,N_19871);
nand U20346 (N_20346,N_19864,N_19687);
or U20347 (N_20347,N_19781,N_19888);
and U20348 (N_20348,N_19936,N_19736);
and U20349 (N_20349,N_19717,N_19903);
xnor U20350 (N_20350,N_19953,N_19973);
and U20351 (N_20351,N_19607,N_19887);
nor U20352 (N_20352,N_19561,N_19774);
nor U20353 (N_20353,N_19805,N_19901);
nor U20354 (N_20354,N_19644,N_19903);
and U20355 (N_20355,N_19601,N_19792);
and U20356 (N_20356,N_19867,N_19505);
and U20357 (N_20357,N_19941,N_19584);
nand U20358 (N_20358,N_19788,N_19674);
and U20359 (N_20359,N_19668,N_19740);
and U20360 (N_20360,N_19924,N_19696);
and U20361 (N_20361,N_19956,N_19652);
xor U20362 (N_20362,N_19987,N_19937);
and U20363 (N_20363,N_19957,N_19527);
and U20364 (N_20364,N_19955,N_19951);
and U20365 (N_20365,N_19698,N_19677);
and U20366 (N_20366,N_19937,N_19605);
nand U20367 (N_20367,N_19749,N_19689);
or U20368 (N_20368,N_19874,N_19795);
and U20369 (N_20369,N_19715,N_19822);
or U20370 (N_20370,N_19670,N_19978);
nor U20371 (N_20371,N_19613,N_19580);
or U20372 (N_20372,N_19854,N_19719);
or U20373 (N_20373,N_19677,N_19708);
and U20374 (N_20374,N_19704,N_19921);
nor U20375 (N_20375,N_19748,N_19536);
nor U20376 (N_20376,N_19900,N_19654);
nand U20377 (N_20377,N_19975,N_19564);
nor U20378 (N_20378,N_19841,N_19614);
or U20379 (N_20379,N_19534,N_19949);
nand U20380 (N_20380,N_19677,N_19743);
xor U20381 (N_20381,N_19788,N_19573);
and U20382 (N_20382,N_19672,N_19990);
nor U20383 (N_20383,N_19734,N_19722);
xor U20384 (N_20384,N_19892,N_19524);
nand U20385 (N_20385,N_19886,N_19636);
nor U20386 (N_20386,N_19539,N_19675);
xnor U20387 (N_20387,N_19586,N_19916);
nor U20388 (N_20388,N_19635,N_19732);
nand U20389 (N_20389,N_19528,N_19633);
nand U20390 (N_20390,N_19729,N_19977);
and U20391 (N_20391,N_19720,N_19608);
nor U20392 (N_20392,N_19759,N_19838);
xnor U20393 (N_20393,N_19950,N_19679);
and U20394 (N_20394,N_19812,N_19765);
or U20395 (N_20395,N_19780,N_19743);
nor U20396 (N_20396,N_19619,N_19929);
xor U20397 (N_20397,N_19987,N_19956);
or U20398 (N_20398,N_19992,N_19559);
and U20399 (N_20399,N_19695,N_19508);
xor U20400 (N_20400,N_19800,N_19901);
or U20401 (N_20401,N_19861,N_19952);
and U20402 (N_20402,N_19817,N_19582);
and U20403 (N_20403,N_19747,N_19712);
and U20404 (N_20404,N_19900,N_19928);
nand U20405 (N_20405,N_19590,N_19744);
and U20406 (N_20406,N_19897,N_19828);
nor U20407 (N_20407,N_19945,N_19556);
and U20408 (N_20408,N_19743,N_19651);
and U20409 (N_20409,N_19525,N_19702);
and U20410 (N_20410,N_19531,N_19895);
xnor U20411 (N_20411,N_19934,N_19738);
and U20412 (N_20412,N_19794,N_19589);
or U20413 (N_20413,N_19607,N_19835);
nor U20414 (N_20414,N_19898,N_19602);
nor U20415 (N_20415,N_19783,N_19577);
or U20416 (N_20416,N_19897,N_19610);
nand U20417 (N_20417,N_19531,N_19672);
xor U20418 (N_20418,N_19899,N_19574);
and U20419 (N_20419,N_19818,N_19756);
or U20420 (N_20420,N_19631,N_19953);
and U20421 (N_20421,N_19934,N_19859);
and U20422 (N_20422,N_19809,N_19646);
xor U20423 (N_20423,N_19812,N_19680);
nand U20424 (N_20424,N_19920,N_19829);
and U20425 (N_20425,N_19653,N_19760);
or U20426 (N_20426,N_19999,N_19606);
or U20427 (N_20427,N_19861,N_19600);
xnor U20428 (N_20428,N_19787,N_19821);
xnor U20429 (N_20429,N_19836,N_19724);
nand U20430 (N_20430,N_19868,N_19879);
and U20431 (N_20431,N_19793,N_19803);
xnor U20432 (N_20432,N_19664,N_19717);
xor U20433 (N_20433,N_19861,N_19997);
and U20434 (N_20434,N_19621,N_19645);
nand U20435 (N_20435,N_19950,N_19583);
and U20436 (N_20436,N_19752,N_19845);
xor U20437 (N_20437,N_19927,N_19792);
xor U20438 (N_20438,N_19887,N_19962);
nand U20439 (N_20439,N_19891,N_19708);
or U20440 (N_20440,N_19745,N_19941);
nand U20441 (N_20441,N_19776,N_19974);
or U20442 (N_20442,N_19504,N_19958);
nand U20443 (N_20443,N_19793,N_19943);
or U20444 (N_20444,N_19984,N_19871);
or U20445 (N_20445,N_19936,N_19813);
and U20446 (N_20446,N_19823,N_19654);
or U20447 (N_20447,N_19996,N_19593);
nand U20448 (N_20448,N_19546,N_19621);
and U20449 (N_20449,N_19784,N_19503);
xnor U20450 (N_20450,N_19970,N_19905);
or U20451 (N_20451,N_19795,N_19858);
or U20452 (N_20452,N_19575,N_19911);
nor U20453 (N_20453,N_19880,N_19875);
nand U20454 (N_20454,N_19973,N_19751);
nor U20455 (N_20455,N_19639,N_19534);
nor U20456 (N_20456,N_19547,N_19693);
or U20457 (N_20457,N_19753,N_19591);
nand U20458 (N_20458,N_19872,N_19889);
nor U20459 (N_20459,N_19835,N_19979);
nor U20460 (N_20460,N_19592,N_19526);
and U20461 (N_20461,N_19621,N_19893);
nand U20462 (N_20462,N_19859,N_19525);
nor U20463 (N_20463,N_19755,N_19948);
or U20464 (N_20464,N_19801,N_19880);
and U20465 (N_20465,N_19791,N_19630);
xor U20466 (N_20466,N_19770,N_19519);
or U20467 (N_20467,N_19946,N_19831);
and U20468 (N_20468,N_19840,N_19972);
and U20469 (N_20469,N_19561,N_19568);
nand U20470 (N_20470,N_19668,N_19684);
or U20471 (N_20471,N_19541,N_19554);
xnor U20472 (N_20472,N_19631,N_19801);
xor U20473 (N_20473,N_19687,N_19897);
nor U20474 (N_20474,N_19819,N_19670);
or U20475 (N_20475,N_19787,N_19724);
and U20476 (N_20476,N_19763,N_19655);
xnor U20477 (N_20477,N_19524,N_19939);
xor U20478 (N_20478,N_19652,N_19673);
nor U20479 (N_20479,N_19537,N_19922);
xor U20480 (N_20480,N_19875,N_19650);
xnor U20481 (N_20481,N_19719,N_19707);
and U20482 (N_20482,N_19666,N_19902);
or U20483 (N_20483,N_19851,N_19515);
xor U20484 (N_20484,N_19970,N_19648);
xnor U20485 (N_20485,N_19722,N_19993);
or U20486 (N_20486,N_19566,N_19867);
nand U20487 (N_20487,N_19566,N_19524);
and U20488 (N_20488,N_19747,N_19694);
or U20489 (N_20489,N_19664,N_19975);
nor U20490 (N_20490,N_19711,N_19916);
or U20491 (N_20491,N_19587,N_19773);
and U20492 (N_20492,N_19979,N_19585);
xnor U20493 (N_20493,N_19972,N_19989);
nor U20494 (N_20494,N_19552,N_19574);
or U20495 (N_20495,N_19618,N_19526);
nand U20496 (N_20496,N_19625,N_19535);
and U20497 (N_20497,N_19592,N_19864);
xor U20498 (N_20498,N_19994,N_19849);
or U20499 (N_20499,N_19748,N_19721);
nand U20500 (N_20500,N_20134,N_20155);
nand U20501 (N_20501,N_20302,N_20394);
nand U20502 (N_20502,N_20236,N_20006);
nor U20503 (N_20503,N_20050,N_20309);
nor U20504 (N_20504,N_20183,N_20335);
or U20505 (N_20505,N_20142,N_20288);
nor U20506 (N_20506,N_20168,N_20170);
or U20507 (N_20507,N_20382,N_20350);
nand U20508 (N_20508,N_20087,N_20274);
nor U20509 (N_20509,N_20258,N_20051);
or U20510 (N_20510,N_20432,N_20189);
and U20511 (N_20511,N_20406,N_20135);
nor U20512 (N_20512,N_20230,N_20348);
and U20513 (N_20513,N_20018,N_20496);
nand U20514 (N_20514,N_20329,N_20402);
and U20515 (N_20515,N_20115,N_20223);
xor U20516 (N_20516,N_20488,N_20017);
xor U20517 (N_20517,N_20352,N_20431);
nand U20518 (N_20518,N_20208,N_20347);
nand U20519 (N_20519,N_20460,N_20298);
and U20520 (N_20520,N_20033,N_20275);
and U20521 (N_20521,N_20069,N_20032);
nor U20522 (N_20522,N_20169,N_20466);
nor U20523 (N_20523,N_20080,N_20222);
xor U20524 (N_20524,N_20372,N_20068);
or U20525 (N_20525,N_20296,N_20340);
or U20526 (N_20526,N_20178,N_20415);
nand U20527 (N_20527,N_20037,N_20196);
nand U20528 (N_20528,N_20081,N_20244);
and U20529 (N_20529,N_20007,N_20445);
nor U20530 (N_20530,N_20127,N_20217);
or U20531 (N_20531,N_20004,N_20425);
or U20532 (N_20532,N_20345,N_20437);
nand U20533 (N_20533,N_20163,N_20088);
nand U20534 (N_20534,N_20011,N_20457);
and U20535 (N_20535,N_20031,N_20359);
or U20536 (N_20536,N_20283,N_20175);
nand U20537 (N_20537,N_20111,N_20143);
nor U20538 (N_20538,N_20167,N_20197);
and U20539 (N_20539,N_20426,N_20240);
and U20540 (N_20540,N_20319,N_20027);
and U20541 (N_20541,N_20130,N_20060);
xnor U20542 (N_20542,N_20003,N_20364);
nor U20543 (N_20543,N_20267,N_20491);
xor U20544 (N_20544,N_20405,N_20164);
nor U20545 (N_20545,N_20366,N_20370);
nand U20546 (N_20546,N_20157,N_20061);
or U20547 (N_20547,N_20278,N_20441);
or U20548 (N_20548,N_20048,N_20424);
nand U20549 (N_20549,N_20328,N_20277);
nand U20550 (N_20550,N_20066,N_20023);
xnor U20551 (N_20551,N_20132,N_20124);
nor U20552 (N_20552,N_20332,N_20318);
nand U20553 (N_20553,N_20138,N_20276);
nor U20554 (N_20554,N_20059,N_20357);
or U20555 (N_20555,N_20290,N_20409);
or U20556 (N_20556,N_20478,N_20213);
xor U20557 (N_20557,N_20246,N_20005);
xnor U20558 (N_20558,N_20131,N_20487);
xor U20559 (N_20559,N_20078,N_20042);
xnor U20560 (N_20560,N_20158,N_20316);
and U20561 (N_20561,N_20243,N_20353);
or U20562 (N_20562,N_20071,N_20362);
nor U20563 (N_20563,N_20133,N_20162);
or U20564 (N_20564,N_20123,N_20417);
or U20565 (N_20565,N_20247,N_20351);
xor U20566 (N_20566,N_20451,N_20248);
xor U20567 (N_20567,N_20024,N_20165);
nor U20568 (N_20568,N_20414,N_20419);
xnor U20569 (N_20569,N_20121,N_20257);
xor U20570 (N_20570,N_20314,N_20054);
nor U20571 (N_20571,N_20303,N_20461);
and U20572 (N_20572,N_20019,N_20373);
nor U20573 (N_20573,N_20263,N_20064);
xnor U20574 (N_20574,N_20304,N_20342);
and U20575 (N_20575,N_20322,N_20021);
xor U20576 (N_20576,N_20376,N_20367);
or U20577 (N_20577,N_20393,N_20447);
xnor U20578 (N_20578,N_20368,N_20210);
or U20579 (N_20579,N_20485,N_20125);
and U20580 (N_20580,N_20079,N_20420);
and U20581 (N_20581,N_20233,N_20300);
xor U20582 (N_20582,N_20324,N_20101);
or U20583 (N_20583,N_20479,N_20379);
xnor U20584 (N_20584,N_20193,N_20205);
xor U20585 (N_20585,N_20105,N_20237);
and U20586 (N_20586,N_20012,N_20295);
nand U20587 (N_20587,N_20471,N_20235);
and U20588 (N_20588,N_20365,N_20336);
and U20589 (N_20589,N_20312,N_20360);
or U20590 (N_20590,N_20390,N_20001);
nor U20591 (N_20591,N_20176,N_20195);
or U20592 (N_20592,N_20057,N_20120);
xor U20593 (N_20593,N_20156,N_20093);
and U20594 (N_20594,N_20442,N_20082);
xor U20595 (N_20595,N_20065,N_20035);
nor U20596 (N_20596,N_20330,N_20077);
or U20597 (N_20597,N_20215,N_20119);
and U20598 (N_20598,N_20483,N_20140);
or U20599 (N_20599,N_20436,N_20200);
xor U20600 (N_20600,N_20467,N_20153);
nor U20601 (N_20601,N_20053,N_20239);
and U20602 (N_20602,N_20022,N_20400);
nand U20603 (N_20603,N_20398,N_20030);
xnor U20604 (N_20604,N_20122,N_20280);
nand U20605 (N_20605,N_20325,N_20286);
nand U20606 (N_20606,N_20076,N_20002);
nand U20607 (N_20607,N_20411,N_20161);
and U20608 (N_20608,N_20070,N_20259);
nor U20609 (N_20609,N_20473,N_20144);
or U20610 (N_20610,N_20049,N_20349);
or U20611 (N_20611,N_20301,N_20034);
nand U20612 (N_20612,N_20427,N_20141);
and U20613 (N_20613,N_20474,N_20421);
or U20614 (N_20614,N_20454,N_20242);
or U20615 (N_20615,N_20270,N_20321);
nand U20616 (N_20616,N_20216,N_20265);
nor U20617 (N_20617,N_20380,N_20046);
or U20618 (N_20618,N_20498,N_20333);
nor U20619 (N_20619,N_20238,N_20305);
and U20620 (N_20620,N_20199,N_20009);
xor U20621 (N_20621,N_20182,N_20391);
nand U20622 (N_20622,N_20245,N_20440);
and U20623 (N_20623,N_20486,N_20449);
or U20624 (N_20624,N_20361,N_20472);
xor U20625 (N_20625,N_20464,N_20084);
xnor U20626 (N_20626,N_20408,N_20202);
and U20627 (N_20627,N_20495,N_20015);
xnor U20628 (N_20628,N_20341,N_20293);
nor U20629 (N_20629,N_20020,N_20413);
or U20630 (N_20630,N_20026,N_20313);
and U20631 (N_20631,N_20085,N_20456);
or U20632 (N_20632,N_20104,N_20294);
and U20633 (N_20633,N_20129,N_20228);
nor U20634 (N_20634,N_20160,N_20090);
nor U20635 (N_20635,N_20067,N_20056);
and U20636 (N_20636,N_20171,N_20261);
or U20637 (N_20637,N_20038,N_20493);
and U20638 (N_20638,N_20102,N_20204);
nor U20639 (N_20639,N_20281,N_20271);
nor U20640 (N_20640,N_20469,N_20180);
nor U20641 (N_20641,N_20455,N_20219);
nand U20642 (N_20642,N_20346,N_20326);
and U20643 (N_20643,N_20430,N_20450);
nand U20644 (N_20644,N_20399,N_20462);
nand U20645 (N_20645,N_20166,N_20494);
and U20646 (N_20646,N_20256,N_20310);
nand U20647 (N_20647,N_20097,N_20331);
and U20648 (N_20648,N_20363,N_20289);
and U20649 (N_20649,N_20126,N_20252);
nor U20650 (N_20650,N_20159,N_20139);
xor U20651 (N_20651,N_20497,N_20315);
nor U20652 (N_20652,N_20098,N_20052);
and U20653 (N_20653,N_20112,N_20181);
nor U20654 (N_20654,N_20291,N_20434);
nor U20655 (N_20655,N_20150,N_20465);
xor U20656 (N_20656,N_20403,N_20386);
or U20657 (N_20657,N_20484,N_20385);
or U20658 (N_20658,N_20186,N_20184);
xnor U20659 (N_20659,N_20279,N_20083);
or U20660 (N_20660,N_20260,N_20106);
nand U20661 (N_20661,N_20377,N_20073);
nor U20662 (N_20662,N_20266,N_20172);
nand U20663 (N_20663,N_20173,N_20418);
nand U20664 (N_20664,N_20475,N_20013);
or U20665 (N_20665,N_20192,N_20401);
xor U20666 (N_20666,N_20369,N_20387);
xnor U20667 (N_20667,N_20422,N_20214);
or U20668 (N_20668,N_20092,N_20152);
and U20669 (N_20669,N_20227,N_20272);
nor U20670 (N_20670,N_20108,N_20014);
or U20671 (N_20671,N_20147,N_20453);
or U20672 (N_20672,N_20095,N_20254);
and U20673 (N_20673,N_20149,N_20397);
and U20674 (N_20674,N_20438,N_20249);
or U20675 (N_20675,N_20389,N_20201);
or U20676 (N_20676,N_20253,N_20458);
nor U20677 (N_20677,N_20358,N_20433);
nand U20678 (N_20678,N_20096,N_20435);
nand U20679 (N_20679,N_20378,N_20194);
and U20680 (N_20680,N_20177,N_20306);
nand U20681 (N_20681,N_20423,N_20452);
and U20682 (N_20682,N_20269,N_20136);
or U20683 (N_20683,N_20174,N_20299);
nor U20684 (N_20684,N_20492,N_20185);
and U20685 (N_20685,N_20187,N_20320);
nand U20686 (N_20686,N_20226,N_20232);
xnor U20687 (N_20687,N_20297,N_20323);
and U20688 (N_20688,N_20407,N_20114);
nand U20689 (N_20689,N_20107,N_20203);
or U20690 (N_20690,N_20327,N_20317);
xor U20691 (N_20691,N_20151,N_20113);
nor U20692 (N_20692,N_20016,N_20499);
and U20693 (N_20693,N_20091,N_20311);
and U20694 (N_20694,N_20028,N_20029);
xor U20695 (N_20695,N_20094,N_20190);
and U20696 (N_20696,N_20392,N_20099);
and U20697 (N_20697,N_20292,N_20481);
or U20698 (N_20698,N_20075,N_20343);
xor U20699 (N_20699,N_20128,N_20356);
and U20700 (N_20700,N_20416,N_20234);
and U20701 (N_20701,N_20250,N_20036);
nor U20702 (N_20702,N_20339,N_20463);
and U20703 (N_20703,N_20118,N_20308);
or U20704 (N_20704,N_20117,N_20148);
or U20705 (N_20705,N_20381,N_20264);
nand U20706 (N_20706,N_20063,N_20116);
nand U20707 (N_20707,N_20448,N_20086);
or U20708 (N_20708,N_20489,N_20355);
nand U20709 (N_20709,N_20262,N_20284);
nand U20710 (N_20710,N_20209,N_20145);
and U20711 (N_20711,N_20251,N_20446);
xnor U20712 (N_20712,N_20137,N_20337);
and U20713 (N_20713,N_20384,N_20410);
or U20714 (N_20714,N_20476,N_20191);
or U20715 (N_20715,N_20282,N_20089);
xor U20716 (N_20716,N_20055,N_20404);
xnor U20717 (N_20717,N_20482,N_20285);
nor U20718 (N_20718,N_20110,N_20109);
and U20719 (N_20719,N_20045,N_20043);
xor U20720 (N_20720,N_20154,N_20490);
and U20721 (N_20721,N_20443,N_20229);
nand U20722 (N_20722,N_20375,N_20255);
nor U20723 (N_20723,N_20354,N_20103);
or U20724 (N_20724,N_20241,N_20072);
or U20725 (N_20725,N_20428,N_20371);
or U20726 (N_20726,N_20383,N_20040);
nand U20727 (N_20727,N_20047,N_20224);
nor U20728 (N_20728,N_20206,N_20338);
or U20729 (N_20729,N_20444,N_20374);
xor U20730 (N_20730,N_20480,N_20395);
nand U20731 (N_20731,N_20429,N_20459);
and U20732 (N_20732,N_20044,N_20211);
nand U20733 (N_20733,N_20439,N_20207);
nand U20734 (N_20734,N_20221,N_20074);
xnor U20735 (N_20735,N_20198,N_20039);
nand U20736 (N_20736,N_20062,N_20388);
nor U20737 (N_20737,N_20100,N_20412);
or U20738 (N_20738,N_20334,N_20010);
xnor U20739 (N_20739,N_20041,N_20470);
nor U20740 (N_20740,N_20231,N_20344);
or U20741 (N_20741,N_20468,N_20008);
nor U20742 (N_20742,N_20268,N_20287);
nand U20743 (N_20743,N_20212,N_20225);
nor U20744 (N_20744,N_20477,N_20396);
and U20745 (N_20745,N_20000,N_20307);
nor U20746 (N_20746,N_20188,N_20058);
or U20747 (N_20747,N_20273,N_20146);
and U20748 (N_20748,N_20218,N_20025);
xor U20749 (N_20749,N_20220,N_20179);
and U20750 (N_20750,N_20409,N_20404);
nand U20751 (N_20751,N_20337,N_20075);
xor U20752 (N_20752,N_20142,N_20486);
nor U20753 (N_20753,N_20101,N_20409);
nor U20754 (N_20754,N_20311,N_20002);
nand U20755 (N_20755,N_20135,N_20144);
xor U20756 (N_20756,N_20413,N_20181);
and U20757 (N_20757,N_20017,N_20121);
and U20758 (N_20758,N_20076,N_20489);
nor U20759 (N_20759,N_20259,N_20141);
or U20760 (N_20760,N_20451,N_20445);
or U20761 (N_20761,N_20489,N_20371);
or U20762 (N_20762,N_20114,N_20350);
and U20763 (N_20763,N_20044,N_20287);
nor U20764 (N_20764,N_20061,N_20028);
nand U20765 (N_20765,N_20054,N_20083);
or U20766 (N_20766,N_20328,N_20046);
nand U20767 (N_20767,N_20334,N_20099);
nor U20768 (N_20768,N_20265,N_20425);
or U20769 (N_20769,N_20454,N_20063);
nor U20770 (N_20770,N_20470,N_20457);
and U20771 (N_20771,N_20492,N_20290);
and U20772 (N_20772,N_20164,N_20032);
and U20773 (N_20773,N_20405,N_20383);
xor U20774 (N_20774,N_20302,N_20188);
or U20775 (N_20775,N_20413,N_20477);
nor U20776 (N_20776,N_20098,N_20157);
nand U20777 (N_20777,N_20358,N_20382);
xor U20778 (N_20778,N_20005,N_20354);
and U20779 (N_20779,N_20272,N_20170);
xor U20780 (N_20780,N_20317,N_20290);
xor U20781 (N_20781,N_20129,N_20429);
nor U20782 (N_20782,N_20295,N_20151);
xor U20783 (N_20783,N_20123,N_20195);
nand U20784 (N_20784,N_20080,N_20057);
and U20785 (N_20785,N_20149,N_20338);
nand U20786 (N_20786,N_20054,N_20395);
and U20787 (N_20787,N_20248,N_20007);
or U20788 (N_20788,N_20049,N_20423);
or U20789 (N_20789,N_20445,N_20011);
nor U20790 (N_20790,N_20369,N_20029);
and U20791 (N_20791,N_20162,N_20391);
or U20792 (N_20792,N_20162,N_20117);
and U20793 (N_20793,N_20163,N_20445);
nor U20794 (N_20794,N_20260,N_20289);
nor U20795 (N_20795,N_20201,N_20363);
and U20796 (N_20796,N_20345,N_20082);
or U20797 (N_20797,N_20103,N_20177);
nor U20798 (N_20798,N_20062,N_20205);
xnor U20799 (N_20799,N_20057,N_20176);
or U20800 (N_20800,N_20047,N_20075);
nor U20801 (N_20801,N_20035,N_20075);
nor U20802 (N_20802,N_20037,N_20221);
nor U20803 (N_20803,N_20374,N_20174);
nor U20804 (N_20804,N_20260,N_20092);
or U20805 (N_20805,N_20020,N_20180);
nand U20806 (N_20806,N_20269,N_20356);
xnor U20807 (N_20807,N_20033,N_20498);
nand U20808 (N_20808,N_20218,N_20157);
and U20809 (N_20809,N_20024,N_20198);
and U20810 (N_20810,N_20321,N_20287);
and U20811 (N_20811,N_20459,N_20166);
or U20812 (N_20812,N_20293,N_20140);
or U20813 (N_20813,N_20130,N_20271);
xor U20814 (N_20814,N_20137,N_20466);
xnor U20815 (N_20815,N_20072,N_20465);
nand U20816 (N_20816,N_20259,N_20359);
xor U20817 (N_20817,N_20111,N_20195);
nor U20818 (N_20818,N_20036,N_20429);
nor U20819 (N_20819,N_20466,N_20429);
and U20820 (N_20820,N_20099,N_20462);
and U20821 (N_20821,N_20087,N_20074);
nand U20822 (N_20822,N_20496,N_20476);
nand U20823 (N_20823,N_20319,N_20347);
nor U20824 (N_20824,N_20097,N_20470);
nor U20825 (N_20825,N_20070,N_20494);
or U20826 (N_20826,N_20295,N_20369);
nor U20827 (N_20827,N_20298,N_20147);
nand U20828 (N_20828,N_20049,N_20150);
and U20829 (N_20829,N_20497,N_20094);
nand U20830 (N_20830,N_20382,N_20083);
and U20831 (N_20831,N_20408,N_20319);
or U20832 (N_20832,N_20117,N_20482);
nand U20833 (N_20833,N_20265,N_20469);
and U20834 (N_20834,N_20174,N_20076);
xnor U20835 (N_20835,N_20334,N_20276);
nand U20836 (N_20836,N_20025,N_20483);
or U20837 (N_20837,N_20293,N_20110);
nand U20838 (N_20838,N_20205,N_20476);
nor U20839 (N_20839,N_20360,N_20468);
or U20840 (N_20840,N_20482,N_20385);
xnor U20841 (N_20841,N_20484,N_20329);
and U20842 (N_20842,N_20081,N_20406);
or U20843 (N_20843,N_20366,N_20423);
nand U20844 (N_20844,N_20006,N_20366);
and U20845 (N_20845,N_20403,N_20304);
nand U20846 (N_20846,N_20448,N_20237);
nand U20847 (N_20847,N_20152,N_20429);
xor U20848 (N_20848,N_20250,N_20432);
xor U20849 (N_20849,N_20321,N_20474);
xnor U20850 (N_20850,N_20304,N_20153);
xnor U20851 (N_20851,N_20349,N_20421);
xnor U20852 (N_20852,N_20069,N_20025);
or U20853 (N_20853,N_20007,N_20481);
and U20854 (N_20854,N_20415,N_20142);
xor U20855 (N_20855,N_20011,N_20274);
nor U20856 (N_20856,N_20393,N_20189);
and U20857 (N_20857,N_20093,N_20033);
xor U20858 (N_20858,N_20312,N_20442);
nand U20859 (N_20859,N_20285,N_20270);
nor U20860 (N_20860,N_20109,N_20032);
nand U20861 (N_20861,N_20365,N_20434);
and U20862 (N_20862,N_20461,N_20380);
xnor U20863 (N_20863,N_20245,N_20078);
xor U20864 (N_20864,N_20140,N_20468);
nor U20865 (N_20865,N_20443,N_20073);
nor U20866 (N_20866,N_20022,N_20376);
xor U20867 (N_20867,N_20193,N_20443);
and U20868 (N_20868,N_20451,N_20280);
or U20869 (N_20869,N_20256,N_20129);
nand U20870 (N_20870,N_20238,N_20306);
and U20871 (N_20871,N_20040,N_20426);
or U20872 (N_20872,N_20400,N_20372);
nor U20873 (N_20873,N_20022,N_20058);
and U20874 (N_20874,N_20105,N_20077);
or U20875 (N_20875,N_20274,N_20414);
nor U20876 (N_20876,N_20236,N_20452);
nor U20877 (N_20877,N_20016,N_20135);
xnor U20878 (N_20878,N_20062,N_20331);
and U20879 (N_20879,N_20070,N_20462);
or U20880 (N_20880,N_20046,N_20160);
or U20881 (N_20881,N_20348,N_20164);
xor U20882 (N_20882,N_20028,N_20458);
or U20883 (N_20883,N_20146,N_20398);
or U20884 (N_20884,N_20138,N_20459);
xor U20885 (N_20885,N_20408,N_20429);
xor U20886 (N_20886,N_20238,N_20490);
xnor U20887 (N_20887,N_20106,N_20422);
and U20888 (N_20888,N_20131,N_20241);
xnor U20889 (N_20889,N_20309,N_20491);
or U20890 (N_20890,N_20201,N_20457);
nor U20891 (N_20891,N_20317,N_20162);
and U20892 (N_20892,N_20314,N_20479);
or U20893 (N_20893,N_20123,N_20238);
and U20894 (N_20894,N_20404,N_20358);
nand U20895 (N_20895,N_20082,N_20336);
nor U20896 (N_20896,N_20189,N_20252);
nor U20897 (N_20897,N_20096,N_20191);
and U20898 (N_20898,N_20277,N_20127);
nand U20899 (N_20899,N_20214,N_20396);
nor U20900 (N_20900,N_20290,N_20009);
or U20901 (N_20901,N_20079,N_20161);
or U20902 (N_20902,N_20415,N_20080);
and U20903 (N_20903,N_20198,N_20472);
nand U20904 (N_20904,N_20019,N_20178);
and U20905 (N_20905,N_20277,N_20336);
xor U20906 (N_20906,N_20195,N_20470);
or U20907 (N_20907,N_20431,N_20112);
xor U20908 (N_20908,N_20197,N_20033);
or U20909 (N_20909,N_20498,N_20183);
nand U20910 (N_20910,N_20248,N_20143);
xnor U20911 (N_20911,N_20415,N_20397);
xnor U20912 (N_20912,N_20177,N_20269);
nor U20913 (N_20913,N_20248,N_20186);
xnor U20914 (N_20914,N_20367,N_20019);
nand U20915 (N_20915,N_20476,N_20210);
nor U20916 (N_20916,N_20166,N_20383);
xnor U20917 (N_20917,N_20286,N_20077);
and U20918 (N_20918,N_20118,N_20284);
nor U20919 (N_20919,N_20182,N_20417);
and U20920 (N_20920,N_20149,N_20272);
or U20921 (N_20921,N_20487,N_20027);
nor U20922 (N_20922,N_20325,N_20327);
nor U20923 (N_20923,N_20117,N_20384);
nor U20924 (N_20924,N_20277,N_20470);
nand U20925 (N_20925,N_20303,N_20126);
nor U20926 (N_20926,N_20332,N_20326);
nor U20927 (N_20927,N_20169,N_20189);
or U20928 (N_20928,N_20323,N_20080);
xor U20929 (N_20929,N_20136,N_20463);
nor U20930 (N_20930,N_20216,N_20475);
and U20931 (N_20931,N_20423,N_20004);
nor U20932 (N_20932,N_20101,N_20122);
and U20933 (N_20933,N_20157,N_20238);
nor U20934 (N_20934,N_20040,N_20097);
xnor U20935 (N_20935,N_20413,N_20385);
and U20936 (N_20936,N_20175,N_20270);
or U20937 (N_20937,N_20008,N_20136);
nand U20938 (N_20938,N_20375,N_20423);
nand U20939 (N_20939,N_20240,N_20242);
xor U20940 (N_20940,N_20250,N_20391);
or U20941 (N_20941,N_20175,N_20408);
and U20942 (N_20942,N_20170,N_20338);
nand U20943 (N_20943,N_20171,N_20097);
xnor U20944 (N_20944,N_20467,N_20171);
or U20945 (N_20945,N_20173,N_20316);
nor U20946 (N_20946,N_20204,N_20038);
xnor U20947 (N_20947,N_20373,N_20374);
nor U20948 (N_20948,N_20375,N_20261);
nor U20949 (N_20949,N_20210,N_20286);
nand U20950 (N_20950,N_20398,N_20086);
and U20951 (N_20951,N_20119,N_20057);
xnor U20952 (N_20952,N_20015,N_20188);
nor U20953 (N_20953,N_20160,N_20093);
and U20954 (N_20954,N_20168,N_20098);
xor U20955 (N_20955,N_20474,N_20043);
and U20956 (N_20956,N_20142,N_20005);
xnor U20957 (N_20957,N_20175,N_20174);
or U20958 (N_20958,N_20435,N_20069);
xor U20959 (N_20959,N_20352,N_20436);
nor U20960 (N_20960,N_20107,N_20446);
nand U20961 (N_20961,N_20259,N_20477);
or U20962 (N_20962,N_20216,N_20039);
xor U20963 (N_20963,N_20378,N_20347);
nor U20964 (N_20964,N_20112,N_20201);
or U20965 (N_20965,N_20129,N_20234);
nand U20966 (N_20966,N_20057,N_20019);
nor U20967 (N_20967,N_20455,N_20027);
and U20968 (N_20968,N_20247,N_20125);
or U20969 (N_20969,N_20256,N_20067);
nor U20970 (N_20970,N_20038,N_20021);
nand U20971 (N_20971,N_20289,N_20234);
nor U20972 (N_20972,N_20285,N_20495);
xor U20973 (N_20973,N_20087,N_20375);
nand U20974 (N_20974,N_20318,N_20406);
nor U20975 (N_20975,N_20303,N_20204);
or U20976 (N_20976,N_20356,N_20057);
nor U20977 (N_20977,N_20200,N_20323);
nor U20978 (N_20978,N_20019,N_20282);
xor U20979 (N_20979,N_20278,N_20143);
and U20980 (N_20980,N_20118,N_20117);
xor U20981 (N_20981,N_20179,N_20397);
nor U20982 (N_20982,N_20105,N_20185);
and U20983 (N_20983,N_20164,N_20162);
nand U20984 (N_20984,N_20336,N_20264);
nand U20985 (N_20985,N_20485,N_20126);
nor U20986 (N_20986,N_20384,N_20321);
nor U20987 (N_20987,N_20219,N_20111);
or U20988 (N_20988,N_20085,N_20024);
nand U20989 (N_20989,N_20165,N_20154);
nand U20990 (N_20990,N_20063,N_20262);
nor U20991 (N_20991,N_20373,N_20361);
or U20992 (N_20992,N_20337,N_20206);
or U20993 (N_20993,N_20381,N_20162);
xnor U20994 (N_20994,N_20136,N_20047);
or U20995 (N_20995,N_20393,N_20431);
nand U20996 (N_20996,N_20356,N_20137);
nand U20997 (N_20997,N_20185,N_20098);
nand U20998 (N_20998,N_20202,N_20190);
and U20999 (N_20999,N_20299,N_20369);
nor U21000 (N_21000,N_20895,N_20782);
nand U21001 (N_21001,N_20863,N_20881);
xor U21002 (N_21002,N_20677,N_20877);
or U21003 (N_21003,N_20565,N_20818);
nor U21004 (N_21004,N_20715,N_20838);
nor U21005 (N_21005,N_20851,N_20774);
nand U21006 (N_21006,N_20972,N_20546);
and U21007 (N_21007,N_20935,N_20945);
or U21008 (N_21008,N_20527,N_20865);
xor U21009 (N_21009,N_20651,N_20650);
or U21010 (N_21010,N_20581,N_20853);
and U21011 (N_21011,N_20634,N_20791);
xor U21012 (N_21012,N_20922,N_20522);
xor U21013 (N_21013,N_20864,N_20684);
and U21014 (N_21014,N_20547,N_20698);
nor U21015 (N_21015,N_20729,N_20513);
nand U21016 (N_21016,N_20883,N_20568);
nor U21017 (N_21017,N_20627,N_20664);
nand U21018 (N_21018,N_20967,N_20887);
xnor U21019 (N_21019,N_20599,N_20716);
nand U21020 (N_21020,N_20825,N_20798);
xnor U21021 (N_21021,N_20893,N_20850);
nand U21022 (N_21022,N_20806,N_20794);
xor U21023 (N_21023,N_20563,N_20997);
nand U21024 (N_21024,N_20544,N_20663);
nor U21025 (N_21025,N_20692,N_20982);
nand U21026 (N_21026,N_20548,N_20847);
or U21027 (N_21027,N_20830,N_20586);
and U21028 (N_21028,N_20585,N_20696);
or U21029 (N_21029,N_20828,N_20552);
xor U21030 (N_21030,N_20783,N_20896);
xnor U21031 (N_21031,N_20977,N_20910);
nor U21032 (N_21032,N_20587,N_20555);
and U21033 (N_21033,N_20758,N_20837);
nand U21034 (N_21034,N_20619,N_20511);
nor U21035 (N_21035,N_20905,N_20719);
or U21036 (N_21036,N_20970,N_20625);
and U21037 (N_21037,N_20916,N_20988);
xnor U21038 (N_21038,N_20593,N_20868);
and U21039 (N_21039,N_20665,N_20960);
xor U21040 (N_21040,N_20582,N_20814);
xnor U21041 (N_21041,N_20860,N_20776);
nand U21042 (N_21042,N_20539,N_20992);
xor U21043 (N_21043,N_20752,N_20870);
nand U21044 (N_21044,N_20605,N_20571);
nor U21045 (N_21045,N_20829,N_20943);
nand U21046 (N_21046,N_20512,N_20801);
or U21047 (N_21047,N_20687,N_20792);
nand U21048 (N_21048,N_20574,N_20562);
and U21049 (N_21049,N_20827,N_20656);
or U21050 (N_21050,N_20950,N_20611);
xnor U21051 (N_21051,N_20869,N_20652);
or U21052 (N_21052,N_20614,N_20983);
xor U21053 (N_21053,N_20842,N_20709);
nor U21054 (N_21054,N_20840,N_20721);
nor U21055 (N_21055,N_20785,N_20816);
nand U21056 (N_21056,N_20841,N_20937);
nor U21057 (N_21057,N_20630,N_20736);
or U21058 (N_21058,N_20787,N_20961);
or U21059 (N_21059,N_20720,N_20525);
xnor U21060 (N_21060,N_20873,N_20956);
and U21061 (N_21061,N_20531,N_20903);
nor U21062 (N_21062,N_20628,N_20508);
xnor U21063 (N_21063,N_20954,N_20631);
and U21064 (N_21064,N_20884,N_20739);
nand U21065 (N_21065,N_20566,N_20671);
xor U21066 (N_21066,N_20749,N_20673);
and U21067 (N_21067,N_20810,N_20510);
nor U21068 (N_21068,N_20995,N_20955);
and U21069 (N_21069,N_20844,N_20748);
and U21070 (N_21070,N_20642,N_20596);
xnor U21071 (N_21071,N_20880,N_20901);
nand U21072 (N_21072,N_20760,N_20660);
and U21073 (N_21073,N_20679,N_20537);
and U21074 (N_21074,N_20608,N_20545);
or U21075 (N_21075,N_20882,N_20770);
or U21076 (N_21076,N_20507,N_20725);
xnor U21077 (N_21077,N_20526,N_20885);
and U21078 (N_21078,N_20570,N_20681);
nor U21079 (N_21079,N_20971,N_20958);
xnor U21080 (N_21080,N_20584,N_20784);
xor U21081 (N_21081,N_20620,N_20824);
nor U21082 (N_21082,N_20558,N_20936);
nand U21083 (N_21083,N_20705,N_20823);
nand U21084 (N_21084,N_20603,N_20606);
nand U21085 (N_21085,N_20849,N_20986);
xor U21086 (N_21086,N_20985,N_20858);
nand U21087 (N_21087,N_20909,N_20676);
or U21088 (N_21088,N_20775,N_20528);
nand U21089 (N_21089,N_20815,N_20598);
nand U21090 (N_21090,N_20848,N_20672);
nand U21091 (N_21091,N_20662,N_20921);
nor U21092 (N_21092,N_20978,N_20668);
xnor U21093 (N_21093,N_20621,N_20949);
nor U21094 (N_21094,N_20649,N_20762);
nor U21095 (N_21095,N_20800,N_20908);
xnor U21096 (N_21096,N_20688,N_20789);
xnor U21097 (N_21097,N_20898,N_20993);
xor U21098 (N_21098,N_20741,N_20900);
nor U21099 (N_21099,N_20811,N_20615);
nand U21100 (N_21100,N_20948,N_20694);
xor U21101 (N_21101,N_20890,N_20894);
xnor U21102 (N_21102,N_20891,N_20561);
nand U21103 (N_21103,N_20533,N_20714);
and U21104 (N_21104,N_20549,N_20808);
nand U21105 (N_21105,N_20521,N_20689);
nand U21106 (N_21106,N_20786,N_20589);
xnor U21107 (N_21107,N_20790,N_20996);
nand U21108 (N_21108,N_20711,N_20722);
nor U21109 (N_21109,N_20999,N_20966);
and U21110 (N_21110,N_20822,N_20889);
and U21111 (N_21111,N_20892,N_20907);
xnor U21112 (N_21112,N_20703,N_20919);
nand U21113 (N_21113,N_20929,N_20503);
or U21114 (N_21114,N_20754,N_20706);
and U21115 (N_21115,N_20796,N_20515);
nor U21116 (N_21116,N_20583,N_20836);
and U21117 (N_21117,N_20540,N_20700);
xor U21118 (N_21118,N_20857,N_20607);
xor U21119 (N_21119,N_20744,N_20831);
and U21120 (N_21120,N_20695,N_20740);
or U21121 (N_21121,N_20832,N_20871);
nor U21122 (N_21122,N_20612,N_20872);
or U21123 (N_21123,N_20579,N_20809);
nand U21124 (N_21124,N_20933,N_20779);
or U21125 (N_21125,N_20707,N_20699);
or U21126 (N_21126,N_20874,N_20718);
and U21127 (N_21127,N_20588,N_20506);
and U21128 (N_21128,N_20538,N_20732);
nand U21129 (N_21129,N_20653,N_20523);
or U21130 (N_21130,N_20536,N_20514);
nor U21131 (N_21131,N_20876,N_20576);
nor U21132 (N_21132,N_20813,N_20728);
nor U21133 (N_21133,N_20622,N_20569);
or U21134 (N_21134,N_20975,N_20553);
or U21135 (N_21135,N_20856,N_20658);
or U21136 (N_21136,N_20980,N_20804);
nor U21137 (N_21137,N_20843,N_20793);
and U21138 (N_21138,N_20633,N_20575);
or U21139 (N_21139,N_20723,N_20670);
nor U21140 (N_21140,N_20987,N_20604);
and U21141 (N_21141,N_20551,N_20644);
nor U21142 (N_21142,N_20738,N_20984);
xor U21143 (N_21143,N_20712,N_20917);
nand U21144 (N_21144,N_20952,N_20964);
nor U21145 (N_21145,N_20686,N_20592);
and U21146 (N_21146,N_20897,N_20654);
nand U21147 (N_21147,N_20685,N_20780);
nand U21148 (N_21148,N_20940,N_20938);
and U21149 (N_21149,N_20500,N_20807);
nor U21150 (N_21150,N_20624,N_20701);
nor U21151 (N_21151,N_20772,N_20852);
nand U21152 (N_21152,N_20519,N_20666);
and U21153 (N_21153,N_20717,N_20990);
and U21154 (N_21154,N_20934,N_20639);
nand U21155 (N_21155,N_20965,N_20918);
and U21156 (N_21156,N_20959,N_20501);
nand U21157 (N_21157,N_20573,N_20683);
and U21158 (N_21158,N_20682,N_20991);
xnor U21159 (N_21159,N_20915,N_20957);
or U21160 (N_21160,N_20866,N_20930);
or U21161 (N_21161,N_20577,N_20963);
xnor U21162 (N_21162,N_20751,N_20733);
xnor U21163 (N_21163,N_20602,N_20618);
xnor U21164 (N_21164,N_20953,N_20632);
nor U21165 (N_21165,N_20636,N_20517);
or U21166 (N_21166,N_20989,N_20661);
nor U21167 (N_21167,N_20973,N_20557);
nor U21168 (N_21168,N_20941,N_20771);
nor U21169 (N_21169,N_20730,N_20839);
or U21170 (N_21170,N_20773,N_20914);
nor U21171 (N_21171,N_20731,N_20926);
nand U21172 (N_21172,N_20591,N_20886);
xor U21173 (N_21173,N_20928,N_20899);
or U21174 (N_21174,N_20502,N_20643);
and U21175 (N_21175,N_20834,N_20845);
nand U21176 (N_21176,N_20743,N_20559);
and U21177 (N_21177,N_20595,N_20710);
nor U21178 (N_21178,N_20659,N_20920);
nand U21179 (N_21179,N_20803,N_20702);
nor U21180 (N_21180,N_20906,N_20704);
or U21181 (N_21181,N_20680,N_20968);
and U21182 (N_21182,N_20931,N_20669);
xor U21183 (N_21183,N_20764,N_20594);
xnor U21184 (N_21184,N_20925,N_20767);
or U21185 (N_21185,N_20805,N_20578);
nand U21186 (N_21186,N_20504,N_20610);
xnor U21187 (N_21187,N_20590,N_20947);
and U21188 (N_21188,N_20724,N_20826);
nand U21189 (N_21189,N_20855,N_20678);
xnor U21190 (N_21190,N_20647,N_20924);
or U21191 (N_21191,N_20623,N_20674);
nor U21192 (N_21192,N_20974,N_20629);
xor U21193 (N_21193,N_20944,N_20769);
and U21194 (N_21194,N_20912,N_20609);
nand U21195 (N_21195,N_20757,N_20726);
nor U21196 (N_21196,N_20761,N_20788);
or U21197 (N_21197,N_20962,N_20600);
and U21198 (N_21198,N_20580,N_20946);
and U21199 (N_21199,N_20613,N_20846);
nand U21200 (N_21200,N_20747,N_20781);
nor U21201 (N_21201,N_20759,N_20904);
or U21202 (N_21202,N_20998,N_20802);
nor U21203 (N_21203,N_20541,N_20572);
or U21204 (N_21204,N_20902,N_20753);
nand U21205 (N_21205,N_20756,N_20861);
xor U21206 (N_21206,N_20835,N_20693);
nor U21207 (N_21207,N_20854,N_20516);
nor U21208 (N_21208,N_20820,N_20878);
nor U21209 (N_21209,N_20969,N_20543);
nor U21210 (N_21210,N_20532,N_20617);
nor U21211 (N_21211,N_20645,N_20667);
xor U21212 (N_21212,N_20534,N_20505);
nor U21213 (N_21213,N_20812,N_20750);
xnor U21214 (N_21214,N_20777,N_20932);
and U21215 (N_21215,N_20737,N_20879);
nor U21216 (N_21216,N_20994,N_20690);
nand U21217 (N_21217,N_20821,N_20939);
or U21218 (N_21218,N_20768,N_20550);
nor U21219 (N_21219,N_20833,N_20859);
nand U21220 (N_21220,N_20979,N_20691);
xnor U21221 (N_21221,N_20951,N_20745);
nor U21222 (N_21222,N_20742,N_20763);
and U21223 (N_21223,N_20535,N_20675);
nand U21224 (N_21224,N_20560,N_20655);
xor U21225 (N_21225,N_20509,N_20520);
xnor U21226 (N_21226,N_20638,N_20616);
and U21227 (N_21227,N_20641,N_20637);
xnor U21228 (N_21228,N_20713,N_20923);
xnor U21229 (N_21229,N_20888,N_20727);
nand U21230 (N_21230,N_20640,N_20518);
or U21231 (N_21231,N_20875,N_20981);
xnor U21232 (N_21232,N_20554,N_20601);
and U21233 (N_21233,N_20635,N_20797);
nand U21234 (N_21234,N_20657,N_20755);
or U21235 (N_21235,N_20697,N_20556);
or U21236 (N_21236,N_20765,N_20626);
and U21237 (N_21237,N_20646,N_20819);
xnor U21238 (N_21238,N_20795,N_20799);
xor U21239 (N_21239,N_20734,N_20913);
xor U21240 (N_21240,N_20766,N_20911);
nor U21241 (N_21241,N_20735,N_20867);
nand U21242 (N_21242,N_20927,N_20746);
xnor U21243 (N_21243,N_20862,N_20530);
nand U21244 (N_21244,N_20708,N_20524);
nor U21245 (N_21245,N_20567,N_20648);
nor U21246 (N_21246,N_20529,N_20942);
or U21247 (N_21247,N_20542,N_20564);
xnor U21248 (N_21248,N_20778,N_20976);
or U21249 (N_21249,N_20817,N_20597);
nand U21250 (N_21250,N_20903,N_20696);
nand U21251 (N_21251,N_20595,N_20754);
nor U21252 (N_21252,N_20941,N_20989);
nand U21253 (N_21253,N_20855,N_20877);
xor U21254 (N_21254,N_20865,N_20755);
and U21255 (N_21255,N_20757,N_20880);
or U21256 (N_21256,N_20615,N_20707);
nor U21257 (N_21257,N_20650,N_20992);
nor U21258 (N_21258,N_20691,N_20779);
nor U21259 (N_21259,N_20588,N_20935);
and U21260 (N_21260,N_20644,N_20589);
nor U21261 (N_21261,N_20584,N_20915);
and U21262 (N_21262,N_20606,N_20912);
nand U21263 (N_21263,N_20986,N_20770);
nor U21264 (N_21264,N_20553,N_20840);
xor U21265 (N_21265,N_20684,N_20619);
xor U21266 (N_21266,N_20960,N_20520);
or U21267 (N_21267,N_20610,N_20593);
or U21268 (N_21268,N_20802,N_20716);
nand U21269 (N_21269,N_20731,N_20767);
nor U21270 (N_21270,N_20635,N_20819);
xor U21271 (N_21271,N_20882,N_20586);
xor U21272 (N_21272,N_20829,N_20997);
or U21273 (N_21273,N_20625,N_20821);
or U21274 (N_21274,N_20993,N_20641);
or U21275 (N_21275,N_20502,N_20637);
xnor U21276 (N_21276,N_20801,N_20584);
nand U21277 (N_21277,N_20832,N_20997);
xnor U21278 (N_21278,N_20795,N_20760);
or U21279 (N_21279,N_20956,N_20787);
xor U21280 (N_21280,N_20561,N_20735);
and U21281 (N_21281,N_20675,N_20944);
xor U21282 (N_21282,N_20938,N_20656);
or U21283 (N_21283,N_20823,N_20693);
and U21284 (N_21284,N_20642,N_20632);
and U21285 (N_21285,N_20709,N_20544);
nand U21286 (N_21286,N_20509,N_20500);
nand U21287 (N_21287,N_20607,N_20606);
xnor U21288 (N_21288,N_20549,N_20510);
or U21289 (N_21289,N_20885,N_20611);
nand U21290 (N_21290,N_20559,N_20564);
nor U21291 (N_21291,N_20502,N_20746);
xnor U21292 (N_21292,N_20531,N_20611);
nor U21293 (N_21293,N_20718,N_20771);
xor U21294 (N_21294,N_20946,N_20795);
nand U21295 (N_21295,N_20984,N_20937);
nand U21296 (N_21296,N_20788,N_20826);
or U21297 (N_21297,N_20926,N_20888);
nor U21298 (N_21298,N_20670,N_20712);
nand U21299 (N_21299,N_20584,N_20953);
and U21300 (N_21300,N_20731,N_20865);
or U21301 (N_21301,N_20536,N_20734);
xnor U21302 (N_21302,N_20597,N_20576);
and U21303 (N_21303,N_20922,N_20994);
and U21304 (N_21304,N_20845,N_20507);
xnor U21305 (N_21305,N_20763,N_20552);
xnor U21306 (N_21306,N_20515,N_20811);
or U21307 (N_21307,N_20794,N_20592);
nor U21308 (N_21308,N_20706,N_20561);
and U21309 (N_21309,N_20728,N_20543);
nand U21310 (N_21310,N_20606,N_20719);
nand U21311 (N_21311,N_20655,N_20961);
or U21312 (N_21312,N_20991,N_20938);
nor U21313 (N_21313,N_20831,N_20976);
xnor U21314 (N_21314,N_20505,N_20736);
or U21315 (N_21315,N_20977,N_20856);
xor U21316 (N_21316,N_20962,N_20841);
xnor U21317 (N_21317,N_20931,N_20735);
and U21318 (N_21318,N_20637,N_20658);
and U21319 (N_21319,N_20624,N_20687);
nor U21320 (N_21320,N_20993,N_20560);
or U21321 (N_21321,N_20614,N_20744);
or U21322 (N_21322,N_20887,N_20525);
and U21323 (N_21323,N_20947,N_20607);
and U21324 (N_21324,N_20855,N_20985);
and U21325 (N_21325,N_20833,N_20552);
and U21326 (N_21326,N_20933,N_20594);
xor U21327 (N_21327,N_20843,N_20825);
nand U21328 (N_21328,N_20559,N_20764);
xor U21329 (N_21329,N_20744,N_20571);
nor U21330 (N_21330,N_20666,N_20729);
and U21331 (N_21331,N_20868,N_20988);
nand U21332 (N_21332,N_20520,N_20925);
nand U21333 (N_21333,N_20772,N_20837);
or U21334 (N_21334,N_20574,N_20850);
and U21335 (N_21335,N_20957,N_20932);
and U21336 (N_21336,N_20581,N_20755);
nor U21337 (N_21337,N_20975,N_20609);
nor U21338 (N_21338,N_20658,N_20821);
and U21339 (N_21339,N_20795,N_20729);
xnor U21340 (N_21340,N_20879,N_20943);
and U21341 (N_21341,N_20504,N_20763);
nor U21342 (N_21342,N_20674,N_20504);
and U21343 (N_21343,N_20898,N_20699);
or U21344 (N_21344,N_20725,N_20874);
or U21345 (N_21345,N_20708,N_20937);
nor U21346 (N_21346,N_20862,N_20805);
nand U21347 (N_21347,N_20603,N_20999);
nand U21348 (N_21348,N_20524,N_20580);
xor U21349 (N_21349,N_20551,N_20850);
or U21350 (N_21350,N_20885,N_20898);
nor U21351 (N_21351,N_20833,N_20712);
or U21352 (N_21352,N_20515,N_20607);
and U21353 (N_21353,N_20843,N_20683);
nand U21354 (N_21354,N_20818,N_20828);
and U21355 (N_21355,N_20720,N_20518);
nand U21356 (N_21356,N_20927,N_20540);
nor U21357 (N_21357,N_20747,N_20531);
and U21358 (N_21358,N_20503,N_20734);
nand U21359 (N_21359,N_20737,N_20936);
and U21360 (N_21360,N_20533,N_20663);
nor U21361 (N_21361,N_20660,N_20842);
nor U21362 (N_21362,N_20766,N_20915);
xor U21363 (N_21363,N_20777,N_20756);
nand U21364 (N_21364,N_20597,N_20863);
or U21365 (N_21365,N_20918,N_20874);
xnor U21366 (N_21366,N_20770,N_20693);
nand U21367 (N_21367,N_20765,N_20658);
or U21368 (N_21368,N_20843,N_20745);
and U21369 (N_21369,N_20564,N_20782);
nand U21370 (N_21370,N_20665,N_20939);
or U21371 (N_21371,N_20959,N_20567);
or U21372 (N_21372,N_20902,N_20798);
nor U21373 (N_21373,N_20910,N_20927);
xor U21374 (N_21374,N_20649,N_20615);
nor U21375 (N_21375,N_20842,N_20744);
nor U21376 (N_21376,N_20689,N_20926);
or U21377 (N_21377,N_20607,N_20635);
or U21378 (N_21378,N_20951,N_20833);
nor U21379 (N_21379,N_20886,N_20877);
nor U21380 (N_21380,N_20580,N_20897);
or U21381 (N_21381,N_20647,N_20979);
or U21382 (N_21382,N_20665,N_20556);
nor U21383 (N_21383,N_20927,N_20757);
nand U21384 (N_21384,N_20574,N_20634);
nand U21385 (N_21385,N_20773,N_20850);
xor U21386 (N_21386,N_20622,N_20728);
xor U21387 (N_21387,N_20815,N_20957);
nand U21388 (N_21388,N_20750,N_20830);
xnor U21389 (N_21389,N_20573,N_20828);
or U21390 (N_21390,N_20976,N_20783);
nor U21391 (N_21391,N_20937,N_20948);
nor U21392 (N_21392,N_20514,N_20755);
nor U21393 (N_21393,N_20570,N_20733);
or U21394 (N_21394,N_20757,N_20982);
or U21395 (N_21395,N_20509,N_20757);
nor U21396 (N_21396,N_20976,N_20769);
and U21397 (N_21397,N_20879,N_20597);
nand U21398 (N_21398,N_20786,N_20701);
or U21399 (N_21399,N_20997,N_20547);
or U21400 (N_21400,N_20822,N_20666);
and U21401 (N_21401,N_20644,N_20960);
and U21402 (N_21402,N_20516,N_20900);
xnor U21403 (N_21403,N_20838,N_20517);
nand U21404 (N_21404,N_20645,N_20627);
nor U21405 (N_21405,N_20829,N_20930);
or U21406 (N_21406,N_20945,N_20572);
and U21407 (N_21407,N_20599,N_20646);
xor U21408 (N_21408,N_20530,N_20585);
nor U21409 (N_21409,N_20839,N_20745);
or U21410 (N_21410,N_20654,N_20521);
nand U21411 (N_21411,N_20626,N_20729);
nor U21412 (N_21412,N_20955,N_20663);
nand U21413 (N_21413,N_20987,N_20969);
nand U21414 (N_21414,N_20593,N_20516);
nand U21415 (N_21415,N_20856,N_20883);
and U21416 (N_21416,N_20535,N_20522);
and U21417 (N_21417,N_20607,N_20866);
nor U21418 (N_21418,N_20828,N_20641);
nor U21419 (N_21419,N_20525,N_20882);
nand U21420 (N_21420,N_20701,N_20872);
nand U21421 (N_21421,N_20790,N_20906);
xnor U21422 (N_21422,N_20824,N_20902);
xor U21423 (N_21423,N_20777,N_20906);
xor U21424 (N_21424,N_20932,N_20939);
xor U21425 (N_21425,N_20918,N_20605);
nand U21426 (N_21426,N_20644,N_20720);
and U21427 (N_21427,N_20579,N_20572);
and U21428 (N_21428,N_20701,N_20673);
xnor U21429 (N_21429,N_20711,N_20595);
xor U21430 (N_21430,N_20952,N_20677);
xnor U21431 (N_21431,N_20562,N_20968);
nand U21432 (N_21432,N_20869,N_20794);
or U21433 (N_21433,N_20756,N_20713);
nand U21434 (N_21434,N_20963,N_20869);
nor U21435 (N_21435,N_20995,N_20935);
nand U21436 (N_21436,N_20794,N_20747);
nand U21437 (N_21437,N_20634,N_20745);
xor U21438 (N_21438,N_20623,N_20836);
nor U21439 (N_21439,N_20633,N_20609);
xnor U21440 (N_21440,N_20732,N_20560);
or U21441 (N_21441,N_20524,N_20774);
nor U21442 (N_21442,N_20881,N_20645);
nor U21443 (N_21443,N_20581,N_20741);
or U21444 (N_21444,N_20978,N_20598);
xor U21445 (N_21445,N_20956,N_20692);
nand U21446 (N_21446,N_20722,N_20743);
nand U21447 (N_21447,N_20933,N_20832);
nor U21448 (N_21448,N_20909,N_20910);
xnor U21449 (N_21449,N_20797,N_20643);
and U21450 (N_21450,N_20552,N_20721);
nor U21451 (N_21451,N_20842,N_20611);
and U21452 (N_21452,N_20957,N_20838);
or U21453 (N_21453,N_20744,N_20996);
nor U21454 (N_21454,N_20923,N_20799);
or U21455 (N_21455,N_20562,N_20981);
nor U21456 (N_21456,N_20816,N_20985);
or U21457 (N_21457,N_20528,N_20937);
and U21458 (N_21458,N_20554,N_20634);
nor U21459 (N_21459,N_20648,N_20847);
or U21460 (N_21460,N_20760,N_20703);
or U21461 (N_21461,N_20945,N_20847);
nand U21462 (N_21462,N_20527,N_20800);
xnor U21463 (N_21463,N_20892,N_20657);
and U21464 (N_21464,N_20692,N_20795);
and U21465 (N_21465,N_20508,N_20834);
nor U21466 (N_21466,N_20603,N_20767);
or U21467 (N_21467,N_20877,N_20604);
or U21468 (N_21468,N_20929,N_20793);
or U21469 (N_21469,N_20875,N_20883);
xnor U21470 (N_21470,N_20692,N_20787);
nand U21471 (N_21471,N_20706,N_20655);
or U21472 (N_21472,N_20943,N_20736);
xor U21473 (N_21473,N_20503,N_20748);
nor U21474 (N_21474,N_20956,N_20774);
nor U21475 (N_21475,N_20573,N_20894);
nand U21476 (N_21476,N_20701,N_20615);
or U21477 (N_21477,N_20965,N_20701);
nor U21478 (N_21478,N_20741,N_20728);
nor U21479 (N_21479,N_20939,N_20996);
xnor U21480 (N_21480,N_20819,N_20663);
nor U21481 (N_21481,N_20505,N_20974);
or U21482 (N_21482,N_20927,N_20741);
or U21483 (N_21483,N_20636,N_20909);
nand U21484 (N_21484,N_20847,N_20851);
xor U21485 (N_21485,N_20983,N_20699);
nand U21486 (N_21486,N_20951,N_20549);
xnor U21487 (N_21487,N_20881,N_20742);
xnor U21488 (N_21488,N_20710,N_20826);
xor U21489 (N_21489,N_20886,N_20876);
or U21490 (N_21490,N_20996,N_20517);
nand U21491 (N_21491,N_20693,N_20750);
and U21492 (N_21492,N_20592,N_20923);
xor U21493 (N_21493,N_20890,N_20990);
or U21494 (N_21494,N_20707,N_20730);
xor U21495 (N_21495,N_20846,N_20783);
nand U21496 (N_21496,N_20536,N_20972);
xor U21497 (N_21497,N_20653,N_20740);
nand U21498 (N_21498,N_20787,N_20746);
nand U21499 (N_21499,N_20594,N_20756);
or U21500 (N_21500,N_21496,N_21456);
or U21501 (N_21501,N_21485,N_21223);
nand U21502 (N_21502,N_21240,N_21470);
and U21503 (N_21503,N_21398,N_21077);
nor U21504 (N_21504,N_21466,N_21012);
nor U21505 (N_21505,N_21126,N_21402);
nand U21506 (N_21506,N_21182,N_21306);
nor U21507 (N_21507,N_21432,N_21028);
nand U21508 (N_21508,N_21053,N_21147);
nor U21509 (N_21509,N_21097,N_21285);
and U21510 (N_21510,N_21139,N_21146);
and U21511 (N_21511,N_21125,N_21294);
nand U21512 (N_21512,N_21277,N_21207);
nor U21513 (N_21513,N_21250,N_21027);
and U21514 (N_21514,N_21368,N_21450);
xor U21515 (N_21515,N_21347,N_21406);
nor U21516 (N_21516,N_21312,N_21313);
and U21517 (N_21517,N_21006,N_21002);
xor U21518 (N_21518,N_21167,N_21117);
or U21519 (N_21519,N_21248,N_21445);
nand U21520 (N_21520,N_21155,N_21314);
or U21521 (N_21521,N_21113,N_21369);
nor U21522 (N_21522,N_21258,N_21441);
nand U21523 (N_21523,N_21089,N_21462);
or U21524 (N_21524,N_21142,N_21279);
nor U21525 (N_21525,N_21290,N_21330);
or U21526 (N_21526,N_21409,N_21246);
nor U21527 (N_21527,N_21032,N_21423);
or U21528 (N_21528,N_21088,N_21080);
nand U21529 (N_21529,N_21137,N_21448);
xor U21530 (N_21530,N_21299,N_21498);
or U21531 (N_21531,N_21245,N_21127);
xnor U21532 (N_21532,N_21220,N_21405);
nor U21533 (N_21533,N_21106,N_21070);
and U21534 (N_21534,N_21394,N_21284);
nor U21535 (N_21535,N_21380,N_21172);
xor U21536 (N_21536,N_21252,N_21309);
nor U21537 (N_21537,N_21046,N_21278);
xnor U21538 (N_21538,N_21339,N_21084);
nand U21539 (N_21539,N_21224,N_21271);
nor U21540 (N_21540,N_21098,N_21192);
nand U21541 (N_21541,N_21283,N_21040);
and U21542 (N_21542,N_21011,N_21363);
nor U21543 (N_21543,N_21030,N_21442);
and U21544 (N_21544,N_21161,N_21204);
xor U21545 (N_21545,N_21103,N_21352);
and U21546 (N_21546,N_21034,N_21232);
xnor U21547 (N_21547,N_21473,N_21397);
or U21548 (N_21548,N_21023,N_21244);
or U21549 (N_21549,N_21020,N_21047);
nand U21550 (N_21550,N_21326,N_21391);
and U21551 (N_21551,N_21014,N_21188);
nor U21552 (N_21552,N_21367,N_21447);
or U21553 (N_21553,N_21395,N_21385);
and U21554 (N_21554,N_21476,N_21428);
and U21555 (N_21555,N_21136,N_21334);
nand U21556 (N_21556,N_21481,N_21381);
xnor U21557 (N_21557,N_21133,N_21486);
nand U21558 (N_21558,N_21375,N_21200);
and U21559 (N_21559,N_21179,N_21067);
nor U21560 (N_21560,N_21357,N_21229);
or U21561 (N_21561,N_21305,N_21256);
and U21562 (N_21562,N_21328,N_21396);
xor U21563 (N_21563,N_21162,N_21453);
xor U21564 (N_21564,N_21490,N_21164);
nand U21565 (N_21565,N_21063,N_21230);
nand U21566 (N_21566,N_21303,N_21355);
or U21567 (N_21567,N_21377,N_21298);
nor U21568 (N_21568,N_21071,N_21425);
nand U21569 (N_21569,N_21109,N_21110);
xnor U21570 (N_21570,N_21132,N_21376);
or U21571 (N_21571,N_21190,N_21181);
xor U21572 (N_21572,N_21078,N_21015);
nor U21573 (N_21573,N_21141,N_21185);
nor U21574 (N_21574,N_21460,N_21083);
nand U21575 (N_21575,N_21482,N_21016);
xor U21576 (N_21576,N_21356,N_21241);
nor U21577 (N_21577,N_21461,N_21079);
nand U21578 (N_21578,N_21307,N_21024);
nor U21579 (N_21579,N_21198,N_21492);
and U21580 (N_21580,N_21493,N_21433);
or U21581 (N_21581,N_21175,N_21327);
nand U21582 (N_21582,N_21050,N_21257);
xor U21583 (N_21583,N_21060,N_21178);
nand U21584 (N_21584,N_21472,N_21003);
or U21585 (N_21585,N_21295,N_21095);
or U21586 (N_21586,N_21411,N_21426);
nand U21587 (N_21587,N_21177,N_21101);
nand U21588 (N_21588,N_21215,N_21051);
and U21589 (N_21589,N_21421,N_21158);
nor U21590 (N_21590,N_21499,N_21238);
and U21591 (N_21591,N_21281,N_21171);
nor U21592 (N_21592,N_21082,N_21276);
nand U21593 (N_21593,N_21350,N_21165);
nand U21594 (N_21594,N_21389,N_21086);
or U21595 (N_21595,N_21297,N_21249);
and U21596 (N_21596,N_21143,N_21388);
xor U21597 (N_21597,N_21324,N_21475);
xnor U21598 (N_21598,N_21316,N_21152);
and U21599 (N_21599,N_21222,N_21173);
or U21600 (N_21600,N_21315,N_21464);
xor U21601 (N_21601,N_21069,N_21438);
or U21602 (N_21602,N_21452,N_21008);
nor U21603 (N_21603,N_21058,N_21302);
and U21604 (N_21604,N_21468,N_21214);
and U21605 (N_21605,N_21065,N_21251);
or U21606 (N_21606,N_21168,N_21081);
nand U21607 (N_21607,N_21203,N_21404);
xnor U21608 (N_21608,N_21189,N_21195);
xnor U21609 (N_21609,N_21123,N_21108);
nor U21610 (N_21610,N_21044,N_21226);
nand U21611 (N_21611,N_21212,N_21427);
nor U21612 (N_21612,N_21231,N_21469);
xor U21613 (N_21613,N_21237,N_21366);
and U21614 (N_21614,N_21094,N_21444);
nor U21615 (N_21615,N_21085,N_21193);
nand U21616 (N_21616,N_21041,N_21134);
nor U21617 (N_21617,N_21009,N_21199);
xnor U21618 (N_21618,N_21340,N_21383);
nand U21619 (N_21619,N_21497,N_21037);
or U21620 (N_21620,N_21112,N_21410);
nand U21621 (N_21621,N_21415,N_21436);
xnor U21622 (N_21622,N_21273,N_21039);
nand U21623 (N_21623,N_21384,N_21268);
and U21624 (N_21624,N_21477,N_21107);
nor U21625 (N_21625,N_21331,N_21194);
nand U21626 (N_21626,N_21122,N_21239);
nor U21627 (N_21627,N_21073,N_21236);
and U21628 (N_21628,N_21036,N_21262);
nor U21629 (N_21629,N_21437,N_21054);
and U21630 (N_21630,N_21004,N_21018);
nor U21631 (N_21631,N_21272,N_21131);
and U21632 (N_21632,N_21035,N_21120);
nand U21633 (N_21633,N_21105,N_21156);
and U21634 (N_21634,N_21337,N_21260);
and U21635 (N_21635,N_21042,N_21099);
or U21636 (N_21636,N_21286,N_21414);
and U21637 (N_21637,N_21412,N_21048);
nor U21638 (N_21638,N_21019,N_21010);
and U21639 (N_21639,N_21234,N_21259);
nand U21640 (N_21640,N_21253,N_21187);
and U21641 (N_21641,N_21225,N_21480);
nand U21642 (N_21642,N_21227,N_21379);
or U21643 (N_21643,N_21254,N_21049);
xnor U21644 (N_21644,N_21293,N_21373);
and U21645 (N_21645,N_21282,N_21043);
xor U21646 (N_21646,N_21184,N_21288);
nor U21647 (N_21647,N_21311,N_21062);
or U21648 (N_21648,N_21364,N_21458);
nor U21649 (N_21649,N_21300,N_21144);
nor U21650 (N_21650,N_21275,N_21341);
nor U21651 (N_21651,N_21055,N_21335);
and U21652 (N_21652,N_21233,N_21361);
and U21653 (N_21653,N_21483,N_21176);
nor U21654 (N_21654,N_21348,N_21209);
nor U21655 (N_21655,N_21093,N_21129);
and U21656 (N_21656,N_21374,N_21145);
nand U21657 (N_21657,N_21066,N_21358);
nand U21658 (N_21658,N_21429,N_21274);
nor U21659 (N_21659,N_21205,N_21333);
nand U21660 (N_21660,N_21180,N_21026);
nor U21661 (N_21661,N_21463,N_21217);
or U21662 (N_21662,N_21296,N_21033);
xor U21663 (N_21663,N_21201,N_21092);
xnor U21664 (N_21664,N_21210,N_21163);
xnor U21665 (N_21665,N_21128,N_21159);
or U21666 (N_21666,N_21045,N_21439);
and U21667 (N_21667,N_21100,N_21074);
xnor U21668 (N_21668,N_21365,N_21455);
xor U21669 (N_21669,N_21243,N_21495);
or U21670 (N_21670,N_21266,N_21301);
xor U21671 (N_21671,N_21076,N_21261);
nand U21672 (N_21672,N_21474,N_21057);
and U21673 (N_21673,N_21321,N_21052);
nor U21674 (N_21674,N_21114,N_21091);
xor U21675 (N_21675,N_21446,N_21005);
or U21676 (N_21676,N_21124,N_21235);
or U21677 (N_21677,N_21007,N_21451);
or U21678 (N_21678,N_21332,N_21135);
nor U21679 (N_21679,N_21216,N_21149);
xnor U21680 (N_21680,N_21292,N_21202);
nor U21681 (N_21681,N_21170,N_21068);
nor U21682 (N_21682,N_21280,N_21401);
xor U21683 (N_21683,N_21443,N_21343);
nor U21684 (N_21684,N_21121,N_21154);
nand U21685 (N_21685,N_21169,N_21319);
xor U21686 (N_21686,N_21387,N_21449);
or U21687 (N_21687,N_21111,N_21392);
nand U21688 (N_21688,N_21420,N_21038);
nand U21689 (N_21689,N_21310,N_21219);
xor U21690 (N_21690,N_21000,N_21064);
and U21691 (N_21691,N_21269,N_21342);
and U21692 (N_21692,N_21228,N_21457);
nand U21693 (N_21693,N_21400,N_21191);
nand U21694 (N_21694,N_21287,N_21072);
nand U21695 (N_21695,N_21317,N_21408);
and U21696 (N_21696,N_21491,N_21403);
nor U21697 (N_21697,N_21407,N_21150);
and U21698 (N_21698,N_21488,N_21075);
or U21699 (N_21699,N_21242,N_21336);
nor U21700 (N_21700,N_21025,N_21160);
nor U21701 (N_21701,N_21130,N_21304);
nand U21702 (N_21702,N_21061,N_21087);
nor U21703 (N_21703,N_21213,N_21265);
or U21704 (N_21704,N_21399,N_21351);
nand U21705 (N_21705,N_21353,N_21386);
nor U21706 (N_21706,N_21320,N_21218);
nand U21707 (N_21707,N_21029,N_21022);
and U21708 (N_21708,N_21056,N_21267);
nor U21709 (N_21709,N_21390,N_21416);
or U21710 (N_21710,N_21489,N_21211);
or U21711 (N_21711,N_21349,N_21354);
or U21712 (N_21712,N_21208,N_21148);
nor U21713 (N_21713,N_21157,N_21440);
xnor U21714 (N_21714,N_21174,N_21059);
nor U21715 (N_21715,N_21318,N_21418);
xor U21716 (N_21716,N_21289,N_21459);
nor U21717 (N_21717,N_21102,N_21494);
and U21718 (N_21718,N_21104,N_21338);
xor U21719 (N_21719,N_21140,N_21291);
nor U21720 (N_21720,N_21153,N_21151);
nand U21721 (N_21721,N_21435,N_21370);
and U21722 (N_21722,N_21308,N_21430);
and U21723 (N_21723,N_21325,N_21345);
or U21724 (N_21724,N_21467,N_21013);
or U21725 (N_21725,N_21479,N_21431);
nor U21726 (N_21726,N_21183,N_21221);
nand U21727 (N_21727,N_21247,N_21264);
and U21728 (N_21728,N_21138,N_21031);
and U21729 (N_21729,N_21001,N_21166);
or U21730 (N_21730,N_21471,N_21362);
nand U21731 (N_21731,N_21413,N_21255);
and U21732 (N_21732,N_21393,N_21454);
or U21733 (N_21733,N_21197,N_21359);
and U21734 (N_21734,N_21382,N_21021);
nand U21735 (N_21735,N_21371,N_21263);
nand U21736 (N_21736,N_21422,N_21478);
nor U21737 (N_21737,N_21419,N_21329);
xor U21738 (N_21738,N_21360,N_21344);
nand U21739 (N_21739,N_21434,N_21346);
or U21740 (N_21740,N_21186,N_21417);
and U21741 (N_21741,N_21323,N_21465);
nand U21742 (N_21742,N_21116,N_21270);
nand U21743 (N_21743,N_21118,N_21372);
xor U21744 (N_21744,N_21424,N_21119);
xnor U21745 (N_21745,N_21206,N_21196);
or U21746 (N_21746,N_21322,N_21115);
nand U21747 (N_21747,N_21487,N_21484);
xnor U21748 (N_21748,N_21017,N_21378);
xor U21749 (N_21749,N_21096,N_21090);
or U21750 (N_21750,N_21384,N_21110);
nor U21751 (N_21751,N_21166,N_21192);
or U21752 (N_21752,N_21020,N_21155);
nor U21753 (N_21753,N_21109,N_21030);
or U21754 (N_21754,N_21291,N_21475);
xnor U21755 (N_21755,N_21034,N_21241);
xor U21756 (N_21756,N_21398,N_21060);
xnor U21757 (N_21757,N_21283,N_21071);
or U21758 (N_21758,N_21022,N_21145);
xor U21759 (N_21759,N_21406,N_21000);
nor U21760 (N_21760,N_21390,N_21344);
and U21761 (N_21761,N_21221,N_21091);
nor U21762 (N_21762,N_21258,N_21233);
nor U21763 (N_21763,N_21023,N_21147);
or U21764 (N_21764,N_21073,N_21445);
nor U21765 (N_21765,N_21256,N_21478);
xnor U21766 (N_21766,N_21333,N_21348);
and U21767 (N_21767,N_21333,N_21365);
nand U21768 (N_21768,N_21349,N_21439);
and U21769 (N_21769,N_21471,N_21185);
xor U21770 (N_21770,N_21300,N_21068);
or U21771 (N_21771,N_21074,N_21194);
and U21772 (N_21772,N_21339,N_21340);
nor U21773 (N_21773,N_21073,N_21377);
nand U21774 (N_21774,N_21412,N_21175);
and U21775 (N_21775,N_21316,N_21320);
nand U21776 (N_21776,N_21406,N_21249);
and U21777 (N_21777,N_21429,N_21276);
nand U21778 (N_21778,N_21090,N_21465);
and U21779 (N_21779,N_21180,N_21137);
nor U21780 (N_21780,N_21154,N_21031);
or U21781 (N_21781,N_21191,N_21423);
nor U21782 (N_21782,N_21210,N_21019);
nor U21783 (N_21783,N_21352,N_21016);
nor U21784 (N_21784,N_21098,N_21410);
or U21785 (N_21785,N_21000,N_21410);
or U21786 (N_21786,N_21205,N_21035);
and U21787 (N_21787,N_21089,N_21012);
xor U21788 (N_21788,N_21394,N_21051);
nor U21789 (N_21789,N_21354,N_21325);
or U21790 (N_21790,N_21454,N_21301);
and U21791 (N_21791,N_21394,N_21428);
or U21792 (N_21792,N_21117,N_21137);
and U21793 (N_21793,N_21174,N_21062);
or U21794 (N_21794,N_21012,N_21122);
xnor U21795 (N_21795,N_21278,N_21115);
nor U21796 (N_21796,N_21295,N_21185);
nand U21797 (N_21797,N_21418,N_21325);
or U21798 (N_21798,N_21076,N_21090);
or U21799 (N_21799,N_21411,N_21473);
nand U21800 (N_21800,N_21378,N_21037);
and U21801 (N_21801,N_21381,N_21288);
and U21802 (N_21802,N_21012,N_21028);
and U21803 (N_21803,N_21308,N_21075);
nand U21804 (N_21804,N_21478,N_21058);
nor U21805 (N_21805,N_21068,N_21375);
nor U21806 (N_21806,N_21331,N_21021);
xor U21807 (N_21807,N_21146,N_21332);
nand U21808 (N_21808,N_21193,N_21307);
xor U21809 (N_21809,N_21145,N_21126);
or U21810 (N_21810,N_21120,N_21476);
nor U21811 (N_21811,N_21409,N_21312);
nor U21812 (N_21812,N_21086,N_21246);
and U21813 (N_21813,N_21265,N_21015);
nand U21814 (N_21814,N_21151,N_21421);
nand U21815 (N_21815,N_21465,N_21369);
and U21816 (N_21816,N_21314,N_21409);
xor U21817 (N_21817,N_21231,N_21318);
nor U21818 (N_21818,N_21451,N_21182);
nor U21819 (N_21819,N_21408,N_21197);
nor U21820 (N_21820,N_21355,N_21109);
xnor U21821 (N_21821,N_21077,N_21034);
nor U21822 (N_21822,N_21121,N_21497);
nor U21823 (N_21823,N_21424,N_21111);
and U21824 (N_21824,N_21146,N_21069);
and U21825 (N_21825,N_21478,N_21297);
xnor U21826 (N_21826,N_21240,N_21227);
nand U21827 (N_21827,N_21106,N_21002);
nand U21828 (N_21828,N_21099,N_21337);
xor U21829 (N_21829,N_21097,N_21253);
xor U21830 (N_21830,N_21493,N_21418);
or U21831 (N_21831,N_21431,N_21370);
nor U21832 (N_21832,N_21383,N_21001);
and U21833 (N_21833,N_21437,N_21035);
nor U21834 (N_21834,N_21015,N_21278);
nand U21835 (N_21835,N_21369,N_21324);
nor U21836 (N_21836,N_21136,N_21243);
nand U21837 (N_21837,N_21060,N_21326);
or U21838 (N_21838,N_21126,N_21355);
and U21839 (N_21839,N_21134,N_21293);
nor U21840 (N_21840,N_21198,N_21130);
or U21841 (N_21841,N_21338,N_21065);
nor U21842 (N_21842,N_21396,N_21305);
nor U21843 (N_21843,N_21035,N_21092);
nor U21844 (N_21844,N_21480,N_21431);
or U21845 (N_21845,N_21232,N_21176);
nand U21846 (N_21846,N_21443,N_21114);
or U21847 (N_21847,N_21403,N_21266);
nand U21848 (N_21848,N_21101,N_21090);
or U21849 (N_21849,N_21457,N_21307);
and U21850 (N_21850,N_21320,N_21390);
or U21851 (N_21851,N_21161,N_21295);
or U21852 (N_21852,N_21212,N_21241);
xor U21853 (N_21853,N_21204,N_21424);
nand U21854 (N_21854,N_21283,N_21233);
or U21855 (N_21855,N_21076,N_21442);
xnor U21856 (N_21856,N_21060,N_21202);
and U21857 (N_21857,N_21442,N_21321);
and U21858 (N_21858,N_21468,N_21262);
nand U21859 (N_21859,N_21259,N_21284);
and U21860 (N_21860,N_21035,N_21401);
or U21861 (N_21861,N_21114,N_21089);
and U21862 (N_21862,N_21309,N_21468);
and U21863 (N_21863,N_21086,N_21253);
or U21864 (N_21864,N_21068,N_21260);
xnor U21865 (N_21865,N_21415,N_21180);
xor U21866 (N_21866,N_21246,N_21385);
nand U21867 (N_21867,N_21265,N_21473);
nor U21868 (N_21868,N_21391,N_21491);
and U21869 (N_21869,N_21191,N_21353);
nor U21870 (N_21870,N_21227,N_21494);
xor U21871 (N_21871,N_21095,N_21277);
xnor U21872 (N_21872,N_21289,N_21061);
nor U21873 (N_21873,N_21038,N_21484);
xnor U21874 (N_21874,N_21368,N_21473);
xnor U21875 (N_21875,N_21382,N_21336);
and U21876 (N_21876,N_21204,N_21178);
or U21877 (N_21877,N_21486,N_21210);
or U21878 (N_21878,N_21118,N_21289);
nor U21879 (N_21879,N_21112,N_21328);
or U21880 (N_21880,N_21055,N_21334);
xor U21881 (N_21881,N_21448,N_21142);
and U21882 (N_21882,N_21038,N_21210);
and U21883 (N_21883,N_21179,N_21483);
or U21884 (N_21884,N_21443,N_21111);
and U21885 (N_21885,N_21178,N_21010);
xor U21886 (N_21886,N_21314,N_21182);
nand U21887 (N_21887,N_21024,N_21317);
or U21888 (N_21888,N_21250,N_21361);
and U21889 (N_21889,N_21121,N_21294);
nor U21890 (N_21890,N_21424,N_21158);
or U21891 (N_21891,N_21298,N_21323);
or U21892 (N_21892,N_21142,N_21020);
nand U21893 (N_21893,N_21397,N_21015);
nand U21894 (N_21894,N_21235,N_21339);
nand U21895 (N_21895,N_21213,N_21363);
nand U21896 (N_21896,N_21064,N_21239);
or U21897 (N_21897,N_21151,N_21095);
or U21898 (N_21898,N_21048,N_21089);
nand U21899 (N_21899,N_21322,N_21208);
xor U21900 (N_21900,N_21264,N_21461);
nor U21901 (N_21901,N_21274,N_21281);
or U21902 (N_21902,N_21152,N_21051);
and U21903 (N_21903,N_21167,N_21229);
or U21904 (N_21904,N_21397,N_21096);
or U21905 (N_21905,N_21208,N_21218);
or U21906 (N_21906,N_21009,N_21263);
xor U21907 (N_21907,N_21028,N_21374);
or U21908 (N_21908,N_21296,N_21423);
or U21909 (N_21909,N_21401,N_21377);
and U21910 (N_21910,N_21151,N_21258);
or U21911 (N_21911,N_21131,N_21242);
or U21912 (N_21912,N_21114,N_21227);
xnor U21913 (N_21913,N_21287,N_21192);
and U21914 (N_21914,N_21116,N_21415);
nand U21915 (N_21915,N_21188,N_21282);
nor U21916 (N_21916,N_21333,N_21020);
nor U21917 (N_21917,N_21201,N_21057);
and U21918 (N_21918,N_21233,N_21043);
and U21919 (N_21919,N_21451,N_21062);
nor U21920 (N_21920,N_21352,N_21415);
xnor U21921 (N_21921,N_21257,N_21132);
nand U21922 (N_21922,N_21308,N_21201);
nand U21923 (N_21923,N_21435,N_21010);
or U21924 (N_21924,N_21269,N_21067);
nand U21925 (N_21925,N_21456,N_21369);
nor U21926 (N_21926,N_21499,N_21422);
nand U21927 (N_21927,N_21216,N_21026);
nor U21928 (N_21928,N_21053,N_21012);
and U21929 (N_21929,N_21415,N_21427);
or U21930 (N_21930,N_21247,N_21346);
nor U21931 (N_21931,N_21035,N_21399);
nand U21932 (N_21932,N_21063,N_21462);
nand U21933 (N_21933,N_21227,N_21201);
nor U21934 (N_21934,N_21484,N_21319);
nor U21935 (N_21935,N_21014,N_21000);
xor U21936 (N_21936,N_21251,N_21075);
nor U21937 (N_21937,N_21491,N_21421);
nor U21938 (N_21938,N_21424,N_21125);
nor U21939 (N_21939,N_21081,N_21334);
nor U21940 (N_21940,N_21062,N_21406);
xnor U21941 (N_21941,N_21184,N_21258);
nand U21942 (N_21942,N_21459,N_21165);
or U21943 (N_21943,N_21220,N_21093);
xnor U21944 (N_21944,N_21413,N_21169);
or U21945 (N_21945,N_21264,N_21177);
xor U21946 (N_21946,N_21282,N_21355);
or U21947 (N_21947,N_21146,N_21349);
nor U21948 (N_21948,N_21018,N_21152);
and U21949 (N_21949,N_21298,N_21122);
and U21950 (N_21950,N_21386,N_21073);
nand U21951 (N_21951,N_21142,N_21375);
or U21952 (N_21952,N_21237,N_21150);
nand U21953 (N_21953,N_21468,N_21027);
or U21954 (N_21954,N_21274,N_21175);
or U21955 (N_21955,N_21364,N_21007);
nand U21956 (N_21956,N_21251,N_21098);
nand U21957 (N_21957,N_21002,N_21295);
nor U21958 (N_21958,N_21280,N_21415);
or U21959 (N_21959,N_21325,N_21080);
nor U21960 (N_21960,N_21324,N_21041);
nor U21961 (N_21961,N_21257,N_21488);
nand U21962 (N_21962,N_21373,N_21026);
nand U21963 (N_21963,N_21027,N_21489);
nand U21964 (N_21964,N_21375,N_21208);
xor U21965 (N_21965,N_21085,N_21331);
nand U21966 (N_21966,N_21253,N_21310);
xor U21967 (N_21967,N_21362,N_21475);
nor U21968 (N_21968,N_21076,N_21415);
and U21969 (N_21969,N_21043,N_21004);
or U21970 (N_21970,N_21355,N_21444);
xor U21971 (N_21971,N_21435,N_21092);
and U21972 (N_21972,N_21131,N_21361);
nor U21973 (N_21973,N_21358,N_21177);
nor U21974 (N_21974,N_21077,N_21056);
nand U21975 (N_21975,N_21235,N_21121);
nor U21976 (N_21976,N_21430,N_21127);
xor U21977 (N_21977,N_21399,N_21023);
nand U21978 (N_21978,N_21282,N_21453);
nand U21979 (N_21979,N_21177,N_21266);
nor U21980 (N_21980,N_21246,N_21411);
xor U21981 (N_21981,N_21241,N_21475);
and U21982 (N_21982,N_21198,N_21412);
nor U21983 (N_21983,N_21140,N_21360);
nand U21984 (N_21984,N_21185,N_21112);
or U21985 (N_21985,N_21346,N_21366);
xnor U21986 (N_21986,N_21126,N_21499);
nand U21987 (N_21987,N_21127,N_21047);
xnor U21988 (N_21988,N_21270,N_21451);
or U21989 (N_21989,N_21352,N_21027);
nand U21990 (N_21990,N_21251,N_21366);
nand U21991 (N_21991,N_21047,N_21194);
and U21992 (N_21992,N_21134,N_21321);
nor U21993 (N_21993,N_21032,N_21049);
nor U21994 (N_21994,N_21138,N_21269);
nand U21995 (N_21995,N_21011,N_21108);
or U21996 (N_21996,N_21396,N_21392);
nand U21997 (N_21997,N_21409,N_21363);
or U21998 (N_21998,N_21408,N_21445);
or U21999 (N_21999,N_21081,N_21373);
xor U22000 (N_22000,N_21657,N_21926);
and U22001 (N_22001,N_21877,N_21928);
nand U22002 (N_22002,N_21943,N_21907);
nor U22003 (N_22003,N_21705,N_21726);
and U22004 (N_22004,N_21909,N_21857);
and U22005 (N_22005,N_21536,N_21760);
and U22006 (N_22006,N_21501,N_21678);
xor U22007 (N_22007,N_21826,N_21790);
or U22008 (N_22008,N_21891,N_21824);
xor U22009 (N_22009,N_21582,N_21889);
nor U22010 (N_22010,N_21597,N_21932);
and U22011 (N_22011,N_21524,N_21915);
or U22012 (N_22012,N_21789,N_21671);
or U22013 (N_22013,N_21893,N_21853);
or U22014 (N_22014,N_21667,N_21776);
nand U22015 (N_22015,N_21908,N_21901);
and U22016 (N_22016,N_21609,N_21700);
and U22017 (N_22017,N_21920,N_21751);
nand U22018 (N_22018,N_21916,N_21995);
nor U22019 (N_22019,N_21814,N_21544);
nor U22020 (N_22020,N_21587,N_21809);
and U22021 (N_22021,N_21565,N_21762);
and U22022 (N_22022,N_21625,N_21757);
or U22023 (N_22023,N_21887,N_21801);
nand U22024 (N_22024,N_21741,N_21845);
or U22025 (N_22025,N_21729,N_21517);
xor U22026 (N_22026,N_21687,N_21799);
nor U22027 (N_22027,N_21500,N_21616);
nand U22028 (N_22028,N_21546,N_21929);
xnor U22029 (N_22029,N_21721,N_21677);
and U22030 (N_22030,N_21764,N_21662);
xnor U22031 (N_22031,N_21882,N_21904);
xor U22032 (N_22032,N_21767,N_21864);
xor U22033 (N_22033,N_21744,N_21993);
or U22034 (N_22034,N_21878,N_21841);
or U22035 (N_22035,N_21532,N_21548);
nor U22036 (N_22036,N_21991,N_21602);
xnor U22037 (N_22037,N_21674,N_21999);
and U22038 (N_22038,N_21795,N_21591);
or U22039 (N_22039,N_21702,N_21676);
and U22040 (N_22040,N_21735,N_21598);
nand U22041 (N_22041,N_21987,N_21545);
xnor U22042 (N_22042,N_21607,N_21569);
nor U22043 (N_22043,N_21634,N_21730);
xor U22044 (N_22044,N_21652,N_21861);
nand U22045 (N_22045,N_21650,N_21525);
nor U22046 (N_22046,N_21781,N_21818);
and U22047 (N_22047,N_21592,N_21577);
nor U22048 (N_22048,N_21879,N_21507);
nor U22049 (N_22049,N_21921,N_21715);
xor U22050 (N_22050,N_21670,N_21549);
nor U22051 (N_22051,N_21686,N_21720);
and U22052 (N_22052,N_21806,N_21732);
or U22053 (N_22053,N_21663,N_21856);
and U22054 (N_22054,N_21843,N_21614);
or U22055 (N_22055,N_21714,N_21881);
nor U22056 (N_22056,N_21977,N_21550);
and U22057 (N_22057,N_21811,N_21945);
xor U22058 (N_22058,N_21573,N_21706);
or U22059 (N_22059,N_21810,N_21838);
nor U22060 (N_22060,N_21738,N_21925);
and U22061 (N_22061,N_21567,N_21871);
or U22062 (N_22062,N_21703,N_21654);
xnor U22063 (N_22063,N_21750,N_21748);
or U22064 (N_22064,N_21967,N_21797);
and U22065 (N_22065,N_21917,N_21745);
or U22066 (N_22066,N_21989,N_21980);
and U22067 (N_22067,N_21533,N_21859);
xor U22068 (N_22068,N_21777,N_21884);
xnor U22069 (N_22069,N_21791,N_21679);
xnor U22070 (N_22070,N_21803,N_21515);
and U22071 (N_22071,N_21656,N_21529);
and U22072 (N_22072,N_21572,N_21561);
or U22073 (N_22073,N_21986,N_21960);
xor U22074 (N_22074,N_21514,N_21900);
nor U22075 (N_22075,N_21802,N_21641);
and U22076 (N_22076,N_21785,N_21880);
and U22077 (N_22077,N_21872,N_21913);
nor U22078 (N_22078,N_21974,N_21761);
nor U22079 (N_22079,N_21825,N_21948);
nor U22080 (N_22080,N_21631,N_21842);
and U22081 (N_22081,N_21771,N_21722);
xor U22082 (N_22082,N_21583,N_21510);
or U22083 (N_22083,N_21635,N_21685);
and U22084 (N_22084,N_21559,N_21905);
nand U22085 (N_22085,N_21638,N_21787);
or U22086 (N_22086,N_21556,N_21890);
xnor U22087 (N_22087,N_21773,N_21794);
nor U22088 (N_22088,N_21672,N_21512);
nor U22089 (N_22089,N_21758,N_21752);
and U22090 (N_22090,N_21769,N_21792);
or U22091 (N_22091,N_21540,N_21832);
and U22092 (N_22092,N_21947,N_21959);
and U22093 (N_22093,N_21938,N_21604);
xor U22094 (N_22094,N_21717,N_21704);
nor U22095 (N_22095,N_21846,N_21903);
or U22096 (N_22096,N_21585,N_21813);
and U22097 (N_22097,N_21593,N_21873);
or U22098 (N_22098,N_21617,N_21504);
xor U22099 (N_22099,N_21847,N_21968);
nand U22100 (N_22100,N_21835,N_21605);
xor U22101 (N_22101,N_21707,N_21973);
nor U22102 (N_22102,N_21855,N_21647);
nor U22103 (N_22103,N_21793,N_21658);
nor U22104 (N_22104,N_21950,N_21990);
and U22105 (N_22105,N_21778,N_21927);
xor U22106 (N_22106,N_21580,N_21731);
nand U22107 (N_22107,N_21581,N_21972);
nand U22108 (N_22108,N_21589,N_21782);
nand U22109 (N_22109,N_21594,N_21552);
nand U22110 (N_22110,N_21516,N_21957);
xor U22111 (N_22111,N_21666,N_21623);
or U22112 (N_22112,N_21754,N_21733);
and U22113 (N_22113,N_21982,N_21911);
nand U22114 (N_22114,N_21914,N_21564);
nor U22115 (N_22115,N_21988,N_21522);
nand U22116 (N_22116,N_21701,N_21840);
nand U22117 (N_22117,N_21958,N_21596);
and U22118 (N_22118,N_21951,N_21940);
and U22119 (N_22119,N_21645,N_21984);
xnor U22120 (N_22120,N_21578,N_21822);
nand U22121 (N_22121,N_21942,N_21865);
nor U22122 (N_22122,N_21981,N_21827);
xnor U22123 (N_22123,N_21590,N_21836);
nor U22124 (N_22124,N_21511,N_21537);
and U22125 (N_22125,N_21883,N_21613);
and U22126 (N_22126,N_21965,N_21770);
xnor U22127 (N_22127,N_21684,N_21772);
or U22128 (N_22128,N_21800,N_21659);
or U22129 (N_22129,N_21543,N_21756);
xor U22130 (N_22130,N_21523,N_21759);
xnor U22131 (N_22131,N_21896,N_21725);
or U22132 (N_22132,N_21521,N_21642);
and U22133 (N_22133,N_21502,N_21553);
nor U22134 (N_22134,N_21723,N_21978);
xor U22135 (N_22135,N_21566,N_21886);
and U22136 (N_22136,N_21775,N_21955);
and U22137 (N_22137,N_21628,N_21503);
or U22138 (N_22138,N_21637,N_21839);
nand U22139 (N_22139,N_21586,N_21994);
or U22140 (N_22140,N_21535,N_21742);
nor U22141 (N_22141,N_21780,N_21530);
xor U22142 (N_22142,N_21817,N_21828);
or U22143 (N_22143,N_21668,N_21557);
nand U22144 (N_22144,N_21719,N_21711);
or U22145 (N_22145,N_21747,N_21520);
xor U22146 (N_22146,N_21620,N_21804);
xor U22147 (N_22147,N_21899,N_21816);
or U22148 (N_22148,N_21830,N_21622);
or U22149 (N_22149,N_21831,N_21610);
and U22150 (N_22150,N_21746,N_21574);
nand U22151 (N_22151,N_21696,N_21858);
or U22152 (N_22152,N_21624,N_21612);
xor U22153 (N_22153,N_21630,N_21985);
nand U22154 (N_22154,N_21576,N_21734);
xor U22155 (N_22155,N_21629,N_21976);
nand U22156 (N_22156,N_21848,N_21956);
nand U22157 (N_22157,N_21874,N_21595);
or U22158 (N_22158,N_21944,N_21639);
xnor U22159 (N_22159,N_21971,N_21615);
nand U22160 (N_22160,N_21588,N_21542);
or U22161 (N_22161,N_21541,N_21692);
xnor U22162 (N_22162,N_21675,N_21681);
nand U22163 (N_22163,N_21788,N_21910);
nand U22164 (N_22164,N_21693,N_21664);
or U22165 (N_22165,N_21560,N_21633);
and U22166 (N_22166,N_21892,N_21718);
or U22167 (N_22167,N_21697,N_21599);
nor U22168 (N_22168,N_21627,N_21755);
nor U22169 (N_22169,N_21563,N_21768);
nor U22170 (N_22170,N_21860,N_21710);
nand U22171 (N_22171,N_21698,N_21661);
nor U22172 (N_22172,N_21689,N_21763);
nand U22173 (N_22173,N_21508,N_21875);
xnor U22174 (N_22174,N_21600,N_21712);
and U22175 (N_22175,N_21834,N_21902);
xor U22176 (N_22176,N_21716,N_21575);
nand U22177 (N_22177,N_21568,N_21680);
and U22178 (N_22178,N_21739,N_21805);
xnor U22179 (N_22179,N_21708,N_21695);
nor U22180 (N_22180,N_21798,N_21966);
or U22181 (N_22181,N_21555,N_21694);
or U22182 (N_22182,N_21998,N_21779);
nor U22183 (N_22183,N_21518,N_21919);
xnor U22184 (N_22184,N_21784,N_21954);
and U22185 (N_22185,N_21937,N_21513);
nor U22186 (N_22186,N_21644,N_21939);
xor U22187 (N_22187,N_21812,N_21979);
nand U22188 (N_22188,N_21866,N_21669);
nor U22189 (N_22189,N_21646,N_21728);
nand U22190 (N_22190,N_21737,N_21934);
or U22191 (N_22191,N_21547,N_21648);
nand U22192 (N_22192,N_21709,N_21531);
nand U22193 (N_22193,N_21946,N_21626);
nand U22194 (N_22194,N_21821,N_21736);
nor U22195 (N_22195,N_21505,N_21961);
nor U22196 (N_22196,N_21796,N_21823);
nand U22197 (N_22197,N_21527,N_21649);
or U22198 (N_22198,N_21894,N_21509);
nand U22199 (N_22199,N_21660,N_21851);
xnor U22200 (N_22200,N_21571,N_21786);
nor U22201 (N_22201,N_21941,N_21888);
or U22202 (N_22202,N_21611,N_21895);
nor U22203 (N_22203,N_21876,N_21808);
and U22204 (N_22204,N_21570,N_21844);
or U22205 (N_22205,N_21727,N_21953);
xnor U22206 (N_22206,N_21551,N_21691);
xnor U22207 (N_22207,N_21743,N_21643);
xnor U22208 (N_22208,N_21618,N_21636);
and U22209 (N_22209,N_21898,N_21952);
nor U22210 (N_22210,N_21765,N_21783);
xor U22211 (N_22211,N_21930,N_21584);
or U22212 (N_22212,N_21562,N_21603);
xnor U22213 (N_22213,N_21606,N_21897);
xnor U22214 (N_22214,N_21713,N_21683);
xnor U22215 (N_22215,N_21753,N_21749);
or U22216 (N_22216,N_21539,N_21554);
xor U22217 (N_22217,N_21740,N_21837);
or U22218 (N_22218,N_21820,N_21601);
nand U22219 (N_22219,N_21534,N_21653);
xor U22220 (N_22220,N_21724,N_21867);
nor U22221 (N_22221,N_21506,N_21870);
or U22222 (N_22222,N_21690,N_21933);
nand U22223 (N_22223,N_21949,N_21558);
xor U22224 (N_22224,N_21970,N_21935);
or U22225 (N_22225,N_21519,N_21774);
or U22226 (N_22226,N_21924,N_21632);
or U22227 (N_22227,N_21969,N_21885);
or U22228 (N_22228,N_21538,N_21608);
xor U22229 (N_22229,N_21983,N_21997);
and U22230 (N_22230,N_21579,N_21829);
nand U22231 (N_22231,N_21963,N_21931);
nand U22232 (N_22232,N_21640,N_21962);
xnor U22233 (N_22233,N_21996,N_21665);
or U22234 (N_22234,N_21619,N_21621);
xnor U22235 (N_22235,N_21655,N_21869);
and U22236 (N_22236,N_21849,N_21699);
xor U22237 (N_22237,N_21854,N_21918);
and U22238 (N_22238,N_21992,N_21673);
nand U22239 (N_22239,N_21833,N_21688);
xnor U22240 (N_22240,N_21852,N_21923);
nor U22241 (N_22241,N_21906,N_21912);
nor U22242 (N_22242,N_21868,N_21682);
nand U22243 (N_22243,N_21863,N_21850);
or U22244 (N_22244,N_21815,N_21936);
or U22245 (N_22245,N_21807,N_21526);
and U22246 (N_22246,N_21922,N_21862);
nor U22247 (N_22247,N_21766,N_21651);
nand U22248 (N_22248,N_21819,N_21528);
nor U22249 (N_22249,N_21964,N_21975);
nand U22250 (N_22250,N_21630,N_21712);
and U22251 (N_22251,N_21967,N_21724);
xor U22252 (N_22252,N_21671,N_21787);
xor U22253 (N_22253,N_21658,N_21513);
xor U22254 (N_22254,N_21527,N_21873);
nor U22255 (N_22255,N_21626,N_21695);
or U22256 (N_22256,N_21780,N_21855);
nor U22257 (N_22257,N_21883,N_21691);
nor U22258 (N_22258,N_21782,N_21689);
nor U22259 (N_22259,N_21875,N_21816);
nor U22260 (N_22260,N_21734,N_21775);
or U22261 (N_22261,N_21635,N_21914);
or U22262 (N_22262,N_21696,N_21730);
or U22263 (N_22263,N_21534,N_21981);
xnor U22264 (N_22264,N_21701,N_21507);
nand U22265 (N_22265,N_21702,N_21621);
nand U22266 (N_22266,N_21736,N_21684);
and U22267 (N_22267,N_21681,N_21955);
nor U22268 (N_22268,N_21736,N_21776);
nand U22269 (N_22269,N_21744,N_21543);
nand U22270 (N_22270,N_21901,N_21824);
nor U22271 (N_22271,N_21971,N_21851);
nor U22272 (N_22272,N_21920,N_21601);
nand U22273 (N_22273,N_21531,N_21705);
or U22274 (N_22274,N_21667,N_21960);
and U22275 (N_22275,N_21887,N_21914);
xnor U22276 (N_22276,N_21750,N_21811);
or U22277 (N_22277,N_21605,N_21916);
nand U22278 (N_22278,N_21575,N_21965);
or U22279 (N_22279,N_21666,N_21934);
or U22280 (N_22280,N_21933,N_21772);
nand U22281 (N_22281,N_21606,N_21546);
nor U22282 (N_22282,N_21675,N_21505);
nor U22283 (N_22283,N_21905,N_21640);
or U22284 (N_22284,N_21701,N_21652);
nand U22285 (N_22285,N_21767,N_21988);
nor U22286 (N_22286,N_21712,N_21744);
and U22287 (N_22287,N_21634,N_21542);
nor U22288 (N_22288,N_21795,N_21848);
or U22289 (N_22289,N_21902,N_21958);
nand U22290 (N_22290,N_21956,N_21613);
nor U22291 (N_22291,N_21696,N_21605);
and U22292 (N_22292,N_21836,N_21710);
nand U22293 (N_22293,N_21890,N_21630);
xor U22294 (N_22294,N_21847,N_21833);
xor U22295 (N_22295,N_21647,N_21595);
nand U22296 (N_22296,N_21754,N_21509);
or U22297 (N_22297,N_21582,N_21927);
xor U22298 (N_22298,N_21631,N_21791);
nand U22299 (N_22299,N_21827,N_21886);
nor U22300 (N_22300,N_21897,N_21690);
or U22301 (N_22301,N_21820,N_21949);
nor U22302 (N_22302,N_21792,N_21565);
nor U22303 (N_22303,N_21836,N_21780);
xor U22304 (N_22304,N_21973,N_21983);
nand U22305 (N_22305,N_21541,N_21629);
xnor U22306 (N_22306,N_21935,N_21926);
nand U22307 (N_22307,N_21521,N_21830);
xor U22308 (N_22308,N_21865,N_21883);
nand U22309 (N_22309,N_21574,N_21975);
and U22310 (N_22310,N_21908,N_21852);
nor U22311 (N_22311,N_21872,N_21685);
or U22312 (N_22312,N_21633,N_21530);
nand U22313 (N_22313,N_21552,N_21821);
nor U22314 (N_22314,N_21653,N_21660);
nor U22315 (N_22315,N_21776,N_21753);
and U22316 (N_22316,N_21697,N_21933);
nor U22317 (N_22317,N_21500,N_21796);
xor U22318 (N_22318,N_21625,N_21703);
nand U22319 (N_22319,N_21814,N_21738);
nand U22320 (N_22320,N_21835,N_21952);
or U22321 (N_22321,N_21613,N_21766);
xnor U22322 (N_22322,N_21570,N_21870);
xnor U22323 (N_22323,N_21963,N_21913);
nor U22324 (N_22324,N_21837,N_21586);
xor U22325 (N_22325,N_21966,N_21828);
nand U22326 (N_22326,N_21810,N_21726);
and U22327 (N_22327,N_21860,N_21991);
nand U22328 (N_22328,N_21628,N_21587);
xnor U22329 (N_22329,N_21797,N_21585);
nand U22330 (N_22330,N_21930,N_21816);
xnor U22331 (N_22331,N_21824,N_21751);
nand U22332 (N_22332,N_21816,N_21608);
nand U22333 (N_22333,N_21802,N_21712);
and U22334 (N_22334,N_21532,N_21850);
and U22335 (N_22335,N_21586,N_21979);
nand U22336 (N_22336,N_21659,N_21720);
nand U22337 (N_22337,N_21838,N_21629);
nand U22338 (N_22338,N_21766,N_21937);
nor U22339 (N_22339,N_21973,N_21910);
nand U22340 (N_22340,N_21952,N_21550);
nand U22341 (N_22341,N_21997,N_21694);
or U22342 (N_22342,N_21651,N_21982);
xor U22343 (N_22343,N_21919,N_21719);
nor U22344 (N_22344,N_21742,N_21600);
or U22345 (N_22345,N_21699,N_21948);
or U22346 (N_22346,N_21622,N_21675);
nand U22347 (N_22347,N_21854,N_21995);
or U22348 (N_22348,N_21532,N_21549);
nand U22349 (N_22349,N_21988,N_21649);
xor U22350 (N_22350,N_21519,N_21643);
nand U22351 (N_22351,N_21529,N_21666);
and U22352 (N_22352,N_21951,N_21850);
nand U22353 (N_22353,N_21820,N_21913);
nor U22354 (N_22354,N_21503,N_21842);
nor U22355 (N_22355,N_21731,N_21764);
nand U22356 (N_22356,N_21873,N_21975);
or U22357 (N_22357,N_21539,N_21974);
or U22358 (N_22358,N_21991,N_21806);
xor U22359 (N_22359,N_21915,N_21691);
or U22360 (N_22360,N_21555,N_21661);
xor U22361 (N_22361,N_21847,N_21527);
and U22362 (N_22362,N_21794,N_21645);
nand U22363 (N_22363,N_21719,N_21899);
or U22364 (N_22364,N_21660,N_21627);
xnor U22365 (N_22365,N_21515,N_21502);
nand U22366 (N_22366,N_21953,N_21514);
nor U22367 (N_22367,N_21891,N_21865);
xnor U22368 (N_22368,N_21995,N_21886);
xor U22369 (N_22369,N_21922,N_21529);
and U22370 (N_22370,N_21675,N_21678);
or U22371 (N_22371,N_21609,N_21600);
or U22372 (N_22372,N_21956,N_21726);
nand U22373 (N_22373,N_21734,N_21984);
nand U22374 (N_22374,N_21923,N_21691);
or U22375 (N_22375,N_21882,N_21736);
or U22376 (N_22376,N_21924,N_21807);
nor U22377 (N_22377,N_21868,N_21797);
and U22378 (N_22378,N_21596,N_21512);
nor U22379 (N_22379,N_21659,N_21697);
nor U22380 (N_22380,N_21700,N_21688);
nand U22381 (N_22381,N_21827,N_21982);
or U22382 (N_22382,N_21789,N_21921);
xnor U22383 (N_22383,N_21512,N_21809);
nand U22384 (N_22384,N_21729,N_21996);
or U22385 (N_22385,N_21545,N_21843);
xnor U22386 (N_22386,N_21512,N_21892);
nand U22387 (N_22387,N_21546,N_21877);
and U22388 (N_22388,N_21754,N_21507);
and U22389 (N_22389,N_21681,N_21657);
xor U22390 (N_22390,N_21884,N_21987);
nand U22391 (N_22391,N_21769,N_21766);
or U22392 (N_22392,N_21695,N_21544);
nand U22393 (N_22393,N_21774,N_21819);
or U22394 (N_22394,N_21971,N_21784);
or U22395 (N_22395,N_21850,N_21959);
xor U22396 (N_22396,N_21704,N_21898);
or U22397 (N_22397,N_21596,N_21785);
or U22398 (N_22398,N_21788,N_21918);
nor U22399 (N_22399,N_21829,N_21808);
xor U22400 (N_22400,N_21675,N_21867);
or U22401 (N_22401,N_21569,N_21963);
or U22402 (N_22402,N_21537,N_21928);
and U22403 (N_22403,N_21806,N_21820);
and U22404 (N_22404,N_21853,N_21655);
and U22405 (N_22405,N_21857,N_21581);
nand U22406 (N_22406,N_21880,N_21654);
nand U22407 (N_22407,N_21837,N_21804);
or U22408 (N_22408,N_21628,N_21683);
nor U22409 (N_22409,N_21769,N_21822);
and U22410 (N_22410,N_21561,N_21952);
and U22411 (N_22411,N_21540,N_21678);
and U22412 (N_22412,N_21522,N_21539);
or U22413 (N_22413,N_21852,N_21949);
and U22414 (N_22414,N_21807,N_21708);
nand U22415 (N_22415,N_21803,N_21833);
xor U22416 (N_22416,N_21600,N_21537);
or U22417 (N_22417,N_21567,N_21560);
nor U22418 (N_22418,N_21793,N_21864);
or U22419 (N_22419,N_21566,N_21680);
nand U22420 (N_22420,N_21835,N_21848);
nor U22421 (N_22421,N_21514,N_21565);
and U22422 (N_22422,N_21586,N_21656);
nand U22423 (N_22423,N_21815,N_21512);
xor U22424 (N_22424,N_21728,N_21605);
and U22425 (N_22425,N_21824,N_21820);
nand U22426 (N_22426,N_21975,N_21847);
or U22427 (N_22427,N_21702,N_21875);
xor U22428 (N_22428,N_21622,N_21559);
nand U22429 (N_22429,N_21532,N_21514);
xnor U22430 (N_22430,N_21573,N_21905);
or U22431 (N_22431,N_21603,N_21869);
xnor U22432 (N_22432,N_21531,N_21846);
and U22433 (N_22433,N_21778,N_21648);
nand U22434 (N_22434,N_21955,N_21961);
or U22435 (N_22435,N_21774,N_21508);
nand U22436 (N_22436,N_21986,N_21512);
nor U22437 (N_22437,N_21865,N_21646);
xor U22438 (N_22438,N_21952,N_21500);
xnor U22439 (N_22439,N_21910,N_21785);
xor U22440 (N_22440,N_21730,N_21651);
or U22441 (N_22441,N_21754,N_21931);
and U22442 (N_22442,N_21806,N_21798);
or U22443 (N_22443,N_21841,N_21660);
nor U22444 (N_22444,N_21909,N_21980);
nand U22445 (N_22445,N_21817,N_21549);
or U22446 (N_22446,N_21796,N_21725);
nand U22447 (N_22447,N_21834,N_21835);
and U22448 (N_22448,N_21776,N_21911);
and U22449 (N_22449,N_21771,N_21550);
xnor U22450 (N_22450,N_21946,N_21662);
and U22451 (N_22451,N_21700,N_21546);
and U22452 (N_22452,N_21987,N_21769);
xnor U22453 (N_22453,N_21643,N_21977);
or U22454 (N_22454,N_21814,N_21844);
nor U22455 (N_22455,N_21801,N_21563);
or U22456 (N_22456,N_21506,N_21820);
nor U22457 (N_22457,N_21560,N_21929);
and U22458 (N_22458,N_21602,N_21592);
xor U22459 (N_22459,N_21649,N_21641);
and U22460 (N_22460,N_21797,N_21706);
nand U22461 (N_22461,N_21531,N_21841);
or U22462 (N_22462,N_21969,N_21799);
nand U22463 (N_22463,N_21528,N_21922);
and U22464 (N_22464,N_21650,N_21917);
nor U22465 (N_22465,N_21891,N_21787);
nand U22466 (N_22466,N_21703,N_21598);
and U22467 (N_22467,N_21667,N_21869);
and U22468 (N_22468,N_21971,N_21548);
or U22469 (N_22469,N_21672,N_21794);
and U22470 (N_22470,N_21578,N_21909);
and U22471 (N_22471,N_21625,N_21622);
and U22472 (N_22472,N_21920,N_21787);
and U22473 (N_22473,N_21968,N_21819);
nor U22474 (N_22474,N_21924,N_21568);
or U22475 (N_22475,N_21698,N_21625);
or U22476 (N_22476,N_21643,N_21869);
nand U22477 (N_22477,N_21893,N_21577);
nand U22478 (N_22478,N_21939,N_21567);
nor U22479 (N_22479,N_21998,N_21903);
and U22480 (N_22480,N_21540,N_21853);
xor U22481 (N_22481,N_21663,N_21849);
nand U22482 (N_22482,N_21842,N_21739);
and U22483 (N_22483,N_21806,N_21545);
and U22484 (N_22484,N_21996,N_21655);
nand U22485 (N_22485,N_21644,N_21522);
nor U22486 (N_22486,N_21650,N_21735);
or U22487 (N_22487,N_21546,N_21519);
xnor U22488 (N_22488,N_21624,N_21738);
or U22489 (N_22489,N_21619,N_21913);
xor U22490 (N_22490,N_21548,N_21879);
nand U22491 (N_22491,N_21503,N_21796);
xnor U22492 (N_22492,N_21552,N_21504);
nand U22493 (N_22493,N_21837,N_21536);
xor U22494 (N_22494,N_21571,N_21588);
xor U22495 (N_22495,N_21514,N_21628);
xnor U22496 (N_22496,N_21586,N_21789);
nand U22497 (N_22497,N_21666,N_21757);
nand U22498 (N_22498,N_21617,N_21999);
nor U22499 (N_22499,N_21628,N_21997);
xnor U22500 (N_22500,N_22092,N_22150);
xor U22501 (N_22501,N_22243,N_22163);
xor U22502 (N_22502,N_22483,N_22405);
nand U22503 (N_22503,N_22285,N_22244);
nand U22504 (N_22504,N_22084,N_22442);
nor U22505 (N_22505,N_22383,N_22110);
or U22506 (N_22506,N_22009,N_22379);
and U22507 (N_22507,N_22202,N_22474);
nand U22508 (N_22508,N_22189,N_22429);
or U22509 (N_22509,N_22021,N_22051);
nand U22510 (N_22510,N_22332,N_22002);
nand U22511 (N_22511,N_22449,N_22000);
nand U22512 (N_22512,N_22470,N_22030);
and U22513 (N_22513,N_22094,N_22065);
nor U22514 (N_22514,N_22329,N_22121);
or U22515 (N_22515,N_22495,N_22378);
xor U22516 (N_22516,N_22486,N_22364);
nand U22517 (N_22517,N_22188,N_22006);
or U22518 (N_22518,N_22415,N_22177);
xor U22519 (N_22519,N_22257,N_22348);
xor U22520 (N_22520,N_22184,N_22220);
or U22521 (N_22521,N_22225,N_22413);
nor U22522 (N_22522,N_22129,N_22386);
xor U22523 (N_22523,N_22450,N_22443);
xnor U22524 (N_22524,N_22180,N_22201);
xor U22525 (N_22525,N_22458,N_22303);
and U22526 (N_22526,N_22161,N_22104);
nand U22527 (N_22527,N_22463,N_22230);
and U22528 (N_22528,N_22290,N_22147);
or U22529 (N_22529,N_22194,N_22295);
xnor U22530 (N_22530,N_22054,N_22434);
nand U22531 (N_22531,N_22428,N_22390);
or U22532 (N_22532,N_22334,N_22081);
nand U22533 (N_22533,N_22440,N_22418);
or U22534 (N_22534,N_22456,N_22060);
xnor U22535 (N_22535,N_22263,N_22254);
xor U22536 (N_22536,N_22077,N_22269);
xnor U22537 (N_22537,N_22176,N_22034);
nor U22538 (N_22538,N_22248,N_22143);
nand U22539 (N_22539,N_22175,N_22420);
and U22540 (N_22540,N_22069,N_22493);
and U22541 (N_22541,N_22144,N_22370);
or U22542 (N_22542,N_22212,N_22361);
and U22543 (N_22543,N_22119,N_22135);
or U22544 (N_22544,N_22242,N_22190);
and U22545 (N_22545,N_22033,N_22130);
and U22546 (N_22546,N_22306,N_22036);
xor U22547 (N_22547,N_22158,N_22446);
xor U22548 (N_22548,N_22337,N_22252);
or U22549 (N_22549,N_22345,N_22462);
nand U22550 (N_22550,N_22102,N_22208);
nor U22551 (N_22551,N_22310,N_22321);
nand U22552 (N_22552,N_22204,N_22120);
xor U22553 (N_22553,N_22430,N_22111);
xnor U22554 (N_22554,N_22437,N_22160);
xor U22555 (N_22555,N_22196,N_22232);
or U22556 (N_22556,N_22497,N_22057);
nor U22557 (N_22557,N_22498,N_22192);
nand U22558 (N_22558,N_22042,N_22480);
xnor U22559 (N_22559,N_22347,N_22424);
nand U22560 (N_22560,N_22426,N_22074);
nand U22561 (N_22561,N_22317,N_22387);
or U22562 (N_22562,N_22289,N_22320);
and U22563 (N_22563,N_22384,N_22344);
nand U22564 (N_22564,N_22479,N_22156);
or U22565 (N_22565,N_22322,N_22088);
and U22566 (N_22566,N_22134,N_22145);
nand U22567 (N_22567,N_22358,N_22432);
xnor U22568 (N_22568,N_22186,N_22234);
nor U22569 (N_22569,N_22411,N_22318);
or U22570 (N_22570,N_22153,N_22423);
nor U22571 (N_22571,N_22284,N_22399);
nor U22572 (N_22572,N_22372,N_22162);
or U22573 (N_22573,N_22445,N_22187);
nand U22574 (N_22574,N_22068,N_22286);
and U22575 (N_22575,N_22078,N_22044);
nand U22576 (N_22576,N_22231,N_22211);
xnor U22577 (N_22577,N_22035,N_22118);
nand U22578 (N_22578,N_22249,N_22251);
nor U22579 (N_22579,N_22408,N_22195);
and U22580 (N_22580,N_22316,N_22441);
xor U22581 (N_22581,N_22311,N_22105);
or U22582 (N_22582,N_22273,N_22086);
or U22583 (N_22583,N_22228,N_22271);
nand U22584 (N_22584,N_22340,N_22182);
and U22585 (N_22585,N_22038,N_22416);
xor U22586 (N_22586,N_22315,N_22059);
nand U22587 (N_22587,N_22001,N_22342);
nand U22588 (N_22588,N_22075,N_22301);
nand U22589 (N_22589,N_22478,N_22014);
xnor U22590 (N_22590,N_22245,N_22266);
nand U22591 (N_22591,N_22116,N_22374);
nor U22592 (N_22592,N_22421,N_22451);
nor U22593 (N_22593,N_22089,N_22298);
xor U22594 (N_22594,N_22373,N_22011);
nor U22595 (N_22595,N_22137,N_22066);
or U22596 (N_22596,N_22327,N_22258);
or U22597 (N_22597,N_22296,N_22359);
nand U22598 (N_22598,N_22123,N_22395);
or U22599 (N_22599,N_22193,N_22235);
nor U22600 (N_22600,N_22159,N_22091);
nand U22601 (N_22601,N_22433,N_22095);
and U22602 (N_22602,N_22064,N_22029);
nor U22603 (N_22603,N_22496,N_22466);
xnor U22604 (N_22604,N_22255,N_22238);
xor U22605 (N_22605,N_22414,N_22114);
nand U22606 (N_22606,N_22328,N_22149);
xor U22607 (N_22607,N_22331,N_22100);
nand U22608 (N_22608,N_22073,N_22490);
or U22609 (N_22609,N_22122,N_22346);
xnor U22610 (N_22610,N_22047,N_22023);
and U22611 (N_22611,N_22302,N_22313);
or U22612 (N_22612,N_22046,N_22319);
and U22613 (N_22613,N_22053,N_22085);
xor U22614 (N_22614,N_22356,N_22056);
and U22615 (N_22615,N_22274,N_22039);
nor U22616 (N_22616,N_22343,N_22216);
nand U22617 (N_22617,N_22008,N_22173);
nor U22618 (N_22618,N_22324,N_22461);
xnor U22619 (N_22619,N_22133,N_22402);
nor U22620 (N_22620,N_22262,N_22063);
xor U22621 (N_22621,N_22219,N_22293);
or U22622 (N_22622,N_22200,N_22012);
or U22623 (N_22623,N_22027,N_22377);
nand U22624 (N_22624,N_22409,N_22357);
or U22625 (N_22625,N_22106,N_22169);
and U22626 (N_22626,N_22097,N_22172);
xor U22627 (N_22627,N_22025,N_22024);
xor U22628 (N_22628,N_22481,N_22492);
nor U22629 (N_22629,N_22157,N_22369);
nand U22630 (N_22630,N_22048,N_22341);
nand U22631 (N_22631,N_22350,N_22491);
xor U22632 (N_22632,N_22107,N_22272);
xor U22633 (N_22633,N_22468,N_22087);
xnor U22634 (N_22634,N_22391,N_22007);
nand U22635 (N_22635,N_22292,N_22325);
and U22636 (N_22636,N_22385,N_22397);
and U22637 (N_22637,N_22224,N_22004);
nor U22638 (N_22638,N_22239,N_22488);
nor U22639 (N_22639,N_22166,N_22139);
and U22640 (N_22640,N_22394,N_22287);
or U22641 (N_22641,N_22256,N_22223);
and U22642 (N_22642,N_22181,N_22406);
nand U22643 (N_22643,N_22467,N_22055);
and U22644 (N_22644,N_22291,N_22407);
xnor U22645 (N_22645,N_22236,N_22032);
nor U22646 (N_22646,N_22401,N_22140);
or U22647 (N_22647,N_22323,N_22452);
nand U22648 (N_22648,N_22233,N_22198);
nor U22649 (N_22649,N_22240,N_22037);
or U22650 (N_22650,N_22412,N_22366);
xnor U22651 (N_22651,N_22015,N_22307);
or U22652 (N_22652,N_22058,N_22098);
xnor U22653 (N_22653,N_22214,N_22473);
xor U22654 (N_22654,N_22131,N_22392);
xnor U22655 (N_22655,N_22022,N_22281);
and U22656 (N_22656,N_22151,N_22448);
or U22657 (N_22657,N_22241,N_22351);
xnor U22658 (N_22658,N_22381,N_22174);
nor U22659 (N_22659,N_22080,N_22339);
and U22660 (N_22660,N_22113,N_22419);
xnor U22661 (N_22661,N_22277,N_22382);
xor U22662 (N_22662,N_22457,N_22270);
or U22663 (N_22663,N_22209,N_22472);
or U22664 (N_22664,N_22375,N_22222);
and U22665 (N_22665,N_22167,N_22203);
or U22666 (N_22666,N_22218,N_22112);
nand U22667 (N_22667,N_22312,N_22132);
nor U22668 (N_22668,N_22380,N_22288);
and U22669 (N_22669,N_22128,N_22265);
and U22670 (N_22670,N_22283,N_22090);
and U22671 (N_22671,N_22020,N_22072);
xnor U22672 (N_22672,N_22197,N_22101);
xor U22673 (N_22673,N_22217,N_22179);
nor U22674 (N_22674,N_22422,N_22431);
nand U22675 (N_22675,N_22469,N_22487);
xor U22676 (N_22676,N_22362,N_22309);
xnor U22677 (N_22677,N_22052,N_22155);
xnor U22678 (N_22678,N_22017,N_22494);
nor U22679 (N_22679,N_22425,N_22304);
xnor U22680 (N_22680,N_22178,N_22314);
or U22681 (N_22681,N_22389,N_22099);
nand U22682 (N_22682,N_22227,N_22125);
and U22683 (N_22683,N_22003,N_22109);
or U22684 (N_22684,N_22124,N_22278);
and U22685 (N_22685,N_22282,N_22349);
nand U22686 (N_22686,N_22326,N_22400);
xor U22687 (N_22687,N_22253,N_22115);
nor U22688 (N_22688,N_22477,N_22185);
nor U22689 (N_22689,N_22018,N_22465);
nand U22690 (N_22690,N_22164,N_22237);
nand U22691 (N_22691,N_22367,N_22096);
and U22692 (N_22692,N_22210,N_22117);
nand U22693 (N_22693,N_22213,N_22050);
xor U22694 (N_22694,N_22082,N_22070);
or U22695 (N_22695,N_22259,N_22028);
nor U22696 (N_22696,N_22205,N_22215);
xnor U22697 (N_22697,N_22404,N_22010);
xor U22698 (N_22698,N_22436,N_22136);
and U22699 (N_22699,N_22294,N_22041);
or U22700 (N_22700,N_22103,N_22247);
xor U22701 (N_22701,N_22335,N_22229);
nand U22702 (N_22702,N_22453,N_22062);
or U22703 (N_22703,N_22019,N_22447);
nor U22704 (N_22704,N_22170,N_22267);
nor U22705 (N_22705,N_22146,N_22045);
and U22706 (N_22706,N_22427,N_22083);
and U22707 (N_22707,N_22031,N_22067);
xor U22708 (N_22708,N_22297,N_22460);
nand U22709 (N_22709,N_22250,N_22154);
nand U22710 (N_22710,N_22299,N_22435);
and U22711 (N_22711,N_22275,N_22471);
xnor U22712 (N_22712,N_22005,N_22264);
xnor U22713 (N_22713,N_22376,N_22016);
and U22714 (N_22714,N_22142,N_22300);
and U22715 (N_22715,N_22268,N_22165);
nor U22716 (N_22716,N_22444,N_22464);
nor U22717 (N_22717,N_22152,N_22459);
nand U22718 (N_22718,N_22191,N_22371);
nand U22719 (N_22719,N_22168,N_22148);
nor U22720 (N_22720,N_22226,N_22485);
and U22721 (N_22721,N_22499,N_22355);
nand U22722 (N_22722,N_22338,N_22206);
and U22723 (N_22723,N_22308,N_22352);
nor U22724 (N_22724,N_22475,N_22454);
nor U22725 (N_22725,N_22439,N_22398);
xnor U22726 (N_22726,N_22261,N_22365);
and U22727 (N_22727,N_22410,N_22127);
and U22728 (N_22728,N_22138,N_22396);
nand U22729 (N_22729,N_22141,N_22360);
nand U22730 (N_22730,N_22076,N_22207);
nor U22731 (N_22731,N_22093,N_22049);
and U22732 (N_22732,N_22363,N_22071);
or U22733 (N_22733,N_22260,N_22353);
or U22734 (N_22734,N_22026,N_22330);
nor U22735 (N_22735,N_22393,N_22279);
or U22736 (N_22736,N_22489,N_22482);
xor U22737 (N_22737,N_22221,N_22108);
nand U22738 (N_22738,N_22043,N_22417);
or U22739 (N_22739,N_22280,N_22013);
nor U22740 (N_22740,N_22484,N_22354);
or U22741 (N_22741,N_22183,N_22061);
nand U22742 (N_22742,N_22438,N_22388);
xor U22743 (N_22743,N_22171,N_22126);
nand U22744 (N_22744,N_22079,N_22455);
xnor U22745 (N_22745,N_22305,N_22040);
xor U22746 (N_22746,N_22333,N_22336);
nor U22747 (N_22747,N_22403,N_22476);
xor U22748 (N_22748,N_22368,N_22199);
or U22749 (N_22749,N_22246,N_22276);
or U22750 (N_22750,N_22192,N_22368);
or U22751 (N_22751,N_22159,N_22477);
nand U22752 (N_22752,N_22483,N_22066);
nand U22753 (N_22753,N_22171,N_22140);
or U22754 (N_22754,N_22401,N_22010);
nor U22755 (N_22755,N_22064,N_22385);
xor U22756 (N_22756,N_22252,N_22365);
nor U22757 (N_22757,N_22149,N_22429);
nand U22758 (N_22758,N_22183,N_22383);
xnor U22759 (N_22759,N_22176,N_22088);
xor U22760 (N_22760,N_22246,N_22050);
xnor U22761 (N_22761,N_22498,N_22496);
and U22762 (N_22762,N_22218,N_22207);
and U22763 (N_22763,N_22283,N_22205);
xnor U22764 (N_22764,N_22132,N_22160);
or U22765 (N_22765,N_22333,N_22054);
xor U22766 (N_22766,N_22223,N_22108);
xor U22767 (N_22767,N_22337,N_22454);
and U22768 (N_22768,N_22461,N_22241);
nor U22769 (N_22769,N_22460,N_22004);
and U22770 (N_22770,N_22435,N_22163);
nor U22771 (N_22771,N_22232,N_22087);
nand U22772 (N_22772,N_22109,N_22121);
xor U22773 (N_22773,N_22431,N_22157);
or U22774 (N_22774,N_22394,N_22452);
xnor U22775 (N_22775,N_22150,N_22203);
and U22776 (N_22776,N_22337,N_22194);
and U22777 (N_22777,N_22434,N_22172);
and U22778 (N_22778,N_22453,N_22468);
and U22779 (N_22779,N_22326,N_22448);
nand U22780 (N_22780,N_22162,N_22077);
xor U22781 (N_22781,N_22468,N_22298);
or U22782 (N_22782,N_22361,N_22484);
and U22783 (N_22783,N_22340,N_22374);
nor U22784 (N_22784,N_22053,N_22431);
nor U22785 (N_22785,N_22303,N_22343);
nand U22786 (N_22786,N_22397,N_22441);
xnor U22787 (N_22787,N_22497,N_22015);
nand U22788 (N_22788,N_22107,N_22158);
xor U22789 (N_22789,N_22273,N_22443);
or U22790 (N_22790,N_22386,N_22322);
xor U22791 (N_22791,N_22237,N_22069);
xor U22792 (N_22792,N_22297,N_22047);
nor U22793 (N_22793,N_22258,N_22443);
xnor U22794 (N_22794,N_22101,N_22067);
nor U22795 (N_22795,N_22384,N_22445);
or U22796 (N_22796,N_22412,N_22163);
nand U22797 (N_22797,N_22288,N_22303);
xnor U22798 (N_22798,N_22064,N_22033);
nor U22799 (N_22799,N_22418,N_22454);
or U22800 (N_22800,N_22194,N_22270);
nand U22801 (N_22801,N_22251,N_22244);
or U22802 (N_22802,N_22476,N_22249);
xnor U22803 (N_22803,N_22353,N_22346);
or U22804 (N_22804,N_22159,N_22276);
xor U22805 (N_22805,N_22094,N_22444);
or U22806 (N_22806,N_22067,N_22363);
nand U22807 (N_22807,N_22058,N_22059);
or U22808 (N_22808,N_22244,N_22143);
nor U22809 (N_22809,N_22481,N_22013);
nand U22810 (N_22810,N_22411,N_22439);
nand U22811 (N_22811,N_22077,N_22220);
nand U22812 (N_22812,N_22101,N_22487);
and U22813 (N_22813,N_22293,N_22372);
xor U22814 (N_22814,N_22382,N_22473);
or U22815 (N_22815,N_22290,N_22037);
nand U22816 (N_22816,N_22128,N_22270);
or U22817 (N_22817,N_22399,N_22371);
and U22818 (N_22818,N_22364,N_22311);
or U22819 (N_22819,N_22231,N_22322);
nor U22820 (N_22820,N_22483,N_22277);
xnor U22821 (N_22821,N_22320,N_22112);
nand U22822 (N_22822,N_22372,N_22309);
nand U22823 (N_22823,N_22166,N_22248);
nor U22824 (N_22824,N_22199,N_22030);
and U22825 (N_22825,N_22415,N_22273);
xor U22826 (N_22826,N_22243,N_22078);
and U22827 (N_22827,N_22074,N_22199);
nor U22828 (N_22828,N_22330,N_22378);
xnor U22829 (N_22829,N_22152,N_22369);
nor U22830 (N_22830,N_22084,N_22403);
nand U22831 (N_22831,N_22291,N_22033);
and U22832 (N_22832,N_22257,N_22057);
xor U22833 (N_22833,N_22269,N_22096);
and U22834 (N_22834,N_22329,N_22440);
nor U22835 (N_22835,N_22005,N_22483);
nand U22836 (N_22836,N_22192,N_22140);
and U22837 (N_22837,N_22231,N_22453);
nor U22838 (N_22838,N_22317,N_22461);
nand U22839 (N_22839,N_22200,N_22285);
xor U22840 (N_22840,N_22490,N_22017);
nor U22841 (N_22841,N_22012,N_22210);
nor U22842 (N_22842,N_22378,N_22108);
and U22843 (N_22843,N_22263,N_22260);
nand U22844 (N_22844,N_22176,N_22083);
nor U22845 (N_22845,N_22089,N_22170);
xnor U22846 (N_22846,N_22036,N_22295);
nand U22847 (N_22847,N_22351,N_22157);
or U22848 (N_22848,N_22245,N_22050);
nor U22849 (N_22849,N_22104,N_22324);
nor U22850 (N_22850,N_22306,N_22013);
or U22851 (N_22851,N_22046,N_22394);
or U22852 (N_22852,N_22446,N_22048);
nor U22853 (N_22853,N_22282,N_22393);
and U22854 (N_22854,N_22238,N_22141);
xor U22855 (N_22855,N_22395,N_22182);
and U22856 (N_22856,N_22251,N_22209);
xor U22857 (N_22857,N_22190,N_22275);
or U22858 (N_22858,N_22382,N_22024);
or U22859 (N_22859,N_22460,N_22437);
or U22860 (N_22860,N_22090,N_22335);
or U22861 (N_22861,N_22263,N_22033);
nor U22862 (N_22862,N_22418,N_22359);
and U22863 (N_22863,N_22106,N_22183);
and U22864 (N_22864,N_22208,N_22489);
nand U22865 (N_22865,N_22202,N_22381);
or U22866 (N_22866,N_22050,N_22089);
nor U22867 (N_22867,N_22167,N_22011);
and U22868 (N_22868,N_22059,N_22253);
or U22869 (N_22869,N_22436,N_22377);
and U22870 (N_22870,N_22025,N_22281);
xnor U22871 (N_22871,N_22188,N_22037);
nor U22872 (N_22872,N_22473,N_22192);
nand U22873 (N_22873,N_22075,N_22236);
and U22874 (N_22874,N_22489,N_22340);
xor U22875 (N_22875,N_22377,N_22090);
or U22876 (N_22876,N_22253,N_22416);
or U22877 (N_22877,N_22018,N_22320);
or U22878 (N_22878,N_22080,N_22170);
xor U22879 (N_22879,N_22168,N_22428);
and U22880 (N_22880,N_22456,N_22335);
or U22881 (N_22881,N_22137,N_22181);
xnor U22882 (N_22882,N_22110,N_22010);
or U22883 (N_22883,N_22215,N_22231);
nor U22884 (N_22884,N_22037,N_22268);
and U22885 (N_22885,N_22401,N_22496);
nand U22886 (N_22886,N_22211,N_22157);
and U22887 (N_22887,N_22464,N_22243);
and U22888 (N_22888,N_22317,N_22307);
or U22889 (N_22889,N_22078,N_22378);
and U22890 (N_22890,N_22079,N_22496);
and U22891 (N_22891,N_22021,N_22227);
nand U22892 (N_22892,N_22208,N_22130);
or U22893 (N_22893,N_22336,N_22299);
nand U22894 (N_22894,N_22254,N_22366);
nor U22895 (N_22895,N_22184,N_22234);
nand U22896 (N_22896,N_22074,N_22160);
and U22897 (N_22897,N_22142,N_22467);
and U22898 (N_22898,N_22326,N_22422);
xnor U22899 (N_22899,N_22352,N_22108);
nor U22900 (N_22900,N_22108,N_22398);
or U22901 (N_22901,N_22450,N_22480);
nand U22902 (N_22902,N_22096,N_22228);
and U22903 (N_22903,N_22053,N_22034);
xor U22904 (N_22904,N_22058,N_22254);
and U22905 (N_22905,N_22053,N_22096);
and U22906 (N_22906,N_22015,N_22366);
nand U22907 (N_22907,N_22318,N_22003);
nor U22908 (N_22908,N_22067,N_22204);
nor U22909 (N_22909,N_22035,N_22439);
xnor U22910 (N_22910,N_22085,N_22282);
nand U22911 (N_22911,N_22403,N_22013);
xor U22912 (N_22912,N_22295,N_22187);
or U22913 (N_22913,N_22322,N_22286);
or U22914 (N_22914,N_22006,N_22003);
or U22915 (N_22915,N_22197,N_22212);
xor U22916 (N_22916,N_22423,N_22180);
xnor U22917 (N_22917,N_22026,N_22318);
nand U22918 (N_22918,N_22085,N_22022);
or U22919 (N_22919,N_22150,N_22194);
and U22920 (N_22920,N_22000,N_22472);
or U22921 (N_22921,N_22022,N_22203);
and U22922 (N_22922,N_22445,N_22158);
nor U22923 (N_22923,N_22339,N_22392);
nand U22924 (N_22924,N_22104,N_22318);
xnor U22925 (N_22925,N_22142,N_22429);
nand U22926 (N_22926,N_22401,N_22077);
and U22927 (N_22927,N_22055,N_22444);
nand U22928 (N_22928,N_22107,N_22197);
nand U22929 (N_22929,N_22404,N_22215);
nor U22930 (N_22930,N_22373,N_22271);
xnor U22931 (N_22931,N_22280,N_22460);
nor U22932 (N_22932,N_22173,N_22183);
nand U22933 (N_22933,N_22359,N_22212);
or U22934 (N_22934,N_22184,N_22189);
nor U22935 (N_22935,N_22144,N_22173);
xor U22936 (N_22936,N_22216,N_22007);
and U22937 (N_22937,N_22051,N_22224);
nand U22938 (N_22938,N_22231,N_22200);
nor U22939 (N_22939,N_22318,N_22305);
and U22940 (N_22940,N_22391,N_22087);
and U22941 (N_22941,N_22340,N_22484);
and U22942 (N_22942,N_22481,N_22101);
nand U22943 (N_22943,N_22021,N_22281);
xnor U22944 (N_22944,N_22399,N_22313);
nor U22945 (N_22945,N_22207,N_22033);
nand U22946 (N_22946,N_22363,N_22377);
and U22947 (N_22947,N_22263,N_22249);
nand U22948 (N_22948,N_22249,N_22217);
and U22949 (N_22949,N_22288,N_22052);
nor U22950 (N_22950,N_22050,N_22091);
nand U22951 (N_22951,N_22007,N_22367);
nor U22952 (N_22952,N_22031,N_22493);
or U22953 (N_22953,N_22227,N_22363);
xor U22954 (N_22954,N_22441,N_22037);
nor U22955 (N_22955,N_22404,N_22259);
and U22956 (N_22956,N_22243,N_22193);
nand U22957 (N_22957,N_22073,N_22366);
xnor U22958 (N_22958,N_22133,N_22400);
or U22959 (N_22959,N_22027,N_22077);
and U22960 (N_22960,N_22100,N_22206);
or U22961 (N_22961,N_22319,N_22441);
nand U22962 (N_22962,N_22453,N_22404);
and U22963 (N_22963,N_22252,N_22223);
and U22964 (N_22964,N_22272,N_22391);
or U22965 (N_22965,N_22344,N_22212);
and U22966 (N_22966,N_22285,N_22188);
or U22967 (N_22967,N_22383,N_22463);
nand U22968 (N_22968,N_22158,N_22423);
nor U22969 (N_22969,N_22111,N_22310);
xor U22970 (N_22970,N_22450,N_22043);
nor U22971 (N_22971,N_22002,N_22494);
xor U22972 (N_22972,N_22170,N_22240);
nor U22973 (N_22973,N_22416,N_22252);
or U22974 (N_22974,N_22053,N_22461);
nor U22975 (N_22975,N_22224,N_22475);
xor U22976 (N_22976,N_22437,N_22089);
nand U22977 (N_22977,N_22391,N_22127);
nor U22978 (N_22978,N_22410,N_22036);
or U22979 (N_22979,N_22246,N_22362);
or U22980 (N_22980,N_22423,N_22065);
nand U22981 (N_22981,N_22156,N_22066);
xor U22982 (N_22982,N_22055,N_22159);
and U22983 (N_22983,N_22452,N_22476);
and U22984 (N_22984,N_22173,N_22313);
nor U22985 (N_22985,N_22212,N_22226);
nor U22986 (N_22986,N_22477,N_22283);
nor U22987 (N_22987,N_22213,N_22042);
or U22988 (N_22988,N_22327,N_22353);
or U22989 (N_22989,N_22087,N_22378);
nor U22990 (N_22990,N_22164,N_22337);
nor U22991 (N_22991,N_22232,N_22003);
or U22992 (N_22992,N_22299,N_22311);
nand U22993 (N_22993,N_22231,N_22173);
nor U22994 (N_22994,N_22057,N_22431);
or U22995 (N_22995,N_22190,N_22335);
or U22996 (N_22996,N_22082,N_22088);
nor U22997 (N_22997,N_22264,N_22006);
and U22998 (N_22998,N_22377,N_22081);
and U22999 (N_22999,N_22035,N_22063);
nand U23000 (N_23000,N_22867,N_22513);
or U23001 (N_23001,N_22924,N_22830);
and U23002 (N_23002,N_22973,N_22877);
or U23003 (N_23003,N_22705,N_22986);
and U23004 (N_23004,N_22645,N_22920);
or U23005 (N_23005,N_22884,N_22788);
and U23006 (N_23006,N_22792,N_22925);
nand U23007 (N_23007,N_22623,N_22827);
or U23008 (N_23008,N_22587,N_22574);
xor U23009 (N_23009,N_22820,N_22807);
and U23010 (N_23010,N_22663,N_22833);
or U23011 (N_23011,N_22941,N_22997);
nand U23012 (N_23012,N_22654,N_22912);
nor U23013 (N_23013,N_22950,N_22904);
or U23014 (N_23014,N_22648,N_22853);
nor U23015 (N_23015,N_22787,N_22710);
xor U23016 (N_23016,N_22745,N_22949);
xor U23017 (N_23017,N_22926,N_22659);
or U23018 (N_23018,N_22693,N_22503);
and U23019 (N_23019,N_22763,N_22982);
and U23020 (N_23020,N_22678,N_22696);
nor U23021 (N_23021,N_22634,N_22768);
and U23022 (N_23022,N_22774,N_22893);
xnor U23023 (N_23023,N_22981,N_22721);
nand U23024 (N_23024,N_22860,N_22551);
or U23025 (N_23025,N_22621,N_22600);
xor U23026 (N_23026,N_22602,N_22773);
nor U23027 (N_23027,N_22980,N_22523);
and U23028 (N_23028,N_22521,N_22501);
and U23029 (N_23029,N_22687,N_22670);
nor U23030 (N_23030,N_22772,N_22970);
and U23031 (N_23031,N_22822,N_22957);
nand U23032 (N_23032,N_22631,N_22714);
nor U23033 (N_23033,N_22847,N_22591);
or U23034 (N_23034,N_22617,N_22979);
xor U23035 (N_23035,N_22756,N_22613);
nor U23036 (N_23036,N_22850,N_22961);
and U23037 (N_23037,N_22858,N_22769);
nor U23038 (N_23038,N_22545,N_22667);
nor U23039 (N_23039,N_22736,N_22895);
nor U23040 (N_23040,N_22878,N_22801);
or U23041 (N_23041,N_22707,N_22864);
nand U23042 (N_23042,N_22798,N_22715);
xor U23043 (N_23043,N_22859,N_22777);
xnor U23044 (N_23044,N_22866,N_22976);
and U23045 (N_23045,N_22977,N_22831);
nand U23046 (N_23046,N_22789,N_22751);
nor U23047 (N_23047,N_22910,N_22594);
xnor U23048 (N_23048,N_22684,N_22532);
nand U23049 (N_23049,N_22557,N_22682);
nor U23050 (N_23050,N_22703,N_22578);
and U23051 (N_23051,N_22708,N_22914);
nand U23052 (N_23052,N_22725,N_22806);
nand U23053 (N_23053,N_22967,N_22996);
and U23054 (N_23054,N_22778,N_22965);
nor U23055 (N_23055,N_22896,N_22985);
and U23056 (N_23056,N_22849,N_22596);
or U23057 (N_23057,N_22731,N_22641);
or U23058 (N_23058,N_22540,N_22931);
and U23059 (N_23059,N_22589,N_22579);
nand U23060 (N_23060,N_22837,N_22702);
nand U23061 (N_23061,N_22507,N_22987);
or U23062 (N_23062,N_22544,N_22894);
nand U23063 (N_23063,N_22658,N_22709);
and U23064 (N_23064,N_22716,N_22584);
or U23065 (N_23065,N_22597,N_22586);
nor U23066 (N_23066,N_22952,N_22771);
xor U23067 (N_23067,N_22585,N_22505);
nor U23068 (N_23068,N_22577,N_22533);
nor U23069 (N_23069,N_22939,N_22560);
nor U23070 (N_23070,N_22992,N_22642);
nand U23071 (N_23071,N_22514,N_22947);
nor U23072 (N_23072,N_22908,N_22516);
or U23073 (N_23073,N_22636,N_22990);
or U23074 (N_23074,N_22828,N_22862);
or U23075 (N_23075,N_22918,N_22512);
or U23076 (N_23076,N_22783,N_22868);
nor U23077 (N_23077,N_22765,N_22601);
or U23078 (N_23078,N_22680,N_22610);
nor U23079 (N_23079,N_22936,N_22564);
xor U23080 (N_23080,N_22762,N_22735);
or U23081 (N_23081,N_22672,N_22741);
or U23082 (N_23082,N_22661,N_22802);
nor U23083 (N_23083,N_22826,N_22846);
nand U23084 (N_23084,N_22842,N_22885);
nor U23085 (N_23085,N_22812,N_22723);
nor U23086 (N_23086,N_22592,N_22993);
and U23087 (N_23087,N_22562,N_22824);
xor U23088 (N_23088,N_22819,N_22852);
xor U23089 (N_23089,N_22500,N_22948);
xnor U23090 (N_23090,N_22711,N_22558);
or U23091 (N_23091,N_22653,N_22886);
or U23092 (N_23092,N_22671,N_22724);
and U23093 (N_23093,N_22882,N_22518);
and U23094 (N_23094,N_22625,N_22855);
nand U23095 (N_23095,N_22938,N_22954);
and U23096 (N_23096,N_22984,N_22757);
or U23097 (N_23097,N_22538,N_22553);
nand U23098 (N_23098,N_22622,N_22676);
xor U23099 (N_23099,N_22836,N_22744);
and U23100 (N_23100,N_22543,N_22699);
nor U23101 (N_23101,N_22835,N_22632);
and U23102 (N_23102,N_22966,N_22962);
nand U23103 (N_23103,N_22905,N_22673);
or U23104 (N_23104,N_22502,N_22999);
and U23105 (N_23105,N_22958,N_22730);
xnor U23106 (N_23106,N_22509,N_22790);
or U23107 (N_23107,N_22548,N_22683);
or U23108 (N_23108,N_22733,N_22616);
and U23109 (N_23109,N_22635,N_22690);
and U23110 (N_23110,N_22619,N_22704);
nor U23111 (N_23111,N_22903,N_22640);
or U23112 (N_23112,N_22732,N_22537);
xor U23113 (N_23113,N_22650,N_22739);
or U23114 (N_23114,N_22565,N_22593);
nand U23115 (N_23115,N_22876,N_22697);
nand U23116 (N_23116,N_22856,N_22701);
and U23117 (N_23117,N_22698,N_22628);
nand U23118 (N_23118,N_22573,N_22655);
xnor U23119 (N_23119,N_22508,N_22604);
nor U23120 (N_23120,N_22590,N_22536);
and U23121 (N_23121,N_22953,N_22688);
xor U23122 (N_23122,N_22529,N_22695);
xnor U23123 (N_23123,N_22898,N_22746);
nor U23124 (N_23124,N_22740,N_22932);
or U23125 (N_23125,N_22607,N_22897);
nor U23126 (N_23126,N_22998,N_22646);
and U23127 (N_23127,N_22825,N_22726);
or U23128 (N_23128,N_22612,N_22720);
nor U23129 (N_23129,N_22764,N_22728);
xnor U23130 (N_23130,N_22951,N_22629);
xnor U23131 (N_23131,N_22840,N_22524);
and U23132 (N_23132,N_22677,N_22839);
nand U23133 (N_23133,N_22813,N_22988);
or U23134 (N_23134,N_22775,N_22566);
or U23135 (N_23135,N_22738,N_22547);
or U23136 (N_23136,N_22916,N_22760);
and U23137 (N_23137,N_22892,N_22517);
nor U23138 (N_23138,N_22755,N_22782);
xnor U23139 (N_23139,N_22615,N_22729);
and U23140 (N_23140,N_22643,N_22575);
or U23141 (N_23141,N_22510,N_22934);
or U23142 (N_23142,N_22700,N_22754);
and U23143 (N_23143,N_22794,N_22972);
nor U23144 (N_23144,N_22675,N_22883);
nor U23145 (N_23145,N_22909,N_22552);
nor U23146 (N_23146,N_22901,N_22656);
nand U23147 (N_23147,N_22913,N_22890);
nor U23148 (N_23148,N_22964,N_22681);
and U23149 (N_23149,N_22861,N_22874);
nor U23150 (N_23150,N_22706,N_22665);
and U23151 (N_23151,N_22571,N_22955);
and U23152 (N_23152,N_22580,N_22569);
or U23153 (N_23153,N_22603,N_22811);
nor U23154 (N_23154,N_22555,N_22821);
nor U23155 (N_23155,N_22791,N_22570);
and U23156 (N_23156,N_22722,N_22804);
nor U23157 (N_23157,N_22823,N_22511);
nand U23158 (N_23158,N_22797,N_22618);
nand U23159 (N_23159,N_22686,N_22749);
nor U23160 (N_23160,N_22857,N_22796);
and U23161 (N_23161,N_22567,N_22525);
nor U23162 (N_23162,N_22546,N_22832);
nor U23163 (N_23163,N_22515,N_22539);
and U23164 (N_23164,N_22759,N_22713);
nand U23165 (N_23165,N_22712,N_22810);
nor U23166 (N_23166,N_22550,N_22679);
xnor U23167 (N_23167,N_22906,N_22968);
nor U23168 (N_23168,N_22556,N_22752);
xnor U23169 (N_23169,N_22753,N_22887);
or U23170 (N_23170,N_22929,N_22814);
nor U23171 (N_23171,N_22803,N_22785);
xor U23172 (N_23172,N_22647,N_22637);
or U23173 (N_23173,N_22917,N_22923);
nand U23174 (N_23174,N_22871,N_22599);
and U23175 (N_23175,N_22776,N_22535);
nand U23176 (N_23176,N_22651,N_22534);
xor U23177 (N_23177,N_22668,N_22624);
nor U23178 (N_23178,N_22638,N_22927);
and U23179 (N_23179,N_22542,N_22626);
nor U23180 (N_23180,N_22800,N_22915);
nand U23181 (N_23181,N_22748,N_22946);
xor U23182 (N_23182,N_22943,N_22719);
or U23183 (N_23183,N_22891,N_22974);
nor U23184 (N_23184,N_22963,N_22660);
nand U23185 (N_23185,N_22817,N_22530);
or U23186 (N_23186,N_22689,N_22921);
and U23187 (N_23187,N_22605,N_22779);
nand U23188 (N_23188,N_22780,N_22971);
and U23189 (N_23189,N_22742,N_22793);
nor U23190 (N_23190,N_22994,N_22956);
nor U23191 (N_23191,N_22899,N_22900);
xnor U23192 (N_23192,N_22843,N_22922);
xor U23193 (N_23193,N_22691,N_22588);
xnor U23194 (N_23194,N_22649,N_22737);
xnor U23195 (N_23195,N_22606,N_22718);
nand U23196 (N_23196,N_22975,N_22944);
nand U23197 (N_23197,N_22863,N_22669);
xor U23198 (N_23198,N_22506,N_22928);
nor U23199 (N_23199,N_22829,N_22657);
or U23200 (N_23200,N_22614,N_22609);
or U23201 (N_23201,N_22834,N_22662);
or U23202 (N_23202,N_22809,N_22784);
xnor U23203 (N_23203,N_22870,N_22630);
or U23204 (N_23204,N_22781,N_22559);
nand U23205 (N_23205,N_22845,N_22945);
xnor U23206 (N_23206,N_22816,N_22937);
and U23207 (N_23207,N_22935,N_22983);
nor U23208 (N_23208,N_22561,N_22750);
or U23209 (N_23209,N_22572,N_22583);
nor U23210 (N_23210,N_22608,N_22865);
nand U23211 (N_23211,N_22881,N_22554);
xnor U23212 (N_23212,N_22611,N_22815);
nor U23213 (N_23213,N_22805,N_22664);
nor U23214 (N_23214,N_22844,N_22519);
nor U23215 (N_23215,N_22879,N_22598);
nor U23216 (N_23216,N_22685,N_22851);
nand U23217 (N_23217,N_22991,N_22727);
xnor U23218 (N_23218,N_22639,N_22902);
xor U23219 (N_23219,N_22989,N_22959);
nand U23220 (N_23220,N_22581,N_22767);
or U23221 (N_23221,N_22869,N_22969);
and U23222 (N_23222,N_22888,N_22854);
and U23223 (N_23223,N_22717,N_22995);
xnor U23224 (N_23224,N_22576,N_22940);
nand U23225 (N_23225,N_22520,N_22549);
nand U23226 (N_23226,N_22582,N_22692);
nand U23227 (N_23227,N_22786,N_22978);
and U23228 (N_23228,N_22531,N_22620);
or U23229 (N_23229,N_22911,N_22522);
xnor U23230 (N_23230,N_22933,N_22528);
and U23231 (N_23231,N_22818,N_22960);
xor U23232 (N_23232,N_22799,N_22541);
and U23233 (N_23233,N_22942,N_22873);
or U23234 (N_23234,N_22644,N_22734);
xnor U23235 (N_23235,N_22568,N_22504);
nand U23236 (N_23236,N_22758,N_22766);
nand U23237 (N_23237,N_22907,N_22674);
xor U23238 (N_23238,N_22880,N_22889);
xnor U23239 (N_23239,N_22808,N_22930);
nor U23240 (N_23240,N_22795,N_22633);
xnor U23241 (N_23241,N_22872,N_22761);
or U23242 (N_23242,N_22848,N_22838);
nor U23243 (N_23243,N_22694,N_22841);
and U23244 (N_23244,N_22563,N_22595);
and U23245 (N_23245,N_22875,N_22526);
and U23246 (N_23246,N_22919,N_22627);
or U23247 (N_23247,N_22666,N_22747);
and U23248 (N_23248,N_22770,N_22527);
nand U23249 (N_23249,N_22652,N_22743);
nor U23250 (N_23250,N_22908,N_22620);
xor U23251 (N_23251,N_22669,N_22743);
or U23252 (N_23252,N_22770,N_22856);
and U23253 (N_23253,N_22627,N_22625);
nor U23254 (N_23254,N_22896,N_22906);
and U23255 (N_23255,N_22731,N_22839);
and U23256 (N_23256,N_22941,N_22979);
or U23257 (N_23257,N_22780,N_22686);
nand U23258 (N_23258,N_22509,N_22590);
nand U23259 (N_23259,N_22528,N_22782);
nor U23260 (N_23260,N_22750,N_22719);
and U23261 (N_23261,N_22599,N_22884);
nor U23262 (N_23262,N_22509,N_22708);
nand U23263 (N_23263,N_22562,N_22589);
and U23264 (N_23264,N_22510,N_22900);
nand U23265 (N_23265,N_22635,N_22876);
nor U23266 (N_23266,N_22606,N_22926);
nor U23267 (N_23267,N_22559,N_22886);
and U23268 (N_23268,N_22774,N_22837);
or U23269 (N_23269,N_22851,N_22773);
and U23270 (N_23270,N_22794,N_22699);
and U23271 (N_23271,N_22803,N_22858);
nor U23272 (N_23272,N_22761,N_22551);
nand U23273 (N_23273,N_22775,N_22888);
and U23274 (N_23274,N_22651,N_22780);
or U23275 (N_23275,N_22968,N_22894);
or U23276 (N_23276,N_22707,N_22936);
nand U23277 (N_23277,N_22509,N_22625);
nand U23278 (N_23278,N_22715,N_22933);
xor U23279 (N_23279,N_22597,N_22830);
nor U23280 (N_23280,N_22754,N_22728);
xor U23281 (N_23281,N_22906,N_22849);
nand U23282 (N_23282,N_22901,N_22629);
xor U23283 (N_23283,N_22970,N_22628);
or U23284 (N_23284,N_22692,N_22753);
nand U23285 (N_23285,N_22652,N_22632);
or U23286 (N_23286,N_22817,N_22887);
or U23287 (N_23287,N_22799,N_22807);
xnor U23288 (N_23288,N_22736,N_22846);
or U23289 (N_23289,N_22869,N_22970);
xor U23290 (N_23290,N_22847,N_22778);
nand U23291 (N_23291,N_22526,N_22580);
nand U23292 (N_23292,N_22655,N_22788);
and U23293 (N_23293,N_22544,N_22875);
and U23294 (N_23294,N_22969,N_22755);
nand U23295 (N_23295,N_22924,N_22951);
or U23296 (N_23296,N_22995,N_22531);
nand U23297 (N_23297,N_22540,N_22684);
and U23298 (N_23298,N_22774,N_22730);
xnor U23299 (N_23299,N_22948,N_22700);
nor U23300 (N_23300,N_22934,N_22546);
nand U23301 (N_23301,N_22584,N_22865);
nand U23302 (N_23302,N_22596,N_22615);
xnor U23303 (N_23303,N_22511,N_22700);
nor U23304 (N_23304,N_22898,N_22703);
xor U23305 (N_23305,N_22563,N_22667);
or U23306 (N_23306,N_22732,N_22947);
nand U23307 (N_23307,N_22835,N_22918);
and U23308 (N_23308,N_22636,N_22846);
xor U23309 (N_23309,N_22830,N_22654);
nor U23310 (N_23310,N_22560,N_22635);
xnor U23311 (N_23311,N_22754,N_22777);
and U23312 (N_23312,N_22650,N_22587);
nor U23313 (N_23313,N_22708,N_22994);
nor U23314 (N_23314,N_22791,N_22793);
xor U23315 (N_23315,N_22757,N_22964);
nand U23316 (N_23316,N_22914,N_22776);
xor U23317 (N_23317,N_22695,N_22835);
or U23318 (N_23318,N_22743,N_22666);
or U23319 (N_23319,N_22979,N_22735);
and U23320 (N_23320,N_22933,N_22802);
and U23321 (N_23321,N_22843,N_22710);
or U23322 (N_23322,N_22864,N_22731);
nor U23323 (N_23323,N_22786,N_22932);
or U23324 (N_23324,N_22795,N_22504);
nand U23325 (N_23325,N_22813,N_22976);
nand U23326 (N_23326,N_22859,N_22689);
xor U23327 (N_23327,N_22786,N_22750);
or U23328 (N_23328,N_22544,N_22824);
xnor U23329 (N_23329,N_22645,N_22997);
and U23330 (N_23330,N_22767,N_22931);
and U23331 (N_23331,N_22538,N_22945);
or U23332 (N_23332,N_22842,N_22742);
xnor U23333 (N_23333,N_22574,N_22968);
nor U23334 (N_23334,N_22502,N_22865);
nor U23335 (N_23335,N_22899,N_22861);
and U23336 (N_23336,N_22978,N_22723);
and U23337 (N_23337,N_22603,N_22939);
and U23338 (N_23338,N_22554,N_22945);
nor U23339 (N_23339,N_22839,N_22858);
and U23340 (N_23340,N_22826,N_22646);
xor U23341 (N_23341,N_22774,N_22975);
xnor U23342 (N_23342,N_22810,N_22559);
nand U23343 (N_23343,N_22641,N_22968);
and U23344 (N_23344,N_22564,N_22506);
xnor U23345 (N_23345,N_22610,N_22554);
and U23346 (N_23346,N_22654,N_22828);
and U23347 (N_23347,N_22814,N_22904);
or U23348 (N_23348,N_22856,N_22532);
or U23349 (N_23349,N_22577,N_22921);
xor U23350 (N_23350,N_22726,N_22988);
or U23351 (N_23351,N_22707,N_22684);
nor U23352 (N_23352,N_22521,N_22716);
and U23353 (N_23353,N_22707,N_22925);
or U23354 (N_23354,N_22691,N_22901);
and U23355 (N_23355,N_22902,N_22845);
nand U23356 (N_23356,N_22898,N_22732);
or U23357 (N_23357,N_22951,N_22838);
nor U23358 (N_23358,N_22979,N_22624);
and U23359 (N_23359,N_22509,N_22959);
xnor U23360 (N_23360,N_22742,N_22817);
and U23361 (N_23361,N_22801,N_22702);
xnor U23362 (N_23362,N_22606,N_22655);
nand U23363 (N_23363,N_22621,N_22884);
nand U23364 (N_23364,N_22958,N_22792);
nor U23365 (N_23365,N_22830,N_22504);
or U23366 (N_23366,N_22514,N_22999);
or U23367 (N_23367,N_22971,N_22683);
xnor U23368 (N_23368,N_22989,N_22751);
or U23369 (N_23369,N_22548,N_22999);
nand U23370 (N_23370,N_22517,N_22580);
and U23371 (N_23371,N_22675,N_22505);
xor U23372 (N_23372,N_22657,N_22806);
nor U23373 (N_23373,N_22977,N_22596);
nor U23374 (N_23374,N_22562,N_22501);
or U23375 (N_23375,N_22769,N_22836);
nand U23376 (N_23376,N_22707,N_22898);
nor U23377 (N_23377,N_22636,N_22750);
or U23378 (N_23378,N_22883,N_22946);
xnor U23379 (N_23379,N_22800,N_22804);
nor U23380 (N_23380,N_22557,N_22567);
xor U23381 (N_23381,N_22954,N_22881);
nand U23382 (N_23382,N_22690,N_22576);
or U23383 (N_23383,N_22904,N_22764);
nor U23384 (N_23384,N_22815,N_22752);
or U23385 (N_23385,N_22580,N_22518);
and U23386 (N_23386,N_22658,N_22987);
or U23387 (N_23387,N_22979,N_22532);
nor U23388 (N_23388,N_22994,N_22974);
nor U23389 (N_23389,N_22849,N_22769);
or U23390 (N_23390,N_22593,N_22878);
or U23391 (N_23391,N_22813,N_22560);
nand U23392 (N_23392,N_22918,N_22529);
or U23393 (N_23393,N_22854,N_22775);
or U23394 (N_23394,N_22692,N_22909);
xnor U23395 (N_23395,N_22509,N_22990);
and U23396 (N_23396,N_22951,N_22531);
nand U23397 (N_23397,N_22851,N_22593);
or U23398 (N_23398,N_22504,N_22752);
or U23399 (N_23399,N_22533,N_22510);
or U23400 (N_23400,N_22892,N_22917);
or U23401 (N_23401,N_22610,N_22877);
and U23402 (N_23402,N_22640,N_22993);
nor U23403 (N_23403,N_22826,N_22877);
and U23404 (N_23404,N_22928,N_22910);
and U23405 (N_23405,N_22804,N_22853);
nand U23406 (N_23406,N_22560,N_22885);
nor U23407 (N_23407,N_22657,N_22763);
or U23408 (N_23408,N_22927,N_22870);
and U23409 (N_23409,N_22813,N_22777);
xor U23410 (N_23410,N_22620,N_22547);
or U23411 (N_23411,N_22978,N_22658);
nor U23412 (N_23412,N_22655,N_22902);
or U23413 (N_23413,N_22880,N_22563);
xnor U23414 (N_23414,N_22866,N_22523);
nand U23415 (N_23415,N_22585,N_22801);
nand U23416 (N_23416,N_22836,N_22914);
nand U23417 (N_23417,N_22788,N_22837);
nand U23418 (N_23418,N_22918,N_22857);
and U23419 (N_23419,N_22765,N_22793);
nand U23420 (N_23420,N_22965,N_22584);
xor U23421 (N_23421,N_22590,N_22581);
and U23422 (N_23422,N_22595,N_22545);
xor U23423 (N_23423,N_22969,N_22984);
xnor U23424 (N_23424,N_22677,N_22997);
and U23425 (N_23425,N_22768,N_22708);
xnor U23426 (N_23426,N_22907,N_22993);
or U23427 (N_23427,N_22709,N_22637);
or U23428 (N_23428,N_22897,N_22518);
xor U23429 (N_23429,N_22727,N_22988);
xnor U23430 (N_23430,N_22805,N_22627);
nor U23431 (N_23431,N_22623,N_22699);
xnor U23432 (N_23432,N_22964,N_22751);
xnor U23433 (N_23433,N_22541,N_22673);
and U23434 (N_23434,N_22621,N_22838);
xor U23435 (N_23435,N_22675,N_22790);
or U23436 (N_23436,N_22684,N_22644);
xor U23437 (N_23437,N_22995,N_22501);
nand U23438 (N_23438,N_22592,N_22703);
nand U23439 (N_23439,N_22819,N_22993);
nor U23440 (N_23440,N_22848,N_22535);
nand U23441 (N_23441,N_22502,N_22776);
or U23442 (N_23442,N_22712,N_22575);
nand U23443 (N_23443,N_22918,N_22873);
and U23444 (N_23444,N_22961,N_22856);
nor U23445 (N_23445,N_22638,N_22579);
nand U23446 (N_23446,N_22815,N_22736);
xnor U23447 (N_23447,N_22982,N_22782);
xnor U23448 (N_23448,N_22508,N_22992);
or U23449 (N_23449,N_22674,N_22603);
or U23450 (N_23450,N_22969,N_22571);
and U23451 (N_23451,N_22898,N_22589);
or U23452 (N_23452,N_22650,N_22910);
xor U23453 (N_23453,N_22875,N_22677);
xor U23454 (N_23454,N_22872,N_22531);
nand U23455 (N_23455,N_22682,N_22627);
nand U23456 (N_23456,N_22555,N_22677);
or U23457 (N_23457,N_22771,N_22832);
and U23458 (N_23458,N_22980,N_22868);
and U23459 (N_23459,N_22693,N_22911);
or U23460 (N_23460,N_22538,N_22846);
or U23461 (N_23461,N_22653,N_22609);
xnor U23462 (N_23462,N_22939,N_22581);
nand U23463 (N_23463,N_22918,N_22604);
xor U23464 (N_23464,N_22705,N_22627);
nor U23465 (N_23465,N_22536,N_22966);
nor U23466 (N_23466,N_22764,N_22518);
nand U23467 (N_23467,N_22509,N_22876);
and U23468 (N_23468,N_22571,N_22915);
nand U23469 (N_23469,N_22532,N_22698);
nor U23470 (N_23470,N_22554,N_22783);
nor U23471 (N_23471,N_22769,N_22639);
or U23472 (N_23472,N_22897,N_22613);
and U23473 (N_23473,N_22791,N_22549);
or U23474 (N_23474,N_22549,N_22505);
xor U23475 (N_23475,N_22674,N_22520);
and U23476 (N_23476,N_22784,N_22543);
xnor U23477 (N_23477,N_22745,N_22814);
nor U23478 (N_23478,N_22849,N_22902);
xor U23479 (N_23479,N_22933,N_22841);
nor U23480 (N_23480,N_22787,N_22861);
and U23481 (N_23481,N_22860,N_22687);
nor U23482 (N_23482,N_22999,N_22762);
and U23483 (N_23483,N_22979,N_22918);
nor U23484 (N_23484,N_22697,N_22546);
or U23485 (N_23485,N_22681,N_22564);
and U23486 (N_23486,N_22786,N_22675);
xnor U23487 (N_23487,N_22630,N_22924);
or U23488 (N_23488,N_22599,N_22925);
nor U23489 (N_23489,N_22852,N_22553);
xor U23490 (N_23490,N_22625,N_22569);
xor U23491 (N_23491,N_22617,N_22646);
xnor U23492 (N_23492,N_22781,N_22901);
or U23493 (N_23493,N_22787,N_22746);
and U23494 (N_23494,N_22755,N_22728);
and U23495 (N_23495,N_22979,N_22670);
xnor U23496 (N_23496,N_22821,N_22559);
and U23497 (N_23497,N_22881,N_22835);
or U23498 (N_23498,N_22934,N_22744);
nor U23499 (N_23499,N_22735,N_22716);
and U23500 (N_23500,N_23133,N_23345);
xor U23501 (N_23501,N_23462,N_23492);
or U23502 (N_23502,N_23113,N_23474);
nand U23503 (N_23503,N_23189,N_23134);
and U23504 (N_23504,N_23114,N_23188);
nor U23505 (N_23505,N_23344,N_23022);
or U23506 (N_23506,N_23318,N_23436);
nand U23507 (N_23507,N_23351,N_23000);
nor U23508 (N_23508,N_23050,N_23235);
nor U23509 (N_23509,N_23300,N_23006);
xor U23510 (N_23510,N_23168,N_23037);
and U23511 (N_23511,N_23288,N_23031);
nor U23512 (N_23512,N_23232,N_23122);
or U23513 (N_23513,N_23417,N_23066);
xor U23514 (N_23514,N_23392,N_23103);
and U23515 (N_23515,N_23098,N_23328);
and U23516 (N_23516,N_23401,N_23322);
nand U23517 (N_23517,N_23280,N_23120);
and U23518 (N_23518,N_23337,N_23061);
xor U23519 (N_23519,N_23316,N_23338);
nor U23520 (N_23520,N_23495,N_23472);
xor U23521 (N_23521,N_23071,N_23083);
nor U23522 (N_23522,N_23175,N_23262);
nand U23523 (N_23523,N_23226,N_23329);
nor U23524 (N_23524,N_23433,N_23258);
xor U23525 (N_23525,N_23424,N_23169);
xnor U23526 (N_23526,N_23397,N_23459);
or U23527 (N_23527,N_23242,N_23172);
or U23528 (N_23528,N_23427,N_23039);
or U23529 (N_23529,N_23295,N_23382);
nand U23530 (N_23530,N_23185,N_23221);
nand U23531 (N_23531,N_23480,N_23135);
nor U23532 (N_23532,N_23278,N_23155);
or U23533 (N_23533,N_23217,N_23012);
xnor U23534 (N_23534,N_23091,N_23241);
nor U23535 (N_23535,N_23391,N_23104);
and U23536 (N_23536,N_23054,N_23115);
nor U23537 (N_23537,N_23149,N_23013);
or U23538 (N_23538,N_23056,N_23180);
and U23539 (N_23539,N_23411,N_23121);
xnor U23540 (N_23540,N_23245,N_23257);
nand U23541 (N_23541,N_23111,N_23036);
nor U23542 (N_23542,N_23171,N_23034);
nor U23543 (N_23543,N_23364,N_23255);
or U23544 (N_23544,N_23100,N_23314);
and U23545 (N_23545,N_23365,N_23461);
and U23546 (N_23546,N_23445,N_23488);
and U23547 (N_23547,N_23279,N_23299);
nor U23548 (N_23548,N_23118,N_23271);
nand U23549 (N_23549,N_23035,N_23192);
nor U23550 (N_23550,N_23044,N_23159);
xor U23551 (N_23551,N_23415,N_23346);
and U23552 (N_23552,N_23307,N_23088);
and U23553 (N_23553,N_23208,N_23440);
nor U23554 (N_23554,N_23116,N_23040);
and U23555 (N_23555,N_23426,N_23306);
xor U23556 (N_23556,N_23292,N_23386);
nor U23557 (N_23557,N_23026,N_23330);
or U23558 (N_23558,N_23482,N_23249);
and U23559 (N_23559,N_23049,N_23222);
nand U23560 (N_23560,N_23231,N_23315);
nand U23561 (N_23561,N_23448,N_23234);
and U23562 (N_23562,N_23290,N_23097);
xor U23563 (N_23563,N_23385,N_23106);
nand U23564 (N_23564,N_23205,N_23112);
xnor U23565 (N_23565,N_23340,N_23124);
xnor U23566 (N_23566,N_23291,N_23261);
or U23567 (N_23567,N_23094,N_23178);
or U23568 (N_23568,N_23442,N_23408);
xnor U23569 (N_23569,N_23407,N_23151);
nand U23570 (N_23570,N_23360,N_23263);
or U23571 (N_23571,N_23047,N_23468);
nor U23572 (N_23572,N_23019,N_23405);
nand U23573 (N_23573,N_23355,N_23005);
and U23574 (N_23574,N_23395,N_23252);
or U23575 (N_23575,N_23033,N_23419);
xor U23576 (N_23576,N_23285,N_23260);
or U23577 (N_23577,N_23313,N_23282);
nand U23578 (N_23578,N_23399,N_23420);
and U23579 (N_23579,N_23493,N_23418);
or U23580 (N_23580,N_23335,N_23020);
or U23581 (N_23581,N_23014,N_23219);
nand U23582 (N_23582,N_23085,N_23238);
or U23583 (N_23583,N_23001,N_23389);
nor U23584 (N_23584,N_23074,N_23491);
nor U23585 (N_23585,N_23007,N_23366);
and U23586 (N_23586,N_23394,N_23177);
and U23587 (N_23587,N_23297,N_23204);
xnor U23588 (N_23588,N_23356,N_23421);
xor U23589 (N_23589,N_23136,N_23131);
xnor U23590 (N_23590,N_23009,N_23494);
nor U23591 (N_23591,N_23464,N_23467);
or U23592 (N_23592,N_23406,N_23368);
nor U23593 (N_23593,N_23473,N_23326);
or U23594 (N_23594,N_23447,N_23072);
nor U23595 (N_23595,N_23293,N_23196);
or U23596 (N_23596,N_23471,N_23281);
nand U23597 (N_23597,N_23361,N_23422);
and U23598 (N_23598,N_23075,N_23287);
nand U23599 (N_23599,N_23150,N_23463);
nand U23600 (N_23600,N_23441,N_23298);
and U23601 (N_23601,N_23230,N_23302);
or U23602 (N_23602,N_23373,N_23450);
nor U23603 (N_23603,N_23046,N_23478);
and U23604 (N_23604,N_23331,N_23080);
xnor U23605 (N_23605,N_23431,N_23224);
or U23606 (N_23606,N_23200,N_23206);
xnor U23607 (N_23607,N_23376,N_23380);
or U23608 (N_23608,N_23324,N_23123);
or U23609 (N_23609,N_23301,N_23455);
nand U23610 (N_23610,N_23030,N_23213);
or U23611 (N_23611,N_23363,N_23065);
xnor U23612 (N_23612,N_23476,N_23430);
or U23613 (N_23613,N_23108,N_23129);
and U23614 (N_23614,N_23244,N_23143);
or U23615 (N_23615,N_23070,N_23349);
xnor U23616 (N_23616,N_23369,N_23400);
and U23617 (N_23617,N_23081,N_23348);
nor U23618 (N_23618,N_23485,N_23449);
nand U23619 (N_23619,N_23225,N_23011);
xor U23620 (N_23620,N_23409,N_23269);
nand U23621 (N_23621,N_23055,N_23381);
nand U23622 (N_23622,N_23499,N_23358);
and U23623 (N_23623,N_23148,N_23038);
or U23624 (N_23624,N_23387,N_23139);
and U23625 (N_23625,N_23132,N_23145);
and U23626 (N_23626,N_23275,N_23021);
nand U23627 (N_23627,N_23157,N_23137);
and U23628 (N_23628,N_23342,N_23119);
xor U23629 (N_23629,N_23062,N_23432);
xor U23630 (N_23630,N_23125,N_23227);
or U23631 (N_23631,N_23203,N_23060);
or U23632 (N_23632,N_23353,N_23460);
nor U23633 (N_23633,N_23439,N_23423);
nor U23634 (N_23634,N_23246,N_23379);
xor U23635 (N_23635,N_23454,N_23265);
nand U23636 (N_23636,N_23105,N_23152);
xor U23637 (N_23637,N_23236,N_23296);
and U23638 (N_23638,N_23087,N_23211);
and U23639 (N_23639,N_23154,N_23190);
nor U23640 (N_23640,N_23174,N_23384);
or U23641 (N_23641,N_23202,N_23248);
xor U23642 (N_23642,N_23179,N_23479);
or U23643 (N_23643,N_23093,N_23414);
xor U23644 (N_23644,N_23220,N_23374);
nand U23645 (N_23645,N_23141,N_23371);
and U23646 (N_23646,N_23194,N_23250);
nand U23647 (N_23647,N_23140,N_23166);
xor U23648 (N_23648,N_23067,N_23308);
xnor U23649 (N_23649,N_23270,N_23429);
xor U23650 (N_23650,N_23048,N_23084);
or U23651 (N_23651,N_23162,N_23210);
xnor U23652 (N_23652,N_23413,N_23333);
nand U23653 (N_23653,N_23023,N_23228);
nor U23654 (N_23654,N_23193,N_23233);
or U23655 (N_23655,N_23195,N_23101);
or U23656 (N_23656,N_23239,N_23216);
xnor U23657 (N_23657,N_23410,N_23069);
and U23658 (N_23658,N_23343,N_23428);
xor U23659 (N_23659,N_23045,N_23486);
nand U23660 (N_23660,N_23041,N_23497);
or U23661 (N_23661,N_23016,N_23332);
or U23662 (N_23662,N_23452,N_23443);
nand U23663 (N_23663,N_23393,N_23465);
or U23664 (N_23664,N_23483,N_23444);
and U23665 (N_23665,N_23187,N_23086);
nor U23666 (N_23666,N_23043,N_23117);
nor U23667 (N_23667,N_23218,N_23456);
or U23668 (N_23668,N_23243,N_23147);
or U23669 (N_23669,N_23289,N_23372);
nor U23670 (N_23670,N_23357,N_23215);
and U23671 (N_23671,N_23490,N_23068);
nand U23672 (N_23672,N_23237,N_23469);
nand U23673 (N_23673,N_23323,N_23176);
xnor U23674 (N_23674,N_23077,N_23303);
or U23675 (N_23675,N_23317,N_23339);
and U23676 (N_23676,N_23453,N_23199);
nor U23677 (N_23677,N_23256,N_23446);
xnor U23678 (N_23678,N_23102,N_23277);
or U23679 (N_23679,N_23063,N_23350);
nand U23680 (N_23680,N_23425,N_23398);
nand U23681 (N_23681,N_23484,N_23027);
or U23682 (N_23682,N_23390,N_23092);
or U23683 (N_23683,N_23017,N_23223);
and U23684 (N_23684,N_23264,N_23470);
and U23685 (N_23685,N_23259,N_23325);
or U23686 (N_23686,N_23286,N_23186);
nand U23687 (N_23687,N_23240,N_23438);
nand U23688 (N_23688,N_23073,N_23367);
and U23689 (N_23689,N_23352,N_23146);
nand U23690 (N_23690,N_23181,N_23434);
nand U23691 (N_23691,N_23251,N_23138);
xor U23692 (N_23692,N_23311,N_23274);
nor U23693 (N_23693,N_23182,N_23008);
or U23694 (N_23694,N_23029,N_23058);
nand U23695 (N_23695,N_23183,N_23128);
xor U23696 (N_23696,N_23018,N_23078);
xnor U23697 (N_23697,N_23321,N_23396);
and U23698 (N_23698,N_23253,N_23403);
or U23699 (N_23699,N_23336,N_23377);
xor U23700 (N_23700,N_23266,N_23082);
xnor U23701 (N_23701,N_23099,N_23341);
and U23702 (N_23702,N_23170,N_23370);
nand U23703 (N_23703,N_23052,N_23109);
nor U23704 (N_23704,N_23003,N_23076);
xnor U23705 (N_23705,N_23327,N_23404);
or U23706 (N_23706,N_23412,N_23004);
nand U23707 (N_23707,N_23028,N_23110);
xnor U23708 (N_23708,N_23229,N_23284);
nand U23709 (N_23709,N_23214,N_23267);
xnor U23710 (N_23710,N_23156,N_23487);
nand U23711 (N_23711,N_23126,N_23362);
nor U23712 (N_23712,N_23184,N_23160);
nand U23713 (N_23713,N_23107,N_23198);
and U23714 (N_23714,N_23466,N_23320);
nand U23715 (N_23715,N_23144,N_23312);
nor U23716 (N_23716,N_23191,N_23359);
or U23717 (N_23717,N_23272,N_23051);
or U23718 (N_23718,N_23207,N_23010);
or U23719 (N_23719,N_23015,N_23304);
and U23720 (N_23720,N_23130,N_23163);
and U23721 (N_23721,N_23276,N_23002);
or U23722 (N_23722,N_23388,N_23153);
nand U23723 (N_23723,N_23212,N_23498);
and U23724 (N_23724,N_23142,N_23268);
and U23725 (N_23725,N_23477,N_23209);
and U23726 (N_23726,N_23095,N_23319);
or U23727 (N_23727,N_23375,N_23247);
nor U23728 (N_23728,N_23057,N_23402);
nor U23729 (N_23729,N_23089,N_23489);
xnor U23730 (N_23730,N_23475,N_23173);
xor U23731 (N_23731,N_23096,N_23053);
xor U23732 (N_23732,N_23334,N_23161);
or U23733 (N_23733,N_23201,N_23294);
and U23734 (N_23734,N_23197,N_23309);
xnor U23735 (N_23735,N_23310,N_23254);
or U23736 (N_23736,N_23024,N_23435);
nand U23737 (N_23737,N_23273,N_23451);
xnor U23738 (N_23738,N_23496,N_23378);
nor U23739 (N_23739,N_23158,N_23437);
nand U23740 (N_23740,N_23458,N_23383);
nor U23741 (N_23741,N_23165,N_23032);
nor U23742 (N_23742,N_23090,N_23481);
or U23743 (N_23743,N_23416,N_23064);
and U23744 (N_23744,N_23025,N_23059);
and U23745 (N_23745,N_23283,N_23042);
nor U23746 (N_23746,N_23347,N_23079);
nand U23747 (N_23747,N_23354,N_23457);
nor U23748 (N_23748,N_23167,N_23164);
or U23749 (N_23749,N_23127,N_23305);
xor U23750 (N_23750,N_23276,N_23026);
nor U23751 (N_23751,N_23079,N_23295);
nand U23752 (N_23752,N_23162,N_23456);
xnor U23753 (N_23753,N_23194,N_23227);
nand U23754 (N_23754,N_23067,N_23395);
nor U23755 (N_23755,N_23169,N_23289);
or U23756 (N_23756,N_23265,N_23151);
nand U23757 (N_23757,N_23461,N_23205);
or U23758 (N_23758,N_23188,N_23231);
and U23759 (N_23759,N_23146,N_23482);
nor U23760 (N_23760,N_23043,N_23006);
xor U23761 (N_23761,N_23144,N_23417);
or U23762 (N_23762,N_23178,N_23047);
or U23763 (N_23763,N_23096,N_23066);
nand U23764 (N_23764,N_23038,N_23104);
xor U23765 (N_23765,N_23062,N_23218);
or U23766 (N_23766,N_23242,N_23294);
nand U23767 (N_23767,N_23423,N_23197);
and U23768 (N_23768,N_23491,N_23272);
nand U23769 (N_23769,N_23217,N_23094);
nand U23770 (N_23770,N_23080,N_23460);
xor U23771 (N_23771,N_23195,N_23187);
and U23772 (N_23772,N_23417,N_23391);
nand U23773 (N_23773,N_23152,N_23430);
xor U23774 (N_23774,N_23005,N_23216);
and U23775 (N_23775,N_23384,N_23385);
nand U23776 (N_23776,N_23329,N_23129);
nand U23777 (N_23777,N_23123,N_23165);
nor U23778 (N_23778,N_23258,N_23391);
nor U23779 (N_23779,N_23335,N_23405);
nand U23780 (N_23780,N_23418,N_23159);
or U23781 (N_23781,N_23064,N_23404);
nor U23782 (N_23782,N_23085,N_23152);
xor U23783 (N_23783,N_23233,N_23088);
nor U23784 (N_23784,N_23372,N_23241);
and U23785 (N_23785,N_23374,N_23016);
xor U23786 (N_23786,N_23113,N_23304);
and U23787 (N_23787,N_23003,N_23444);
or U23788 (N_23788,N_23298,N_23036);
nor U23789 (N_23789,N_23205,N_23032);
nand U23790 (N_23790,N_23006,N_23306);
and U23791 (N_23791,N_23350,N_23422);
xnor U23792 (N_23792,N_23041,N_23168);
nand U23793 (N_23793,N_23258,N_23264);
nand U23794 (N_23794,N_23369,N_23066);
nor U23795 (N_23795,N_23194,N_23212);
nor U23796 (N_23796,N_23266,N_23466);
nor U23797 (N_23797,N_23265,N_23307);
nand U23798 (N_23798,N_23443,N_23127);
and U23799 (N_23799,N_23177,N_23063);
xnor U23800 (N_23800,N_23026,N_23239);
or U23801 (N_23801,N_23435,N_23151);
nor U23802 (N_23802,N_23261,N_23368);
and U23803 (N_23803,N_23399,N_23086);
xnor U23804 (N_23804,N_23373,N_23006);
nor U23805 (N_23805,N_23364,N_23292);
nand U23806 (N_23806,N_23334,N_23162);
nor U23807 (N_23807,N_23492,N_23192);
xnor U23808 (N_23808,N_23297,N_23085);
nand U23809 (N_23809,N_23155,N_23170);
or U23810 (N_23810,N_23214,N_23414);
and U23811 (N_23811,N_23241,N_23240);
and U23812 (N_23812,N_23024,N_23098);
nor U23813 (N_23813,N_23486,N_23154);
nor U23814 (N_23814,N_23286,N_23455);
nand U23815 (N_23815,N_23077,N_23112);
xnor U23816 (N_23816,N_23061,N_23249);
and U23817 (N_23817,N_23477,N_23364);
nor U23818 (N_23818,N_23258,N_23450);
xnor U23819 (N_23819,N_23447,N_23304);
nand U23820 (N_23820,N_23398,N_23121);
and U23821 (N_23821,N_23054,N_23088);
or U23822 (N_23822,N_23286,N_23335);
or U23823 (N_23823,N_23195,N_23203);
nor U23824 (N_23824,N_23024,N_23458);
xor U23825 (N_23825,N_23407,N_23461);
xnor U23826 (N_23826,N_23162,N_23480);
xor U23827 (N_23827,N_23051,N_23425);
xnor U23828 (N_23828,N_23062,N_23398);
and U23829 (N_23829,N_23281,N_23314);
or U23830 (N_23830,N_23425,N_23142);
and U23831 (N_23831,N_23443,N_23187);
or U23832 (N_23832,N_23433,N_23295);
xor U23833 (N_23833,N_23416,N_23304);
and U23834 (N_23834,N_23380,N_23404);
or U23835 (N_23835,N_23452,N_23312);
nor U23836 (N_23836,N_23111,N_23307);
xnor U23837 (N_23837,N_23395,N_23459);
and U23838 (N_23838,N_23290,N_23149);
nor U23839 (N_23839,N_23286,N_23493);
nor U23840 (N_23840,N_23458,N_23054);
nand U23841 (N_23841,N_23375,N_23093);
or U23842 (N_23842,N_23274,N_23106);
xnor U23843 (N_23843,N_23179,N_23056);
nor U23844 (N_23844,N_23102,N_23224);
nor U23845 (N_23845,N_23473,N_23096);
xnor U23846 (N_23846,N_23306,N_23401);
nor U23847 (N_23847,N_23259,N_23314);
nand U23848 (N_23848,N_23089,N_23354);
nor U23849 (N_23849,N_23418,N_23073);
nand U23850 (N_23850,N_23385,N_23362);
or U23851 (N_23851,N_23147,N_23470);
or U23852 (N_23852,N_23424,N_23050);
nand U23853 (N_23853,N_23213,N_23388);
nand U23854 (N_23854,N_23442,N_23373);
or U23855 (N_23855,N_23342,N_23375);
or U23856 (N_23856,N_23284,N_23198);
xor U23857 (N_23857,N_23464,N_23468);
xnor U23858 (N_23858,N_23132,N_23031);
and U23859 (N_23859,N_23421,N_23289);
nand U23860 (N_23860,N_23344,N_23411);
and U23861 (N_23861,N_23179,N_23481);
nor U23862 (N_23862,N_23046,N_23225);
and U23863 (N_23863,N_23405,N_23016);
or U23864 (N_23864,N_23097,N_23335);
nor U23865 (N_23865,N_23262,N_23275);
nand U23866 (N_23866,N_23053,N_23173);
and U23867 (N_23867,N_23225,N_23344);
nand U23868 (N_23868,N_23275,N_23302);
and U23869 (N_23869,N_23497,N_23151);
xnor U23870 (N_23870,N_23078,N_23027);
xor U23871 (N_23871,N_23129,N_23161);
nor U23872 (N_23872,N_23382,N_23288);
and U23873 (N_23873,N_23108,N_23214);
or U23874 (N_23874,N_23412,N_23011);
nor U23875 (N_23875,N_23348,N_23483);
or U23876 (N_23876,N_23096,N_23309);
and U23877 (N_23877,N_23218,N_23294);
nor U23878 (N_23878,N_23354,N_23170);
or U23879 (N_23879,N_23199,N_23133);
xor U23880 (N_23880,N_23056,N_23052);
nand U23881 (N_23881,N_23000,N_23448);
nor U23882 (N_23882,N_23070,N_23252);
nor U23883 (N_23883,N_23315,N_23009);
nand U23884 (N_23884,N_23149,N_23428);
nand U23885 (N_23885,N_23231,N_23244);
xor U23886 (N_23886,N_23108,N_23252);
xnor U23887 (N_23887,N_23167,N_23193);
nand U23888 (N_23888,N_23397,N_23080);
or U23889 (N_23889,N_23412,N_23294);
or U23890 (N_23890,N_23228,N_23387);
xor U23891 (N_23891,N_23158,N_23328);
and U23892 (N_23892,N_23282,N_23221);
nor U23893 (N_23893,N_23068,N_23425);
nor U23894 (N_23894,N_23001,N_23170);
nand U23895 (N_23895,N_23364,N_23191);
xnor U23896 (N_23896,N_23388,N_23125);
or U23897 (N_23897,N_23064,N_23227);
nand U23898 (N_23898,N_23265,N_23444);
xnor U23899 (N_23899,N_23482,N_23479);
xor U23900 (N_23900,N_23487,N_23187);
and U23901 (N_23901,N_23014,N_23444);
or U23902 (N_23902,N_23016,N_23440);
or U23903 (N_23903,N_23221,N_23028);
nand U23904 (N_23904,N_23365,N_23145);
nor U23905 (N_23905,N_23245,N_23481);
and U23906 (N_23906,N_23154,N_23038);
xor U23907 (N_23907,N_23005,N_23360);
and U23908 (N_23908,N_23107,N_23225);
or U23909 (N_23909,N_23057,N_23093);
nor U23910 (N_23910,N_23350,N_23351);
xnor U23911 (N_23911,N_23475,N_23292);
nor U23912 (N_23912,N_23486,N_23058);
nor U23913 (N_23913,N_23432,N_23389);
xor U23914 (N_23914,N_23410,N_23385);
nand U23915 (N_23915,N_23453,N_23356);
or U23916 (N_23916,N_23398,N_23163);
nand U23917 (N_23917,N_23395,N_23280);
and U23918 (N_23918,N_23452,N_23186);
and U23919 (N_23919,N_23296,N_23021);
xor U23920 (N_23920,N_23067,N_23045);
or U23921 (N_23921,N_23205,N_23215);
nor U23922 (N_23922,N_23450,N_23045);
nand U23923 (N_23923,N_23006,N_23477);
nand U23924 (N_23924,N_23488,N_23407);
xor U23925 (N_23925,N_23354,N_23133);
or U23926 (N_23926,N_23411,N_23207);
or U23927 (N_23927,N_23075,N_23468);
nand U23928 (N_23928,N_23251,N_23116);
or U23929 (N_23929,N_23041,N_23437);
nor U23930 (N_23930,N_23017,N_23427);
nor U23931 (N_23931,N_23041,N_23471);
nand U23932 (N_23932,N_23449,N_23010);
and U23933 (N_23933,N_23304,N_23183);
or U23934 (N_23934,N_23118,N_23112);
or U23935 (N_23935,N_23355,N_23499);
xor U23936 (N_23936,N_23293,N_23155);
nand U23937 (N_23937,N_23355,N_23425);
nand U23938 (N_23938,N_23149,N_23044);
and U23939 (N_23939,N_23198,N_23050);
nand U23940 (N_23940,N_23121,N_23439);
nand U23941 (N_23941,N_23344,N_23433);
nand U23942 (N_23942,N_23369,N_23471);
xnor U23943 (N_23943,N_23206,N_23182);
nand U23944 (N_23944,N_23458,N_23261);
nand U23945 (N_23945,N_23079,N_23065);
nor U23946 (N_23946,N_23417,N_23000);
and U23947 (N_23947,N_23407,N_23214);
nor U23948 (N_23948,N_23194,N_23319);
or U23949 (N_23949,N_23464,N_23085);
or U23950 (N_23950,N_23389,N_23092);
and U23951 (N_23951,N_23006,N_23005);
nor U23952 (N_23952,N_23019,N_23029);
and U23953 (N_23953,N_23454,N_23091);
or U23954 (N_23954,N_23008,N_23420);
nor U23955 (N_23955,N_23424,N_23221);
nor U23956 (N_23956,N_23366,N_23280);
nand U23957 (N_23957,N_23043,N_23205);
xnor U23958 (N_23958,N_23067,N_23030);
xor U23959 (N_23959,N_23421,N_23056);
nand U23960 (N_23960,N_23260,N_23435);
nand U23961 (N_23961,N_23270,N_23220);
xor U23962 (N_23962,N_23011,N_23397);
or U23963 (N_23963,N_23461,N_23310);
nor U23964 (N_23964,N_23139,N_23082);
or U23965 (N_23965,N_23046,N_23008);
or U23966 (N_23966,N_23111,N_23472);
nor U23967 (N_23967,N_23041,N_23266);
nand U23968 (N_23968,N_23344,N_23446);
xor U23969 (N_23969,N_23241,N_23329);
and U23970 (N_23970,N_23372,N_23470);
and U23971 (N_23971,N_23367,N_23478);
nand U23972 (N_23972,N_23029,N_23014);
nor U23973 (N_23973,N_23280,N_23451);
nand U23974 (N_23974,N_23336,N_23075);
or U23975 (N_23975,N_23182,N_23308);
xor U23976 (N_23976,N_23311,N_23187);
and U23977 (N_23977,N_23313,N_23458);
nor U23978 (N_23978,N_23224,N_23304);
and U23979 (N_23979,N_23460,N_23413);
and U23980 (N_23980,N_23402,N_23261);
nor U23981 (N_23981,N_23399,N_23249);
nand U23982 (N_23982,N_23351,N_23062);
and U23983 (N_23983,N_23373,N_23412);
xor U23984 (N_23984,N_23094,N_23314);
xnor U23985 (N_23985,N_23234,N_23411);
and U23986 (N_23986,N_23025,N_23245);
nor U23987 (N_23987,N_23107,N_23397);
xor U23988 (N_23988,N_23222,N_23142);
and U23989 (N_23989,N_23186,N_23053);
and U23990 (N_23990,N_23388,N_23481);
nand U23991 (N_23991,N_23490,N_23446);
or U23992 (N_23992,N_23278,N_23096);
or U23993 (N_23993,N_23408,N_23028);
nor U23994 (N_23994,N_23213,N_23214);
nand U23995 (N_23995,N_23032,N_23252);
and U23996 (N_23996,N_23436,N_23191);
or U23997 (N_23997,N_23149,N_23000);
xnor U23998 (N_23998,N_23421,N_23395);
xnor U23999 (N_23999,N_23346,N_23491);
nor U24000 (N_24000,N_23711,N_23657);
and U24001 (N_24001,N_23887,N_23529);
nand U24002 (N_24002,N_23930,N_23628);
or U24003 (N_24003,N_23883,N_23703);
xnor U24004 (N_24004,N_23666,N_23846);
xor U24005 (N_24005,N_23557,N_23639);
nand U24006 (N_24006,N_23689,N_23881);
and U24007 (N_24007,N_23756,N_23927);
nand U24008 (N_24008,N_23630,N_23848);
xor U24009 (N_24009,N_23692,N_23794);
or U24010 (N_24010,N_23698,N_23747);
nor U24011 (N_24011,N_23514,N_23580);
nor U24012 (N_24012,N_23560,N_23549);
and U24013 (N_24013,N_23578,N_23901);
nor U24014 (N_24014,N_23530,N_23502);
xor U24015 (N_24015,N_23825,N_23800);
and U24016 (N_24016,N_23873,N_23551);
nor U24017 (N_24017,N_23660,N_23590);
nor U24018 (N_24018,N_23500,N_23627);
or U24019 (N_24019,N_23774,N_23798);
nand U24020 (N_24020,N_23909,N_23712);
nor U24021 (N_24021,N_23928,N_23793);
nor U24022 (N_24022,N_23884,N_23776);
nand U24023 (N_24023,N_23737,N_23979);
xnor U24024 (N_24024,N_23576,N_23746);
nand U24025 (N_24025,N_23690,N_23541);
nor U24026 (N_24026,N_23618,N_23650);
nor U24027 (N_24027,N_23841,N_23987);
nand U24028 (N_24028,N_23516,N_23852);
and U24029 (N_24029,N_23603,N_23519);
nand U24030 (N_24030,N_23687,N_23625);
or U24031 (N_24031,N_23587,N_23545);
or U24032 (N_24032,N_23658,N_23681);
nand U24033 (N_24033,N_23527,N_23934);
or U24034 (N_24034,N_23907,N_23862);
and U24035 (N_24035,N_23685,N_23836);
and U24036 (N_24036,N_23732,N_23568);
or U24037 (N_24037,N_23693,N_23786);
nand U24038 (N_24038,N_23614,N_23569);
xor U24039 (N_24039,N_23608,N_23989);
nor U24040 (N_24040,N_23912,N_23750);
xnor U24041 (N_24041,N_23937,N_23763);
nor U24042 (N_24042,N_23914,N_23634);
nand U24043 (N_24043,N_23577,N_23880);
xor U24044 (N_24044,N_23816,N_23762);
and U24045 (N_24045,N_23758,N_23949);
and U24046 (N_24046,N_23531,N_23840);
and U24047 (N_24047,N_23645,N_23702);
xor U24048 (N_24048,N_23931,N_23809);
nand U24049 (N_24049,N_23697,N_23775);
xor U24050 (N_24050,N_23575,N_23801);
xor U24051 (N_24051,N_23503,N_23612);
nor U24052 (N_24052,N_23954,N_23688);
nor U24053 (N_24053,N_23957,N_23643);
and U24054 (N_24054,N_23594,N_23921);
nand U24055 (N_24055,N_23923,N_23865);
nor U24056 (N_24056,N_23749,N_23992);
or U24057 (N_24057,N_23651,N_23906);
and U24058 (N_24058,N_23559,N_23673);
or U24059 (N_24059,N_23581,N_23790);
or U24060 (N_24060,N_23999,N_23609);
xnor U24061 (N_24061,N_23891,N_23785);
and U24062 (N_24062,N_23769,N_23695);
nand U24063 (N_24063,N_23879,N_23829);
or U24064 (N_24064,N_23858,N_23871);
nand U24065 (N_24065,N_23694,N_23726);
nor U24066 (N_24066,N_23772,N_23561);
nor U24067 (N_24067,N_23853,N_23538);
and U24068 (N_24068,N_23970,N_23742);
nand U24069 (N_24069,N_23622,N_23550);
nor U24070 (N_24070,N_23504,N_23908);
nor U24071 (N_24071,N_23547,N_23570);
and U24072 (N_24072,N_23913,N_23704);
or U24073 (N_24073,N_23669,N_23574);
xnor U24074 (N_24074,N_23579,N_23866);
nand U24075 (N_24075,N_23636,N_23566);
nor U24076 (N_24076,N_23599,N_23876);
or U24077 (N_24077,N_23562,N_23915);
nand U24078 (N_24078,N_23696,N_23926);
and U24079 (N_24079,N_23882,N_23683);
nand U24080 (N_24080,N_23617,N_23986);
nor U24081 (N_24081,N_23997,N_23713);
nand U24082 (N_24082,N_23827,N_23739);
and U24083 (N_24083,N_23918,N_23546);
and U24084 (N_24084,N_23822,N_23721);
nand U24085 (N_24085,N_23782,N_23616);
nand U24086 (N_24086,N_23610,N_23832);
and U24087 (N_24087,N_23679,N_23585);
nor U24088 (N_24088,N_23571,N_23735);
nand U24089 (N_24089,N_23602,N_23837);
nor U24090 (N_24090,N_23637,N_23802);
nor U24091 (N_24091,N_23935,N_23864);
nor U24092 (N_24092,N_23933,N_23626);
or U24093 (N_24093,N_23905,N_23761);
or U24094 (N_24094,N_23552,N_23813);
nor U24095 (N_24095,N_23572,N_23936);
xnor U24096 (N_24096,N_23993,N_23856);
xor U24097 (N_24097,N_23854,N_23861);
nor U24098 (N_24098,N_23642,N_23819);
xnor U24099 (N_24099,N_23640,N_23944);
nor U24100 (N_24100,N_23648,N_23564);
nand U24101 (N_24101,N_23520,N_23605);
or U24102 (N_24102,N_23661,N_23952);
xor U24103 (N_24103,N_23667,N_23535);
nand U24104 (N_24104,N_23733,N_23788);
nor U24105 (N_24105,N_23615,N_23902);
xor U24106 (N_24106,N_23613,N_23893);
xor U24107 (N_24107,N_23972,N_23973);
nand U24108 (N_24108,N_23911,N_23528);
nand U24109 (N_24109,N_23730,N_23606);
or U24110 (N_24110,N_23515,N_23674);
and U24111 (N_24111,N_23592,N_23682);
nand U24112 (N_24112,N_23596,N_23565);
nand U24113 (N_24113,N_23998,N_23611);
nand U24114 (N_24114,N_23960,N_23863);
and U24115 (N_24115,N_23939,N_23718);
nor U24116 (N_24116,N_23595,N_23719);
xnor U24117 (N_24117,N_23878,N_23525);
nor U24118 (N_24118,N_23983,N_23760);
xor U24119 (N_24119,N_23966,N_23795);
or U24120 (N_24120,N_23767,N_23765);
xnor U24121 (N_24121,N_23728,N_23955);
nor U24122 (N_24122,N_23924,N_23818);
nand U24123 (N_24123,N_23898,N_23787);
and U24124 (N_24124,N_23991,N_23723);
or U24125 (N_24125,N_23875,N_23620);
nand U24126 (N_24126,N_23870,N_23812);
or U24127 (N_24127,N_23722,N_23641);
nand U24128 (N_24128,N_23833,N_23994);
or U24129 (N_24129,N_23623,N_23544);
and U24130 (N_24130,N_23830,N_23505);
or U24131 (N_24131,N_23962,N_23981);
xnor U24132 (N_24132,N_23976,N_23586);
or U24133 (N_24133,N_23951,N_23647);
nand U24134 (N_24134,N_23676,N_23900);
xor U24135 (N_24135,N_23821,N_23633);
nor U24136 (N_24136,N_23707,N_23895);
or U24137 (N_24137,N_23654,N_23517);
nor U24138 (N_24138,N_23542,N_23532);
nor U24139 (N_24139,N_23563,N_23662);
xnor U24140 (N_24140,N_23932,N_23946);
nor U24141 (N_24141,N_23539,N_23664);
xor U24142 (N_24142,N_23850,N_23554);
xor U24143 (N_24143,N_23867,N_23600);
or U24144 (N_24144,N_23675,N_23736);
xnor U24145 (N_24145,N_23963,N_23584);
xnor U24146 (N_24146,N_23709,N_23598);
nor U24147 (N_24147,N_23556,N_23548);
and U24148 (N_24148,N_23656,N_23834);
and U24149 (N_24149,N_23740,N_23555);
and U24150 (N_24150,N_23894,N_23512);
nand U24151 (N_24151,N_23537,N_23824);
nand U24152 (N_24152,N_23948,N_23806);
nor U24153 (N_24153,N_23965,N_23638);
xor U24154 (N_24154,N_23872,N_23971);
nor U24155 (N_24155,N_23859,N_23671);
and U24156 (N_24156,N_23567,N_23810);
nand U24157 (N_24157,N_23714,N_23844);
and U24158 (N_24158,N_23885,N_23984);
and U24159 (N_24159,N_23588,N_23757);
or U24160 (N_24160,N_23773,N_23734);
nor U24161 (N_24161,N_23591,N_23518);
nor U24162 (N_24162,N_23593,N_23890);
xnor U24163 (N_24163,N_23899,N_23843);
nor U24164 (N_24164,N_23791,N_23803);
and U24165 (N_24165,N_23978,N_23526);
xnor U24166 (N_24166,N_23838,N_23956);
or U24167 (N_24167,N_23950,N_23943);
nor U24168 (N_24168,N_23982,N_23701);
nand U24169 (N_24169,N_23699,N_23583);
nor U24170 (N_24170,N_23513,N_23748);
nor U24171 (N_24171,N_23521,N_23892);
nor U24172 (N_24172,N_23534,N_23869);
or U24173 (N_24173,N_23835,N_23938);
nor U24174 (N_24174,N_23889,N_23753);
or U24175 (N_24175,N_23644,N_23509);
or U24176 (N_24176,N_23919,N_23621);
and U24177 (N_24177,N_23959,N_23705);
xor U24178 (N_24178,N_23977,N_23823);
xor U24179 (N_24179,N_23652,N_23635);
nand U24180 (N_24180,N_23817,N_23573);
nor U24181 (N_24181,N_23783,N_23868);
xnor U24182 (N_24182,N_23855,N_23764);
xor U24183 (N_24183,N_23796,N_23508);
or U24184 (N_24184,N_23745,N_23511);
or U24185 (N_24185,N_23670,N_23896);
or U24186 (N_24186,N_23738,N_23731);
xor U24187 (N_24187,N_23780,N_23710);
and U24188 (N_24188,N_23826,N_23706);
xnor U24189 (N_24189,N_23789,N_23649);
nor U24190 (N_24190,N_23831,N_23589);
xor U24191 (N_24191,N_23888,N_23533);
nor U24192 (N_24192,N_23877,N_23631);
nor U24193 (N_24193,N_23624,N_23607);
xnor U24194 (N_24194,N_23849,N_23799);
and U24195 (N_24195,N_23604,N_23672);
xor U24196 (N_24196,N_23536,N_23668);
nand U24197 (N_24197,N_23792,N_23820);
xnor U24198 (N_24198,N_23700,N_23808);
xnor U24199 (N_24199,N_23543,N_23540);
nor U24200 (N_24200,N_23916,N_23842);
nor U24201 (N_24201,N_23632,N_23845);
or U24202 (N_24202,N_23629,N_23797);
and U24203 (N_24203,N_23969,N_23715);
or U24204 (N_24204,N_23727,N_23751);
nand U24205 (N_24205,N_23655,N_23851);
or U24206 (N_24206,N_23910,N_23558);
nand U24207 (N_24207,N_23807,N_23729);
nor U24208 (N_24208,N_23759,N_23886);
nor U24209 (N_24209,N_23925,N_23523);
and U24210 (N_24210,N_23874,N_23975);
nand U24211 (N_24211,N_23968,N_23922);
nand U24212 (N_24212,N_23725,N_23619);
or U24213 (N_24213,N_23678,N_23684);
nand U24214 (N_24214,N_23501,N_23720);
or U24215 (N_24215,N_23929,N_23805);
nor U24216 (N_24216,N_23777,N_23961);
nor U24217 (N_24217,N_23964,N_23917);
nand U24218 (N_24218,N_23847,N_23768);
and U24219 (N_24219,N_23724,N_23814);
nand U24220 (N_24220,N_23897,N_23743);
xnor U24221 (N_24221,N_23990,N_23940);
xor U24222 (N_24222,N_23665,N_23781);
xnor U24223 (N_24223,N_23980,N_23646);
and U24224 (N_24224,N_23766,N_23686);
or U24225 (N_24225,N_23680,N_23659);
or U24226 (N_24226,N_23967,N_23953);
nand U24227 (N_24227,N_23677,N_23510);
or U24228 (N_24228,N_23708,N_23601);
and U24229 (N_24229,N_23815,N_23996);
or U24230 (N_24230,N_23904,N_23974);
nor U24231 (N_24231,N_23811,N_23507);
nor U24232 (N_24232,N_23958,N_23754);
nand U24233 (N_24233,N_23522,N_23828);
or U24234 (N_24234,N_23985,N_23771);
nor U24235 (N_24235,N_23597,N_23663);
nor U24236 (N_24236,N_23716,N_23691);
or U24237 (N_24237,N_23784,N_23779);
and U24238 (N_24238,N_23506,N_23945);
or U24239 (N_24239,N_23717,N_23741);
nand U24240 (N_24240,N_23903,N_23770);
nand U24241 (N_24241,N_23995,N_23804);
nand U24242 (N_24242,N_23582,N_23755);
nor U24243 (N_24243,N_23920,N_23744);
xor U24244 (N_24244,N_23947,N_23553);
xnor U24245 (N_24245,N_23778,N_23941);
xor U24246 (N_24246,N_23857,N_23524);
nand U24247 (N_24247,N_23988,N_23860);
nand U24248 (N_24248,N_23942,N_23653);
nor U24249 (N_24249,N_23752,N_23839);
or U24250 (N_24250,N_23677,N_23717);
xor U24251 (N_24251,N_23635,N_23750);
or U24252 (N_24252,N_23968,N_23674);
or U24253 (N_24253,N_23994,N_23738);
nor U24254 (N_24254,N_23697,N_23611);
nor U24255 (N_24255,N_23816,N_23653);
xor U24256 (N_24256,N_23998,N_23829);
nor U24257 (N_24257,N_23949,N_23579);
and U24258 (N_24258,N_23794,N_23674);
xnor U24259 (N_24259,N_23703,N_23501);
xnor U24260 (N_24260,N_23739,N_23702);
nor U24261 (N_24261,N_23981,N_23832);
and U24262 (N_24262,N_23775,N_23823);
nand U24263 (N_24263,N_23533,N_23703);
or U24264 (N_24264,N_23707,N_23810);
and U24265 (N_24265,N_23901,N_23758);
nor U24266 (N_24266,N_23573,N_23860);
or U24267 (N_24267,N_23843,N_23921);
and U24268 (N_24268,N_23923,N_23976);
and U24269 (N_24269,N_23845,N_23685);
xor U24270 (N_24270,N_23939,N_23826);
and U24271 (N_24271,N_23582,N_23809);
nor U24272 (N_24272,N_23663,N_23754);
nor U24273 (N_24273,N_23823,N_23703);
or U24274 (N_24274,N_23771,N_23588);
xor U24275 (N_24275,N_23769,N_23964);
xor U24276 (N_24276,N_23621,N_23916);
or U24277 (N_24277,N_23509,N_23859);
xor U24278 (N_24278,N_23846,N_23797);
or U24279 (N_24279,N_23566,N_23544);
nor U24280 (N_24280,N_23895,N_23715);
nor U24281 (N_24281,N_23807,N_23816);
and U24282 (N_24282,N_23539,N_23653);
and U24283 (N_24283,N_23559,N_23612);
and U24284 (N_24284,N_23688,N_23873);
or U24285 (N_24285,N_23924,N_23757);
xnor U24286 (N_24286,N_23617,N_23967);
and U24287 (N_24287,N_23902,N_23896);
nand U24288 (N_24288,N_23610,N_23895);
xor U24289 (N_24289,N_23734,N_23560);
nor U24290 (N_24290,N_23666,N_23684);
or U24291 (N_24291,N_23784,N_23814);
xor U24292 (N_24292,N_23578,N_23596);
and U24293 (N_24293,N_23502,N_23738);
and U24294 (N_24294,N_23922,N_23770);
or U24295 (N_24295,N_23838,N_23793);
and U24296 (N_24296,N_23605,N_23959);
nor U24297 (N_24297,N_23997,N_23917);
or U24298 (N_24298,N_23714,N_23696);
nand U24299 (N_24299,N_23678,N_23685);
nand U24300 (N_24300,N_23907,N_23744);
and U24301 (N_24301,N_23554,N_23867);
nand U24302 (N_24302,N_23765,N_23801);
nor U24303 (N_24303,N_23652,N_23993);
nand U24304 (N_24304,N_23924,N_23583);
nor U24305 (N_24305,N_23580,N_23610);
or U24306 (N_24306,N_23991,N_23568);
nand U24307 (N_24307,N_23988,N_23972);
nor U24308 (N_24308,N_23843,N_23761);
nand U24309 (N_24309,N_23526,N_23804);
and U24310 (N_24310,N_23772,N_23942);
nand U24311 (N_24311,N_23683,N_23781);
xnor U24312 (N_24312,N_23754,N_23919);
nand U24313 (N_24313,N_23656,N_23641);
nor U24314 (N_24314,N_23594,N_23814);
xor U24315 (N_24315,N_23687,N_23551);
and U24316 (N_24316,N_23576,N_23971);
nor U24317 (N_24317,N_23694,N_23922);
nand U24318 (N_24318,N_23577,N_23907);
and U24319 (N_24319,N_23881,N_23673);
and U24320 (N_24320,N_23937,N_23782);
or U24321 (N_24321,N_23587,N_23537);
nor U24322 (N_24322,N_23649,N_23695);
and U24323 (N_24323,N_23991,N_23572);
xor U24324 (N_24324,N_23835,N_23676);
xnor U24325 (N_24325,N_23704,N_23699);
and U24326 (N_24326,N_23636,N_23857);
xor U24327 (N_24327,N_23729,N_23967);
and U24328 (N_24328,N_23917,N_23815);
nand U24329 (N_24329,N_23642,N_23887);
and U24330 (N_24330,N_23922,N_23816);
nor U24331 (N_24331,N_23637,N_23894);
nand U24332 (N_24332,N_23964,N_23825);
xnor U24333 (N_24333,N_23685,N_23764);
xor U24334 (N_24334,N_23944,N_23556);
and U24335 (N_24335,N_23744,N_23592);
xnor U24336 (N_24336,N_23768,N_23960);
nor U24337 (N_24337,N_23980,N_23773);
nor U24338 (N_24338,N_23616,N_23747);
nand U24339 (N_24339,N_23550,N_23879);
or U24340 (N_24340,N_23995,N_23689);
or U24341 (N_24341,N_23695,N_23617);
xnor U24342 (N_24342,N_23757,N_23585);
or U24343 (N_24343,N_23801,N_23996);
or U24344 (N_24344,N_23972,N_23551);
xor U24345 (N_24345,N_23794,N_23736);
and U24346 (N_24346,N_23876,N_23665);
xnor U24347 (N_24347,N_23842,N_23616);
nor U24348 (N_24348,N_23513,N_23699);
nor U24349 (N_24349,N_23963,N_23848);
xnor U24350 (N_24350,N_23885,N_23803);
nand U24351 (N_24351,N_23721,N_23934);
and U24352 (N_24352,N_23800,N_23827);
xor U24353 (N_24353,N_23991,N_23807);
xnor U24354 (N_24354,N_23881,N_23872);
or U24355 (N_24355,N_23741,N_23829);
and U24356 (N_24356,N_23893,N_23652);
or U24357 (N_24357,N_23840,N_23640);
nand U24358 (N_24358,N_23683,N_23858);
nand U24359 (N_24359,N_23847,N_23940);
and U24360 (N_24360,N_23737,N_23892);
nand U24361 (N_24361,N_23743,N_23946);
nand U24362 (N_24362,N_23881,N_23888);
and U24363 (N_24363,N_23646,N_23806);
and U24364 (N_24364,N_23728,N_23794);
nor U24365 (N_24365,N_23619,N_23922);
nor U24366 (N_24366,N_23774,N_23884);
or U24367 (N_24367,N_23960,N_23586);
and U24368 (N_24368,N_23506,N_23984);
or U24369 (N_24369,N_23697,N_23744);
nand U24370 (N_24370,N_23897,N_23980);
xnor U24371 (N_24371,N_23533,N_23977);
nor U24372 (N_24372,N_23715,N_23728);
and U24373 (N_24373,N_23786,N_23623);
nand U24374 (N_24374,N_23551,N_23527);
nor U24375 (N_24375,N_23510,N_23708);
xnor U24376 (N_24376,N_23857,N_23837);
xor U24377 (N_24377,N_23533,N_23989);
nor U24378 (N_24378,N_23738,N_23566);
xnor U24379 (N_24379,N_23853,N_23658);
nor U24380 (N_24380,N_23511,N_23851);
xor U24381 (N_24381,N_23895,N_23802);
nand U24382 (N_24382,N_23685,N_23642);
nor U24383 (N_24383,N_23544,N_23556);
nor U24384 (N_24384,N_23560,N_23987);
and U24385 (N_24385,N_23879,N_23815);
and U24386 (N_24386,N_23692,N_23748);
nand U24387 (N_24387,N_23650,N_23703);
and U24388 (N_24388,N_23893,N_23712);
and U24389 (N_24389,N_23981,N_23525);
xor U24390 (N_24390,N_23649,N_23612);
and U24391 (N_24391,N_23868,N_23724);
or U24392 (N_24392,N_23739,N_23758);
nor U24393 (N_24393,N_23870,N_23582);
or U24394 (N_24394,N_23957,N_23525);
nand U24395 (N_24395,N_23862,N_23998);
and U24396 (N_24396,N_23609,N_23758);
and U24397 (N_24397,N_23559,N_23615);
and U24398 (N_24398,N_23924,N_23518);
xor U24399 (N_24399,N_23892,N_23884);
and U24400 (N_24400,N_23673,N_23546);
nand U24401 (N_24401,N_23767,N_23956);
or U24402 (N_24402,N_23651,N_23964);
nand U24403 (N_24403,N_23500,N_23940);
xor U24404 (N_24404,N_23568,N_23847);
or U24405 (N_24405,N_23867,N_23710);
xnor U24406 (N_24406,N_23638,N_23784);
xnor U24407 (N_24407,N_23644,N_23941);
or U24408 (N_24408,N_23727,N_23602);
xnor U24409 (N_24409,N_23761,N_23940);
nand U24410 (N_24410,N_23703,N_23985);
xnor U24411 (N_24411,N_23885,N_23591);
or U24412 (N_24412,N_23683,N_23997);
or U24413 (N_24413,N_23864,N_23658);
nor U24414 (N_24414,N_23965,N_23760);
xnor U24415 (N_24415,N_23648,N_23647);
or U24416 (N_24416,N_23711,N_23780);
or U24417 (N_24417,N_23608,N_23595);
nand U24418 (N_24418,N_23742,N_23886);
nor U24419 (N_24419,N_23868,N_23810);
and U24420 (N_24420,N_23773,N_23675);
xnor U24421 (N_24421,N_23848,N_23577);
nor U24422 (N_24422,N_23614,N_23670);
xnor U24423 (N_24423,N_23947,N_23777);
nand U24424 (N_24424,N_23799,N_23730);
nand U24425 (N_24425,N_23925,N_23728);
nor U24426 (N_24426,N_23708,N_23646);
xnor U24427 (N_24427,N_23763,N_23658);
and U24428 (N_24428,N_23538,N_23838);
xnor U24429 (N_24429,N_23940,N_23742);
or U24430 (N_24430,N_23885,N_23764);
or U24431 (N_24431,N_23761,N_23747);
nor U24432 (N_24432,N_23583,N_23835);
nand U24433 (N_24433,N_23738,N_23670);
nand U24434 (N_24434,N_23645,N_23954);
nand U24435 (N_24435,N_23977,N_23701);
nor U24436 (N_24436,N_23889,N_23816);
or U24437 (N_24437,N_23976,N_23963);
or U24438 (N_24438,N_23899,N_23583);
nor U24439 (N_24439,N_23555,N_23534);
xnor U24440 (N_24440,N_23510,N_23719);
nor U24441 (N_24441,N_23886,N_23641);
nand U24442 (N_24442,N_23678,N_23875);
or U24443 (N_24443,N_23733,N_23883);
or U24444 (N_24444,N_23602,N_23822);
nand U24445 (N_24445,N_23910,N_23702);
or U24446 (N_24446,N_23758,N_23564);
or U24447 (N_24447,N_23936,N_23584);
or U24448 (N_24448,N_23685,N_23548);
nor U24449 (N_24449,N_23635,N_23840);
and U24450 (N_24450,N_23669,N_23743);
nand U24451 (N_24451,N_23642,N_23641);
or U24452 (N_24452,N_23621,N_23559);
and U24453 (N_24453,N_23697,N_23752);
nor U24454 (N_24454,N_23850,N_23839);
xnor U24455 (N_24455,N_23874,N_23554);
and U24456 (N_24456,N_23764,N_23597);
or U24457 (N_24457,N_23738,N_23830);
xnor U24458 (N_24458,N_23934,N_23935);
xor U24459 (N_24459,N_23578,N_23860);
and U24460 (N_24460,N_23964,N_23856);
nor U24461 (N_24461,N_23713,N_23842);
xnor U24462 (N_24462,N_23727,N_23806);
or U24463 (N_24463,N_23581,N_23833);
nor U24464 (N_24464,N_23674,N_23983);
or U24465 (N_24465,N_23806,N_23599);
xnor U24466 (N_24466,N_23986,N_23509);
nor U24467 (N_24467,N_23969,N_23601);
or U24468 (N_24468,N_23819,N_23666);
xnor U24469 (N_24469,N_23815,N_23636);
nor U24470 (N_24470,N_23888,N_23767);
and U24471 (N_24471,N_23680,N_23619);
and U24472 (N_24472,N_23945,N_23574);
nor U24473 (N_24473,N_23633,N_23973);
and U24474 (N_24474,N_23588,N_23863);
and U24475 (N_24475,N_23581,N_23820);
or U24476 (N_24476,N_23752,N_23920);
nor U24477 (N_24477,N_23517,N_23897);
nor U24478 (N_24478,N_23731,N_23764);
nand U24479 (N_24479,N_23926,N_23720);
xnor U24480 (N_24480,N_23627,N_23900);
xnor U24481 (N_24481,N_23562,N_23748);
and U24482 (N_24482,N_23554,N_23717);
or U24483 (N_24483,N_23739,N_23820);
nor U24484 (N_24484,N_23804,N_23646);
or U24485 (N_24485,N_23965,N_23822);
or U24486 (N_24486,N_23693,N_23618);
nand U24487 (N_24487,N_23547,N_23835);
nand U24488 (N_24488,N_23541,N_23808);
and U24489 (N_24489,N_23535,N_23529);
nor U24490 (N_24490,N_23713,N_23728);
or U24491 (N_24491,N_23629,N_23613);
and U24492 (N_24492,N_23790,N_23948);
or U24493 (N_24493,N_23697,N_23966);
xor U24494 (N_24494,N_23727,N_23697);
nor U24495 (N_24495,N_23964,N_23894);
xor U24496 (N_24496,N_23825,N_23615);
xnor U24497 (N_24497,N_23772,N_23963);
or U24498 (N_24498,N_23504,N_23796);
nor U24499 (N_24499,N_23980,N_23644);
or U24500 (N_24500,N_24309,N_24198);
xor U24501 (N_24501,N_24450,N_24386);
nand U24502 (N_24502,N_24275,N_24432);
nand U24503 (N_24503,N_24026,N_24126);
nor U24504 (N_24504,N_24497,N_24188);
or U24505 (N_24505,N_24042,N_24241);
and U24506 (N_24506,N_24059,N_24127);
nor U24507 (N_24507,N_24474,N_24005);
xnor U24508 (N_24508,N_24023,N_24212);
and U24509 (N_24509,N_24134,N_24380);
or U24510 (N_24510,N_24123,N_24251);
nand U24511 (N_24511,N_24051,N_24219);
and U24512 (N_24512,N_24192,N_24265);
xor U24513 (N_24513,N_24046,N_24053);
xor U24514 (N_24514,N_24366,N_24151);
or U24515 (N_24515,N_24112,N_24461);
or U24516 (N_24516,N_24224,N_24490);
and U24517 (N_24517,N_24245,N_24458);
or U24518 (N_24518,N_24365,N_24261);
nand U24519 (N_24519,N_24253,N_24434);
xnor U24520 (N_24520,N_24471,N_24300);
xnor U24521 (N_24521,N_24164,N_24273);
or U24522 (N_24522,N_24246,N_24489);
xnor U24523 (N_24523,N_24463,N_24286);
nor U24524 (N_24524,N_24327,N_24371);
or U24525 (N_24525,N_24495,N_24338);
nand U24526 (N_24526,N_24021,N_24311);
xor U24527 (N_24527,N_24289,N_24211);
and U24528 (N_24528,N_24141,N_24284);
nand U24529 (N_24529,N_24230,N_24235);
and U24530 (N_24530,N_24105,N_24295);
or U24531 (N_24531,N_24416,N_24177);
or U24532 (N_24532,N_24499,N_24285);
nor U24533 (N_24533,N_24006,N_24031);
or U24534 (N_24534,N_24207,N_24063);
nand U24535 (N_24535,N_24390,N_24299);
nor U24536 (N_24536,N_24190,N_24218);
nor U24537 (N_24537,N_24444,N_24435);
nor U24538 (N_24538,N_24479,N_24247);
nand U24539 (N_24539,N_24248,N_24131);
xnor U24540 (N_24540,N_24167,N_24076);
xor U24541 (N_24541,N_24028,N_24341);
xnor U24542 (N_24542,N_24157,N_24339);
and U24543 (N_24543,N_24406,N_24020);
xor U24544 (N_24544,N_24173,N_24152);
or U24545 (N_24545,N_24209,N_24359);
and U24546 (N_24546,N_24159,N_24003);
xor U24547 (N_24547,N_24290,N_24057);
xor U24548 (N_24548,N_24122,N_24364);
nand U24549 (N_24549,N_24140,N_24029);
nand U24550 (N_24550,N_24037,N_24121);
or U24551 (N_24551,N_24018,N_24119);
or U24552 (N_24552,N_24050,N_24475);
and U24553 (N_24553,N_24111,N_24405);
or U24554 (N_24554,N_24217,N_24130);
and U24555 (N_24555,N_24153,N_24070);
xnor U24556 (N_24556,N_24473,N_24162);
and U24557 (N_24557,N_24436,N_24414);
nand U24558 (N_24558,N_24472,N_24387);
and U24559 (N_24559,N_24457,N_24236);
and U24560 (N_24560,N_24370,N_24039);
and U24561 (N_24561,N_24454,N_24013);
and U24562 (N_24562,N_24197,N_24221);
nor U24563 (N_24563,N_24388,N_24120);
or U24564 (N_24564,N_24482,N_24361);
nor U24565 (N_24565,N_24208,N_24225);
nor U24566 (N_24566,N_24049,N_24168);
nor U24567 (N_24567,N_24348,N_24445);
nor U24568 (N_24568,N_24250,N_24079);
and U24569 (N_24569,N_24081,N_24147);
and U24570 (N_24570,N_24194,N_24417);
or U24571 (N_24571,N_24408,N_24086);
or U24572 (N_24572,N_24085,N_24351);
and U24573 (N_24573,N_24316,N_24452);
nand U24574 (N_24574,N_24389,N_24038);
or U24575 (N_24575,N_24484,N_24419);
or U24576 (N_24576,N_24174,N_24082);
and U24577 (N_24577,N_24143,N_24329);
nand U24578 (N_24578,N_24424,N_24137);
and U24579 (N_24579,N_24277,N_24437);
xor U24580 (N_24580,N_24342,N_24220);
nand U24581 (N_24581,N_24106,N_24447);
nor U24582 (N_24582,N_24008,N_24090);
nand U24583 (N_24583,N_24462,N_24396);
or U24584 (N_24584,N_24045,N_24179);
nand U24585 (N_24585,N_24293,N_24056);
nor U24586 (N_24586,N_24492,N_24158);
and U24587 (N_24587,N_24315,N_24401);
nor U24588 (N_24588,N_24460,N_24075);
xnor U24589 (N_24589,N_24421,N_24428);
xor U24590 (N_24590,N_24100,N_24128);
nand U24591 (N_24591,N_24234,N_24430);
and U24592 (N_24592,N_24000,N_24360);
nor U24593 (N_24593,N_24054,N_24047);
and U24594 (N_24594,N_24093,N_24249);
xor U24595 (N_24595,N_24165,N_24302);
and U24596 (N_24596,N_24259,N_24017);
nand U24597 (N_24597,N_24233,N_24080);
nand U24598 (N_24598,N_24097,N_24478);
and U24599 (N_24599,N_24014,N_24203);
nor U24600 (N_24600,N_24335,N_24308);
nor U24601 (N_24601,N_24496,N_24296);
or U24602 (N_24602,N_24071,N_24292);
xnor U24603 (N_24603,N_24160,N_24262);
nor U24604 (N_24604,N_24092,N_24161);
and U24605 (N_24605,N_24375,N_24010);
nor U24606 (N_24606,N_24096,N_24135);
xor U24607 (N_24607,N_24318,N_24349);
or U24608 (N_24608,N_24114,N_24468);
xor U24609 (N_24609,N_24287,N_24266);
xnor U24610 (N_24610,N_24288,N_24303);
and U24611 (N_24611,N_24422,N_24263);
nand U24612 (N_24612,N_24398,N_24024);
nor U24613 (N_24613,N_24324,N_24073);
or U24614 (N_24614,N_24238,N_24078);
xor U24615 (N_24615,N_24015,N_24352);
nand U24616 (N_24616,N_24367,N_24117);
and U24617 (N_24617,N_24493,N_24058);
xor U24618 (N_24618,N_24466,N_24115);
xnor U24619 (N_24619,N_24226,N_24169);
xnor U24620 (N_24620,N_24483,N_24146);
nand U24621 (N_24621,N_24283,N_24439);
nor U24622 (N_24622,N_24354,N_24215);
nand U24623 (N_24623,N_24155,N_24442);
nor U24624 (N_24624,N_24477,N_24260);
or U24625 (N_24625,N_24362,N_24269);
or U24626 (N_24626,N_24423,N_24291);
or U24627 (N_24627,N_24068,N_24016);
nand U24628 (N_24628,N_24425,N_24310);
nand U24629 (N_24629,N_24464,N_24343);
nand U24630 (N_24630,N_24195,N_24229);
nor U24631 (N_24631,N_24069,N_24089);
or U24632 (N_24632,N_24200,N_24313);
or U24633 (N_24633,N_24184,N_24205);
nand U24634 (N_24634,N_24274,N_24084);
nand U24635 (N_24635,N_24353,N_24369);
nor U24636 (N_24636,N_24107,N_24002);
nor U24637 (N_24637,N_24098,N_24007);
xnor U24638 (N_24638,N_24376,N_24124);
nor U24639 (N_24639,N_24171,N_24346);
or U24640 (N_24640,N_24382,N_24465);
nand U24641 (N_24641,N_24334,N_24487);
nor U24642 (N_24642,N_24377,N_24022);
xor U24643 (N_24643,N_24418,N_24032);
xnor U24644 (N_24644,N_24138,N_24358);
and U24645 (N_24645,N_24108,N_24061);
nand U24646 (N_24646,N_24040,N_24228);
or U24647 (N_24647,N_24453,N_24301);
or U24648 (N_24648,N_24297,N_24257);
and U24649 (N_24649,N_24095,N_24488);
xnor U24650 (N_24650,N_24223,N_24103);
nand U24651 (N_24651,N_24149,N_24427);
nand U24652 (N_24652,N_24163,N_24456);
nand U24653 (N_24653,N_24041,N_24252);
or U24654 (N_24654,N_24196,N_24467);
or U24655 (N_24655,N_24116,N_24443);
xnor U24656 (N_24656,N_24144,N_24088);
nand U24657 (N_24657,N_24065,N_24320);
nor U24658 (N_24658,N_24317,N_24044);
nand U24659 (N_24659,N_24214,N_24133);
xor U24660 (N_24660,N_24404,N_24231);
nand U24661 (N_24661,N_24321,N_24438);
nor U24662 (N_24662,N_24270,N_24363);
and U24663 (N_24663,N_24239,N_24411);
nand U24664 (N_24664,N_24048,N_24383);
nand U24665 (N_24665,N_24373,N_24368);
nor U24666 (N_24666,N_24412,N_24305);
nor U24667 (N_24667,N_24176,N_24113);
nand U24668 (N_24668,N_24441,N_24175);
nor U24669 (N_24669,N_24001,N_24172);
and U24670 (N_24670,N_24276,N_24244);
nor U24671 (N_24671,N_24400,N_24227);
nand U24672 (N_24672,N_24307,N_24099);
nor U24673 (N_24673,N_24280,N_24480);
and U24674 (N_24674,N_24268,N_24344);
nand U24675 (N_24675,N_24136,N_24110);
xor U24676 (N_24676,N_24181,N_24298);
and U24677 (N_24677,N_24381,N_24402);
nor U24678 (N_24678,N_24395,N_24199);
nand U24679 (N_24679,N_24148,N_24333);
and U24680 (N_24680,N_24448,N_24429);
xnor U24681 (N_24681,N_24204,N_24118);
xnor U24682 (N_24682,N_24420,N_24470);
and U24683 (N_24683,N_24030,N_24271);
or U24684 (N_24684,N_24072,N_24446);
nor U24685 (N_24685,N_24356,N_24403);
nor U24686 (N_24686,N_24355,N_24449);
or U24687 (N_24687,N_24415,N_24350);
xnor U24688 (N_24688,N_24347,N_24399);
nor U24689 (N_24689,N_24319,N_24440);
xor U24690 (N_24690,N_24469,N_24009);
xor U24691 (N_24691,N_24393,N_24156);
or U24692 (N_24692,N_24378,N_24272);
and U24693 (N_24693,N_24256,N_24187);
or U24694 (N_24694,N_24459,N_24232);
nand U24695 (N_24695,N_24237,N_24064);
and U24696 (N_24696,N_24498,N_24258);
or U24697 (N_24697,N_24222,N_24332);
nor U24698 (N_24698,N_24340,N_24264);
and U24699 (N_24699,N_24189,N_24035);
and U24700 (N_24700,N_24240,N_24043);
xnor U24701 (N_24701,N_24306,N_24036);
nand U24702 (N_24702,N_24077,N_24102);
or U24703 (N_24703,N_24004,N_24142);
xnor U24704 (N_24704,N_24433,N_24379);
and U24705 (N_24705,N_24336,N_24314);
nor U24706 (N_24706,N_24060,N_24201);
xor U24707 (N_24707,N_24410,N_24034);
nand U24708 (N_24708,N_24426,N_24385);
xnor U24709 (N_24709,N_24182,N_24087);
nor U24710 (N_24710,N_24392,N_24325);
nor U24711 (N_24711,N_24074,N_24322);
xnor U24712 (N_24712,N_24331,N_24067);
or U24713 (N_24713,N_24357,N_24094);
and U24714 (N_24714,N_24323,N_24154);
nand U24715 (N_24715,N_24372,N_24374);
nand U24716 (N_24716,N_24213,N_24278);
nand U24717 (N_24717,N_24312,N_24407);
xnor U24718 (N_24718,N_24191,N_24185);
and U24719 (N_24719,N_24413,N_24485);
nand U24720 (N_24720,N_24019,N_24281);
and U24721 (N_24721,N_24206,N_24326);
nor U24722 (N_24722,N_24170,N_24255);
nor U24723 (N_24723,N_24337,N_24052);
nand U24724 (N_24724,N_24062,N_24025);
nand U24725 (N_24725,N_24125,N_24216);
and U24726 (N_24726,N_24166,N_24104);
or U24727 (N_24727,N_24476,N_24101);
and U24728 (N_24728,N_24294,N_24012);
and U24729 (N_24729,N_24486,N_24397);
xor U24730 (N_24730,N_24145,N_24083);
nand U24731 (N_24731,N_24384,N_24186);
xnor U24732 (N_24732,N_24451,N_24494);
or U24733 (N_24733,N_24394,N_24491);
nor U24734 (N_24734,N_24243,N_24033);
nand U24735 (N_24735,N_24027,N_24254);
xnor U24736 (N_24736,N_24202,N_24193);
xnor U24737 (N_24737,N_24279,N_24066);
nor U24738 (N_24738,N_24242,N_24267);
and U24739 (N_24739,N_24431,N_24091);
and U24740 (N_24740,N_24304,N_24129);
nand U24741 (N_24741,N_24345,N_24139);
nand U24742 (N_24742,N_24330,N_24282);
and U24743 (N_24743,N_24178,N_24328);
xor U24744 (N_24744,N_24055,N_24109);
nand U24745 (N_24745,N_24481,N_24183);
nand U24746 (N_24746,N_24132,N_24210);
xnor U24747 (N_24747,N_24180,N_24011);
and U24748 (N_24748,N_24409,N_24150);
xnor U24749 (N_24749,N_24391,N_24455);
or U24750 (N_24750,N_24056,N_24385);
and U24751 (N_24751,N_24113,N_24400);
and U24752 (N_24752,N_24396,N_24279);
xor U24753 (N_24753,N_24378,N_24382);
xor U24754 (N_24754,N_24036,N_24149);
xor U24755 (N_24755,N_24457,N_24298);
or U24756 (N_24756,N_24113,N_24301);
nand U24757 (N_24757,N_24280,N_24450);
nor U24758 (N_24758,N_24048,N_24050);
nand U24759 (N_24759,N_24361,N_24062);
xor U24760 (N_24760,N_24190,N_24040);
xnor U24761 (N_24761,N_24114,N_24293);
and U24762 (N_24762,N_24245,N_24018);
nor U24763 (N_24763,N_24295,N_24212);
nand U24764 (N_24764,N_24499,N_24031);
and U24765 (N_24765,N_24168,N_24007);
and U24766 (N_24766,N_24251,N_24364);
or U24767 (N_24767,N_24445,N_24400);
or U24768 (N_24768,N_24287,N_24191);
nor U24769 (N_24769,N_24441,N_24203);
xnor U24770 (N_24770,N_24307,N_24448);
xor U24771 (N_24771,N_24492,N_24087);
and U24772 (N_24772,N_24062,N_24387);
nor U24773 (N_24773,N_24266,N_24365);
and U24774 (N_24774,N_24255,N_24430);
and U24775 (N_24775,N_24269,N_24262);
xor U24776 (N_24776,N_24313,N_24090);
nand U24777 (N_24777,N_24353,N_24342);
nand U24778 (N_24778,N_24233,N_24357);
xnor U24779 (N_24779,N_24091,N_24457);
nand U24780 (N_24780,N_24075,N_24162);
nand U24781 (N_24781,N_24129,N_24178);
xor U24782 (N_24782,N_24185,N_24034);
or U24783 (N_24783,N_24156,N_24192);
nand U24784 (N_24784,N_24195,N_24040);
and U24785 (N_24785,N_24202,N_24473);
nor U24786 (N_24786,N_24432,N_24237);
and U24787 (N_24787,N_24081,N_24121);
xor U24788 (N_24788,N_24070,N_24125);
or U24789 (N_24789,N_24247,N_24378);
xnor U24790 (N_24790,N_24206,N_24121);
xor U24791 (N_24791,N_24170,N_24307);
and U24792 (N_24792,N_24417,N_24228);
xnor U24793 (N_24793,N_24074,N_24105);
or U24794 (N_24794,N_24211,N_24054);
or U24795 (N_24795,N_24338,N_24466);
or U24796 (N_24796,N_24138,N_24480);
xor U24797 (N_24797,N_24426,N_24228);
or U24798 (N_24798,N_24472,N_24307);
nand U24799 (N_24799,N_24102,N_24163);
nand U24800 (N_24800,N_24311,N_24134);
xor U24801 (N_24801,N_24440,N_24393);
xor U24802 (N_24802,N_24134,N_24384);
nor U24803 (N_24803,N_24141,N_24496);
and U24804 (N_24804,N_24166,N_24260);
or U24805 (N_24805,N_24274,N_24037);
nand U24806 (N_24806,N_24492,N_24130);
xnor U24807 (N_24807,N_24470,N_24033);
and U24808 (N_24808,N_24403,N_24225);
or U24809 (N_24809,N_24279,N_24190);
xor U24810 (N_24810,N_24199,N_24273);
xor U24811 (N_24811,N_24002,N_24362);
nand U24812 (N_24812,N_24059,N_24239);
nand U24813 (N_24813,N_24105,N_24385);
and U24814 (N_24814,N_24108,N_24303);
nand U24815 (N_24815,N_24296,N_24417);
or U24816 (N_24816,N_24222,N_24324);
xnor U24817 (N_24817,N_24006,N_24007);
or U24818 (N_24818,N_24280,N_24318);
xor U24819 (N_24819,N_24142,N_24468);
and U24820 (N_24820,N_24454,N_24364);
and U24821 (N_24821,N_24424,N_24207);
or U24822 (N_24822,N_24454,N_24265);
xnor U24823 (N_24823,N_24151,N_24067);
and U24824 (N_24824,N_24083,N_24141);
xnor U24825 (N_24825,N_24349,N_24094);
and U24826 (N_24826,N_24488,N_24281);
and U24827 (N_24827,N_24410,N_24191);
nor U24828 (N_24828,N_24098,N_24324);
or U24829 (N_24829,N_24250,N_24377);
or U24830 (N_24830,N_24194,N_24302);
and U24831 (N_24831,N_24282,N_24038);
nor U24832 (N_24832,N_24202,N_24275);
and U24833 (N_24833,N_24376,N_24070);
and U24834 (N_24834,N_24120,N_24104);
nor U24835 (N_24835,N_24344,N_24101);
nor U24836 (N_24836,N_24082,N_24409);
or U24837 (N_24837,N_24022,N_24321);
nor U24838 (N_24838,N_24494,N_24496);
nor U24839 (N_24839,N_24205,N_24292);
nor U24840 (N_24840,N_24326,N_24314);
or U24841 (N_24841,N_24102,N_24116);
nand U24842 (N_24842,N_24262,N_24274);
nor U24843 (N_24843,N_24057,N_24124);
xor U24844 (N_24844,N_24405,N_24273);
and U24845 (N_24845,N_24191,N_24333);
and U24846 (N_24846,N_24322,N_24287);
xnor U24847 (N_24847,N_24402,N_24157);
or U24848 (N_24848,N_24294,N_24042);
nand U24849 (N_24849,N_24136,N_24253);
nor U24850 (N_24850,N_24186,N_24044);
and U24851 (N_24851,N_24466,N_24164);
nand U24852 (N_24852,N_24244,N_24225);
nand U24853 (N_24853,N_24338,N_24086);
nand U24854 (N_24854,N_24342,N_24337);
xnor U24855 (N_24855,N_24154,N_24299);
nor U24856 (N_24856,N_24288,N_24236);
and U24857 (N_24857,N_24253,N_24018);
and U24858 (N_24858,N_24359,N_24283);
or U24859 (N_24859,N_24023,N_24429);
nand U24860 (N_24860,N_24147,N_24192);
nand U24861 (N_24861,N_24165,N_24170);
and U24862 (N_24862,N_24352,N_24194);
or U24863 (N_24863,N_24146,N_24118);
nand U24864 (N_24864,N_24406,N_24027);
nand U24865 (N_24865,N_24461,N_24285);
xnor U24866 (N_24866,N_24099,N_24047);
or U24867 (N_24867,N_24042,N_24043);
xnor U24868 (N_24868,N_24295,N_24156);
or U24869 (N_24869,N_24136,N_24382);
xnor U24870 (N_24870,N_24444,N_24096);
or U24871 (N_24871,N_24246,N_24296);
xnor U24872 (N_24872,N_24247,N_24244);
nor U24873 (N_24873,N_24141,N_24044);
nor U24874 (N_24874,N_24200,N_24479);
or U24875 (N_24875,N_24338,N_24333);
xor U24876 (N_24876,N_24452,N_24093);
nor U24877 (N_24877,N_24175,N_24160);
nor U24878 (N_24878,N_24064,N_24141);
xnor U24879 (N_24879,N_24005,N_24342);
nand U24880 (N_24880,N_24460,N_24409);
xor U24881 (N_24881,N_24145,N_24444);
or U24882 (N_24882,N_24005,N_24450);
nor U24883 (N_24883,N_24405,N_24045);
and U24884 (N_24884,N_24218,N_24134);
nand U24885 (N_24885,N_24163,N_24327);
and U24886 (N_24886,N_24136,N_24249);
xnor U24887 (N_24887,N_24194,N_24381);
nor U24888 (N_24888,N_24336,N_24141);
nor U24889 (N_24889,N_24309,N_24488);
nand U24890 (N_24890,N_24151,N_24126);
nand U24891 (N_24891,N_24078,N_24385);
and U24892 (N_24892,N_24456,N_24426);
and U24893 (N_24893,N_24332,N_24295);
nand U24894 (N_24894,N_24439,N_24125);
xor U24895 (N_24895,N_24098,N_24122);
nor U24896 (N_24896,N_24207,N_24256);
xnor U24897 (N_24897,N_24059,N_24078);
or U24898 (N_24898,N_24361,N_24239);
nand U24899 (N_24899,N_24180,N_24450);
and U24900 (N_24900,N_24389,N_24226);
and U24901 (N_24901,N_24087,N_24405);
xor U24902 (N_24902,N_24446,N_24496);
xnor U24903 (N_24903,N_24269,N_24232);
nand U24904 (N_24904,N_24065,N_24257);
and U24905 (N_24905,N_24360,N_24483);
or U24906 (N_24906,N_24088,N_24018);
or U24907 (N_24907,N_24006,N_24124);
or U24908 (N_24908,N_24194,N_24131);
nor U24909 (N_24909,N_24248,N_24296);
and U24910 (N_24910,N_24154,N_24001);
xnor U24911 (N_24911,N_24453,N_24404);
nor U24912 (N_24912,N_24194,N_24208);
and U24913 (N_24913,N_24348,N_24031);
or U24914 (N_24914,N_24377,N_24208);
and U24915 (N_24915,N_24313,N_24027);
nand U24916 (N_24916,N_24417,N_24400);
nor U24917 (N_24917,N_24462,N_24028);
nand U24918 (N_24918,N_24480,N_24467);
and U24919 (N_24919,N_24229,N_24401);
or U24920 (N_24920,N_24423,N_24369);
nor U24921 (N_24921,N_24397,N_24383);
nor U24922 (N_24922,N_24445,N_24304);
or U24923 (N_24923,N_24274,N_24488);
and U24924 (N_24924,N_24314,N_24113);
and U24925 (N_24925,N_24127,N_24021);
and U24926 (N_24926,N_24287,N_24497);
nor U24927 (N_24927,N_24014,N_24493);
and U24928 (N_24928,N_24221,N_24229);
xnor U24929 (N_24929,N_24384,N_24415);
and U24930 (N_24930,N_24160,N_24455);
nor U24931 (N_24931,N_24259,N_24055);
and U24932 (N_24932,N_24035,N_24336);
and U24933 (N_24933,N_24166,N_24362);
and U24934 (N_24934,N_24080,N_24121);
or U24935 (N_24935,N_24203,N_24007);
or U24936 (N_24936,N_24411,N_24098);
nand U24937 (N_24937,N_24163,N_24495);
or U24938 (N_24938,N_24490,N_24060);
nor U24939 (N_24939,N_24149,N_24406);
and U24940 (N_24940,N_24028,N_24445);
xor U24941 (N_24941,N_24414,N_24168);
nor U24942 (N_24942,N_24384,N_24483);
nand U24943 (N_24943,N_24165,N_24121);
or U24944 (N_24944,N_24247,N_24154);
nand U24945 (N_24945,N_24045,N_24244);
or U24946 (N_24946,N_24166,N_24198);
nand U24947 (N_24947,N_24395,N_24293);
nand U24948 (N_24948,N_24360,N_24160);
nor U24949 (N_24949,N_24433,N_24026);
or U24950 (N_24950,N_24016,N_24193);
nor U24951 (N_24951,N_24170,N_24309);
xor U24952 (N_24952,N_24416,N_24227);
nor U24953 (N_24953,N_24452,N_24184);
and U24954 (N_24954,N_24259,N_24241);
and U24955 (N_24955,N_24477,N_24460);
and U24956 (N_24956,N_24000,N_24436);
or U24957 (N_24957,N_24114,N_24285);
or U24958 (N_24958,N_24330,N_24324);
or U24959 (N_24959,N_24451,N_24069);
nor U24960 (N_24960,N_24448,N_24087);
and U24961 (N_24961,N_24222,N_24337);
nand U24962 (N_24962,N_24155,N_24170);
or U24963 (N_24963,N_24097,N_24314);
nor U24964 (N_24964,N_24095,N_24373);
xnor U24965 (N_24965,N_24395,N_24361);
nand U24966 (N_24966,N_24445,N_24059);
xnor U24967 (N_24967,N_24141,N_24089);
nand U24968 (N_24968,N_24087,N_24271);
and U24969 (N_24969,N_24110,N_24200);
nand U24970 (N_24970,N_24100,N_24124);
or U24971 (N_24971,N_24265,N_24317);
xor U24972 (N_24972,N_24184,N_24445);
nor U24973 (N_24973,N_24297,N_24160);
and U24974 (N_24974,N_24200,N_24470);
nor U24975 (N_24975,N_24378,N_24096);
and U24976 (N_24976,N_24336,N_24073);
xor U24977 (N_24977,N_24329,N_24352);
or U24978 (N_24978,N_24174,N_24153);
or U24979 (N_24979,N_24194,N_24071);
nand U24980 (N_24980,N_24038,N_24152);
or U24981 (N_24981,N_24126,N_24150);
nor U24982 (N_24982,N_24351,N_24127);
nand U24983 (N_24983,N_24403,N_24440);
and U24984 (N_24984,N_24261,N_24428);
nor U24985 (N_24985,N_24351,N_24217);
xor U24986 (N_24986,N_24270,N_24105);
nand U24987 (N_24987,N_24173,N_24132);
xnor U24988 (N_24988,N_24340,N_24263);
and U24989 (N_24989,N_24040,N_24061);
xor U24990 (N_24990,N_24211,N_24103);
nand U24991 (N_24991,N_24160,N_24443);
and U24992 (N_24992,N_24084,N_24083);
or U24993 (N_24993,N_24180,N_24384);
and U24994 (N_24994,N_24367,N_24032);
and U24995 (N_24995,N_24089,N_24307);
nand U24996 (N_24996,N_24436,N_24443);
nand U24997 (N_24997,N_24112,N_24136);
xnor U24998 (N_24998,N_24027,N_24122);
nand U24999 (N_24999,N_24186,N_24124);
nor U25000 (N_25000,N_24878,N_24994);
or U25001 (N_25001,N_24528,N_24943);
nand U25002 (N_25002,N_24643,N_24588);
and U25003 (N_25003,N_24745,N_24567);
nand U25004 (N_25004,N_24999,N_24713);
and U25005 (N_25005,N_24992,N_24852);
or U25006 (N_25006,N_24502,N_24654);
xnor U25007 (N_25007,N_24947,N_24846);
nor U25008 (N_25008,N_24792,N_24694);
and U25009 (N_25009,N_24904,N_24711);
nor U25010 (N_25010,N_24923,N_24721);
or U25011 (N_25011,N_24700,N_24996);
nor U25012 (N_25012,N_24738,N_24599);
xnor U25013 (N_25013,N_24801,N_24608);
or U25014 (N_25014,N_24649,N_24749);
xor U25015 (N_25015,N_24642,N_24916);
xnor U25016 (N_25016,N_24618,N_24979);
nor U25017 (N_25017,N_24803,N_24504);
nand U25018 (N_25018,N_24744,N_24731);
xnor U25019 (N_25019,N_24962,N_24871);
or U25020 (N_25020,N_24714,N_24593);
or U25021 (N_25021,N_24679,N_24733);
nand U25022 (N_25022,N_24970,N_24676);
or U25023 (N_25023,N_24816,N_24865);
xnor U25024 (N_25024,N_24836,N_24837);
nor U25025 (N_25025,N_24685,N_24965);
xor U25026 (N_25026,N_24977,N_24578);
or U25027 (N_25027,N_24523,N_24555);
xor U25028 (N_25028,N_24840,N_24696);
nand U25029 (N_25029,N_24921,N_24531);
or U25030 (N_25030,N_24814,N_24621);
xnor U25031 (N_25031,N_24874,N_24625);
and U25032 (N_25032,N_24752,N_24762);
xor U25033 (N_25033,N_24791,N_24520);
xnor U25034 (N_25034,N_24628,N_24632);
or U25035 (N_25035,N_24764,N_24688);
nand U25036 (N_25036,N_24712,N_24845);
or U25037 (N_25037,N_24842,N_24532);
xor U25038 (N_25038,N_24748,N_24760);
and U25039 (N_25039,N_24701,N_24975);
or U25040 (N_25040,N_24615,N_24873);
nand U25041 (N_25041,N_24849,N_24674);
xnor U25042 (N_25042,N_24743,N_24561);
nand U25043 (N_25043,N_24716,N_24747);
nand U25044 (N_25044,N_24880,N_24525);
and U25045 (N_25045,N_24751,N_24899);
and U25046 (N_25046,N_24914,N_24927);
nand U25047 (N_25047,N_24956,N_24972);
nand U25048 (N_25048,N_24834,N_24683);
or U25049 (N_25049,N_24919,N_24690);
or U25050 (N_25050,N_24997,N_24945);
xnor U25051 (N_25051,N_24856,N_24802);
or U25052 (N_25052,N_24828,N_24663);
nor U25053 (N_25053,N_24825,N_24616);
or U25054 (N_25054,N_24887,N_24510);
xnor U25055 (N_25055,N_24551,N_24785);
and U25056 (N_25056,N_24987,N_24798);
or U25057 (N_25057,N_24544,N_24854);
xnor U25058 (N_25058,N_24793,N_24967);
or U25059 (N_25059,N_24838,N_24547);
xor U25060 (N_25060,N_24960,N_24895);
xor U25061 (N_25061,N_24583,N_24860);
nand U25062 (N_25062,N_24613,N_24804);
and U25063 (N_25063,N_24824,N_24682);
xor U25064 (N_25064,N_24884,N_24806);
xnor U25065 (N_25065,N_24678,N_24695);
and U25066 (N_25066,N_24991,N_24641);
nor U25067 (N_25067,N_24783,N_24777);
nor U25068 (N_25068,N_24626,N_24560);
and U25069 (N_25069,N_24835,N_24570);
and U25070 (N_25070,N_24697,N_24565);
and U25071 (N_25071,N_24766,N_24848);
nor U25072 (N_25072,N_24993,N_24647);
nand U25073 (N_25073,N_24867,N_24774);
and U25074 (N_25074,N_24959,N_24844);
nor U25075 (N_25075,N_24732,N_24581);
and U25076 (N_25076,N_24754,N_24717);
and U25077 (N_25077,N_24763,N_24596);
and U25078 (N_25078,N_24557,N_24981);
nand U25079 (N_25079,N_24589,N_24818);
or U25080 (N_25080,N_24590,N_24522);
and U25081 (N_25081,N_24984,N_24868);
nand U25082 (N_25082,N_24724,N_24808);
and U25083 (N_25083,N_24820,N_24709);
nand U25084 (N_25084,N_24636,N_24656);
nand U25085 (N_25085,N_24909,N_24897);
and U25086 (N_25086,N_24813,N_24668);
nand U25087 (N_25087,N_24669,N_24817);
nand U25088 (N_25088,N_24646,N_24657);
and U25089 (N_25089,N_24794,N_24910);
xor U25090 (N_25090,N_24689,N_24508);
nor U25091 (N_25091,N_24603,N_24841);
nand U25092 (N_25092,N_24526,N_24638);
and U25093 (N_25093,N_24619,N_24606);
or U25094 (N_25094,N_24660,N_24926);
nand U25095 (N_25095,N_24637,N_24799);
and U25096 (N_25096,N_24549,N_24604);
nand U25097 (N_25097,N_24784,N_24976);
xnor U25098 (N_25098,N_24903,N_24985);
nor U25099 (N_25099,N_24753,N_24807);
or U25100 (N_25100,N_24719,N_24691);
nand U25101 (N_25101,N_24958,N_24624);
nand U25102 (N_25102,N_24986,N_24995);
nand U25103 (N_25103,N_24584,N_24595);
nor U25104 (N_25104,N_24827,N_24915);
nor U25105 (N_25105,N_24750,N_24586);
or U25106 (N_25106,N_24514,N_24665);
nand U25107 (N_25107,N_24969,N_24759);
xor U25108 (N_25108,N_24574,N_24545);
xnor U25109 (N_25109,N_24662,N_24866);
nor U25110 (N_25110,N_24773,N_24853);
nor U25111 (N_25111,N_24964,N_24500);
or U25112 (N_25112,N_24631,N_24672);
xor U25113 (N_25113,N_24515,N_24881);
xor U25114 (N_25114,N_24609,N_24620);
or U25115 (N_25115,N_24861,N_24851);
xnor U25116 (N_25116,N_24907,N_24686);
or U25117 (N_25117,N_24896,N_24612);
and U25118 (N_25118,N_24534,N_24627);
or U25119 (N_25119,N_24829,N_24629);
or U25120 (N_25120,N_24571,N_24894);
nand U25121 (N_25121,N_24790,N_24651);
nor U25122 (N_25122,N_24601,N_24602);
nand U25123 (N_25123,N_24772,N_24706);
nand U25124 (N_25124,N_24537,N_24891);
and U25125 (N_25125,N_24900,N_24901);
xor U25126 (N_25126,N_24677,N_24902);
and U25127 (N_25127,N_24684,N_24832);
or U25128 (N_25128,N_24811,N_24533);
and U25129 (N_25129,N_24670,N_24779);
or U25130 (N_25130,N_24558,N_24756);
nor U25131 (N_25131,N_24862,N_24710);
and U25132 (N_25132,N_24890,N_24505);
or U25133 (N_25133,N_24990,N_24585);
nor U25134 (N_25134,N_24587,N_24704);
nor U25135 (N_25135,N_24623,N_24591);
xor U25136 (N_25136,N_24847,N_24725);
xor U25137 (N_25137,N_24573,N_24575);
or U25138 (N_25138,N_24973,N_24889);
or U25139 (N_25139,N_24949,N_24998);
nor U25140 (N_25140,N_24776,N_24529);
nand U25141 (N_25141,N_24611,N_24705);
and U25142 (N_25142,N_24942,N_24655);
xor U25143 (N_25143,N_24800,N_24506);
and U25144 (N_25144,N_24550,N_24918);
nand U25145 (N_25145,N_24727,N_24906);
nor U25146 (N_25146,N_24644,N_24607);
and U25147 (N_25147,N_24989,N_24518);
nand U25148 (N_25148,N_24519,N_24787);
and U25149 (N_25149,N_24703,N_24680);
or U25150 (N_25150,N_24730,N_24786);
nor U25151 (N_25151,N_24513,N_24941);
or U25152 (N_25152,N_24598,N_24737);
nor U25153 (N_25153,N_24931,N_24815);
nor U25154 (N_25154,N_24592,N_24819);
xnor U25155 (N_25155,N_24564,N_24671);
nor U25156 (N_25156,N_24938,N_24857);
and U25157 (N_25157,N_24954,N_24882);
nor U25158 (N_25158,N_24940,N_24877);
and U25159 (N_25159,N_24582,N_24610);
nand U25160 (N_25160,N_24934,N_24501);
nor U25161 (N_25161,N_24512,N_24830);
or U25162 (N_25162,N_24864,N_24952);
nor U25163 (N_25163,N_24707,N_24594);
and U25164 (N_25164,N_24755,N_24600);
xnor U25165 (N_25165,N_24666,N_24963);
and U25166 (N_25166,N_24879,N_24980);
nor U25167 (N_25167,N_24734,N_24988);
xor U25168 (N_25168,N_24948,N_24635);
nor U25169 (N_25169,N_24539,N_24722);
nand U25170 (N_25170,N_24516,N_24950);
or U25171 (N_25171,N_24870,N_24805);
or U25172 (N_25172,N_24645,N_24788);
nand U25173 (N_25173,N_24729,N_24661);
and U25174 (N_25174,N_24576,N_24823);
nor U25175 (N_25175,N_24568,N_24780);
nand U25176 (N_25176,N_24978,N_24524);
or U25177 (N_25177,N_24653,N_24789);
and U25178 (N_25178,N_24634,N_24968);
or U25179 (N_25179,N_24546,N_24888);
nor U25180 (N_25180,N_24858,N_24863);
or U25181 (N_25181,N_24886,N_24767);
and U25182 (N_25182,N_24742,N_24920);
nand U25183 (N_25183,N_24859,N_24698);
and U25184 (N_25184,N_24699,N_24933);
nor U25185 (N_25185,N_24892,N_24809);
and U25186 (N_25186,N_24944,N_24736);
xor U25187 (N_25187,N_24869,N_24741);
xor U25188 (N_25188,N_24775,N_24580);
xnor U25189 (N_25189,N_24702,N_24530);
nor U25190 (N_25190,N_24850,N_24511);
nor U25191 (N_25191,N_24681,N_24553);
and U25192 (N_25192,N_24566,N_24739);
nor U25193 (N_25193,N_24687,N_24912);
and U25194 (N_25194,N_24572,N_24543);
and U25195 (N_25195,N_24843,N_24821);
and U25196 (N_25196,N_24936,N_24778);
or U25197 (N_25197,N_24548,N_24939);
nand U25198 (N_25198,N_24839,N_24723);
nand U25199 (N_25199,N_24652,N_24810);
nor U25200 (N_25200,N_24639,N_24893);
or U25201 (N_25201,N_24708,N_24605);
nand U25202 (N_25202,N_24913,N_24633);
nand U25203 (N_25203,N_24872,N_24535);
nand U25204 (N_25204,N_24797,N_24795);
nand U25205 (N_25205,N_24517,N_24664);
xnor U25206 (N_25206,N_24951,N_24740);
xor U25207 (N_25207,N_24957,N_24768);
nand U25208 (N_25208,N_24930,N_24982);
nand U25209 (N_25209,N_24782,N_24536);
and U25210 (N_25210,N_24735,N_24559);
nand U25211 (N_25211,N_24855,N_24971);
nor U25212 (N_25212,N_24563,N_24746);
xnor U25213 (N_25213,N_24761,N_24715);
or U25214 (N_25214,N_24720,N_24577);
or U25215 (N_25215,N_24922,N_24507);
or U25216 (N_25216,N_24614,N_24503);
or U25217 (N_25217,N_24728,N_24579);
and U25218 (N_25218,N_24781,N_24883);
and U25219 (N_25219,N_24554,N_24898);
xnor U25220 (N_25220,N_24667,N_24974);
nand U25221 (N_25221,N_24961,N_24552);
or U25222 (N_25222,N_24833,N_24812);
nor U25223 (N_25223,N_24648,N_24932);
nand U25224 (N_25224,N_24765,N_24675);
nor U25225 (N_25225,N_24630,N_24538);
xnor U25226 (N_25226,N_24540,N_24928);
and U25227 (N_25227,N_24541,N_24718);
or U25228 (N_25228,N_24692,N_24562);
nor U25229 (N_25229,N_24769,N_24796);
nand U25230 (N_25230,N_24831,N_24946);
nor U25231 (N_25231,N_24955,N_24924);
xnor U25232 (N_25232,N_24650,N_24509);
xnor U25233 (N_25233,N_24521,N_24659);
nand U25234 (N_25234,N_24597,N_24771);
nor U25235 (N_25235,N_24673,N_24929);
or U25236 (N_25236,N_24726,N_24617);
or U25237 (N_25237,N_24826,N_24556);
nand U25238 (N_25238,N_24966,N_24770);
nor U25239 (N_25239,N_24905,N_24640);
nand U25240 (N_25240,N_24757,N_24542);
nand U25241 (N_25241,N_24658,N_24876);
nand U25242 (N_25242,N_24527,N_24983);
nor U25243 (N_25243,N_24953,N_24937);
nor U25244 (N_25244,N_24917,N_24693);
nor U25245 (N_25245,N_24758,N_24569);
nand U25246 (N_25246,N_24885,N_24911);
nor U25247 (N_25247,N_24935,N_24925);
xor U25248 (N_25248,N_24908,N_24822);
nand U25249 (N_25249,N_24875,N_24622);
or U25250 (N_25250,N_24893,N_24922);
xor U25251 (N_25251,N_24598,N_24980);
xor U25252 (N_25252,N_24649,N_24789);
nor U25253 (N_25253,N_24622,N_24606);
xor U25254 (N_25254,N_24584,N_24649);
and U25255 (N_25255,N_24586,N_24615);
xnor U25256 (N_25256,N_24917,N_24514);
and U25257 (N_25257,N_24791,N_24807);
xnor U25258 (N_25258,N_24640,N_24695);
or U25259 (N_25259,N_24862,N_24723);
or U25260 (N_25260,N_24733,N_24584);
nand U25261 (N_25261,N_24559,N_24914);
nor U25262 (N_25262,N_24645,N_24950);
and U25263 (N_25263,N_24617,N_24930);
xor U25264 (N_25264,N_24557,N_24735);
or U25265 (N_25265,N_24889,N_24813);
or U25266 (N_25266,N_24932,N_24720);
nor U25267 (N_25267,N_24615,N_24560);
or U25268 (N_25268,N_24865,N_24748);
xor U25269 (N_25269,N_24808,N_24924);
or U25270 (N_25270,N_24521,N_24853);
or U25271 (N_25271,N_24947,N_24784);
or U25272 (N_25272,N_24834,N_24792);
or U25273 (N_25273,N_24652,N_24944);
xor U25274 (N_25274,N_24701,N_24534);
nor U25275 (N_25275,N_24691,N_24511);
nand U25276 (N_25276,N_24845,N_24502);
or U25277 (N_25277,N_24755,N_24695);
xnor U25278 (N_25278,N_24672,N_24742);
or U25279 (N_25279,N_24805,N_24544);
nor U25280 (N_25280,N_24734,N_24586);
nor U25281 (N_25281,N_24969,N_24689);
xnor U25282 (N_25282,N_24716,N_24738);
nand U25283 (N_25283,N_24818,N_24736);
nand U25284 (N_25284,N_24939,N_24974);
and U25285 (N_25285,N_24567,N_24560);
or U25286 (N_25286,N_24523,N_24547);
and U25287 (N_25287,N_24562,N_24553);
xor U25288 (N_25288,N_24961,N_24956);
nand U25289 (N_25289,N_24747,N_24914);
xnor U25290 (N_25290,N_24766,N_24542);
and U25291 (N_25291,N_24720,N_24796);
nand U25292 (N_25292,N_24998,N_24644);
nor U25293 (N_25293,N_24916,N_24657);
nor U25294 (N_25294,N_24758,N_24869);
and U25295 (N_25295,N_24580,N_24539);
nor U25296 (N_25296,N_24886,N_24623);
xnor U25297 (N_25297,N_24832,N_24815);
nor U25298 (N_25298,N_24946,N_24740);
nor U25299 (N_25299,N_24975,N_24757);
nand U25300 (N_25300,N_24747,N_24707);
nand U25301 (N_25301,N_24876,N_24634);
xnor U25302 (N_25302,N_24891,N_24751);
nor U25303 (N_25303,N_24710,N_24539);
or U25304 (N_25304,N_24828,N_24952);
or U25305 (N_25305,N_24873,N_24824);
nand U25306 (N_25306,N_24671,N_24666);
nand U25307 (N_25307,N_24903,N_24566);
or U25308 (N_25308,N_24736,N_24651);
xor U25309 (N_25309,N_24760,N_24571);
nor U25310 (N_25310,N_24786,N_24992);
nand U25311 (N_25311,N_24972,N_24980);
nor U25312 (N_25312,N_24756,N_24929);
xnor U25313 (N_25313,N_24803,N_24569);
nor U25314 (N_25314,N_24822,N_24528);
nor U25315 (N_25315,N_24562,N_24539);
nor U25316 (N_25316,N_24572,N_24544);
xor U25317 (N_25317,N_24826,N_24896);
or U25318 (N_25318,N_24944,N_24833);
and U25319 (N_25319,N_24887,N_24679);
or U25320 (N_25320,N_24602,N_24966);
and U25321 (N_25321,N_24796,N_24835);
or U25322 (N_25322,N_24812,N_24596);
and U25323 (N_25323,N_24891,N_24566);
nor U25324 (N_25324,N_24551,N_24676);
nand U25325 (N_25325,N_24750,N_24774);
nand U25326 (N_25326,N_24664,N_24653);
xnor U25327 (N_25327,N_24535,N_24793);
xor U25328 (N_25328,N_24926,N_24636);
xnor U25329 (N_25329,N_24904,N_24901);
nor U25330 (N_25330,N_24615,N_24598);
nand U25331 (N_25331,N_24787,N_24504);
xnor U25332 (N_25332,N_24906,N_24883);
nand U25333 (N_25333,N_24928,N_24578);
xnor U25334 (N_25334,N_24729,N_24634);
xnor U25335 (N_25335,N_24697,N_24708);
nand U25336 (N_25336,N_24990,N_24538);
nand U25337 (N_25337,N_24605,N_24777);
and U25338 (N_25338,N_24993,N_24639);
nand U25339 (N_25339,N_24842,N_24544);
and U25340 (N_25340,N_24607,N_24551);
xor U25341 (N_25341,N_24540,N_24920);
and U25342 (N_25342,N_24790,N_24738);
nand U25343 (N_25343,N_24605,N_24698);
and U25344 (N_25344,N_24667,N_24852);
and U25345 (N_25345,N_24820,N_24586);
or U25346 (N_25346,N_24793,N_24805);
xor U25347 (N_25347,N_24952,N_24626);
nand U25348 (N_25348,N_24783,N_24771);
and U25349 (N_25349,N_24531,N_24872);
or U25350 (N_25350,N_24558,N_24512);
xnor U25351 (N_25351,N_24513,N_24633);
and U25352 (N_25352,N_24869,N_24780);
and U25353 (N_25353,N_24530,N_24742);
and U25354 (N_25354,N_24616,N_24719);
nor U25355 (N_25355,N_24763,N_24958);
xnor U25356 (N_25356,N_24670,N_24664);
nand U25357 (N_25357,N_24762,N_24523);
or U25358 (N_25358,N_24780,N_24654);
or U25359 (N_25359,N_24580,N_24869);
nand U25360 (N_25360,N_24927,N_24711);
nor U25361 (N_25361,N_24855,N_24706);
nor U25362 (N_25362,N_24809,N_24850);
and U25363 (N_25363,N_24939,N_24664);
xor U25364 (N_25364,N_24577,N_24525);
nor U25365 (N_25365,N_24802,N_24991);
xor U25366 (N_25366,N_24786,N_24864);
and U25367 (N_25367,N_24683,N_24546);
xnor U25368 (N_25368,N_24863,N_24848);
and U25369 (N_25369,N_24547,N_24735);
nor U25370 (N_25370,N_24829,N_24882);
nand U25371 (N_25371,N_24798,N_24896);
nor U25372 (N_25372,N_24513,N_24891);
nor U25373 (N_25373,N_24629,N_24631);
or U25374 (N_25374,N_24688,N_24713);
and U25375 (N_25375,N_24825,N_24943);
and U25376 (N_25376,N_24784,N_24600);
nor U25377 (N_25377,N_24876,N_24612);
or U25378 (N_25378,N_24956,N_24527);
nor U25379 (N_25379,N_24951,N_24864);
nand U25380 (N_25380,N_24785,N_24748);
or U25381 (N_25381,N_24990,N_24721);
nor U25382 (N_25382,N_24817,N_24780);
nand U25383 (N_25383,N_24624,N_24917);
and U25384 (N_25384,N_24929,N_24780);
or U25385 (N_25385,N_24710,N_24838);
nand U25386 (N_25386,N_24607,N_24969);
nor U25387 (N_25387,N_24858,N_24905);
or U25388 (N_25388,N_24927,N_24557);
nor U25389 (N_25389,N_24895,N_24715);
nand U25390 (N_25390,N_24535,N_24578);
and U25391 (N_25391,N_24623,N_24583);
xor U25392 (N_25392,N_24543,N_24582);
nor U25393 (N_25393,N_24505,N_24656);
xnor U25394 (N_25394,N_24545,N_24865);
nand U25395 (N_25395,N_24849,N_24898);
and U25396 (N_25396,N_24554,N_24728);
or U25397 (N_25397,N_24627,N_24699);
nand U25398 (N_25398,N_24757,N_24907);
or U25399 (N_25399,N_24822,N_24727);
xnor U25400 (N_25400,N_24863,N_24685);
nand U25401 (N_25401,N_24706,N_24702);
or U25402 (N_25402,N_24586,N_24873);
or U25403 (N_25403,N_24622,N_24952);
or U25404 (N_25404,N_24806,N_24658);
nor U25405 (N_25405,N_24552,N_24957);
or U25406 (N_25406,N_24885,N_24881);
nor U25407 (N_25407,N_24569,N_24538);
and U25408 (N_25408,N_24658,N_24666);
xor U25409 (N_25409,N_24829,N_24520);
nor U25410 (N_25410,N_24638,N_24944);
xor U25411 (N_25411,N_24627,N_24600);
xor U25412 (N_25412,N_24693,N_24761);
or U25413 (N_25413,N_24855,N_24670);
and U25414 (N_25414,N_24591,N_24725);
nand U25415 (N_25415,N_24559,N_24951);
xnor U25416 (N_25416,N_24886,N_24677);
and U25417 (N_25417,N_24835,N_24549);
xnor U25418 (N_25418,N_24630,N_24675);
and U25419 (N_25419,N_24515,N_24878);
and U25420 (N_25420,N_24693,N_24819);
or U25421 (N_25421,N_24589,N_24820);
or U25422 (N_25422,N_24973,N_24502);
or U25423 (N_25423,N_24611,N_24677);
nor U25424 (N_25424,N_24572,N_24745);
and U25425 (N_25425,N_24725,N_24646);
nand U25426 (N_25426,N_24828,N_24931);
and U25427 (N_25427,N_24627,N_24894);
nand U25428 (N_25428,N_24621,N_24749);
or U25429 (N_25429,N_24820,N_24608);
nand U25430 (N_25430,N_24584,N_24634);
or U25431 (N_25431,N_24714,N_24881);
nor U25432 (N_25432,N_24556,N_24586);
nor U25433 (N_25433,N_24742,N_24651);
nand U25434 (N_25434,N_24743,N_24718);
xnor U25435 (N_25435,N_24648,N_24514);
or U25436 (N_25436,N_24727,N_24639);
nor U25437 (N_25437,N_24605,N_24822);
or U25438 (N_25438,N_24796,N_24773);
nand U25439 (N_25439,N_24898,N_24826);
nor U25440 (N_25440,N_24947,N_24808);
and U25441 (N_25441,N_24641,N_24637);
or U25442 (N_25442,N_24506,N_24912);
or U25443 (N_25443,N_24842,N_24968);
nand U25444 (N_25444,N_24973,N_24722);
and U25445 (N_25445,N_24906,N_24783);
nor U25446 (N_25446,N_24515,N_24527);
nand U25447 (N_25447,N_24574,N_24536);
and U25448 (N_25448,N_24562,N_24832);
and U25449 (N_25449,N_24988,N_24659);
nor U25450 (N_25450,N_24568,N_24934);
nand U25451 (N_25451,N_24545,N_24635);
xor U25452 (N_25452,N_24731,N_24876);
nand U25453 (N_25453,N_24759,N_24930);
and U25454 (N_25454,N_24574,N_24522);
xnor U25455 (N_25455,N_24754,N_24512);
nand U25456 (N_25456,N_24580,N_24753);
or U25457 (N_25457,N_24609,N_24716);
and U25458 (N_25458,N_24537,N_24919);
or U25459 (N_25459,N_24556,N_24682);
or U25460 (N_25460,N_24718,N_24841);
or U25461 (N_25461,N_24618,N_24889);
nor U25462 (N_25462,N_24583,N_24972);
xnor U25463 (N_25463,N_24855,N_24836);
xnor U25464 (N_25464,N_24935,N_24608);
nand U25465 (N_25465,N_24822,N_24658);
nand U25466 (N_25466,N_24832,N_24809);
or U25467 (N_25467,N_24896,N_24905);
xor U25468 (N_25468,N_24623,N_24566);
or U25469 (N_25469,N_24725,N_24778);
xnor U25470 (N_25470,N_24856,N_24598);
or U25471 (N_25471,N_24559,N_24529);
nand U25472 (N_25472,N_24665,N_24786);
or U25473 (N_25473,N_24700,N_24725);
or U25474 (N_25474,N_24649,N_24691);
nor U25475 (N_25475,N_24828,N_24629);
xor U25476 (N_25476,N_24607,N_24564);
or U25477 (N_25477,N_24582,N_24558);
nand U25478 (N_25478,N_24801,N_24926);
or U25479 (N_25479,N_24799,N_24851);
nand U25480 (N_25480,N_24517,N_24648);
and U25481 (N_25481,N_24678,N_24732);
xor U25482 (N_25482,N_24801,N_24931);
or U25483 (N_25483,N_24506,N_24854);
and U25484 (N_25484,N_24989,N_24686);
nor U25485 (N_25485,N_24849,N_24699);
nor U25486 (N_25486,N_24522,N_24518);
or U25487 (N_25487,N_24888,N_24532);
or U25488 (N_25488,N_24534,N_24522);
xor U25489 (N_25489,N_24871,N_24659);
xor U25490 (N_25490,N_24554,N_24524);
nand U25491 (N_25491,N_24561,N_24667);
nor U25492 (N_25492,N_24981,N_24814);
nor U25493 (N_25493,N_24588,N_24957);
nand U25494 (N_25494,N_24963,N_24555);
nor U25495 (N_25495,N_24939,N_24638);
nor U25496 (N_25496,N_24734,N_24805);
or U25497 (N_25497,N_24641,N_24858);
nor U25498 (N_25498,N_24613,N_24825);
xnor U25499 (N_25499,N_24514,N_24818);
or U25500 (N_25500,N_25012,N_25025);
and U25501 (N_25501,N_25114,N_25305);
and U25502 (N_25502,N_25095,N_25386);
and U25503 (N_25503,N_25091,N_25082);
and U25504 (N_25504,N_25120,N_25262);
xor U25505 (N_25505,N_25182,N_25209);
or U25506 (N_25506,N_25045,N_25158);
or U25507 (N_25507,N_25469,N_25108);
nand U25508 (N_25508,N_25499,N_25018);
nor U25509 (N_25509,N_25276,N_25044);
nor U25510 (N_25510,N_25171,N_25477);
nand U25511 (N_25511,N_25401,N_25273);
nor U25512 (N_25512,N_25010,N_25349);
nand U25513 (N_25513,N_25041,N_25079);
nor U25514 (N_25514,N_25133,N_25419);
and U25515 (N_25515,N_25465,N_25433);
nand U25516 (N_25516,N_25314,N_25301);
nor U25517 (N_25517,N_25294,N_25358);
nor U25518 (N_25518,N_25284,N_25493);
nor U25519 (N_25519,N_25008,N_25255);
or U25520 (N_25520,N_25107,N_25420);
nor U25521 (N_25521,N_25020,N_25156);
or U25522 (N_25522,N_25054,N_25212);
nor U25523 (N_25523,N_25405,N_25221);
nor U25524 (N_25524,N_25444,N_25080);
nor U25525 (N_25525,N_25023,N_25462);
nand U25526 (N_25526,N_25382,N_25222);
or U25527 (N_25527,N_25103,N_25119);
nand U25528 (N_25528,N_25056,N_25085);
or U25529 (N_25529,N_25388,N_25202);
xnor U25530 (N_25530,N_25347,N_25004);
nand U25531 (N_25531,N_25352,N_25363);
and U25532 (N_25532,N_25243,N_25063);
or U25533 (N_25533,N_25105,N_25367);
and U25534 (N_25534,N_25278,N_25261);
or U25535 (N_25535,N_25205,N_25192);
nor U25536 (N_25536,N_25373,N_25092);
xor U25537 (N_25537,N_25183,N_25207);
nor U25538 (N_25538,N_25142,N_25193);
or U25539 (N_25539,N_25365,N_25001);
or U25540 (N_25540,N_25286,N_25140);
nand U25541 (N_25541,N_25005,N_25011);
nand U25542 (N_25542,N_25459,N_25332);
nand U25543 (N_25543,N_25200,N_25123);
or U25544 (N_25544,N_25225,N_25246);
or U25545 (N_25545,N_25149,N_25135);
or U25546 (N_25546,N_25344,N_25280);
xnor U25547 (N_25547,N_25293,N_25190);
and U25548 (N_25548,N_25113,N_25453);
and U25549 (N_25549,N_25152,N_25109);
nand U25550 (N_25550,N_25320,N_25403);
or U25551 (N_25551,N_25297,N_25154);
nor U25552 (N_25552,N_25498,N_25089);
xor U25553 (N_25553,N_25308,N_25351);
and U25554 (N_25554,N_25224,N_25185);
xor U25555 (N_25555,N_25300,N_25425);
xor U25556 (N_25556,N_25464,N_25307);
and U25557 (N_25557,N_25443,N_25309);
xnor U25558 (N_25558,N_25368,N_25027);
nand U25559 (N_25559,N_25125,N_25328);
and U25560 (N_25560,N_25413,N_25239);
nand U25561 (N_25561,N_25399,N_25042);
nand U25562 (N_25562,N_25093,N_25326);
nand U25563 (N_25563,N_25484,N_25483);
or U25564 (N_25564,N_25395,N_25245);
and U25565 (N_25565,N_25129,N_25478);
nor U25566 (N_25566,N_25219,N_25440);
nor U25567 (N_25567,N_25298,N_25371);
nand U25568 (N_25568,N_25227,N_25168);
nand U25569 (N_25569,N_25026,N_25260);
nor U25570 (N_25570,N_25176,N_25350);
or U25571 (N_25571,N_25069,N_25241);
nand U25572 (N_25572,N_25148,N_25354);
and U25573 (N_25573,N_25355,N_25270);
nor U25574 (N_25574,N_25177,N_25429);
or U25575 (N_25575,N_25060,N_25451);
xnor U25576 (N_25576,N_25238,N_25240);
nor U25577 (N_25577,N_25046,N_25461);
and U25578 (N_25578,N_25218,N_25242);
nor U25579 (N_25579,N_25251,N_25492);
and U25580 (N_25580,N_25009,N_25163);
nand U25581 (N_25581,N_25417,N_25311);
and U25582 (N_25582,N_25160,N_25393);
or U25583 (N_25583,N_25043,N_25104);
or U25584 (N_25584,N_25166,N_25057);
xnor U25585 (N_25585,N_25384,N_25460);
and U25586 (N_25586,N_25064,N_25488);
nor U25587 (N_25587,N_25254,N_25007);
nor U25588 (N_25588,N_25400,N_25272);
nand U25589 (N_25589,N_25283,N_25256);
xnor U25590 (N_25590,N_25128,N_25345);
or U25591 (N_25591,N_25172,N_25013);
nor U25592 (N_25592,N_25252,N_25035);
and U25593 (N_25593,N_25122,N_25189);
xnor U25594 (N_25594,N_25147,N_25017);
or U25595 (N_25595,N_25385,N_25002);
nor U25596 (N_25596,N_25333,N_25466);
xnor U25597 (N_25597,N_25145,N_25331);
or U25598 (N_25598,N_25383,N_25281);
or U25599 (N_25599,N_25100,N_25475);
nand U25600 (N_25600,N_25290,N_25141);
nand U25601 (N_25601,N_25366,N_25404);
nand U25602 (N_25602,N_25394,N_25051);
or U25603 (N_25603,N_25277,N_25235);
xor U25604 (N_25604,N_25282,N_25423);
and U25605 (N_25605,N_25445,N_25111);
xor U25606 (N_25606,N_25402,N_25426);
or U25607 (N_25607,N_25410,N_25144);
or U25608 (N_25608,N_25430,N_25310);
or U25609 (N_25609,N_25039,N_25077);
xor U25610 (N_25610,N_25428,N_25204);
or U25611 (N_25611,N_25447,N_25340);
or U25612 (N_25612,N_25237,N_25369);
and U25613 (N_25613,N_25047,N_25067);
and U25614 (N_25614,N_25438,N_25315);
xor U25615 (N_25615,N_25247,N_25132);
nor U25616 (N_25616,N_25357,N_25442);
nand U25617 (N_25617,N_25186,N_25486);
or U25618 (N_25618,N_25296,N_25397);
and U25619 (N_25619,N_25374,N_25343);
and U25620 (N_25620,N_25034,N_25415);
and U25621 (N_25621,N_25096,N_25471);
xor U25622 (N_25622,N_25101,N_25076);
nor U25623 (N_25623,N_25169,N_25361);
xnor U25624 (N_25624,N_25031,N_25329);
or U25625 (N_25625,N_25179,N_25220);
nand U25626 (N_25626,N_25234,N_25304);
xor U25627 (N_25627,N_25275,N_25303);
xnor U25628 (N_25628,N_25421,N_25263);
nand U25629 (N_25629,N_25016,N_25375);
nand U25630 (N_25630,N_25248,N_25479);
nand U25631 (N_25631,N_25407,N_25267);
xor U25632 (N_25632,N_25110,N_25233);
and U25633 (N_25633,N_25431,N_25292);
and U25634 (N_25634,N_25372,N_25159);
and U25635 (N_25635,N_25230,N_25151);
nand U25636 (N_25636,N_25086,N_25195);
or U25637 (N_25637,N_25223,N_25130);
and U25638 (N_25638,N_25161,N_25409);
and U25639 (N_25639,N_25335,N_25019);
and U25640 (N_25640,N_25143,N_25482);
and U25641 (N_25641,N_25274,N_25138);
nor U25642 (N_25642,N_25115,N_25131);
xor U25643 (N_25643,N_25434,N_25253);
nand U25644 (N_25644,N_25124,N_25049);
and U25645 (N_25645,N_25491,N_25066);
and U25646 (N_25646,N_25048,N_25055);
or U25647 (N_25647,N_25319,N_25106);
xor U25648 (N_25648,N_25061,N_25435);
and U25649 (N_25649,N_25370,N_25380);
and U25650 (N_25650,N_25032,N_25037);
and U25651 (N_25651,N_25287,N_25487);
nor U25652 (N_25652,N_25244,N_25436);
nor U25653 (N_25653,N_25422,N_25083);
or U25654 (N_25654,N_25029,N_25208);
nand U25655 (N_25655,N_25336,N_25014);
or U25656 (N_25656,N_25452,N_25181);
and U25657 (N_25657,N_25164,N_25213);
nand U25658 (N_25658,N_25053,N_25050);
xnor U25659 (N_25659,N_25389,N_25090);
nand U25660 (N_25660,N_25424,N_25341);
nand U25661 (N_25661,N_25153,N_25289);
and U25662 (N_25662,N_25325,N_25059);
and U25663 (N_25663,N_25097,N_25199);
xor U25664 (N_25664,N_25338,N_25454);
and U25665 (N_25665,N_25450,N_25150);
and U25666 (N_25666,N_25075,N_25188);
nand U25667 (N_25667,N_25302,N_25494);
and U25668 (N_25668,N_25265,N_25228);
or U25669 (N_25669,N_25117,N_25021);
xnor U25670 (N_25670,N_25448,N_25006);
and U25671 (N_25671,N_25036,N_25378);
and U25672 (N_25672,N_25362,N_25216);
nand U25673 (N_25673,N_25157,N_25206);
nand U25674 (N_25674,N_25446,N_25194);
nor U25675 (N_25675,N_25364,N_25467);
and U25676 (N_25676,N_25078,N_25203);
or U25677 (N_25677,N_25285,N_25330);
nor U25678 (N_25678,N_25268,N_25264);
or U25679 (N_25679,N_25348,N_25327);
xor U25680 (N_25680,N_25271,N_25071);
xor U25681 (N_25681,N_25196,N_25170);
xnor U25682 (N_25682,N_25377,N_25102);
nand U25683 (N_25683,N_25038,N_25088);
nand U25684 (N_25684,N_25392,N_25187);
nand U25685 (N_25685,N_25481,N_25058);
nand U25686 (N_25686,N_25458,N_25198);
and U25687 (N_25687,N_25473,N_25406);
or U25688 (N_25688,N_25342,N_25000);
or U25689 (N_25689,N_25455,N_25210);
or U25690 (N_25690,N_25353,N_25229);
xor U25691 (N_25691,N_25441,N_25312);
and U25692 (N_25692,N_25266,N_25074);
xor U25693 (N_25693,N_25184,N_25250);
nor U25694 (N_25694,N_25288,N_25073);
and U25695 (N_25695,N_25098,N_25418);
and U25696 (N_25696,N_25360,N_25359);
and U25697 (N_25697,N_25191,N_25211);
nand U25698 (N_25698,N_25249,N_25313);
or U25699 (N_25699,N_25231,N_25356);
or U25700 (N_25700,N_25062,N_25180);
nor U25701 (N_25701,N_25173,N_25391);
and U25702 (N_25702,N_25379,N_25121);
xnor U25703 (N_25703,N_25236,N_25087);
and U25704 (N_25704,N_25390,N_25449);
nor U25705 (N_25705,N_25306,N_25259);
xor U25706 (N_25706,N_25174,N_25099);
xor U25707 (N_25707,N_25197,N_25030);
nand U25708 (N_25708,N_25334,N_25028);
or U25709 (N_25709,N_25472,N_25068);
and U25710 (N_25710,N_25457,N_25416);
xor U25711 (N_25711,N_25411,N_25497);
nand U25712 (N_25712,N_25490,N_25162);
xnor U25713 (N_25713,N_25201,N_25412);
and U25714 (N_25714,N_25094,N_25474);
xnor U25715 (N_25715,N_25072,N_25127);
or U25716 (N_25716,N_25414,N_25258);
nor U25717 (N_25717,N_25387,N_25084);
xnor U25718 (N_25718,N_25065,N_25024);
xnor U25719 (N_25719,N_25485,N_25337);
xnor U25720 (N_25720,N_25324,N_25316);
nand U25721 (N_25721,N_25480,N_25015);
xor U25722 (N_25722,N_25476,N_25022);
nand U25723 (N_25723,N_25033,N_25439);
xor U25724 (N_25724,N_25214,N_25217);
nand U25725 (N_25725,N_25322,N_25295);
nand U25726 (N_25726,N_25139,N_25134);
nor U25727 (N_25727,N_25321,N_25470);
nand U25728 (N_25728,N_25081,N_25175);
and U25729 (N_25729,N_25126,N_25112);
nor U25730 (N_25730,N_25003,N_25489);
nor U25731 (N_25731,N_25437,N_25070);
xnor U25732 (N_25732,N_25323,N_25040);
nand U25733 (N_25733,N_25215,N_25456);
nor U25734 (N_25734,N_25116,N_25165);
or U25735 (N_25735,N_25137,N_25317);
and U25736 (N_25736,N_25291,N_25167);
nand U25737 (N_25737,N_25146,N_25463);
or U25738 (N_25738,N_25346,N_25381);
nor U25739 (N_25739,N_25432,N_25408);
and U25740 (N_25740,N_25468,N_25257);
xor U25741 (N_25741,N_25427,N_25279);
nor U25742 (N_25742,N_25118,N_25052);
and U25743 (N_25743,N_25299,N_25398);
nand U25744 (N_25744,N_25376,N_25232);
nor U25745 (N_25745,N_25269,N_25495);
nor U25746 (N_25746,N_25178,N_25226);
or U25747 (N_25747,N_25318,N_25136);
or U25748 (N_25748,N_25339,N_25155);
or U25749 (N_25749,N_25496,N_25396);
nand U25750 (N_25750,N_25137,N_25441);
and U25751 (N_25751,N_25366,N_25069);
nand U25752 (N_25752,N_25298,N_25440);
and U25753 (N_25753,N_25445,N_25275);
nand U25754 (N_25754,N_25232,N_25093);
nor U25755 (N_25755,N_25407,N_25198);
xnor U25756 (N_25756,N_25478,N_25409);
or U25757 (N_25757,N_25065,N_25117);
nand U25758 (N_25758,N_25370,N_25126);
nor U25759 (N_25759,N_25203,N_25480);
nor U25760 (N_25760,N_25360,N_25027);
nand U25761 (N_25761,N_25163,N_25477);
nor U25762 (N_25762,N_25285,N_25020);
and U25763 (N_25763,N_25280,N_25357);
and U25764 (N_25764,N_25044,N_25098);
or U25765 (N_25765,N_25127,N_25312);
nor U25766 (N_25766,N_25310,N_25317);
and U25767 (N_25767,N_25434,N_25431);
or U25768 (N_25768,N_25143,N_25322);
and U25769 (N_25769,N_25004,N_25337);
or U25770 (N_25770,N_25361,N_25232);
nand U25771 (N_25771,N_25055,N_25178);
or U25772 (N_25772,N_25320,N_25296);
xnor U25773 (N_25773,N_25239,N_25185);
and U25774 (N_25774,N_25439,N_25434);
and U25775 (N_25775,N_25414,N_25059);
xnor U25776 (N_25776,N_25114,N_25112);
nor U25777 (N_25777,N_25189,N_25401);
or U25778 (N_25778,N_25499,N_25253);
xnor U25779 (N_25779,N_25357,N_25413);
nand U25780 (N_25780,N_25317,N_25067);
nor U25781 (N_25781,N_25084,N_25487);
xnor U25782 (N_25782,N_25409,N_25343);
or U25783 (N_25783,N_25083,N_25030);
xnor U25784 (N_25784,N_25051,N_25407);
nand U25785 (N_25785,N_25384,N_25452);
xor U25786 (N_25786,N_25460,N_25078);
xnor U25787 (N_25787,N_25322,N_25481);
nand U25788 (N_25788,N_25295,N_25172);
and U25789 (N_25789,N_25190,N_25284);
nand U25790 (N_25790,N_25292,N_25007);
nor U25791 (N_25791,N_25114,N_25302);
xnor U25792 (N_25792,N_25457,N_25058);
nor U25793 (N_25793,N_25040,N_25157);
xor U25794 (N_25794,N_25054,N_25281);
or U25795 (N_25795,N_25010,N_25343);
xor U25796 (N_25796,N_25413,N_25341);
or U25797 (N_25797,N_25026,N_25484);
and U25798 (N_25798,N_25276,N_25343);
nor U25799 (N_25799,N_25424,N_25269);
or U25800 (N_25800,N_25042,N_25176);
xnor U25801 (N_25801,N_25047,N_25377);
or U25802 (N_25802,N_25323,N_25436);
and U25803 (N_25803,N_25348,N_25118);
nor U25804 (N_25804,N_25459,N_25231);
nand U25805 (N_25805,N_25059,N_25256);
or U25806 (N_25806,N_25098,N_25107);
and U25807 (N_25807,N_25093,N_25223);
or U25808 (N_25808,N_25498,N_25079);
and U25809 (N_25809,N_25380,N_25009);
nand U25810 (N_25810,N_25160,N_25436);
or U25811 (N_25811,N_25436,N_25235);
or U25812 (N_25812,N_25319,N_25181);
nand U25813 (N_25813,N_25069,N_25268);
nor U25814 (N_25814,N_25048,N_25206);
and U25815 (N_25815,N_25131,N_25429);
and U25816 (N_25816,N_25170,N_25306);
nand U25817 (N_25817,N_25269,N_25036);
and U25818 (N_25818,N_25430,N_25268);
nor U25819 (N_25819,N_25174,N_25091);
nand U25820 (N_25820,N_25315,N_25044);
and U25821 (N_25821,N_25395,N_25110);
nor U25822 (N_25822,N_25236,N_25283);
xnor U25823 (N_25823,N_25158,N_25263);
and U25824 (N_25824,N_25406,N_25128);
or U25825 (N_25825,N_25042,N_25132);
nand U25826 (N_25826,N_25233,N_25115);
and U25827 (N_25827,N_25083,N_25130);
xor U25828 (N_25828,N_25036,N_25258);
nor U25829 (N_25829,N_25099,N_25262);
xnor U25830 (N_25830,N_25485,N_25403);
nand U25831 (N_25831,N_25097,N_25049);
nor U25832 (N_25832,N_25087,N_25431);
or U25833 (N_25833,N_25090,N_25121);
xor U25834 (N_25834,N_25472,N_25058);
or U25835 (N_25835,N_25422,N_25148);
nand U25836 (N_25836,N_25015,N_25350);
and U25837 (N_25837,N_25141,N_25176);
and U25838 (N_25838,N_25284,N_25332);
nand U25839 (N_25839,N_25297,N_25398);
nand U25840 (N_25840,N_25283,N_25223);
nand U25841 (N_25841,N_25018,N_25359);
nor U25842 (N_25842,N_25289,N_25052);
and U25843 (N_25843,N_25141,N_25085);
or U25844 (N_25844,N_25186,N_25461);
and U25845 (N_25845,N_25235,N_25288);
nand U25846 (N_25846,N_25183,N_25271);
or U25847 (N_25847,N_25277,N_25411);
xor U25848 (N_25848,N_25485,N_25449);
and U25849 (N_25849,N_25125,N_25302);
nand U25850 (N_25850,N_25420,N_25379);
nor U25851 (N_25851,N_25016,N_25022);
nor U25852 (N_25852,N_25010,N_25357);
nand U25853 (N_25853,N_25398,N_25350);
or U25854 (N_25854,N_25354,N_25142);
and U25855 (N_25855,N_25384,N_25224);
xnor U25856 (N_25856,N_25275,N_25465);
and U25857 (N_25857,N_25456,N_25461);
or U25858 (N_25858,N_25033,N_25180);
xor U25859 (N_25859,N_25427,N_25321);
and U25860 (N_25860,N_25439,N_25374);
nand U25861 (N_25861,N_25092,N_25170);
or U25862 (N_25862,N_25076,N_25295);
nor U25863 (N_25863,N_25221,N_25363);
nor U25864 (N_25864,N_25119,N_25284);
nand U25865 (N_25865,N_25342,N_25201);
and U25866 (N_25866,N_25089,N_25443);
or U25867 (N_25867,N_25468,N_25018);
nor U25868 (N_25868,N_25160,N_25227);
nor U25869 (N_25869,N_25255,N_25232);
nor U25870 (N_25870,N_25283,N_25341);
and U25871 (N_25871,N_25038,N_25106);
or U25872 (N_25872,N_25013,N_25005);
and U25873 (N_25873,N_25127,N_25275);
and U25874 (N_25874,N_25075,N_25325);
nand U25875 (N_25875,N_25060,N_25033);
nand U25876 (N_25876,N_25419,N_25000);
nor U25877 (N_25877,N_25128,N_25170);
nand U25878 (N_25878,N_25345,N_25047);
or U25879 (N_25879,N_25186,N_25455);
nor U25880 (N_25880,N_25375,N_25065);
and U25881 (N_25881,N_25432,N_25087);
nand U25882 (N_25882,N_25047,N_25098);
xnor U25883 (N_25883,N_25444,N_25430);
and U25884 (N_25884,N_25007,N_25366);
nor U25885 (N_25885,N_25053,N_25387);
nand U25886 (N_25886,N_25087,N_25294);
and U25887 (N_25887,N_25288,N_25051);
or U25888 (N_25888,N_25481,N_25347);
or U25889 (N_25889,N_25192,N_25225);
xnor U25890 (N_25890,N_25156,N_25499);
nor U25891 (N_25891,N_25425,N_25330);
xnor U25892 (N_25892,N_25422,N_25190);
xor U25893 (N_25893,N_25373,N_25185);
and U25894 (N_25894,N_25204,N_25437);
nor U25895 (N_25895,N_25023,N_25078);
nor U25896 (N_25896,N_25400,N_25111);
xor U25897 (N_25897,N_25060,N_25223);
or U25898 (N_25898,N_25317,N_25209);
and U25899 (N_25899,N_25321,N_25011);
and U25900 (N_25900,N_25109,N_25198);
xor U25901 (N_25901,N_25080,N_25103);
or U25902 (N_25902,N_25021,N_25189);
xnor U25903 (N_25903,N_25093,N_25487);
nor U25904 (N_25904,N_25315,N_25296);
nor U25905 (N_25905,N_25206,N_25210);
nand U25906 (N_25906,N_25291,N_25300);
nor U25907 (N_25907,N_25335,N_25264);
and U25908 (N_25908,N_25179,N_25452);
xnor U25909 (N_25909,N_25288,N_25216);
nor U25910 (N_25910,N_25464,N_25181);
or U25911 (N_25911,N_25417,N_25328);
nand U25912 (N_25912,N_25051,N_25417);
nand U25913 (N_25913,N_25279,N_25454);
or U25914 (N_25914,N_25101,N_25184);
or U25915 (N_25915,N_25348,N_25259);
nand U25916 (N_25916,N_25312,N_25023);
xnor U25917 (N_25917,N_25467,N_25307);
nand U25918 (N_25918,N_25209,N_25223);
nand U25919 (N_25919,N_25249,N_25457);
and U25920 (N_25920,N_25037,N_25330);
nor U25921 (N_25921,N_25191,N_25226);
nor U25922 (N_25922,N_25016,N_25056);
and U25923 (N_25923,N_25054,N_25430);
nor U25924 (N_25924,N_25377,N_25116);
nor U25925 (N_25925,N_25026,N_25412);
nor U25926 (N_25926,N_25428,N_25367);
nand U25927 (N_25927,N_25106,N_25142);
or U25928 (N_25928,N_25109,N_25352);
nor U25929 (N_25929,N_25281,N_25415);
xnor U25930 (N_25930,N_25172,N_25307);
or U25931 (N_25931,N_25313,N_25316);
xnor U25932 (N_25932,N_25254,N_25306);
and U25933 (N_25933,N_25008,N_25038);
xnor U25934 (N_25934,N_25472,N_25142);
xor U25935 (N_25935,N_25121,N_25208);
xor U25936 (N_25936,N_25346,N_25111);
nor U25937 (N_25937,N_25476,N_25079);
nor U25938 (N_25938,N_25141,N_25054);
or U25939 (N_25939,N_25086,N_25456);
nor U25940 (N_25940,N_25262,N_25397);
or U25941 (N_25941,N_25400,N_25093);
and U25942 (N_25942,N_25318,N_25416);
or U25943 (N_25943,N_25221,N_25222);
or U25944 (N_25944,N_25000,N_25132);
nand U25945 (N_25945,N_25499,N_25239);
nand U25946 (N_25946,N_25337,N_25259);
and U25947 (N_25947,N_25391,N_25443);
nand U25948 (N_25948,N_25140,N_25087);
or U25949 (N_25949,N_25258,N_25353);
and U25950 (N_25950,N_25420,N_25476);
or U25951 (N_25951,N_25449,N_25436);
xor U25952 (N_25952,N_25389,N_25061);
nand U25953 (N_25953,N_25132,N_25307);
nand U25954 (N_25954,N_25296,N_25091);
nand U25955 (N_25955,N_25473,N_25462);
or U25956 (N_25956,N_25016,N_25036);
xor U25957 (N_25957,N_25364,N_25292);
nand U25958 (N_25958,N_25349,N_25340);
xnor U25959 (N_25959,N_25257,N_25102);
or U25960 (N_25960,N_25052,N_25022);
nor U25961 (N_25961,N_25147,N_25065);
nand U25962 (N_25962,N_25468,N_25469);
and U25963 (N_25963,N_25253,N_25323);
or U25964 (N_25964,N_25432,N_25411);
nand U25965 (N_25965,N_25163,N_25231);
nor U25966 (N_25966,N_25473,N_25222);
xor U25967 (N_25967,N_25115,N_25469);
xnor U25968 (N_25968,N_25299,N_25283);
nor U25969 (N_25969,N_25324,N_25200);
nor U25970 (N_25970,N_25315,N_25415);
xnor U25971 (N_25971,N_25412,N_25317);
nand U25972 (N_25972,N_25242,N_25013);
xnor U25973 (N_25973,N_25457,N_25011);
or U25974 (N_25974,N_25430,N_25415);
nor U25975 (N_25975,N_25426,N_25100);
xnor U25976 (N_25976,N_25269,N_25391);
xor U25977 (N_25977,N_25472,N_25097);
and U25978 (N_25978,N_25395,N_25290);
or U25979 (N_25979,N_25199,N_25378);
nand U25980 (N_25980,N_25008,N_25045);
nand U25981 (N_25981,N_25348,N_25046);
nand U25982 (N_25982,N_25115,N_25130);
nor U25983 (N_25983,N_25060,N_25164);
and U25984 (N_25984,N_25128,N_25094);
and U25985 (N_25985,N_25210,N_25329);
nor U25986 (N_25986,N_25020,N_25420);
and U25987 (N_25987,N_25110,N_25010);
nor U25988 (N_25988,N_25430,N_25495);
or U25989 (N_25989,N_25188,N_25460);
nor U25990 (N_25990,N_25498,N_25343);
xor U25991 (N_25991,N_25458,N_25081);
xor U25992 (N_25992,N_25185,N_25270);
nand U25993 (N_25993,N_25032,N_25370);
nor U25994 (N_25994,N_25197,N_25187);
xor U25995 (N_25995,N_25309,N_25372);
nand U25996 (N_25996,N_25296,N_25476);
xor U25997 (N_25997,N_25073,N_25168);
xor U25998 (N_25998,N_25111,N_25481);
and U25999 (N_25999,N_25362,N_25307);
or U26000 (N_26000,N_25689,N_25946);
nand U26001 (N_26001,N_25875,N_25986);
or U26002 (N_26002,N_25863,N_25751);
or U26003 (N_26003,N_25865,N_25830);
xor U26004 (N_26004,N_25658,N_25614);
and U26005 (N_26005,N_25980,N_25564);
xnor U26006 (N_26006,N_25697,N_25687);
xnor U26007 (N_26007,N_25522,N_25790);
and U26008 (N_26008,N_25671,N_25638);
nand U26009 (N_26009,N_25855,N_25909);
xor U26010 (N_26010,N_25698,N_25512);
and U26011 (N_26011,N_25926,N_25668);
nand U26012 (N_26012,N_25913,N_25539);
and U26013 (N_26013,N_25623,N_25703);
or U26014 (N_26014,N_25730,N_25930);
xnor U26015 (N_26015,N_25905,N_25544);
xor U26016 (N_26016,N_25916,N_25938);
xor U26017 (N_26017,N_25919,N_25872);
xnor U26018 (N_26018,N_25957,N_25890);
and U26019 (N_26019,N_25871,N_25887);
nand U26020 (N_26020,N_25649,N_25620);
xor U26021 (N_26021,N_25610,N_25768);
xnor U26022 (N_26022,N_25766,N_25604);
xor U26023 (N_26023,N_25551,N_25912);
xor U26024 (N_26024,N_25633,N_25888);
or U26025 (N_26025,N_25534,N_25677);
nor U26026 (N_26026,N_25796,N_25617);
nand U26027 (N_26027,N_25991,N_25673);
or U26028 (N_26028,N_25669,N_25883);
nand U26029 (N_26029,N_25867,N_25805);
or U26030 (N_26030,N_25793,N_25982);
and U26031 (N_26031,N_25842,N_25981);
nand U26032 (N_26032,N_25901,N_25914);
nor U26033 (N_26033,N_25779,N_25941);
or U26034 (N_26034,N_25840,N_25533);
or U26035 (N_26035,N_25932,N_25776);
or U26036 (N_26036,N_25624,N_25993);
and U26037 (N_26037,N_25746,N_25627);
nand U26038 (N_26038,N_25903,N_25688);
nor U26039 (N_26039,N_25802,N_25812);
nand U26040 (N_26040,N_25613,N_25744);
and U26041 (N_26041,N_25813,N_25977);
and U26042 (N_26042,N_25970,N_25950);
xor U26043 (N_26043,N_25723,N_25735);
or U26044 (N_26044,N_25920,N_25552);
nor U26045 (N_26045,N_25657,N_25710);
xor U26046 (N_26046,N_25737,N_25788);
nand U26047 (N_26047,N_25729,N_25794);
nand U26048 (N_26048,N_25721,N_25515);
or U26049 (N_26049,N_25876,N_25739);
nand U26050 (N_26050,N_25715,N_25672);
nor U26051 (N_26051,N_25616,N_25750);
nand U26052 (N_26052,N_25720,N_25741);
or U26053 (N_26053,N_25956,N_25811);
and U26054 (N_26054,N_25814,N_25700);
nand U26055 (N_26055,N_25719,N_25954);
nor U26056 (N_26056,N_25806,N_25860);
xor U26057 (N_26057,N_25690,N_25763);
nand U26058 (N_26058,N_25747,N_25716);
nor U26059 (N_26059,N_25877,N_25847);
and U26060 (N_26060,N_25824,N_25749);
xor U26061 (N_26061,N_25635,N_25984);
nand U26062 (N_26062,N_25583,N_25574);
nor U26063 (N_26063,N_25519,N_25661);
xnor U26064 (N_26064,N_25902,N_25569);
or U26065 (N_26065,N_25546,N_25791);
or U26066 (N_26066,N_25857,N_25611);
or U26067 (N_26067,N_25797,N_25820);
nor U26068 (N_26068,N_25645,N_25590);
nand U26069 (N_26069,N_25765,N_25640);
or U26070 (N_26070,N_25896,N_25622);
xor U26071 (N_26071,N_25892,N_25667);
xor U26072 (N_26072,N_25540,N_25670);
or U26073 (N_26073,N_25935,N_25816);
and U26074 (N_26074,N_25898,N_25618);
xor U26075 (N_26075,N_25608,N_25748);
or U26076 (N_26076,N_25844,N_25997);
xnor U26077 (N_26077,N_25528,N_25940);
xor U26078 (N_26078,N_25740,N_25949);
or U26079 (N_26079,N_25761,N_25808);
and U26080 (N_26080,N_25800,N_25769);
or U26081 (N_26081,N_25778,N_25502);
nand U26082 (N_26082,N_25937,N_25714);
nor U26083 (N_26083,N_25771,N_25680);
or U26084 (N_26084,N_25835,N_25702);
xnor U26085 (N_26085,N_25707,N_25849);
and U26086 (N_26086,N_25725,N_25848);
xnor U26087 (N_26087,N_25738,N_25567);
or U26088 (N_26088,N_25626,N_25566);
and U26089 (N_26089,N_25555,N_25885);
xor U26090 (N_26090,N_25939,N_25577);
nor U26091 (N_26091,N_25724,N_25601);
or U26092 (N_26092,N_25647,N_25757);
xnor U26093 (N_26093,N_25979,N_25520);
nand U26094 (N_26094,N_25833,N_25609);
nor U26095 (N_26095,N_25948,N_25807);
nor U26096 (N_26096,N_25642,N_25530);
xnor U26097 (N_26097,N_25782,N_25581);
or U26098 (N_26098,N_25952,N_25600);
nand U26099 (N_26099,N_25582,N_25631);
and U26100 (N_26100,N_25586,N_25643);
or U26101 (N_26101,N_25679,N_25545);
xnor U26102 (N_26102,N_25910,N_25861);
and U26103 (N_26103,N_25728,N_25535);
xor U26104 (N_26104,N_25942,N_25795);
xor U26105 (N_26105,N_25711,N_25928);
and U26106 (N_26106,N_25968,N_25961);
nor U26107 (N_26107,N_25962,N_25850);
xnor U26108 (N_26108,N_25606,N_25506);
nor U26109 (N_26109,N_25879,N_25509);
nand U26110 (N_26110,N_25559,N_25517);
and U26111 (N_26111,N_25696,N_25557);
xnor U26112 (N_26112,N_25742,N_25595);
nand U26113 (N_26113,N_25588,N_25501);
nor U26114 (N_26114,N_25662,N_25708);
xor U26115 (N_26115,N_25996,N_25911);
nor U26116 (N_26116,N_25676,N_25718);
or U26117 (N_26117,N_25500,N_25615);
and U26118 (N_26118,N_25752,N_25770);
xor U26119 (N_26119,N_25918,N_25641);
and U26120 (N_26120,N_25925,N_25584);
nor U26121 (N_26121,N_25674,N_25634);
xor U26122 (N_26122,N_25958,N_25505);
or U26123 (N_26123,N_25599,N_25934);
xor U26124 (N_26124,N_25554,N_25772);
nor U26125 (N_26125,N_25691,N_25894);
xnor U26126 (N_26126,N_25525,N_25831);
or U26127 (N_26127,N_25541,N_25666);
and U26128 (N_26128,N_25607,N_25862);
nor U26129 (N_26129,N_25924,N_25699);
nand U26130 (N_26130,N_25843,N_25637);
or U26131 (N_26131,N_25834,N_25683);
xnor U26132 (N_26132,N_25960,N_25503);
nand U26133 (N_26133,N_25838,N_25644);
nand U26134 (N_26134,N_25931,N_25989);
or U26135 (N_26135,N_25787,N_25514);
and U26136 (N_26136,N_25775,N_25823);
and U26137 (N_26137,N_25851,N_25784);
nor U26138 (N_26138,N_25602,N_25652);
nand U26139 (N_26139,N_25895,N_25598);
and U26140 (N_26140,N_25976,N_25908);
and U26141 (N_26141,N_25945,N_25929);
nand U26142 (N_26142,N_25891,N_25659);
xnor U26143 (N_26143,N_25999,N_25656);
nor U26144 (N_26144,N_25510,N_25783);
nand U26145 (N_26145,N_25759,N_25755);
or U26146 (N_26146,N_25907,N_25992);
or U26147 (N_26147,N_25731,N_25648);
or U26148 (N_26148,N_25704,N_25774);
nor U26149 (N_26149,N_25636,N_25874);
nand U26150 (N_26150,N_25837,N_25578);
xor U26151 (N_26151,N_25511,N_25563);
nand U26152 (N_26152,N_25560,N_25959);
nand U26153 (N_26153,N_25589,N_25536);
nand U26154 (N_26154,N_25754,N_25821);
nor U26155 (N_26155,N_25936,N_25665);
nor U26156 (N_26156,N_25504,N_25605);
nor U26157 (N_26157,N_25568,N_25592);
or U26158 (N_26158,N_25839,N_25786);
or U26159 (N_26159,N_25818,N_25974);
and U26160 (N_26160,N_25734,N_25694);
and U26161 (N_26161,N_25881,N_25596);
or U26162 (N_26162,N_25869,N_25884);
or U26163 (N_26163,N_25693,N_25518);
or U26164 (N_26164,N_25927,N_25587);
and U26165 (N_26165,N_25998,N_25822);
nand U26166 (N_26166,N_25827,N_25651);
nand U26167 (N_26167,N_25864,N_25653);
nand U26168 (N_26168,N_25966,N_25985);
xnor U26169 (N_26169,N_25915,N_25889);
nor U26170 (N_26170,N_25675,N_25801);
and U26171 (N_26171,N_25899,N_25681);
xor U26172 (N_26172,N_25994,N_25706);
or U26173 (N_26173,N_25819,N_25900);
nor U26174 (N_26174,N_25524,N_25870);
and U26175 (N_26175,N_25995,N_25523);
nand U26176 (N_26176,N_25701,N_25619);
and U26177 (N_26177,N_25969,N_25799);
nand U26178 (N_26178,N_25580,N_25743);
or U26179 (N_26179,N_25785,N_25562);
xnor U26180 (N_26180,N_25859,N_25953);
and U26181 (N_26181,N_25829,N_25815);
or U26182 (N_26182,N_25964,N_25955);
xor U26183 (N_26183,N_25603,N_25709);
nor U26184 (N_26184,N_25712,N_25886);
xnor U26185 (N_26185,N_25527,N_25722);
or U26186 (N_26186,N_25921,N_25682);
nand U26187 (N_26187,N_25650,N_25753);
nand U26188 (N_26188,N_25917,N_25856);
and U26189 (N_26189,N_25508,N_25943);
nor U26190 (N_26190,N_25773,N_25978);
nor U26191 (N_26191,N_25972,N_25570);
xor U26192 (N_26192,N_25556,N_25858);
nor U26193 (N_26193,N_25591,N_25764);
nor U26194 (N_26194,N_25561,N_25573);
xor U26195 (N_26195,N_25780,N_25987);
nand U26196 (N_26196,N_25678,N_25893);
nor U26197 (N_26197,N_25542,N_25758);
and U26198 (N_26198,N_25558,N_25904);
or U26199 (N_26199,N_25663,N_25594);
and U26200 (N_26200,N_25922,N_25548);
nand U26201 (N_26201,N_25951,N_25836);
or U26202 (N_26202,N_25507,N_25726);
xnor U26203 (N_26203,N_25695,N_25947);
xnor U26204 (N_26204,N_25629,N_25736);
and U26205 (N_26205,N_25628,N_25803);
or U26206 (N_26206,N_25792,N_25762);
nor U26207 (N_26207,N_25732,N_25537);
nor U26208 (N_26208,N_25593,N_25878);
or U26209 (N_26209,N_25575,N_25630);
nand U26210 (N_26210,N_25828,N_25990);
nor U26211 (N_26211,N_25897,N_25717);
xnor U26212 (N_26212,N_25692,N_25809);
nor U26213 (N_26213,N_25852,N_25646);
nor U26214 (N_26214,N_25550,N_25971);
and U26215 (N_26215,N_25933,N_25906);
xor U26216 (N_26216,N_25845,N_25713);
and U26217 (N_26217,N_25767,N_25781);
or U26218 (N_26218,N_25868,N_25549);
and U26219 (N_26219,N_25854,N_25685);
nand U26220 (N_26220,N_25882,N_25846);
and U26221 (N_26221,N_25654,N_25543);
nand U26222 (N_26222,N_25553,N_25866);
or U26223 (N_26223,N_25547,N_25516);
or U26224 (N_26224,N_25621,N_25853);
nor U26225 (N_26225,N_25789,N_25756);
nand U26226 (N_26226,N_25576,N_25810);
or U26227 (N_26227,N_25684,N_25571);
and U26228 (N_26228,N_25612,N_25973);
and U26229 (N_26229,N_25880,N_25825);
nor U26230 (N_26230,N_25526,N_25975);
and U26231 (N_26231,N_25963,N_25760);
nor U26232 (N_26232,N_25529,N_25513);
nand U26233 (N_26233,N_25639,N_25983);
nor U26234 (N_26234,N_25826,N_25625);
nor U26235 (N_26235,N_25632,N_25832);
or U26236 (N_26236,N_25705,N_25841);
nand U26237 (N_26237,N_25579,N_25873);
or U26238 (N_26238,N_25727,N_25745);
nor U26239 (N_26239,N_25655,N_25817);
xnor U26240 (N_26240,N_25585,N_25988);
nor U26241 (N_26241,N_25538,N_25660);
nand U26242 (N_26242,N_25686,N_25965);
nand U26243 (N_26243,N_25923,N_25521);
nand U26244 (N_26244,N_25967,N_25733);
nor U26245 (N_26245,N_25804,N_25664);
nand U26246 (N_26246,N_25565,N_25944);
xor U26247 (N_26247,N_25597,N_25798);
or U26248 (N_26248,N_25532,N_25531);
xor U26249 (N_26249,N_25572,N_25777);
nand U26250 (N_26250,N_25905,N_25552);
nand U26251 (N_26251,N_25578,N_25698);
nand U26252 (N_26252,N_25560,N_25794);
xor U26253 (N_26253,N_25751,N_25657);
xnor U26254 (N_26254,N_25501,N_25991);
and U26255 (N_26255,N_25554,N_25820);
xor U26256 (N_26256,N_25926,N_25652);
or U26257 (N_26257,N_25727,N_25827);
xor U26258 (N_26258,N_25962,N_25700);
xor U26259 (N_26259,N_25847,N_25811);
and U26260 (N_26260,N_25628,N_25608);
xnor U26261 (N_26261,N_25587,N_25919);
and U26262 (N_26262,N_25878,N_25883);
xnor U26263 (N_26263,N_25931,N_25709);
nor U26264 (N_26264,N_25902,N_25671);
nand U26265 (N_26265,N_25970,N_25546);
nor U26266 (N_26266,N_25864,N_25822);
or U26267 (N_26267,N_25869,N_25563);
nand U26268 (N_26268,N_25852,N_25844);
and U26269 (N_26269,N_25744,N_25562);
xor U26270 (N_26270,N_25805,N_25654);
xnor U26271 (N_26271,N_25916,N_25771);
nand U26272 (N_26272,N_25902,N_25851);
xnor U26273 (N_26273,N_25738,N_25928);
and U26274 (N_26274,N_25608,N_25862);
and U26275 (N_26275,N_25853,N_25647);
and U26276 (N_26276,N_25917,N_25711);
nand U26277 (N_26277,N_25985,N_25790);
or U26278 (N_26278,N_25687,N_25772);
and U26279 (N_26279,N_25810,N_25901);
and U26280 (N_26280,N_25604,N_25942);
nand U26281 (N_26281,N_25629,N_25767);
nand U26282 (N_26282,N_25765,N_25961);
nand U26283 (N_26283,N_25611,N_25626);
and U26284 (N_26284,N_25846,N_25962);
and U26285 (N_26285,N_25581,N_25771);
and U26286 (N_26286,N_25595,N_25578);
xor U26287 (N_26287,N_25942,N_25997);
nand U26288 (N_26288,N_25975,N_25694);
nand U26289 (N_26289,N_25723,N_25960);
nand U26290 (N_26290,N_25586,N_25940);
nand U26291 (N_26291,N_25761,N_25803);
xnor U26292 (N_26292,N_25578,N_25536);
or U26293 (N_26293,N_25915,N_25526);
xor U26294 (N_26294,N_25797,N_25867);
and U26295 (N_26295,N_25571,N_25774);
nor U26296 (N_26296,N_25644,N_25758);
nand U26297 (N_26297,N_25718,N_25827);
nor U26298 (N_26298,N_25586,N_25946);
or U26299 (N_26299,N_25563,N_25639);
and U26300 (N_26300,N_25648,N_25857);
xor U26301 (N_26301,N_25662,N_25527);
and U26302 (N_26302,N_25980,N_25539);
xnor U26303 (N_26303,N_25558,N_25659);
xor U26304 (N_26304,N_25692,N_25604);
and U26305 (N_26305,N_25866,N_25710);
and U26306 (N_26306,N_25612,N_25538);
nand U26307 (N_26307,N_25526,N_25533);
nor U26308 (N_26308,N_25662,N_25561);
nand U26309 (N_26309,N_25742,N_25717);
nor U26310 (N_26310,N_25923,N_25856);
nor U26311 (N_26311,N_25952,N_25993);
or U26312 (N_26312,N_25730,N_25707);
xnor U26313 (N_26313,N_25838,N_25797);
or U26314 (N_26314,N_25820,N_25629);
and U26315 (N_26315,N_25864,N_25967);
nor U26316 (N_26316,N_25803,N_25554);
nand U26317 (N_26317,N_25847,N_25780);
nand U26318 (N_26318,N_25505,N_25655);
nor U26319 (N_26319,N_25625,N_25599);
and U26320 (N_26320,N_25956,N_25759);
or U26321 (N_26321,N_25531,N_25815);
nor U26322 (N_26322,N_25763,N_25792);
xor U26323 (N_26323,N_25746,N_25593);
nor U26324 (N_26324,N_25946,N_25637);
nand U26325 (N_26325,N_25998,N_25611);
and U26326 (N_26326,N_25717,N_25782);
xor U26327 (N_26327,N_25662,N_25939);
nand U26328 (N_26328,N_25771,N_25694);
nor U26329 (N_26329,N_25935,N_25653);
nor U26330 (N_26330,N_25726,N_25551);
and U26331 (N_26331,N_25883,N_25722);
nor U26332 (N_26332,N_25691,N_25718);
nor U26333 (N_26333,N_25830,N_25570);
nand U26334 (N_26334,N_25541,N_25740);
nand U26335 (N_26335,N_25839,N_25726);
nor U26336 (N_26336,N_25817,N_25594);
and U26337 (N_26337,N_25713,N_25694);
nor U26338 (N_26338,N_25857,N_25570);
nor U26339 (N_26339,N_25955,N_25515);
nor U26340 (N_26340,N_25963,N_25905);
and U26341 (N_26341,N_25654,N_25723);
and U26342 (N_26342,N_25608,N_25802);
or U26343 (N_26343,N_25861,N_25632);
or U26344 (N_26344,N_25641,N_25896);
xor U26345 (N_26345,N_25692,N_25870);
nor U26346 (N_26346,N_25866,N_25779);
or U26347 (N_26347,N_25951,N_25633);
nor U26348 (N_26348,N_25969,N_25620);
and U26349 (N_26349,N_25814,N_25904);
nor U26350 (N_26350,N_25611,N_25559);
nand U26351 (N_26351,N_25669,N_25876);
xor U26352 (N_26352,N_25809,N_25748);
nand U26353 (N_26353,N_25571,N_25653);
or U26354 (N_26354,N_25778,N_25891);
and U26355 (N_26355,N_25855,N_25702);
nor U26356 (N_26356,N_25810,N_25530);
and U26357 (N_26357,N_25644,N_25800);
xnor U26358 (N_26358,N_25982,N_25666);
nand U26359 (N_26359,N_25886,N_25618);
and U26360 (N_26360,N_25500,N_25564);
xnor U26361 (N_26361,N_25695,N_25641);
nor U26362 (N_26362,N_25829,N_25547);
nor U26363 (N_26363,N_25628,N_25774);
xnor U26364 (N_26364,N_25911,N_25845);
and U26365 (N_26365,N_25822,N_25940);
or U26366 (N_26366,N_25949,N_25777);
xnor U26367 (N_26367,N_25901,N_25934);
or U26368 (N_26368,N_25890,N_25686);
xor U26369 (N_26369,N_25913,N_25534);
and U26370 (N_26370,N_25516,N_25706);
nand U26371 (N_26371,N_25762,N_25998);
and U26372 (N_26372,N_25626,N_25571);
nand U26373 (N_26373,N_25807,N_25882);
nor U26374 (N_26374,N_25595,N_25953);
nor U26375 (N_26375,N_25929,N_25784);
xor U26376 (N_26376,N_25909,N_25895);
and U26377 (N_26377,N_25509,N_25687);
or U26378 (N_26378,N_25888,N_25987);
nand U26379 (N_26379,N_25522,N_25948);
nand U26380 (N_26380,N_25719,N_25965);
nor U26381 (N_26381,N_25680,N_25740);
and U26382 (N_26382,N_25996,N_25547);
or U26383 (N_26383,N_25853,N_25806);
or U26384 (N_26384,N_25845,N_25891);
or U26385 (N_26385,N_25792,N_25635);
xnor U26386 (N_26386,N_25799,N_25744);
nand U26387 (N_26387,N_25516,N_25780);
nor U26388 (N_26388,N_25798,N_25823);
nand U26389 (N_26389,N_25516,N_25896);
xor U26390 (N_26390,N_25816,N_25989);
nor U26391 (N_26391,N_25747,N_25783);
nor U26392 (N_26392,N_25975,N_25554);
nor U26393 (N_26393,N_25787,N_25716);
or U26394 (N_26394,N_25766,N_25840);
or U26395 (N_26395,N_25926,N_25678);
nor U26396 (N_26396,N_25723,N_25779);
nand U26397 (N_26397,N_25762,N_25866);
and U26398 (N_26398,N_25516,N_25904);
xnor U26399 (N_26399,N_25765,N_25899);
and U26400 (N_26400,N_25826,N_25875);
or U26401 (N_26401,N_25890,N_25869);
or U26402 (N_26402,N_25613,N_25995);
or U26403 (N_26403,N_25513,N_25553);
and U26404 (N_26404,N_25576,N_25683);
nand U26405 (N_26405,N_25676,N_25989);
nor U26406 (N_26406,N_25620,N_25548);
nand U26407 (N_26407,N_25702,N_25551);
and U26408 (N_26408,N_25757,N_25943);
nand U26409 (N_26409,N_25776,N_25767);
nor U26410 (N_26410,N_25922,N_25537);
nand U26411 (N_26411,N_25786,N_25605);
xor U26412 (N_26412,N_25619,N_25809);
nor U26413 (N_26413,N_25702,N_25789);
nand U26414 (N_26414,N_25954,N_25997);
nand U26415 (N_26415,N_25952,N_25971);
nor U26416 (N_26416,N_25737,N_25608);
xor U26417 (N_26417,N_25613,N_25864);
xor U26418 (N_26418,N_25940,N_25807);
or U26419 (N_26419,N_25939,N_25581);
and U26420 (N_26420,N_25846,N_25613);
nand U26421 (N_26421,N_25515,N_25807);
and U26422 (N_26422,N_25972,N_25639);
or U26423 (N_26423,N_25861,N_25526);
nand U26424 (N_26424,N_25900,N_25766);
xor U26425 (N_26425,N_25654,N_25927);
nor U26426 (N_26426,N_25762,N_25686);
or U26427 (N_26427,N_25519,N_25949);
xor U26428 (N_26428,N_25935,N_25769);
xnor U26429 (N_26429,N_25721,N_25898);
or U26430 (N_26430,N_25686,N_25737);
or U26431 (N_26431,N_25829,N_25957);
or U26432 (N_26432,N_25941,N_25613);
nand U26433 (N_26433,N_25844,N_25939);
and U26434 (N_26434,N_25822,N_25616);
nor U26435 (N_26435,N_25631,N_25861);
or U26436 (N_26436,N_25810,N_25956);
nand U26437 (N_26437,N_25618,N_25770);
nor U26438 (N_26438,N_25892,N_25935);
nor U26439 (N_26439,N_25709,N_25642);
nand U26440 (N_26440,N_25875,N_25979);
nor U26441 (N_26441,N_25792,N_25925);
or U26442 (N_26442,N_25766,N_25539);
or U26443 (N_26443,N_25567,N_25602);
xnor U26444 (N_26444,N_25929,N_25953);
or U26445 (N_26445,N_25728,N_25851);
nand U26446 (N_26446,N_25991,N_25687);
or U26447 (N_26447,N_25620,N_25963);
nor U26448 (N_26448,N_25833,N_25930);
nor U26449 (N_26449,N_25718,N_25717);
or U26450 (N_26450,N_25574,N_25937);
nor U26451 (N_26451,N_25651,N_25993);
xnor U26452 (N_26452,N_25614,N_25756);
xnor U26453 (N_26453,N_25793,N_25842);
or U26454 (N_26454,N_25846,N_25592);
xnor U26455 (N_26455,N_25772,N_25551);
and U26456 (N_26456,N_25590,N_25801);
or U26457 (N_26457,N_25502,N_25794);
or U26458 (N_26458,N_25658,N_25512);
nand U26459 (N_26459,N_25931,N_25752);
and U26460 (N_26460,N_25850,N_25718);
and U26461 (N_26461,N_25604,N_25696);
and U26462 (N_26462,N_25945,N_25914);
xor U26463 (N_26463,N_25952,N_25975);
nor U26464 (N_26464,N_25819,N_25519);
and U26465 (N_26465,N_25894,N_25533);
or U26466 (N_26466,N_25768,N_25502);
and U26467 (N_26467,N_25533,N_25698);
nor U26468 (N_26468,N_25921,N_25750);
nand U26469 (N_26469,N_25788,N_25839);
xnor U26470 (N_26470,N_25508,N_25616);
or U26471 (N_26471,N_25906,N_25822);
nand U26472 (N_26472,N_25504,N_25571);
xor U26473 (N_26473,N_25704,N_25533);
nor U26474 (N_26474,N_25797,N_25628);
and U26475 (N_26475,N_25932,N_25517);
nand U26476 (N_26476,N_25926,N_25695);
nand U26477 (N_26477,N_25692,N_25545);
nor U26478 (N_26478,N_25731,N_25923);
nand U26479 (N_26479,N_25805,N_25659);
xor U26480 (N_26480,N_25531,N_25875);
nand U26481 (N_26481,N_25884,N_25537);
or U26482 (N_26482,N_25757,N_25988);
nor U26483 (N_26483,N_25743,N_25701);
and U26484 (N_26484,N_25630,N_25758);
and U26485 (N_26485,N_25618,N_25675);
xnor U26486 (N_26486,N_25926,N_25572);
and U26487 (N_26487,N_25678,N_25611);
nand U26488 (N_26488,N_25595,N_25591);
nand U26489 (N_26489,N_25884,N_25816);
or U26490 (N_26490,N_25723,N_25975);
nor U26491 (N_26491,N_25886,N_25800);
or U26492 (N_26492,N_25601,N_25866);
xnor U26493 (N_26493,N_25693,N_25866);
and U26494 (N_26494,N_25854,N_25500);
or U26495 (N_26495,N_25853,N_25885);
xnor U26496 (N_26496,N_25544,N_25606);
xor U26497 (N_26497,N_25813,N_25620);
or U26498 (N_26498,N_25754,N_25791);
nor U26499 (N_26499,N_25520,N_25550);
nor U26500 (N_26500,N_26131,N_26448);
xor U26501 (N_26501,N_26146,N_26422);
nand U26502 (N_26502,N_26257,N_26114);
nor U26503 (N_26503,N_26302,N_26446);
nand U26504 (N_26504,N_26174,N_26037);
and U26505 (N_26505,N_26228,N_26339);
and U26506 (N_26506,N_26371,N_26351);
and U26507 (N_26507,N_26074,N_26135);
or U26508 (N_26508,N_26452,N_26327);
or U26509 (N_26509,N_26071,N_26009);
and U26510 (N_26510,N_26070,N_26349);
xor U26511 (N_26511,N_26436,N_26319);
nand U26512 (N_26512,N_26304,N_26210);
nor U26513 (N_26513,N_26283,N_26193);
nor U26514 (N_26514,N_26031,N_26063);
or U26515 (N_26515,N_26384,N_26399);
or U26516 (N_26516,N_26247,N_26077);
nor U26517 (N_26517,N_26083,N_26175);
or U26518 (N_26518,N_26222,N_26150);
xor U26519 (N_26519,N_26494,N_26321);
nor U26520 (N_26520,N_26005,N_26151);
xor U26521 (N_26521,N_26167,N_26062);
and U26522 (N_26522,N_26482,N_26216);
nor U26523 (N_26523,N_26342,N_26237);
xor U26524 (N_26524,N_26363,N_26055);
nor U26525 (N_26525,N_26292,N_26110);
xnor U26526 (N_26526,N_26359,N_26218);
nand U26527 (N_26527,N_26068,N_26061);
and U26528 (N_26528,N_26407,N_26153);
nor U26529 (N_26529,N_26138,N_26030);
or U26530 (N_26530,N_26271,N_26236);
xnor U26531 (N_26531,N_26212,N_26129);
nor U26532 (N_26532,N_26187,N_26059);
xor U26533 (N_26533,N_26015,N_26289);
nand U26534 (N_26534,N_26326,N_26299);
nand U26535 (N_26535,N_26343,N_26113);
xor U26536 (N_26536,N_26258,N_26166);
or U26537 (N_26537,N_26232,N_26233);
and U26538 (N_26538,N_26393,N_26312);
nor U26539 (N_26539,N_26435,N_26177);
xnor U26540 (N_26540,N_26159,N_26298);
nor U26541 (N_26541,N_26400,N_26365);
nor U26542 (N_26542,N_26473,N_26344);
xor U26543 (N_26543,N_26239,N_26211);
or U26544 (N_26544,N_26185,N_26488);
and U26545 (N_26545,N_26333,N_26352);
nor U26546 (N_26546,N_26388,N_26081);
and U26547 (N_26547,N_26214,N_26097);
xnor U26548 (N_26548,N_26119,N_26161);
nor U26549 (N_26549,N_26054,N_26242);
nand U26550 (N_26550,N_26396,N_26000);
xor U26551 (N_26551,N_26417,N_26140);
xnor U26552 (N_26552,N_26378,N_26092);
nand U26553 (N_26553,N_26035,N_26389);
and U26554 (N_26554,N_26294,N_26291);
and U26555 (N_26555,N_26290,N_26335);
and U26556 (N_26556,N_26002,N_26191);
nor U26557 (N_26557,N_26421,N_26476);
nand U26558 (N_26558,N_26282,N_26186);
nor U26559 (N_26559,N_26226,N_26367);
and U26560 (N_26560,N_26453,N_26330);
xor U26561 (N_26561,N_26273,N_26356);
xor U26562 (N_26562,N_26188,N_26065);
nand U26563 (N_26563,N_26460,N_26109);
xnor U26564 (N_26564,N_26047,N_26042);
or U26565 (N_26565,N_26230,N_26284);
or U26566 (N_26566,N_26178,N_26480);
nand U26567 (N_26567,N_26263,N_26457);
nor U26568 (N_26568,N_26267,N_26464);
nand U26569 (N_26569,N_26353,N_26145);
nand U26570 (N_26570,N_26204,N_26118);
nand U26571 (N_26571,N_26385,N_26038);
nand U26572 (N_26572,N_26034,N_26358);
xnor U26573 (N_26573,N_26391,N_26139);
xnor U26574 (N_26574,N_26004,N_26025);
nand U26575 (N_26575,N_26484,N_26424);
nor U26576 (N_26576,N_26456,N_26149);
nor U26577 (N_26577,N_26449,N_26366);
xnor U26578 (N_26578,N_26324,N_26137);
and U26579 (N_26579,N_26225,N_26102);
nand U26580 (N_26580,N_26433,N_26415);
or U26581 (N_26581,N_26231,N_26397);
nand U26582 (N_26582,N_26332,N_26171);
xor U26583 (N_26583,N_26308,N_26277);
and U26584 (N_26584,N_26437,N_26091);
and U26585 (N_26585,N_26314,N_26027);
or U26586 (N_26586,N_26348,N_26305);
or U26587 (N_26587,N_26136,N_26165);
nand U26588 (N_26588,N_26033,N_26440);
or U26589 (N_26589,N_26049,N_26338);
and U26590 (N_26590,N_26334,N_26147);
nor U26591 (N_26591,N_26196,N_26411);
and U26592 (N_26592,N_26219,N_26126);
nor U26593 (N_26593,N_26079,N_26316);
nand U26594 (N_26594,N_26280,N_26076);
or U26595 (N_26595,N_26429,N_26380);
or U26596 (N_26596,N_26197,N_26434);
nand U26597 (N_26597,N_26101,N_26200);
and U26598 (N_26598,N_26125,N_26229);
nand U26599 (N_26599,N_26016,N_26395);
and U26600 (N_26600,N_26360,N_26479);
nor U26601 (N_26601,N_26279,N_26084);
nor U26602 (N_26602,N_26450,N_26419);
or U26603 (N_26603,N_26007,N_26128);
nand U26604 (N_26604,N_26322,N_26491);
and U26605 (N_26605,N_26160,N_26148);
nand U26606 (N_26606,N_26100,N_26227);
nor U26607 (N_26607,N_26087,N_26439);
nand U26608 (N_26608,N_26072,N_26328);
and U26609 (N_26609,N_26022,N_26336);
and U26610 (N_26610,N_26431,N_26265);
nand U26611 (N_26611,N_26459,N_26379);
nand U26612 (N_26612,N_26454,N_26123);
or U26613 (N_26613,N_26181,N_26408);
or U26614 (N_26614,N_26203,N_26340);
and U26615 (N_26615,N_26492,N_26011);
nand U26616 (N_26616,N_26274,N_26423);
nand U26617 (N_26617,N_26155,N_26272);
and U26618 (N_26618,N_26402,N_26486);
or U26619 (N_26619,N_26205,N_26116);
nor U26620 (N_26620,N_26487,N_26288);
xor U26621 (N_26621,N_26078,N_26192);
nand U26622 (N_26622,N_26368,N_26472);
and U26623 (N_26623,N_26387,N_26040);
or U26624 (N_26624,N_26130,N_26414);
and U26625 (N_26625,N_26451,N_26221);
or U26626 (N_26626,N_26104,N_26194);
and U26627 (N_26627,N_26127,N_26286);
nand U26628 (N_26628,N_26354,N_26154);
or U26629 (N_26629,N_26318,N_26427);
or U26630 (N_26630,N_26382,N_26481);
or U26631 (N_26631,N_26207,N_26066);
and U26632 (N_26632,N_26347,N_26401);
xor U26633 (N_26633,N_26169,N_26093);
xor U26634 (N_26634,N_26303,N_26086);
xnor U26635 (N_26635,N_26412,N_26041);
or U26636 (N_26636,N_26310,N_26253);
xnor U26637 (N_26637,N_26471,N_26003);
xnor U26638 (N_26638,N_26478,N_26162);
nor U26639 (N_26639,N_26133,N_26013);
xnor U26640 (N_26640,N_26323,N_26141);
xor U26641 (N_26641,N_26018,N_26075);
nor U26642 (N_26642,N_26485,N_26331);
or U26643 (N_26643,N_26120,N_26264);
nor U26644 (N_26644,N_26021,N_26262);
or U26645 (N_26645,N_26498,N_26105);
nand U26646 (N_26646,N_26094,N_26409);
nand U26647 (N_26647,N_26251,N_26039);
nor U26648 (N_26648,N_26060,N_26096);
or U26649 (N_26649,N_26179,N_26202);
xnor U26650 (N_26650,N_26483,N_26469);
and U26651 (N_26651,N_26362,N_26489);
xor U26652 (N_26652,N_26244,N_26143);
nand U26653 (N_26653,N_26090,N_26019);
nor U26654 (N_26654,N_26088,N_26441);
or U26655 (N_26655,N_26381,N_26058);
nand U26656 (N_26656,N_26173,N_26325);
xnor U26657 (N_26657,N_26103,N_26275);
or U26658 (N_26658,N_26369,N_26495);
nor U26659 (N_26659,N_26142,N_26345);
and U26660 (N_26660,N_26067,N_26350);
nor U26661 (N_26661,N_26405,N_26132);
or U26662 (N_26662,N_26235,N_26099);
xnor U26663 (N_26663,N_26006,N_26455);
or U26664 (N_26664,N_26108,N_26241);
or U26665 (N_26665,N_26043,N_26050);
and U26666 (N_26666,N_26364,N_26240);
nor U26667 (N_26667,N_26377,N_26410);
or U26668 (N_26668,N_26438,N_26156);
nor U26669 (N_26669,N_26357,N_26246);
nor U26670 (N_26670,N_26445,N_26317);
or U26671 (N_26671,N_26152,N_26180);
xor U26672 (N_26672,N_26425,N_26172);
nor U26673 (N_26673,N_26248,N_26164);
nand U26674 (N_26674,N_26053,N_26069);
nor U26675 (N_26675,N_26144,N_26499);
xnor U26676 (N_26676,N_26028,N_26373);
or U26677 (N_26677,N_26493,N_26297);
nand U26678 (N_26678,N_26008,N_26117);
nand U26679 (N_26679,N_26122,N_26107);
or U26680 (N_26680,N_26458,N_26296);
or U26681 (N_26681,N_26406,N_26320);
or U26682 (N_26682,N_26080,N_26490);
xor U26683 (N_26683,N_26315,N_26183);
xor U26684 (N_26684,N_26256,N_26223);
nor U26685 (N_26685,N_26098,N_26255);
or U26686 (N_26686,N_26209,N_26361);
xor U26687 (N_26687,N_26026,N_26468);
nand U26688 (N_26688,N_26300,N_26287);
xnor U26689 (N_26689,N_26442,N_26112);
xor U26690 (N_26690,N_26010,N_26355);
or U26691 (N_26691,N_26046,N_26269);
xnor U26692 (N_26692,N_26121,N_26184);
xnor U26693 (N_26693,N_26346,N_26462);
and U26694 (N_26694,N_26158,N_26217);
nand U26695 (N_26695,N_26311,N_26386);
nor U26696 (N_26696,N_26443,N_26115);
and U26697 (N_26697,N_26374,N_26111);
nor U26698 (N_26698,N_26383,N_26313);
and U26699 (N_26699,N_26270,N_26259);
and U26700 (N_26700,N_26012,N_26134);
and U26701 (N_26701,N_26428,N_26190);
xnor U26702 (N_26702,N_26163,N_26260);
or U26703 (N_26703,N_26392,N_26001);
nor U26704 (N_26704,N_26461,N_26052);
nor U26705 (N_26705,N_26224,N_26467);
xnor U26706 (N_26706,N_26250,N_26278);
nor U26707 (N_26707,N_26045,N_26020);
xor U26708 (N_26708,N_26199,N_26466);
xor U26709 (N_26709,N_26238,N_26032);
nand U26710 (N_26710,N_26168,N_26249);
nor U26711 (N_26711,N_26176,N_26089);
or U26712 (N_26712,N_26157,N_26444);
nor U26713 (N_26713,N_26208,N_26293);
nand U26714 (N_26714,N_26475,N_26341);
nor U26715 (N_26715,N_26254,N_26375);
nand U26716 (N_26716,N_26309,N_26215);
or U26717 (N_26717,N_26394,N_26029);
xor U26718 (N_26718,N_26268,N_26370);
nand U26719 (N_26719,N_26044,N_26170);
nor U26720 (N_26720,N_26432,N_26082);
and U26721 (N_26721,N_26306,N_26403);
xnor U26722 (N_26722,N_26189,N_26420);
and U26723 (N_26723,N_26474,N_26497);
xor U26724 (N_26724,N_26404,N_26266);
or U26725 (N_26725,N_26261,N_26496);
or U26726 (N_26726,N_26206,N_26418);
nand U26727 (N_26727,N_26234,N_26036);
nor U26728 (N_26728,N_26295,N_26426);
xor U26729 (N_26729,N_26198,N_26276);
xor U26730 (N_26730,N_26220,N_26051);
or U26731 (N_26731,N_26017,N_26463);
xnor U26732 (N_26732,N_26477,N_26376);
or U26733 (N_26733,N_26095,N_26057);
xnor U26734 (N_26734,N_26023,N_26416);
nor U26735 (N_26735,N_26285,N_26252);
nor U26736 (N_26736,N_26243,N_26048);
nand U26737 (N_26737,N_26182,N_26372);
or U26738 (N_26738,N_26124,N_26073);
xor U26739 (N_26739,N_26301,N_26447);
or U26740 (N_26740,N_26329,N_26281);
or U26741 (N_26741,N_26064,N_26201);
or U26742 (N_26742,N_26195,N_26470);
nor U26743 (N_26743,N_26390,N_26465);
or U26744 (N_26744,N_26024,N_26307);
nor U26745 (N_26745,N_26398,N_26106);
nand U26746 (N_26746,N_26245,N_26085);
xor U26747 (N_26747,N_26430,N_26337);
or U26748 (N_26748,N_26413,N_26014);
nand U26749 (N_26749,N_26056,N_26213);
nand U26750 (N_26750,N_26453,N_26236);
and U26751 (N_26751,N_26094,N_26167);
nand U26752 (N_26752,N_26058,N_26355);
nand U26753 (N_26753,N_26498,N_26351);
xnor U26754 (N_26754,N_26327,N_26080);
or U26755 (N_26755,N_26378,N_26449);
xor U26756 (N_26756,N_26208,N_26376);
and U26757 (N_26757,N_26410,N_26311);
nand U26758 (N_26758,N_26281,N_26104);
nor U26759 (N_26759,N_26361,N_26135);
and U26760 (N_26760,N_26049,N_26258);
nor U26761 (N_26761,N_26183,N_26229);
nand U26762 (N_26762,N_26091,N_26492);
xnor U26763 (N_26763,N_26235,N_26061);
or U26764 (N_26764,N_26388,N_26023);
nand U26765 (N_26765,N_26260,N_26299);
or U26766 (N_26766,N_26206,N_26465);
and U26767 (N_26767,N_26358,N_26339);
and U26768 (N_26768,N_26232,N_26473);
nor U26769 (N_26769,N_26220,N_26196);
or U26770 (N_26770,N_26206,N_26126);
xor U26771 (N_26771,N_26147,N_26481);
and U26772 (N_26772,N_26433,N_26219);
or U26773 (N_26773,N_26226,N_26395);
nor U26774 (N_26774,N_26466,N_26215);
or U26775 (N_26775,N_26344,N_26205);
and U26776 (N_26776,N_26427,N_26310);
xnor U26777 (N_26777,N_26154,N_26447);
nor U26778 (N_26778,N_26300,N_26062);
and U26779 (N_26779,N_26237,N_26477);
or U26780 (N_26780,N_26397,N_26052);
nand U26781 (N_26781,N_26046,N_26000);
or U26782 (N_26782,N_26483,N_26477);
or U26783 (N_26783,N_26062,N_26111);
xor U26784 (N_26784,N_26130,N_26312);
nand U26785 (N_26785,N_26345,N_26365);
or U26786 (N_26786,N_26211,N_26462);
or U26787 (N_26787,N_26456,N_26461);
nand U26788 (N_26788,N_26092,N_26209);
and U26789 (N_26789,N_26077,N_26043);
or U26790 (N_26790,N_26483,N_26079);
and U26791 (N_26791,N_26151,N_26142);
nor U26792 (N_26792,N_26043,N_26081);
and U26793 (N_26793,N_26074,N_26086);
nor U26794 (N_26794,N_26186,N_26355);
nor U26795 (N_26795,N_26194,N_26198);
or U26796 (N_26796,N_26163,N_26259);
and U26797 (N_26797,N_26243,N_26465);
and U26798 (N_26798,N_26299,N_26332);
nor U26799 (N_26799,N_26084,N_26356);
xnor U26800 (N_26800,N_26178,N_26163);
nand U26801 (N_26801,N_26048,N_26051);
nand U26802 (N_26802,N_26389,N_26097);
xnor U26803 (N_26803,N_26040,N_26317);
nand U26804 (N_26804,N_26329,N_26258);
nor U26805 (N_26805,N_26484,N_26194);
xor U26806 (N_26806,N_26193,N_26223);
xnor U26807 (N_26807,N_26125,N_26122);
nand U26808 (N_26808,N_26355,N_26424);
and U26809 (N_26809,N_26305,N_26330);
xnor U26810 (N_26810,N_26331,N_26156);
or U26811 (N_26811,N_26103,N_26359);
nand U26812 (N_26812,N_26138,N_26035);
or U26813 (N_26813,N_26219,N_26370);
nor U26814 (N_26814,N_26334,N_26141);
nand U26815 (N_26815,N_26331,N_26403);
nor U26816 (N_26816,N_26386,N_26345);
nor U26817 (N_26817,N_26151,N_26013);
xor U26818 (N_26818,N_26175,N_26058);
xor U26819 (N_26819,N_26385,N_26485);
nor U26820 (N_26820,N_26231,N_26291);
or U26821 (N_26821,N_26109,N_26155);
or U26822 (N_26822,N_26471,N_26067);
nor U26823 (N_26823,N_26455,N_26080);
nor U26824 (N_26824,N_26185,N_26074);
nand U26825 (N_26825,N_26028,N_26360);
and U26826 (N_26826,N_26043,N_26052);
and U26827 (N_26827,N_26049,N_26063);
and U26828 (N_26828,N_26318,N_26039);
nand U26829 (N_26829,N_26347,N_26072);
nand U26830 (N_26830,N_26194,N_26424);
nand U26831 (N_26831,N_26081,N_26481);
and U26832 (N_26832,N_26070,N_26115);
xor U26833 (N_26833,N_26206,N_26463);
nor U26834 (N_26834,N_26295,N_26264);
nor U26835 (N_26835,N_26046,N_26291);
nand U26836 (N_26836,N_26021,N_26201);
nand U26837 (N_26837,N_26306,N_26254);
nor U26838 (N_26838,N_26151,N_26025);
nand U26839 (N_26839,N_26485,N_26039);
xor U26840 (N_26840,N_26461,N_26194);
nand U26841 (N_26841,N_26314,N_26038);
nand U26842 (N_26842,N_26155,N_26319);
xor U26843 (N_26843,N_26471,N_26147);
nor U26844 (N_26844,N_26015,N_26469);
nor U26845 (N_26845,N_26210,N_26456);
xnor U26846 (N_26846,N_26464,N_26463);
or U26847 (N_26847,N_26237,N_26323);
nand U26848 (N_26848,N_26156,N_26276);
xnor U26849 (N_26849,N_26330,N_26383);
xnor U26850 (N_26850,N_26198,N_26115);
xor U26851 (N_26851,N_26053,N_26042);
and U26852 (N_26852,N_26155,N_26150);
and U26853 (N_26853,N_26444,N_26148);
nand U26854 (N_26854,N_26319,N_26309);
or U26855 (N_26855,N_26091,N_26031);
or U26856 (N_26856,N_26241,N_26497);
and U26857 (N_26857,N_26092,N_26414);
nand U26858 (N_26858,N_26123,N_26422);
nor U26859 (N_26859,N_26400,N_26388);
nand U26860 (N_26860,N_26384,N_26033);
nor U26861 (N_26861,N_26252,N_26246);
or U26862 (N_26862,N_26444,N_26435);
and U26863 (N_26863,N_26310,N_26281);
or U26864 (N_26864,N_26128,N_26076);
xnor U26865 (N_26865,N_26098,N_26060);
and U26866 (N_26866,N_26177,N_26024);
xor U26867 (N_26867,N_26483,N_26305);
or U26868 (N_26868,N_26249,N_26095);
nand U26869 (N_26869,N_26193,N_26385);
or U26870 (N_26870,N_26083,N_26028);
or U26871 (N_26871,N_26322,N_26402);
nand U26872 (N_26872,N_26178,N_26126);
nand U26873 (N_26873,N_26489,N_26235);
and U26874 (N_26874,N_26013,N_26086);
or U26875 (N_26875,N_26176,N_26126);
or U26876 (N_26876,N_26263,N_26345);
xnor U26877 (N_26877,N_26254,N_26427);
nand U26878 (N_26878,N_26453,N_26129);
nor U26879 (N_26879,N_26440,N_26227);
and U26880 (N_26880,N_26296,N_26263);
nor U26881 (N_26881,N_26285,N_26464);
nor U26882 (N_26882,N_26345,N_26141);
nand U26883 (N_26883,N_26255,N_26055);
and U26884 (N_26884,N_26251,N_26164);
or U26885 (N_26885,N_26370,N_26346);
and U26886 (N_26886,N_26421,N_26146);
and U26887 (N_26887,N_26242,N_26020);
or U26888 (N_26888,N_26068,N_26337);
or U26889 (N_26889,N_26410,N_26468);
nor U26890 (N_26890,N_26141,N_26264);
nor U26891 (N_26891,N_26224,N_26416);
nor U26892 (N_26892,N_26224,N_26064);
xnor U26893 (N_26893,N_26050,N_26340);
or U26894 (N_26894,N_26484,N_26159);
nor U26895 (N_26895,N_26032,N_26122);
or U26896 (N_26896,N_26013,N_26278);
nor U26897 (N_26897,N_26237,N_26136);
nor U26898 (N_26898,N_26185,N_26268);
and U26899 (N_26899,N_26412,N_26413);
and U26900 (N_26900,N_26458,N_26003);
nand U26901 (N_26901,N_26035,N_26432);
xor U26902 (N_26902,N_26028,N_26064);
and U26903 (N_26903,N_26442,N_26211);
nor U26904 (N_26904,N_26153,N_26113);
or U26905 (N_26905,N_26386,N_26200);
or U26906 (N_26906,N_26116,N_26370);
and U26907 (N_26907,N_26005,N_26246);
and U26908 (N_26908,N_26120,N_26163);
nand U26909 (N_26909,N_26468,N_26371);
nand U26910 (N_26910,N_26448,N_26141);
or U26911 (N_26911,N_26306,N_26393);
nor U26912 (N_26912,N_26169,N_26274);
nor U26913 (N_26913,N_26241,N_26072);
and U26914 (N_26914,N_26392,N_26331);
or U26915 (N_26915,N_26230,N_26301);
and U26916 (N_26916,N_26187,N_26325);
or U26917 (N_26917,N_26156,N_26183);
and U26918 (N_26918,N_26369,N_26214);
and U26919 (N_26919,N_26426,N_26355);
or U26920 (N_26920,N_26144,N_26259);
nor U26921 (N_26921,N_26309,N_26383);
and U26922 (N_26922,N_26370,N_26126);
and U26923 (N_26923,N_26245,N_26473);
and U26924 (N_26924,N_26310,N_26214);
and U26925 (N_26925,N_26022,N_26434);
xnor U26926 (N_26926,N_26104,N_26204);
xnor U26927 (N_26927,N_26019,N_26089);
or U26928 (N_26928,N_26006,N_26499);
nor U26929 (N_26929,N_26439,N_26164);
nor U26930 (N_26930,N_26172,N_26203);
or U26931 (N_26931,N_26133,N_26302);
nand U26932 (N_26932,N_26018,N_26099);
and U26933 (N_26933,N_26190,N_26291);
xnor U26934 (N_26934,N_26294,N_26402);
or U26935 (N_26935,N_26116,N_26326);
or U26936 (N_26936,N_26361,N_26225);
nand U26937 (N_26937,N_26028,N_26044);
nand U26938 (N_26938,N_26181,N_26044);
xor U26939 (N_26939,N_26049,N_26311);
or U26940 (N_26940,N_26012,N_26079);
nor U26941 (N_26941,N_26267,N_26263);
xnor U26942 (N_26942,N_26337,N_26088);
or U26943 (N_26943,N_26142,N_26334);
xnor U26944 (N_26944,N_26251,N_26195);
and U26945 (N_26945,N_26232,N_26108);
nand U26946 (N_26946,N_26093,N_26261);
and U26947 (N_26947,N_26427,N_26062);
or U26948 (N_26948,N_26058,N_26203);
nand U26949 (N_26949,N_26239,N_26204);
nand U26950 (N_26950,N_26135,N_26029);
or U26951 (N_26951,N_26198,N_26131);
nand U26952 (N_26952,N_26086,N_26151);
xor U26953 (N_26953,N_26330,N_26156);
and U26954 (N_26954,N_26424,N_26187);
xnor U26955 (N_26955,N_26426,N_26473);
and U26956 (N_26956,N_26451,N_26160);
nor U26957 (N_26957,N_26053,N_26029);
nand U26958 (N_26958,N_26417,N_26273);
and U26959 (N_26959,N_26040,N_26265);
and U26960 (N_26960,N_26151,N_26465);
nand U26961 (N_26961,N_26291,N_26341);
nand U26962 (N_26962,N_26284,N_26117);
or U26963 (N_26963,N_26215,N_26176);
and U26964 (N_26964,N_26137,N_26441);
nor U26965 (N_26965,N_26355,N_26307);
or U26966 (N_26966,N_26163,N_26326);
nand U26967 (N_26967,N_26241,N_26372);
nand U26968 (N_26968,N_26000,N_26436);
nor U26969 (N_26969,N_26487,N_26260);
or U26970 (N_26970,N_26413,N_26037);
nor U26971 (N_26971,N_26256,N_26090);
and U26972 (N_26972,N_26152,N_26278);
and U26973 (N_26973,N_26097,N_26184);
xor U26974 (N_26974,N_26356,N_26309);
xnor U26975 (N_26975,N_26071,N_26364);
and U26976 (N_26976,N_26172,N_26309);
xnor U26977 (N_26977,N_26136,N_26131);
or U26978 (N_26978,N_26260,N_26011);
or U26979 (N_26979,N_26333,N_26005);
xor U26980 (N_26980,N_26190,N_26327);
and U26981 (N_26981,N_26127,N_26107);
and U26982 (N_26982,N_26064,N_26442);
nand U26983 (N_26983,N_26271,N_26101);
nor U26984 (N_26984,N_26082,N_26449);
nand U26985 (N_26985,N_26276,N_26071);
or U26986 (N_26986,N_26449,N_26311);
xnor U26987 (N_26987,N_26202,N_26125);
nand U26988 (N_26988,N_26399,N_26287);
and U26989 (N_26989,N_26354,N_26092);
and U26990 (N_26990,N_26072,N_26269);
nor U26991 (N_26991,N_26085,N_26083);
nand U26992 (N_26992,N_26053,N_26180);
and U26993 (N_26993,N_26199,N_26389);
nand U26994 (N_26994,N_26009,N_26243);
and U26995 (N_26995,N_26448,N_26342);
nor U26996 (N_26996,N_26332,N_26286);
xor U26997 (N_26997,N_26051,N_26098);
and U26998 (N_26998,N_26137,N_26035);
nor U26999 (N_26999,N_26205,N_26121);
nand U27000 (N_27000,N_26708,N_26612);
and U27001 (N_27001,N_26517,N_26920);
or U27002 (N_27002,N_26873,N_26667);
or U27003 (N_27003,N_26826,N_26809);
xor U27004 (N_27004,N_26638,N_26796);
and U27005 (N_27005,N_26524,N_26872);
nand U27006 (N_27006,N_26684,N_26795);
or U27007 (N_27007,N_26545,N_26541);
or U27008 (N_27008,N_26665,N_26516);
or U27009 (N_27009,N_26553,N_26648);
nor U27010 (N_27010,N_26771,N_26882);
nor U27011 (N_27011,N_26519,N_26959);
nor U27012 (N_27012,N_26570,N_26767);
xor U27013 (N_27013,N_26556,N_26677);
nor U27014 (N_27014,N_26861,N_26670);
nor U27015 (N_27015,N_26792,N_26569);
nor U27016 (N_27016,N_26789,N_26555);
nand U27017 (N_27017,N_26544,N_26835);
or U27018 (N_27018,N_26950,N_26986);
nand U27019 (N_27019,N_26803,N_26630);
nand U27020 (N_27020,N_26855,N_26913);
nor U27021 (N_27021,N_26790,N_26995);
xnor U27022 (N_27022,N_26894,N_26543);
xor U27023 (N_27023,N_26983,N_26916);
and U27024 (N_27024,N_26940,N_26720);
and U27025 (N_27025,N_26586,N_26689);
or U27026 (N_27026,N_26699,N_26899);
nor U27027 (N_27027,N_26726,N_26534);
xor U27028 (N_27028,N_26674,N_26664);
xnor U27029 (N_27029,N_26863,N_26752);
and U27030 (N_27030,N_26999,N_26504);
xor U27031 (N_27031,N_26691,N_26818);
xnor U27032 (N_27032,N_26822,N_26778);
xor U27033 (N_27033,N_26906,N_26837);
and U27034 (N_27034,N_26653,N_26693);
or U27035 (N_27035,N_26565,N_26714);
nand U27036 (N_27036,N_26770,N_26881);
or U27037 (N_27037,N_26785,N_26783);
xnor U27038 (N_27038,N_26523,N_26994);
or U27039 (N_27039,N_26907,N_26529);
nor U27040 (N_27040,N_26814,N_26585);
nand U27041 (N_27041,N_26614,N_26522);
xnor U27042 (N_27042,N_26997,N_26696);
and U27043 (N_27043,N_26563,N_26942);
or U27044 (N_27044,N_26633,N_26948);
xor U27045 (N_27045,N_26635,N_26853);
nor U27046 (N_27046,N_26824,N_26890);
nor U27047 (N_27047,N_26686,N_26905);
xnor U27048 (N_27048,N_26954,N_26632);
xnor U27049 (N_27049,N_26690,N_26596);
xor U27050 (N_27050,N_26535,N_26589);
nand U27051 (N_27051,N_26548,N_26911);
nand U27052 (N_27052,N_26582,N_26839);
and U27053 (N_27053,N_26636,N_26564);
or U27054 (N_27054,N_26955,N_26870);
nor U27055 (N_27055,N_26869,N_26801);
or U27056 (N_27056,N_26985,N_26926);
or U27057 (N_27057,N_26979,N_26981);
nand U27058 (N_27058,N_26896,N_26511);
nand U27059 (N_27059,N_26729,N_26918);
nand U27060 (N_27060,N_26845,N_26990);
xnor U27061 (N_27061,N_26634,N_26876);
or U27062 (N_27062,N_26977,N_26937);
and U27063 (N_27063,N_26935,N_26827);
and U27064 (N_27064,N_26859,N_26621);
and U27065 (N_27065,N_26807,N_26668);
nor U27066 (N_27066,N_26965,N_26603);
xor U27067 (N_27067,N_26850,N_26908);
and U27068 (N_27068,N_26788,N_26888);
and U27069 (N_27069,N_26625,N_26804);
xnor U27070 (N_27070,N_26904,N_26846);
nor U27071 (N_27071,N_26622,N_26542);
xor U27072 (N_27072,N_26927,N_26520);
and U27073 (N_27073,N_26551,N_26830);
nor U27074 (N_27074,N_26507,N_26787);
xor U27075 (N_27075,N_26838,N_26685);
or U27076 (N_27076,N_26640,N_26760);
or U27077 (N_27077,N_26949,N_26660);
or U27078 (N_27078,N_26738,N_26525);
and U27079 (N_27079,N_26521,N_26834);
xnor U27080 (N_27080,N_26610,N_26607);
and U27081 (N_27081,N_26680,N_26731);
and U27082 (N_27082,N_26641,N_26799);
and U27083 (N_27083,N_26812,N_26750);
or U27084 (N_27084,N_26597,N_26931);
xnor U27085 (N_27085,N_26619,N_26700);
nand U27086 (N_27086,N_26945,N_26879);
nor U27087 (N_27087,N_26806,N_26895);
nor U27088 (N_27088,N_26975,N_26584);
or U27089 (N_27089,N_26620,N_26898);
and U27090 (N_27090,N_26580,N_26592);
nand U27091 (N_27091,N_26503,N_26518);
nor U27092 (N_27092,N_26793,N_26832);
nand U27093 (N_27093,N_26721,N_26813);
nand U27094 (N_27094,N_26887,N_26891);
nor U27095 (N_27095,N_26688,N_26577);
or U27096 (N_27096,N_26669,N_26774);
nor U27097 (N_27097,N_26746,N_26854);
or U27098 (N_27098,N_26909,N_26657);
xnor U27099 (N_27099,N_26958,N_26559);
nor U27100 (N_27100,N_26591,N_26572);
xor U27101 (N_27101,N_26704,N_26533);
nor U27102 (N_27102,N_26903,N_26718);
and U27103 (N_27103,N_26605,N_26831);
and U27104 (N_27104,N_26647,N_26840);
nand U27105 (N_27105,N_26659,N_26849);
xnor U27106 (N_27106,N_26554,N_26836);
nand U27107 (N_27107,N_26514,N_26593);
and U27108 (N_27108,N_26505,N_26772);
or U27109 (N_27109,N_26594,N_26815);
xnor U27110 (N_27110,N_26971,N_26627);
nand U27111 (N_27111,N_26515,N_26765);
xor U27112 (N_27112,N_26956,N_26736);
or U27113 (N_27113,N_26848,N_26650);
xnor U27114 (N_27114,N_26805,N_26600);
or U27115 (N_27115,N_26780,N_26698);
xnor U27116 (N_27116,N_26724,N_26877);
nor U27117 (N_27117,N_26508,N_26912);
nand U27118 (N_27118,N_26744,N_26679);
xnor U27119 (N_27119,N_26947,N_26961);
xor U27120 (N_27120,N_26856,N_26798);
or U27121 (N_27121,N_26811,N_26784);
or U27122 (N_27122,N_26722,N_26973);
or U27123 (N_27123,N_26536,N_26883);
or U27124 (N_27124,N_26711,N_26590);
and U27125 (N_27125,N_26506,N_26509);
nor U27126 (N_27126,N_26512,N_26616);
and U27127 (N_27127,N_26637,N_26531);
nand U27128 (N_27128,N_26917,N_26867);
nand U27129 (N_27129,N_26719,N_26609);
and U27130 (N_27130,N_26751,N_26957);
and U27131 (N_27131,N_26608,N_26741);
and U27132 (N_27132,N_26715,N_26930);
and U27133 (N_27133,N_26651,N_26725);
nor U27134 (N_27134,N_26702,N_26847);
nor U27135 (N_27135,N_26717,N_26547);
or U27136 (N_27136,N_26989,N_26860);
or U27137 (N_27137,N_26921,N_26993);
nor U27138 (N_27138,N_26819,N_26695);
xnor U27139 (N_27139,N_26510,N_26540);
and U27140 (N_27140,N_26893,N_26655);
nor U27141 (N_27141,N_26742,N_26578);
and U27142 (N_27142,N_26694,N_26841);
nand U27143 (N_27143,N_26552,N_26528);
xnor U27144 (N_27144,N_26967,N_26623);
nand U27145 (N_27145,N_26713,N_26968);
xnor U27146 (N_27146,N_26966,N_26573);
nand U27147 (N_27147,N_26773,N_26723);
and U27148 (N_27148,N_26757,N_26661);
or U27149 (N_27149,N_26932,N_26735);
and U27150 (N_27150,N_26759,N_26617);
nor U27151 (N_27151,N_26755,N_26558);
nor U27152 (N_27152,N_26864,N_26939);
or U27153 (N_27153,N_26922,N_26613);
and U27154 (N_27154,N_26706,N_26579);
xor U27155 (N_27155,N_26781,N_26575);
or U27156 (N_27156,N_26568,N_26978);
nor U27157 (N_27157,N_26996,N_26892);
nor U27158 (N_27158,N_26962,N_26566);
and U27159 (N_27159,N_26923,N_26933);
nand U27160 (N_27160,N_26902,N_26987);
and U27161 (N_27161,N_26513,N_26952);
nand U27162 (N_27162,N_26502,N_26754);
or U27163 (N_27163,N_26546,N_26972);
nand U27164 (N_27164,N_26743,N_26749);
xor U27165 (N_27165,N_26758,N_26914);
and U27166 (N_27166,N_26823,N_26762);
nand U27167 (N_27167,N_26797,N_26576);
nor U27168 (N_27168,N_26642,N_26557);
xor U27169 (N_27169,N_26526,N_26745);
nor U27170 (N_27170,N_26763,N_26560);
and U27171 (N_27171,N_26969,N_26676);
nand U27172 (N_27172,N_26992,N_26712);
or U27173 (N_27173,N_26984,N_26951);
nor U27174 (N_27174,N_26808,N_26618);
nor U27175 (N_27175,N_26656,N_26733);
nor U27176 (N_27176,N_26875,N_26739);
nor U27177 (N_27177,N_26730,N_26889);
nand U27178 (N_27178,N_26862,N_26764);
nor U27179 (N_27179,N_26943,N_26588);
nand U27180 (N_27180,N_26761,N_26727);
nor U27181 (N_27181,N_26925,N_26606);
or U27182 (N_27182,N_26734,N_26800);
xor U27183 (N_27183,N_26732,N_26756);
xnor U27184 (N_27184,N_26611,N_26550);
or U27185 (N_27185,N_26631,N_26705);
and U27186 (N_27186,N_26598,N_26897);
nor U27187 (N_27187,N_26595,N_26915);
nor U27188 (N_27188,N_26645,N_26938);
nand U27189 (N_27189,N_26581,N_26709);
xnor U27190 (N_27190,N_26615,N_26865);
xnor U27191 (N_27191,N_26946,N_26976);
and U27192 (N_27192,N_26960,N_26782);
or U27193 (N_27193,N_26768,N_26500);
xor U27194 (N_27194,N_26766,N_26639);
and U27195 (N_27195,N_26924,N_26626);
or U27196 (N_27196,N_26681,N_26624);
or U27197 (N_27197,N_26928,N_26777);
nor U27198 (N_27198,N_26666,N_26530);
nand U27199 (N_27199,N_26716,N_26821);
nand U27200 (N_27200,N_26874,N_26786);
or U27201 (N_27201,N_26843,N_26779);
or U27202 (N_27202,N_26697,N_26866);
nor U27203 (N_27203,N_26791,N_26878);
or U27204 (N_27204,N_26682,N_26885);
and U27205 (N_27205,N_26748,N_26549);
nor U27206 (N_27206,N_26934,N_26858);
nand U27207 (N_27207,N_26662,N_26816);
xor U27208 (N_27208,N_26654,N_26663);
nand U27209 (N_27209,N_26941,N_26601);
and U27210 (N_27210,N_26871,N_26672);
and U27211 (N_27211,N_26991,N_26562);
nor U27212 (N_27212,N_26775,N_26658);
and U27213 (N_27213,N_26628,N_26644);
and U27214 (N_27214,N_26629,N_26910);
nand U27215 (N_27215,N_26919,N_26988);
or U27216 (N_27216,N_26820,N_26646);
or U27217 (N_27217,N_26728,N_26737);
or U27218 (N_27218,N_26880,N_26671);
nor U27219 (N_27219,N_26810,N_26740);
nand U27220 (N_27220,N_26687,N_26538);
xnor U27221 (N_27221,N_26936,N_26501);
nand U27222 (N_27222,N_26901,N_26587);
xor U27223 (N_27223,N_26884,N_26817);
nor U27224 (N_27224,N_26794,N_26852);
nor U27225 (N_27225,N_26537,N_26829);
or U27226 (N_27226,N_26900,N_26982);
and U27227 (N_27227,N_26970,N_26802);
or U27228 (N_27228,N_26833,N_26844);
xnor U27229 (N_27229,N_26675,N_26604);
xor U27230 (N_27230,N_26964,N_26998);
or U27231 (N_27231,N_26963,N_26953);
and U27232 (N_27232,N_26673,N_26707);
or U27233 (N_27233,N_26583,N_26851);
or U27234 (N_27234,N_26747,N_26652);
nor U27235 (N_27235,N_26527,N_26842);
nand U27236 (N_27236,N_26532,N_26944);
xnor U27237 (N_27237,N_26776,N_26599);
and U27238 (N_27238,N_26980,N_26567);
nor U27239 (N_27239,N_26857,N_26886);
nand U27240 (N_27240,N_26828,N_26710);
nor U27241 (N_27241,N_26678,N_26692);
nor U27242 (N_27242,N_26929,N_26974);
xnor U27243 (N_27243,N_26703,N_26868);
xor U27244 (N_27244,N_26643,N_26649);
and U27245 (N_27245,N_26602,N_26701);
nor U27246 (N_27246,N_26825,N_26561);
nand U27247 (N_27247,N_26683,N_26574);
nor U27248 (N_27248,N_26539,N_26571);
and U27249 (N_27249,N_26753,N_26769);
xnor U27250 (N_27250,N_26607,N_26776);
xnor U27251 (N_27251,N_26810,N_26508);
and U27252 (N_27252,N_26685,N_26936);
nor U27253 (N_27253,N_26973,N_26905);
or U27254 (N_27254,N_26974,N_26947);
xor U27255 (N_27255,N_26666,N_26971);
xnor U27256 (N_27256,N_26511,N_26923);
nand U27257 (N_27257,N_26510,N_26872);
xnor U27258 (N_27258,N_26779,N_26799);
xnor U27259 (N_27259,N_26702,N_26513);
nand U27260 (N_27260,N_26793,N_26924);
nor U27261 (N_27261,N_26715,N_26753);
nor U27262 (N_27262,N_26619,N_26719);
nor U27263 (N_27263,N_26930,N_26932);
nor U27264 (N_27264,N_26758,N_26959);
xor U27265 (N_27265,N_26799,N_26580);
nand U27266 (N_27266,N_26716,N_26765);
nand U27267 (N_27267,N_26767,N_26757);
and U27268 (N_27268,N_26836,N_26995);
xnor U27269 (N_27269,N_26765,N_26734);
xnor U27270 (N_27270,N_26947,N_26965);
nand U27271 (N_27271,N_26594,N_26889);
nand U27272 (N_27272,N_26740,N_26530);
xor U27273 (N_27273,N_26627,N_26563);
or U27274 (N_27274,N_26692,N_26576);
nor U27275 (N_27275,N_26909,N_26613);
nand U27276 (N_27276,N_26633,N_26593);
nor U27277 (N_27277,N_26716,N_26598);
nor U27278 (N_27278,N_26576,N_26800);
or U27279 (N_27279,N_26982,N_26591);
or U27280 (N_27280,N_26500,N_26584);
nand U27281 (N_27281,N_26679,N_26711);
nand U27282 (N_27282,N_26792,N_26954);
or U27283 (N_27283,N_26644,N_26669);
or U27284 (N_27284,N_26933,N_26767);
nor U27285 (N_27285,N_26716,N_26603);
or U27286 (N_27286,N_26534,N_26537);
xor U27287 (N_27287,N_26534,N_26540);
xor U27288 (N_27288,N_26918,N_26820);
and U27289 (N_27289,N_26980,N_26928);
nor U27290 (N_27290,N_26890,N_26804);
or U27291 (N_27291,N_26629,N_26799);
or U27292 (N_27292,N_26515,N_26773);
xor U27293 (N_27293,N_26594,N_26696);
or U27294 (N_27294,N_26779,N_26829);
nor U27295 (N_27295,N_26527,N_26875);
and U27296 (N_27296,N_26710,N_26518);
or U27297 (N_27297,N_26922,N_26693);
nor U27298 (N_27298,N_26971,N_26536);
and U27299 (N_27299,N_26534,N_26813);
nor U27300 (N_27300,N_26512,N_26577);
or U27301 (N_27301,N_26733,N_26865);
nand U27302 (N_27302,N_26980,N_26806);
xor U27303 (N_27303,N_26775,N_26777);
xnor U27304 (N_27304,N_26777,N_26905);
xnor U27305 (N_27305,N_26989,N_26819);
and U27306 (N_27306,N_26731,N_26871);
and U27307 (N_27307,N_26702,N_26657);
and U27308 (N_27308,N_26914,N_26817);
and U27309 (N_27309,N_26692,N_26856);
nor U27310 (N_27310,N_26511,N_26613);
or U27311 (N_27311,N_26671,N_26924);
xor U27312 (N_27312,N_26781,N_26620);
or U27313 (N_27313,N_26746,N_26596);
nor U27314 (N_27314,N_26636,N_26907);
nand U27315 (N_27315,N_26601,N_26574);
xor U27316 (N_27316,N_26664,N_26685);
nand U27317 (N_27317,N_26765,N_26565);
or U27318 (N_27318,N_26601,N_26801);
or U27319 (N_27319,N_26760,N_26715);
nand U27320 (N_27320,N_26787,N_26886);
nor U27321 (N_27321,N_26966,N_26944);
and U27322 (N_27322,N_26871,N_26512);
or U27323 (N_27323,N_26904,N_26956);
and U27324 (N_27324,N_26761,N_26724);
and U27325 (N_27325,N_26678,N_26551);
nor U27326 (N_27326,N_26685,N_26622);
nand U27327 (N_27327,N_26510,N_26550);
nand U27328 (N_27328,N_26623,N_26729);
xor U27329 (N_27329,N_26635,N_26591);
or U27330 (N_27330,N_26655,N_26638);
xnor U27331 (N_27331,N_26929,N_26748);
nor U27332 (N_27332,N_26907,N_26696);
or U27333 (N_27333,N_26898,N_26963);
xor U27334 (N_27334,N_26653,N_26579);
nand U27335 (N_27335,N_26856,N_26869);
nor U27336 (N_27336,N_26631,N_26938);
nand U27337 (N_27337,N_26566,N_26854);
xor U27338 (N_27338,N_26959,N_26540);
nor U27339 (N_27339,N_26606,N_26530);
nand U27340 (N_27340,N_26752,N_26719);
xnor U27341 (N_27341,N_26738,N_26873);
and U27342 (N_27342,N_26637,N_26773);
nand U27343 (N_27343,N_26614,N_26774);
nand U27344 (N_27344,N_26998,N_26722);
or U27345 (N_27345,N_26980,N_26617);
or U27346 (N_27346,N_26792,N_26959);
nor U27347 (N_27347,N_26844,N_26974);
nand U27348 (N_27348,N_26556,N_26528);
nand U27349 (N_27349,N_26895,N_26831);
nor U27350 (N_27350,N_26592,N_26640);
and U27351 (N_27351,N_26722,N_26602);
nor U27352 (N_27352,N_26694,N_26842);
and U27353 (N_27353,N_26977,N_26696);
xnor U27354 (N_27354,N_26535,N_26869);
xnor U27355 (N_27355,N_26511,N_26912);
and U27356 (N_27356,N_26504,N_26533);
nand U27357 (N_27357,N_26837,N_26985);
nand U27358 (N_27358,N_26636,N_26566);
nand U27359 (N_27359,N_26711,N_26532);
nand U27360 (N_27360,N_26503,N_26535);
and U27361 (N_27361,N_26544,N_26898);
nand U27362 (N_27362,N_26775,N_26712);
nor U27363 (N_27363,N_26552,N_26779);
nor U27364 (N_27364,N_26643,N_26818);
and U27365 (N_27365,N_26755,N_26846);
nor U27366 (N_27366,N_26868,N_26693);
and U27367 (N_27367,N_26806,N_26741);
and U27368 (N_27368,N_26567,N_26748);
nand U27369 (N_27369,N_26702,N_26781);
and U27370 (N_27370,N_26738,N_26767);
nand U27371 (N_27371,N_26773,N_26798);
xnor U27372 (N_27372,N_26748,N_26756);
nor U27373 (N_27373,N_26942,N_26615);
xnor U27374 (N_27374,N_26725,N_26924);
and U27375 (N_27375,N_26872,N_26717);
nor U27376 (N_27376,N_26700,N_26771);
and U27377 (N_27377,N_26650,N_26917);
or U27378 (N_27378,N_26737,N_26618);
xnor U27379 (N_27379,N_26704,N_26667);
xor U27380 (N_27380,N_26677,N_26559);
or U27381 (N_27381,N_26685,N_26536);
nand U27382 (N_27382,N_26526,N_26516);
and U27383 (N_27383,N_26674,N_26793);
nor U27384 (N_27384,N_26750,N_26796);
and U27385 (N_27385,N_26709,N_26616);
xnor U27386 (N_27386,N_26797,N_26857);
or U27387 (N_27387,N_26706,N_26690);
nand U27388 (N_27388,N_26577,N_26518);
and U27389 (N_27389,N_26817,N_26743);
nor U27390 (N_27390,N_26641,N_26902);
nand U27391 (N_27391,N_26585,N_26607);
nor U27392 (N_27392,N_26522,N_26581);
or U27393 (N_27393,N_26963,N_26628);
nand U27394 (N_27394,N_26937,N_26575);
nor U27395 (N_27395,N_26878,N_26838);
and U27396 (N_27396,N_26679,N_26528);
nor U27397 (N_27397,N_26678,N_26834);
xor U27398 (N_27398,N_26708,N_26521);
nor U27399 (N_27399,N_26750,N_26919);
and U27400 (N_27400,N_26750,N_26999);
and U27401 (N_27401,N_26975,N_26606);
or U27402 (N_27402,N_26526,N_26720);
xor U27403 (N_27403,N_26723,N_26760);
xnor U27404 (N_27404,N_26614,N_26658);
and U27405 (N_27405,N_26732,N_26547);
nor U27406 (N_27406,N_26806,N_26793);
xnor U27407 (N_27407,N_26801,N_26620);
and U27408 (N_27408,N_26854,N_26988);
or U27409 (N_27409,N_26702,N_26517);
or U27410 (N_27410,N_26942,N_26720);
and U27411 (N_27411,N_26776,N_26602);
or U27412 (N_27412,N_26683,N_26658);
or U27413 (N_27413,N_26527,N_26973);
xnor U27414 (N_27414,N_26871,N_26852);
nor U27415 (N_27415,N_26618,N_26578);
nand U27416 (N_27416,N_26935,N_26985);
or U27417 (N_27417,N_26603,N_26959);
nand U27418 (N_27418,N_26852,N_26933);
xor U27419 (N_27419,N_26541,N_26613);
xor U27420 (N_27420,N_26667,N_26644);
and U27421 (N_27421,N_26813,N_26799);
nor U27422 (N_27422,N_26879,N_26855);
nand U27423 (N_27423,N_26704,N_26558);
nand U27424 (N_27424,N_26801,N_26762);
nor U27425 (N_27425,N_26591,N_26791);
and U27426 (N_27426,N_26793,N_26969);
nand U27427 (N_27427,N_26735,N_26606);
and U27428 (N_27428,N_26587,N_26841);
nand U27429 (N_27429,N_26509,N_26712);
nand U27430 (N_27430,N_26778,N_26555);
or U27431 (N_27431,N_26969,N_26567);
xor U27432 (N_27432,N_26885,N_26929);
xor U27433 (N_27433,N_26540,N_26861);
and U27434 (N_27434,N_26788,N_26677);
nor U27435 (N_27435,N_26944,N_26562);
and U27436 (N_27436,N_26651,N_26658);
and U27437 (N_27437,N_26521,N_26758);
nor U27438 (N_27438,N_26746,N_26904);
nor U27439 (N_27439,N_26715,N_26605);
nor U27440 (N_27440,N_26828,N_26764);
or U27441 (N_27441,N_26534,N_26743);
and U27442 (N_27442,N_26719,N_26540);
xnor U27443 (N_27443,N_26739,N_26931);
or U27444 (N_27444,N_26702,N_26603);
xor U27445 (N_27445,N_26643,N_26907);
nand U27446 (N_27446,N_26583,N_26527);
or U27447 (N_27447,N_26690,N_26946);
xnor U27448 (N_27448,N_26938,N_26521);
and U27449 (N_27449,N_26622,N_26938);
xor U27450 (N_27450,N_26506,N_26783);
and U27451 (N_27451,N_26553,N_26637);
or U27452 (N_27452,N_26939,N_26758);
nand U27453 (N_27453,N_26942,N_26571);
xor U27454 (N_27454,N_26983,N_26658);
nand U27455 (N_27455,N_26713,N_26647);
and U27456 (N_27456,N_26517,N_26695);
and U27457 (N_27457,N_26599,N_26829);
nor U27458 (N_27458,N_26676,N_26957);
xnor U27459 (N_27459,N_26535,N_26554);
nand U27460 (N_27460,N_26843,N_26840);
or U27461 (N_27461,N_26705,N_26902);
xnor U27462 (N_27462,N_26703,N_26680);
nor U27463 (N_27463,N_26837,N_26650);
xor U27464 (N_27464,N_26712,N_26525);
nand U27465 (N_27465,N_26675,N_26718);
or U27466 (N_27466,N_26533,N_26706);
or U27467 (N_27467,N_26928,N_26891);
and U27468 (N_27468,N_26787,N_26878);
and U27469 (N_27469,N_26621,N_26907);
nand U27470 (N_27470,N_26799,N_26951);
and U27471 (N_27471,N_26500,N_26760);
and U27472 (N_27472,N_26984,N_26825);
or U27473 (N_27473,N_26863,N_26704);
xor U27474 (N_27474,N_26748,N_26705);
and U27475 (N_27475,N_26930,N_26711);
nor U27476 (N_27476,N_26673,N_26633);
nand U27477 (N_27477,N_26974,N_26807);
and U27478 (N_27478,N_26975,N_26878);
nand U27479 (N_27479,N_26775,N_26532);
nor U27480 (N_27480,N_26972,N_26958);
and U27481 (N_27481,N_26562,N_26830);
and U27482 (N_27482,N_26600,N_26727);
nand U27483 (N_27483,N_26587,N_26789);
nor U27484 (N_27484,N_26807,N_26703);
nor U27485 (N_27485,N_26791,N_26782);
nor U27486 (N_27486,N_26856,N_26608);
and U27487 (N_27487,N_26852,N_26805);
or U27488 (N_27488,N_26928,N_26760);
nand U27489 (N_27489,N_26748,N_26689);
or U27490 (N_27490,N_26852,N_26774);
and U27491 (N_27491,N_26562,N_26508);
nand U27492 (N_27492,N_26631,N_26680);
or U27493 (N_27493,N_26596,N_26910);
or U27494 (N_27494,N_26795,N_26906);
nor U27495 (N_27495,N_26893,N_26615);
xor U27496 (N_27496,N_26669,N_26967);
nand U27497 (N_27497,N_26574,N_26755);
xnor U27498 (N_27498,N_26818,N_26614);
and U27499 (N_27499,N_26737,N_26731);
nor U27500 (N_27500,N_27076,N_27294);
nor U27501 (N_27501,N_27266,N_27068);
or U27502 (N_27502,N_27232,N_27041);
or U27503 (N_27503,N_27421,N_27058);
nand U27504 (N_27504,N_27044,N_27430);
or U27505 (N_27505,N_27243,N_27022);
nand U27506 (N_27506,N_27316,N_27252);
or U27507 (N_27507,N_27340,N_27194);
or U27508 (N_27508,N_27391,N_27300);
nand U27509 (N_27509,N_27495,N_27173);
nand U27510 (N_27510,N_27370,N_27347);
nor U27511 (N_27511,N_27008,N_27464);
xor U27512 (N_27512,N_27496,N_27428);
or U27513 (N_27513,N_27024,N_27477);
xor U27514 (N_27514,N_27234,N_27062);
nor U27515 (N_27515,N_27450,N_27147);
nor U27516 (N_27516,N_27480,N_27124);
and U27517 (N_27517,N_27100,N_27228);
nand U27518 (N_27518,N_27424,N_27112);
or U27519 (N_27519,N_27235,N_27321);
or U27520 (N_27520,N_27431,N_27134);
xor U27521 (N_27521,N_27172,N_27113);
and U27522 (N_27522,N_27237,N_27333);
nor U27523 (N_27523,N_27186,N_27334);
and U27524 (N_27524,N_27407,N_27077);
and U27525 (N_27525,N_27032,N_27258);
or U27526 (N_27526,N_27141,N_27011);
xnor U27527 (N_27527,N_27305,N_27109);
nor U27528 (N_27528,N_27073,N_27225);
xnor U27529 (N_27529,N_27362,N_27295);
or U27530 (N_27530,N_27217,N_27314);
and U27531 (N_27531,N_27248,N_27196);
nor U27532 (N_27532,N_27129,N_27440);
and U27533 (N_27533,N_27467,N_27215);
and U27534 (N_27534,N_27045,N_27396);
nand U27535 (N_27535,N_27329,N_27437);
nor U27536 (N_27536,N_27455,N_27063);
and U27537 (N_27537,N_27048,N_27222);
or U27538 (N_27538,N_27326,N_27239);
nor U27539 (N_27539,N_27101,N_27142);
nand U27540 (N_27540,N_27102,N_27031);
nor U27541 (N_27541,N_27473,N_27274);
and U27542 (N_27542,N_27357,N_27490);
and U27543 (N_27543,N_27138,N_27488);
or U27544 (N_27544,N_27187,N_27303);
nand U27545 (N_27545,N_27461,N_27271);
and U27546 (N_27546,N_27210,N_27415);
and U27547 (N_27547,N_27259,N_27249);
or U27548 (N_27548,N_27349,N_27298);
or U27549 (N_27549,N_27075,N_27297);
and U27550 (N_27550,N_27290,N_27175);
nand U27551 (N_27551,N_27317,N_27111);
and U27552 (N_27552,N_27251,N_27498);
and U27553 (N_27553,N_27261,N_27449);
xor U27554 (N_27554,N_27443,N_27025);
and U27555 (N_27555,N_27016,N_27414);
and U27556 (N_27556,N_27466,N_27307);
xor U27557 (N_27557,N_27352,N_27148);
or U27558 (N_27558,N_27462,N_27264);
xnor U27559 (N_27559,N_27236,N_27154);
nor U27560 (N_27560,N_27398,N_27131);
nand U27561 (N_27561,N_27103,N_27468);
nor U27562 (N_27562,N_27211,N_27390);
and U27563 (N_27563,N_27474,N_27319);
nor U27564 (N_27564,N_27409,N_27465);
xor U27565 (N_27565,N_27074,N_27238);
xnor U27566 (N_27566,N_27007,N_27214);
and U27567 (N_27567,N_27284,N_27056);
and U27568 (N_27568,N_27345,N_27223);
nand U27569 (N_27569,N_27156,N_27192);
and U27570 (N_27570,N_27209,N_27489);
nand U27571 (N_27571,N_27050,N_27218);
or U27572 (N_27572,N_27085,N_27036);
nor U27573 (N_27573,N_27081,N_27272);
and U27574 (N_27574,N_27145,N_27023);
nor U27575 (N_27575,N_27402,N_27339);
and U27576 (N_27576,N_27393,N_27457);
xor U27577 (N_27577,N_27379,N_27166);
or U27578 (N_27578,N_27318,N_27312);
and U27579 (N_27579,N_27019,N_27481);
or U27580 (N_27580,N_27230,N_27342);
xor U27581 (N_27581,N_27372,N_27286);
and U27582 (N_27582,N_27091,N_27373);
and U27583 (N_27583,N_27220,N_27322);
nor U27584 (N_27584,N_27219,N_27446);
or U27585 (N_27585,N_27479,N_27423);
nor U27586 (N_27586,N_27400,N_27323);
nand U27587 (N_27587,N_27184,N_27163);
nor U27588 (N_27588,N_27009,N_27208);
and U27589 (N_27589,N_27207,N_27039);
nand U27590 (N_27590,N_27201,N_27010);
nor U27591 (N_27591,N_27059,N_27348);
and U27592 (N_27592,N_27486,N_27065);
nand U27593 (N_27593,N_27277,N_27253);
nand U27594 (N_27594,N_27199,N_27283);
nand U27595 (N_27595,N_27090,N_27381);
nand U27596 (N_27596,N_27397,N_27389);
nand U27597 (N_27597,N_27125,N_27497);
nand U27598 (N_27598,N_27399,N_27313);
nand U27599 (N_27599,N_27107,N_27463);
and U27600 (N_27600,N_27046,N_27188);
and U27601 (N_27601,N_27374,N_27089);
nand U27602 (N_27602,N_27365,N_27469);
or U27603 (N_27603,N_27263,N_27247);
xor U27604 (N_27604,N_27320,N_27413);
nand U27605 (N_27605,N_27071,N_27012);
and U27606 (N_27606,N_27123,N_27441);
or U27607 (N_27607,N_27351,N_27086);
and U27608 (N_27608,N_27080,N_27136);
nand U27609 (N_27609,N_27038,N_27110);
nand U27610 (N_27610,N_27296,N_27410);
nand U27611 (N_27611,N_27132,N_27191);
nand U27612 (N_27612,N_27387,N_27478);
and U27613 (N_27613,N_27030,N_27151);
nand U27614 (N_27614,N_27057,N_27096);
or U27615 (N_27615,N_27176,N_27120);
nor U27616 (N_27616,N_27422,N_27097);
xor U27617 (N_27617,N_27419,N_27162);
xnor U27618 (N_27618,N_27435,N_27104);
nand U27619 (N_27619,N_27153,N_27203);
nand U27620 (N_27620,N_27354,N_27310);
xor U27621 (N_27621,N_27161,N_27099);
and U27622 (N_27622,N_27335,N_27447);
xnor U27623 (N_27623,N_27426,N_27105);
xnor U27624 (N_27624,N_27279,N_27233);
xnor U27625 (N_27625,N_27051,N_27137);
or U27626 (N_27626,N_27392,N_27020);
or U27627 (N_27627,N_27336,N_27287);
nand U27628 (N_27628,N_27382,N_27492);
or U27629 (N_27629,N_27453,N_27052);
nor U27630 (N_27630,N_27363,N_27257);
nor U27631 (N_27631,N_27325,N_27043);
nor U27632 (N_27632,N_27241,N_27394);
or U27633 (N_27633,N_27405,N_27360);
xor U27634 (N_27634,N_27119,N_27002);
xnor U27635 (N_27635,N_27427,N_27017);
nor U27636 (N_27636,N_27343,N_27353);
and U27637 (N_27637,N_27088,N_27095);
or U27638 (N_27638,N_27484,N_27282);
xnor U27639 (N_27639,N_27164,N_27406);
xnor U27640 (N_27640,N_27106,N_27037);
and U27641 (N_27641,N_27006,N_27311);
nand U27642 (N_27642,N_27338,N_27122);
nor U27643 (N_27643,N_27448,N_27491);
and U27644 (N_27644,N_27344,N_27130);
xor U27645 (N_27645,N_27281,N_27383);
xnor U27646 (N_27646,N_27371,N_27035);
nand U27647 (N_27647,N_27034,N_27047);
and U27648 (N_27648,N_27359,N_27304);
xnor U27649 (N_27649,N_27231,N_27366);
nand U27650 (N_27650,N_27337,N_27451);
and U27651 (N_27651,N_27028,N_27053);
or U27652 (N_27652,N_27180,N_27302);
or U27653 (N_27653,N_27289,N_27254);
xnor U27654 (N_27654,N_27408,N_27301);
and U27655 (N_27655,N_27412,N_27442);
nor U27656 (N_27656,N_27270,N_27395);
and U27657 (N_27657,N_27168,N_27240);
or U27658 (N_27658,N_27380,N_27471);
nor U27659 (N_27659,N_27499,N_27268);
and U27660 (N_27660,N_27149,N_27079);
or U27661 (N_27661,N_27386,N_27309);
and U27662 (N_27662,N_27403,N_27157);
nor U27663 (N_27663,N_27328,N_27355);
nand U27664 (N_27664,N_27139,N_27346);
and U27665 (N_27665,N_27143,N_27385);
nand U27666 (N_27666,N_27055,N_27278);
xnor U27667 (N_27667,N_27388,N_27434);
xnor U27668 (N_27668,N_27367,N_27364);
or U27669 (N_27669,N_27144,N_27072);
xor U27670 (N_27670,N_27273,N_27444);
or U27671 (N_27671,N_27021,N_27299);
xor U27672 (N_27672,N_27064,N_27356);
nand U27673 (N_27673,N_27256,N_27040);
or U27674 (N_27674,N_27061,N_27094);
nand U27675 (N_27675,N_27146,N_27160);
and U27676 (N_27676,N_27418,N_27001);
nand U27677 (N_27677,N_27350,N_27202);
nand U27678 (N_27678,N_27369,N_27093);
or U27679 (N_27679,N_27229,N_27114);
xnor U27680 (N_27680,N_27221,N_27165);
nor U27681 (N_27681,N_27375,N_27368);
xor U27682 (N_27682,N_27190,N_27330);
nor U27683 (N_27683,N_27005,N_27445);
or U27684 (N_27684,N_27004,N_27429);
xnor U27685 (N_27685,N_27332,N_27262);
and U27686 (N_27686,N_27452,N_27027);
and U27687 (N_27687,N_27476,N_27069);
nand U27688 (N_27688,N_27015,N_27331);
nor U27689 (N_27689,N_27432,N_27033);
xnor U27690 (N_27690,N_27060,N_27189);
and U27691 (N_27691,N_27459,N_27018);
nand U27692 (N_27692,N_27242,N_27378);
and U27693 (N_27693,N_27205,N_27288);
and U27694 (N_27694,N_27460,N_27159);
xor U27695 (N_27695,N_27185,N_27197);
nand U27696 (N_27696,N_27000,N_27250);
xnor U27697 (N_27697,N_27438,N_27003);
and U27698 (N_27698,N_27275,N_27485);
and U27699 (N_27699,N_27054,N_27026);
nand U27700 (N_27700,N_27170,N_27013);
nand U27701 (N_27701,N_27133,N_27384);
nand U27702 (N_27702,N_27265,N_27245);
nand U27703 (N_27703,N_27127,N_27226);
nor U27704 (N_27704,N_27213,N_27483);
nand U27705 (N_27705,N_27494,N_27315);
nor U27706 (N_27706,N_27292,N_27014);
nand U27707 (N_27707,N_27291,N_27183);
xnor U27708 (N_27708,N_27404,N_27126);
nor U27709 (N_27709,N_27082,N_27327);
nand U27710 (N_27710,N_27193,N_27195);
nand U27711 (N_27711,N_27482,N_27285);
and U27712 (N_27712,N_27216,N_27493);
or U27713 (N_27713,N_27420,N_27454);
nand U27714 (N_27714,N_27084,N_27425);
or U27715 (N_27715,N_27198,N_27260);
nand U27716 (N_27716,N_27377,N_27150);
nor U27717 (N_27717,N_27152,N_27411);
nand U27718 (N_27718,N_27135,N_27181);
xnor U27719 (N_27719,N_27171,N_27244);
or U27720 (N_27720,N_27155,N_27224);
and U27721 (N_27721,N_27049,N_27456);
and U27722 (N_27722,N_27174,N_27115);
nand U27723 (N_27723,N_27341,N_27066);
or U27724 (N_27724,N_27255,N_27167);
nand U27725 (N_27725,N_27267,N_27269);
or U27726 (N_27726,N_27179,N_27361);
or U27727 (N_27727,N_27116,N_27070);
xnor U27728 (N_27728,N_27472,N_27293);
nor U27729 (N_27729,N_27324,N_27087);
or U27730 (N_27730,N_27458,N_27308);
or U27731 (N_27731,N_27475,N_27276);
nor U27732 (N_27732,N_27067,N_27487);
nand U27733 (N_27733,N_27092,N_27169);
nor U27734 (N_27734,N_27121,N_27433);
nor U27735 (N_27735,N_27439,N_27140);
nand U27736 (N_27736,N_27470,N_27246);
xnor U27737 (N_27737,N_27306,N_27083);
and U27738 (N_27738,N_27280,N_27436);
nor U27739 (N_27739,N_27376,N_27128);
or U27740 (N_27740,N_27212,N_27042);
nor U27741 (N_27741,N_27178,N_27098);
nor U27742 (N_27742,N_27078,N_27417);
nand U27743 (N_27743,N_27177,N_27401);
nor U27744 (N_27744,N_27227,N_27117);
xnor U27745 (N_27745,N_27358,N_27158);
nor U27746 (N_27746,N_27416,N_27200);
or U27747 (N_27747,N_27206,N_27182);
nor U27748 (N_27748,N_27204,N_27108);
xnor U27749 (N_27749,N_27029,N_27118);
nand U27750 (N_27750,N_27231,N_27380);
and U27751 (N_27751,N_27404,N_27186);
nand U27752 (N_27752,N_27083,N_27402);
xnor U27753 (N_27753,N_27162,N_27305);
and U27754 (N_27754,N_27105,N_27182);
or U27755 (N_27755,N_27406,N_27370);
and U27756 (N_27756,N_27432,N_27330);
nand U27757 (N_27757,N_27304,N_27417);
and U27758 (N_27758,N_27291,N_27437);
nor U27759 (N_27759,N_27482,N_27215);
xnor U27760 (N_27760,N_27383,N_27176);
nand U27761 (N_27761,N_27425,N_27445);
xor U27762 (N_27762,N_27331,N_27171);
nor U27763 (N_27763,N_27385,N_27270);
and U27764 (N_27764,N_27332,N_27057);
and U27765 (N_27765,N_27333,N_27098);
xnor U27766 (N_27766,N_27195,N_27140);
nor U27767 (N_27767,N_27086,N_27312);
and U27768 (N_27768,N_27498,N_27329);
nand U27769 (N_27769,N_27418,N_27197);
and U27770 (N_27770,N_27094,N_27376);
or U27771 (N_27771,N_27425,N_27346);
xnor U27772 (N_27772,N_27219,N_27398);
nand U27773 (N_27773,N_27341,N_27387);
nor U27774 (N_27774,N_27302,N_27204);
nor U27775 (N_27775,N_27053,N_27058);
or U27776 (N_27776,N_27147,N_27117);
nor U27777 (N_27777,N_27431,N_27035);
and U27778 (N_27778,N_27058,N_27129);
xor U27779 (N_27779,N_27132,N_27291);
xor U27780 (N_27780,N_27279,N_27113);
nor U27781 (N_27781,N_27052,N_27472);
or U27782 (N_27782,N_27294,N_27081);
xor U27783 (N_27783,N_27158,N_27023);
nand U27784 (N_27784,N_27166,N_27128);
and U27785 (N_27785,N_27342,N_27365);
and U27786 (N_27786,N_27413,N_27493);
xor U27787 (N_27787,N_27118,N_27285);
or U27788 (N_27788,N_27404,N_27271);
xnor U27789 (N_27789,N_27046,N_27458);
or U27790 (N_27790,N_27003,N_27317);
nand U27791 (N_27791,N_27440,N_27486);
xnor U27792 (N_27792,N_27055,N_27320);
xnor U27793 (N_27793,N_27034,N_27348);
or U27794 (N_27794,N_27355,N_27200);
and U27795 (N_27795,N_27199,N_27438);
nand U27796 (N_27796,N_27179,N_27216);
xnor U27797 (N_27797,N_27446,N_27288);
nand U27798 (N_27798,N_27327,N_27354);
or U27799 (N_27799,N_27372,N_27183);
or U27800 (N_27800,N_27264,N_27239);
nor U27801 (N_27801,N_27063,N_27143);
and U27802 (N_27802,N_27109,N_27205);
nand U27803 (N_27803,N_27235,N_27074);
nor U27804 (N_27804,N_27077,N_27494);
nand U27805 (N_27805,N_27384,N_27089);
and U27806 (N_27806,N_27103,N_27362);
or U27807 (N_27807,N_27429,N_27252);
or U27808 (N_27808,N_27381,N_27276);
or U27809 (N_27809,N_27222,N_27011);
nor U27810 (N_27810,N_27463,N_27231);
nor U27811 (N_27811,N_27205,N_27417);
nor U27812 (N_27812,N_27176,N_27195);
xnor U27813 (N_27813,N_27136,N_27305);
nand U27814 (N_27814,N_27383,N_27155);
nand U27815 (N_27815,N_27225,N_27280);
and U27816 (N_27816,N_27193,N_27276);
xnor U27817 (N_27817,N_27389,N_27266);
or U27818 (N_27818,N_27341,N_27082);
or U27819 (N_27819,N_27443,N_27100);
or U27820 (N_27820,N_27290,N_27292);
and U27821 (N_27821,N_27098,N_27225);
nand U27822 (N_27822,N_27416,N_27387);
and U27823 (N_27823,N_27347,N_27489);
or U27824 (N_27824,N_27130,N_27380);
nand U27825 (N_27825,N_27353,N_27481);
xnor U27826 (N_27826,N_27407,N_27356);
nor U27827 (N_27827,N_27275,N_27144);
xnor U27828 (N_27828,N_27357,N_27437);
xnor U27829 (N_27829,N_27270,N_27179);
xnor U27830 (N_27830,N_27018,N_27353);
xor U27831 (N_27831,N_27425,N_27188);
xnor U27832 (N_27832,N_27394,N_27486);
xor U27833 (N_27833,N_27291,N_27104);
and U27834 (N_27834,N_27010,N_27184);
nor U27835 (N_27835,N_27267,N_27035);
xor U27836 (N_27836,N_27448,N_27094);
nand U27837 (N_27837,N_27477,N_27396);
and U27838 (N_27838,N_27338,N_27045);
and U27839 (N_27839,N_27053,N_27061);
nand U27840 (N_27840,N_27153,N_27482);
nor U27841 (N_27841,N_27179,N_27124);
nor U27842 (N_27842,N_27166,N_27292);
nand U27843 (N_27843,N_27358,N_27116);
or U27844 (N_27844,N_27048,N_27497);
nor U27845 (N_27845,N_27429,N_27363);
nand U27846 (N_27846,N_27161,N_27209);
and U27847 (N_27847,N_27399,N_27153);
nand U27848 (N_27848,N_27061,N_27273);
xnor U27849 (N_27849,N_27413,N_27411);
xnor U27850 (N_27850,N_27342,N_27160);
and U27851 (N_27851,N_27458,N_27480);
and U27852 (N_27852,N_27094,N_27371);
nor U27853 (N_27853,N_27245,N_27145);
or U27854 (N_27854,N_27208,N_27019);
or U27855 (N_27855,N_27433,N_27031);
xor U27856 (N_27856,N_27299,N_27040);
nand U27857 (N_27857,N_27135,N_27068);
nand U27858 (N_27858,N_27373,N_27311);
nor U27859 (N_27859,N_27012,N_27354);
and U27860 (N_27860,N_27333,N_27145);
nand U27861 (N_27861,N_27335,N_27310);
or U27862 (N_27862,N_27125,N_27349);
xor U27863 (N_27863,N_27222,N_27128);
xor U27864 (N_27864,N_27187,N_27130);
xnor U27865 (N_27865,N_27330,N_27425);
xor U27866 (N_27866,N_27140,N_27147);
xor U27867 (N_27867,N_27208,N_27265);
nor U27868 (N_27868,N_27251,N_27438);
nor U27869 (N_27869,N_27183,N_27095);
and U27870 (N_27870,N_27371,N_27191);
xor U27871 (N_27871,N_27385,N_27414);
nand U27872 (N_27872,N_27324,N_27241);
nor U27873 (N_27873,N_27074,N_27451);
nor U27874 (N_27874,N_27382,N_27370);
or U27875 (N_27875,N_27064,N_27122);
xnor U27876 (N_27876,N_27200,N_27226);
xnor U27877 (N_27877,N_27011,N_27157);
nor U27878 (N_27878,N_27044,N_27250);
nor U27879 (N_27879,N_27237,N_27053);
and U27880 (N_27880,N_27124,N_27319);
nor U27881 (N_27881,N_27400,N_27303);
and U27882 (N_27882,N_27411,N_27190);
nand U27883 (N_27883,N_27366,N_27159);
nand U27884 (N_27884,N_27055,N_27152);
xnor U27885 (N_27885,N_27136,N_27249);
nand U27886 (N_27886,N_27271,N_27024);
or U27887 (N_27887,N_27070,N_27198);
nor U27888 (N_27888,N_27461,N_27169);
nor U27889 (N_27889,N_27168,N_27104);
xnor U27890 (N_27890,N_27068,N_27295);
xnor U27891 (N_27891,N_27378,N_27112);
nand U27892 (N_27892,N_27122,N_27381);
or U27893 (N_27893,N_27439,N_27119);
nand U27894 (N_27894,N_27391,N_27375);
or U27895 (N_27895,N_27337,N_27424);
or U27896 (N_27896,N_27487,N_27011);
or U27897 (N_27897,N_27463,N_27235);
and U27898 (N_27898,N_27136,N_27213);
and U27899 (N_27899,N_27461,N_27198);
nand U27900 (N_27900,N_27475,N_27251);
and U27901 (N_27901,N_27363,N_27139);
xnor U27902 (N_27902,N_27257,N_27322);
xnor U27903 (N_27903,N_27137,N_27223);
or U27904 (N_27904,N_27236,N_27320);
nor U27905 (N_27905,N_27197,N_27449);
and U27906 (N_27906,N_27271,N_27052);
nand U27907 (N_27907,N_27029,N_27079);
nand U27908 (N_27908,N_27264,N_27087);
xnor U27909 (N_27909,N_27251,N_27083);
nor U27910 (N_27910,N_27442,N_27213);
nor U27911 (N_27911,N_27425,N_27490);
or U27912 (N_27912,N_27306,N_27209);
or U27913 (N_27913,N_27375,N_27321);
xnor U27914 (N_27914,N_27316,N_27447);
or U27915 (N_27915,N_27492,N_27226);
nand U27916 (N_27916,N_27291,N_27266);
and U27917 (N_27917,N_27329,N_27190);
and U27918 (N_27918,N_27456,N_27211);
or U27919 (N_27919,N_27166,N_27022);
and U27920 (N_27920,N_27211,N_27162);
and U27921 (N_27921,N_27029,N_27157);
and U27922 (N_27922,N_27464,N_27051);
nor U27923 (N_27923,N_27023,N_27294);
nand U27924 (N_27924,N_27451,N_27291);
nand U27925 (N_27925,N_27497,N_27115);
and U27926 (N_27926,N_27419,N_27038);
nand U27927 (N_27927,N_27287,N_27144);
or U27928 (N_27928,N_27390,N_27397);
and U27929 (N_27929,N_27275,N_27220);
and U27930 (N_27930,N_27234,N_27179);
nand U27931 (N_27931,N_27473,N_27498);
xor U27932 (N_27932,N_27291,N_27233);
nand U27933 (N_27933,N_27416,N_27251);
nand U27934 (N_27934,N_27338,N_27252);
nand U27935 (N_27935,N_27343,N_27454);
and U27936 (N_27936,N_27074,N_27224);
nor U27937 (N_27937,N_27162,N_27260);
xor U27938 (N_27938,N_27385,N_27338);
nand U27939 (N_27939,N_27385,N_27483);
and U27940 (N_27940,N_27299,N_27093);
nand U27941 (N_27941,N_27453,N_27498);
and U27942 (N_27942,N_27199,N_27317);
and U27943 (N_27943,N_27420,N_27199);
or U27944 (N_27944,N_27450,N_27127);
nor U27945 (N_27945,N_27434,N_27064);
or U27946 (N_27946,N_27261,N_27107);
nor U27947 (N_27947,N_27047,N_27344);
or U27948 (N_27948,N_27413,N_27265);
and U27949 (N_27949,N_27133,N_27167);
nor U27950 (N_27950,N_27086,N_27180);
nor U27951 (N_27951,N_27455,N_27338);
nor U27952 (N_27952,N_27422,N_27150);
nand U27953 (N_27953,N_27042,N_27245);
or U27954 (N_27954,N_27256,N_27438);
nand U27955 (N_27955,N_27076,N_27015);
nand U27956 (N_27956,N_27419,N_27354);
nor U27957 (N_27957,N_27290,N_27418);
nor U27958 (N_27958,N_27275,N_27161);
or U27959 (N_27959,N_27317,N_27268);
and U27960 (N_27960,N_27112,N_27380);
nor U27961 (N_27961,N_27320,N_27336);
nor U27962 (N_27962,N_27026,N_27419);
or U27963 (N_27963,N_27298,N_27161);
nand U27964 (N_27964,N_27396,N_27439);
or U27965 (N_27965,N_27391,N_27004);
and U27966 (N_27966,N_27415,N_27342);
nand U27967 (N_27967,N_27279,N_27182);
xnor U27968 (N_27968,N_27092,N_27460);
xor U27969 (N_27969,N_27487,N_27127);
nand U27970 (N_27970,N_27199,N_27001);
nand U27971 (N_27971,N_27372,N_27411);
nor U27972 (N_27972,N_27181,N_27308);
xor U27973 (N_27973,N_27457,N_27301);
or U27974 (N_27974,N_27369,N_27120);
nand U27975 (N_27975,N_27268,N_27091);
nand U27976 (N_27976,N_27472,N_27073);
or U27977 (N_27977,N_27242,N_27425);
xor U27978 (N_27978,N_27352,N_27460);
and U27979 (N_27979,N_27211,N_27143);
nor U27980 (N_27980,N_27002,N_27026);
xor U27981 (N_27981,N_27094,N_27003);
and U27982 (N_27982,N_27219,N_27273);
nor U27983 (N_27983,N_27180,N_27285);
nor U27984 (N_27984,N_27366,N_27052);
nor U27985 (N_27985,N_27149,N_27481);
nor U27986 (N_27986,N_27093,N_27363);
or U27987 (N_27987,N_27011,N_27276);
and U27988 (N_27988,N_27368,N_27086);
or U27989 (N_27989,N_27490,N_27106);
nand U27990 (N_27990,N_27008,N_27425);
nor U27991 (N_27991,N_27457,N_27007);
nand U27992 (N_27992,N_27182,N_27034);
and U27993 (N_27993,N_27035,N_27395);
nor U27994 (N_27994,N_27264,N_27410);
xnor U27995 (N_27995,N_27435,N_27192);
xnor U27996 (N_27996,N_27263,N_27472);
or U27997 (N_27997,N_27459,N_27082);
or U27998 (N_27998,N_27114,N_27275);
or U27999 (N_27999,N_27043,N_27060);
and U28000 (N_28000,N_27604,N_27795);
or U28001 (N_28001,N_27890,N_27928);
xnor U28002 (N_28002,N_27689,N_27757);
and U28003 (N_28003,N_27512,N_27977);
nand U28004 (N_28004,N_27916,N_27637);
nor U28005 (N_28005,N_27675,N_27834);
nor U28006 (N_28006,N_27550,N_27628);
or U28007 (N_28007,N_27863,N_27558);
xnor U28008 (N_28008,N_27679,N_27816);
nor U28009 (N_28009,N_27656,N_27930);
or U28010 (N_28010,N_27767,N_27555);
nor U28011 (N_28011,N_27784,N_27931);
or U28012 (N_28012,N_27765,N_27773);
or U28013 (N_28013,N_27941,N_27501);
xnor U28014 (N_28014,N_27542,N_27797);
and U28015 (N_28015,N_27812,N_27715);
or U28016 (N_28016,N_27774,N_27838);
nand U28017 (N_28017,N_27859,N_27900);
or U28018 (N_28018,N_27504,N_27731);
or U28019 (N_28019,N_27877,N_27851);
xnor U28020 (N_28020,N_27578,N_27721);
nand U28021 (N_28021,N_27945,N_27948);
or U28022 (N_28022,N_27623,N_27577);
xor U28023 (N_28023,N_27821,N_27580);
nand U28024 (N_28024,N_27707,N_27647);
and U28025 (N_28025,N_27989,N_27994);
and U28026 (N_28026,N_27673,N_27665);
nand U28027 (N_28027,N_27563,N_27828);
xnor U28028 (N_28028,N_27841,N_27925);
or U28029 (N_28029,N_27714,N_27786);
and U28030 (N_28030,N_27984,N_27964);
and U28031 (N_28031,N_27858,N_27734);
nor U28032 (N_28032,N_27852,N_27516);
xor U28033 (N_28033,N_27571,N_27593);
nand U28034 (N_28034,N_27870,N_27617);
xor U28035 (N_28035,N_27547,N_27719);
and U28036 (N_28036,N_27517,N_27789);
nor U28037 (N_28037,N_27680,N_27947);
xor U28038 (N_28038,N_27832,N_27836);
nand U28039 (N_28039,N_27709,N_27760);
or U28040 (N_28040,N_27692,N_27686);
and U28041 (N_28041,N_27521,N_27750);
xnor U28042 (N_28042,N_27701,N_27942);
nand U28043 (N_28043,N_27531,N_27515);
nor U28044 (N_28044,N_27952,N_27729);
nor U28045 (N_28045,N_27581,N_27813);
or U28046 (N_28046,N_27988,N_27597);
or U28047 (N_28047,N_27728,N_27814);
or U28048 (N_28048,N_27724,N_27579);
nand U28049 (N_28049,N_27658,N_27536);
and U28050 (N_28050,N_27929,N_27857);
or U28051 (N_28051,N_27888,N_27557);
nand U28052 (N_28052,N_27969,N_27749);
or U28053 (N_28053,N_27631,N_27599);
nor U28054 (N_28054,N_27741,N_27520);
xor U28055 (N_28055,N_27856,N_27509);
nor U28056 (N_28056,N_27913,N_27766);
nand U28057 (N_28057,N_27510,N_27798);
and U28058 (N_28058,N_27691,N_27817);
xnor U28059 (N_28059,N_27533,N_27668);
nor U28060 (N_28060,N_27848,N_27576);
xnor U28061 (N_28061,N_27583,N_27666);
nor U28062 (N_28062,N_27763,N_27805);
or U28063 (N_28063,N_27960,N_27950);
nand U28064 (N_28064,N_27730,N_27713);
or U28065 (N_28065,N_27602,N_27867);
nor U28066 (N_28066,N_27825,N_27582);
nor U28067 (N_28067,N_27710,N_27985);
nor U28068 (N_28068,N_27847,N_27955);
or U28069 (N_28069,N_27899,N_27869);
nor U28070 (N_28070,N_27954,N_27683);
nand U28071 (N_28071,N_27585,N_27840);
and U28072 (N_28072,N_27589,N_27824);
and U28073 (N_28073,N_27973,N_27635);
and U28074 (N_28074,N_27733,N_27562);
xor U28075 (N_28075,N_27905,N_27785);
and U28076 (N_28076,N_27561,N_27554);
or U28077 (N_28077,N_27829,N_27712);
nand U28078 (N_28078,N_27755,N_27696);
xor U28079 (N_28079,N_27779,N_27999);
xnor U28080 (N_28080,N_27541,N_27747);
and U28081 (N_28081,N_27826,N_27519);
nand U28082 (N_28082,N_27889,N_27539);
and U28083 (N_28083,N_27971,N_27986);
nand U28084 (N_28084,N_27753,N_27921);
nor U28085 (N_28085,N_27634,N_27803);
nor U28086 (N_28086,N_27914,N_27564);
and U28087 (N_28087,N_27574,N_27670);
or U28088 (N_28088,N_27871,N_27792);
and U28089 (N_28089,N_27968,N_27982);
and U28090 (N_28090,N_27855,N_27887);
nor U28091 (N_28091,N_27804,N_27746);
or U28092 (N_28092,N_27743,N_27874);
nand U28093 (N_28093,N_27983,N_27676);
and U28094 (N_28094,N_27860,N_27892);
or U28095 (N_28095,N_27752,N_27891);
and U28096 (N_28096,N_27638,N_27782);
or U28097 (N_28097,N_27565,N_27646);
nor U28098 (N_28098,N_27671,N_27991);
or U28099 (N_28099,N_27917,N_27791);
nor U28100 (N_28100,N_27944,N_27610);
or U28101 (N_28101,N_27970,N_27567);
and U28102 (N_28102,N_27699,N_27551);
or U28103 (N_28103,N_27837,N_27649);
xnor U28104 (N_28104,N_27653,N_27961);
and U28105 (N_28105,N_27500,N_27875);
nand U28106 (N_28106,N_27695,N_27811);
or U28107 (N_28107,N_27807,N_27920);
nor U28108 (N_28108,N_27936,N_27919);
nand U28109 (N_28109,N_27976,N_27559);
nand U28110 (N_28110,N_27702,N_27842);
and U28111 (N_28111,N_27513,N_27768);
nand U28112 (N_28112,N_27600,N_27967);
xnor U28113 (N_28113,N_27619,N_27636);
nand U28114 (N_28114,N_27725,N_27940);
xor U28115 (N_28115,N_27751,N_27595);
nor U28116 (N_28116,N_27980,N_27775);
nor U28117 (N_28117,N_27934,N_27885);
xnor U28118 (N_28118,N_27831,N_27962);
nor U28119 (N_28119,N_27545,N_27737);
nand U28120 (N_28120,N_27607,N_27758);
and U28121 (N_28121,N_27932,N_27735);
or U28122 (N_28122,N_27681,N_27528);
or U28123 (N_28123,N_27606,N_27690);
and U28124 (N_28124,N_27896,N_27915);
nor U28125 (N_28125,N_27839,N_27981);
nor U28126 (N_28126,N_27800,N_27845);
nand U28127 (N_28127,N_27663,N_27759);
nor U28128 (N_28128,N_27639,N_27902);
nand U28129 (N_28129,N_27548,N_27694);
nor U28130 (N_28130,N_27793,N_27939);
or U28131 (N_28131,N_27998,N_27777);
xor U28132 (N_28132,N_27864,N_27909);
nor U28133 (N_28133,N_27727,N_27799);
nand U28134 (N_28134,N_27861,N_27553);
xnor U28135 (N_28135,N_27878,N_27620);
xnor U28136 (N_28136,N_27544,N_27951);
nor U28137 (N_28137,N_27794,N_27873);
nor U28138 (N_28138,N_27972,N_27966);
and U28139 (N_28139,N_27632,N_27505);
xor U28140 (N_28140,N_27661,N_27537);
xor U28141 (N_28141,N_27503,N_27996);
and U28142 (N_28142,N_27876,N_27979);
xor U28143 (N_28143,N_27720,N_27990);
or U28144 (N_28144,N_27657,N_27872);
nand U28145 (N_28145,N_27995,N_27974);
and U28146 (N_28146,N_27933,N_27570);
and U28147 (N_28147,N_27953,N_27823);
nand U28148 (N_28148,N_27808,N_27640);
nor U28149 (N_28149,N_27608,N_27862);
nor U28150 (N_28150,N_27687,N_27693);
nor U28151 (N_28151,N_27927,N_27527);
and U28152 (N_28152,N_27802,N_27609);
nor U28153 (N_28153,N_27522,N_27624);
xnor U28154 (N_28154,N_27601,N_27901);
and U28155 (N_28155,N_27603,N_27506);
and U28156 (N_28156,N_27588,N_27507);
or U28157 (N_28157,N_27654,N_27780);
nand U28158 (N_28158,N_27820,N_27771);
nor U28159 (N_28159,N_27770,N_27854);
nand U28160 (N_28160,N_27822,N_27987);
nand U28161 (N_28161,N_27659,N_27810);
or U28162 (N_28162,N_27672,N_27756);
and U28163 (N_28163,N_27651,N_27534);
or U28164 (N_28164,N_27796,N_27575);
nand U28165 (N_28165,N_27778,N_27844);
nand U28166 (N_28166,N_27963,N_27716);
nand U28167 (N_28167,N_27612,N_27833);
nand U28168 (N_28168,N_27865,N_27903);
or U28169 (N_28169,N_27573,N_27523);
nor U28170 (N_28170,N_27879,N_27662);
or U28171 (N_28171,N_27627,N_27697);
nor U28172 (N_28172,N_27742,N_27809);
xor U28173 (N_28173,N_27641,N_27868);
xnor U28174 (N_28174,N_27776,N_27700);
or U28175 (N_28175,N_27764,N_27884);
nand U28176 (N_28176,N_27508,N_27723);
or U28177 (N_28177,N_27738,N_27846);
or U28178 (N_28178,N_27529,N_27975);
and U28179 (N_28179,N_27898,N_27806);
nand U28180 (N_28180,N_27978,N_27586);
nor U28181 (N_28181,N_27923,N_27655);
or U28182 (N_28182,N_27605,N_27590);
or U28183 (N_28183,N_27938,N_27530);
nand U28184 (N_28184,N_27706,N_27918);
and U28185 (N_28185,N_27664,N_27748);
and U28186 (N_28186,N_27788,N_27642);
or U28187 (N_28187,N_27790,N_27678);
or U28188 (N_28188,N_27815,N_27698);
xnor U28189 (N_28189,N_27549,N_27611);
xor U28190 (N_28190,N_27880,N_27912);
xor U28191 (N_28191,N_27532,N_27621);
nand U28192 (N_28192,N_27625,N_27958);
and U28193 (N_28193,N_27568,N_27943);
xor U28194 (N_28194,N_27897,N_27959);
nand U28195 (N_28195,N_27946,N_27911);
or U28196 (N_28196,N_27652,N_27907);
nor U28197 (N_28197,N_27540,N_27718);
nand U28198 (N_28198,N_27740,N_27924);
xnor U28199 (N_28199,N_27626,N_27717);
or U28200 (N_28200,N_27783,N_27648);
or U28201 (N_28201,N_27922,N_27524);
or U28202 (N_28202,N_27704,N_27643);
and U28203 (N_28203,N_27592,N_27937);
and U28204 (N_28204,N_27615,N_27881);
nor U28205 (N_28205,N_27630,N_27965);
nor U28206 (N_28206,N_27762,N_27525);
nand U28207 (N_28207,N_27739,N_27883);
xor U28208 (N_28208,N_27526,N_27732);
or U28209 (N_28209,N_27801,N_27781);
nor U28210 (N_28210,N_27674,N_27556);
and U28211 (N_28211,N_27787,N_27598);
nand U28212 (N_28212,N_27514,N_27853);
nand U28213 (N_28213,N_27761,N_27518);
and U28214 (N_28214,N_27849,N_27754);
nand U28215 (N_28215,N_27895,N_27682);
xnor U28216 (N_28216,N_27543,N_27669);
and U28217 (N_28217,N_27622,N_27818);
and U28218 (N_28218,N_27722,N_27629);
nand U28219 (N_28219,N_27584,N_27819);
nand U28220 (N_28220,N_27502,N_27618);
nand U28221 (N_28221,N_27906,N_27957);
nor U28222 (N_28222,N_27511,N_27935);
xnor U28223 (N_28223,N_27736,N_27908);
or U28224 (N_28224,N_27616,N_27614);
and U28225 (N_28225,N_27745,N_27546);
or U28226 (N_28226,N_27769,N_27882);
or U28227 (N_28227,N_27910,N_27850);
or U28228 (N_28228,N_27667,N_27572);
nand U28229 (N_28229,N_27685,N_27949);
or U28230 (N_28230,N_27830,N_27744);
xnor U28231 (N_28231,N_27591,N_27644);
and U28232 (N_28232,N_27535,N_27569);
nor U28233 (N_28233,N_27660,N_27726);
or U28234 (N_28234,N_27587,N_27538);
xor U28235 (N_28235,N_27866,N_27708);
and U28236 (N_28236,N_27711,N_27677);
and U28237 (N_28237,N_27566,N_27893);
and U28238 (N_28238,N_27992,N_27993);
nor U28239 (N_28239,N_27596,N_27835);
nand U28240 (N_28240,N_27633,N_27703);
xor U28241 (N_28241,N_27688,N_27827);
or U28242 (N_28242,N_27772,N_27552);
and U28243 (N_28243,N_27650,N_27997);
or U28244 (N_28244,N_27705,N_27560);
and U28245 (N_28245,N_27843,N_27926);
or U28246 (N_28246,N_27894,N_27886);
nand U28247 (N_28247,N_27613,N_27904);
or U28248 (N_28248,N_27684,N_27956);
and U28249 (N_28249,N_27645,N_27594);
and U28250 (N_28250,N_27893,N_27530);
and U28251 (N_28251,N_27784,N_27971);
nand U28252 (N_28252,N_27574,N_27933);
xnor U28253 (N_28253,N_27821,N_27750);
xnor U28254 (N_28254,N_27807,N_27921);
and U28255 (N_28255,N_27673,N_27586);
nor U28256 (N_28256,N_27945,N_27887);
or U28257 (N_28257,N_27816,N_27702);
nor U28258 (N_28258,N_27770,N_27910);
xnor U28259 (N_28259,N_27653,N_27548);
or U28260 (N_28260,N_27568,N_27910);
and U28261 (N_28261,N_27696,N_27565);
and U28262 (N_28262,N_27818,N_27704);
nand U28263 (N_28263,N_27995,N_27778);
and U28264 (N_28264,N_27513,N_27781);
xnor U28265 (N_28265,N_27854,N_27989);
nand U28266 (N_28266,N_27713,N_27855);
and U28267 (N_28267,N_27668,N_27743);
nand U28268 (N_28268,N_27632,N_27667);
nor U28269 (N_28269,N_27830,N_27771);
nor U28270 (N_28270,N_27584,N_27802);
nand U28271 (N_28271,N_27970,N_27702);
and U28272 (N_28272,N_27901,N_27849);
and U28273 (N_28273,N_27937,N_27635);
or U28274 (N_28274,N_27672,N_27651);
nor U28275 (N_28275,N_27676,N_27826);
nor U28276 (N_28276,N_27728,N_27889);
nand U28277 (N_28277,N_27716,N_27627);
or U28278 (N_28278,N_27602,N_27562);
xnor U28279 (N_28279,N_27916,N_27989);
nand U28280 (N_28280,N_27847,N_27894);
nand U28281 (N_28281,N_27897,N_27978);
xnor U28282 (N_28282,N_27545,N_27710);
or U28283 (N_28283,N_27831,N_27877);
or U28284 (N_28284,N_27717,N_27951);
nor U28285 (N_28285,N_27684,N_27537);
nor U28286 (N_28286,N_27835,N_27873);
or U28287 (N_28287,N_27880,N_27816);
nor U28288 (N_28288,N_27979,N_27944);
or U28289 (N_28289,N_27757,N_27768);
nor U28290 (N_28290,N_27729,N_27674);
and U28291 (N_28291,N_27924,N_27958);
and U28292 (N_28292,N_27536,N_27785);
nand U28293 (N_28293,N_27536,N_27553);
and U28294 (N_28294,N_27926,N_27811);
and U28295 (N_28295,N_27836,N_27542);
and U28296 (N_28296,N_27824,N_27662);
xor U28297 (N_28297,N_27865,N_27800);
and U28298 (N_28298,N_27945,N_27742);
nor U28299 (N_28299,N_27625,N_27730);
and U28300 (N_28300,N_27537,N_27859);
xnor U28301 (N_28301,N_27805,N_27838);
nor U28302 (N_28302,N_27516,N_27810);
nor U28303 (N_28303,N_27793,N_27779);
or U28304 (N_28304,N_27768,N_27761);
nor U28305 (N_28305,N_27952,N_27987);
or U28306 (N_28306,N_27687,N_27576);
or U28307 (N_28307,N_27952,N_27505);
xnor U28308 (N_28308,N_27945,N_27831);
nor U28309 (N_28309,N_27730,N_27886);
or U28310 (N_28310,N_27787,N_27732);
and U28311 (N_28311,N_27947,N_27998);
nand U28312 (N_28312,N_27648,N_27830);
nor U28313 (N_28313,N_27978,N_27890);
nand U28314 (N_28314,N_27912,N_27772);
nand U28315 (N_28315,N_27628,N_27916);
and U28316 (N_28316,N_27787,N_27554);
nor U28317 (N_28317,N_27962,N_27913);
xnor U28318 (N_28318,N_27649,N_27656);
or U28319 (N_28319,N_27773,N_27768);
or U28320 (N_28320,N_27500,N_27663);
nor U28321 (N_28321,N_27790,N_27811);
nor U28322 (N_28322,N_27817,N_27729);
xor U28323 (N_28323,N_27851,N_27721);
or U28324 (N_28324,N_27701,N_27768);
xor U28325 (N_28325,N_27891,N_27827);
nor U28326 (N_28326,N_27535,N_27861);
or U28327 (N_28327,N_27738,N_27691);
and U28328 (N_28328,N_27581,N_27935);
xor U28329 (N_28329,N_27866,N_27645);
nand U28330 (N_28330,N_27632,N_27841);
nand U28331 (N_28331,N_27905,N_27972);
xnor U28332 (N_28332,N_27964,N_27679);
nand U28333 (N_28333,N_27608,N_27739);
nor U28334 (N_28334,N_27747,N_27885);
or U28335 (N_28335,N_27676,N_27806);
nand U28336 (N_28336,N_27520,N_27969);
and U28337 (N_28337,N_27892,N_27960);
xnor U28338 (N_28338,N_27812,N_27794);
xnor U28339 (N_28339,N_27826,N_27685);
xnor U28340 (N_28340,N_27957,N_27645);
xnor U28341 (N_28341,N_27929,N_27547);
nor U28342 (N_28342,N_27775,N_27974);
nor U28343 (N_28343,N_27514,N_27658);
xor U28344 (N_28344,N_27682,N_27761);
and U28345 (N_28345,N_27864,N_27821);
or U28346 (N_28346,N_27566,N_27646);
nor U28347 (N_28347,N_27669,N_27894);
nand U28348 (N_28348,N_27889,N_27633);
and U28349 (N_28349,N_27830,N_27723);
nor U28350 (N_28350,N_27745,N_27633);
and U28351 (N_28351,N_27961,N_27533);
xor U28352 (N_28352,N_27743,N_27853);
nand U28353 (N_28353,N_27583,N_27981);
and U28354 (N_28354,N_27645,N_27551);
xor U28355 (N_28355,N_27920,N_27760);
nand U28356 (N_28356,N_27848,N_27643);
nor U28357 (N_28357,N_27600,N_27505);
and U28358 (N_28358,N_27728,N_27862);
xnor U28359 (N_28359,N_27788,N_27673);
nor U28360 (N_28360,N_27983,N_27518);
or U28361 (N_28361,N_27598,N_27974);
or U28362 (N_28362,N_27563,N_27704);
or U28363 (N_28363,N_27548,N_27979);
and U28364 (N_28364,N_27663,N_27862);
nand U28365 (N_28365,N_27698,N_27737);
or U28366 (N_28366,N_27942,N_27681);
xnor U28367 (N_28367,N_27883,N_27673);
and U28368 (N_28368,N_27833,N_27528);
and U28369 (N_28369,N_27915,N_27529);
and U28370 (N_28370,N_27645,N_27710);
xnor U28371 (N_28371,N_27761,N_27903);
or U28372 (N_28372,N_27543,N_27679);
and U28373 (N_28373,N_27898,N_27651);
or U28374 (N_28374,N_27883,N_27977);
or U28375 (N_28375,N_27525,N_27761);
and U28376 (N_28376,N_27956,N_27510);
nand U28377 (N_28377,N_27910,N_27890);
nor U28378 (N_28378,N_27810,N_27813);
xnor U28379 (N_28379,N_27820,N_27776);
nor U28380 (N_28380,N_27656,N_27757);
or U28381 (N_28381,N_27644,N_27769);
nand U28382 (N_28382,N_27674,N_27904);
nand U28383 (N_28383,N_27701,N_27593);
and U28384 (N_28384,N_27811,N_27798);
or U28385 (N_28385,N_27561,N_27814);
or U28386 (N_28386,N_27631,N_27827);
xnor U28387 (N_28387,N_27550,N_27980);
xor U28388 (N_28388,N_27551,N_27831);
nand U28389 (N_28389,N_27859,N_27923);
xnor U28390 (N_28390,N_27530,N_27527);
xnor U28391 (N_28391,N_27850,N_27874);
nor U28392 (N_28392,N_27928,N_27510);
and U28393 (N_28393,N_27977,N_27649);
xnor U28394 (N_28394,N_27599,N_27503);
and U28395 (N_28395,N_27614,N_27692);
xnor U28396 (N_28396,N_27943,N_27703);
xnor U28397 (N_28397,N_27584,N_27994);
nand U28398 (N_28398,N_27755,N_27795);
nor U28399 (N_28399,N_27885,N_27756);
nand U28400 (N_28400,N_27662,N_27806);
and U28401 (N_28401,N_27752,N_27847);
and U28402 (N_28402,N_27707,N_27841);
xnor U28403 (N_28403,N_27517,N_27579);
and U28404 (N_28404,N_27859,N_27762);
nand U28405 (N_28405,N_27835,N_27892);
and U28406 (N_28406,N_27678,N_27837);
nor U28407 (N_28407,N_27698,N_27515);
and U28408 (N_28408,N_27524,N_27735);
and U28409 (N_28409,N_27922,N_27904);
or U28410 (N_28410,N_27579,N_27950);
nand U28411 (N_28411,N_27522,N_27659);
nand U28412 (N_28412,N_27571,N_27545);
nor U28413 (N_28413,N_27859,N_27599);
or U28414 (N_28414,N_27932,N_27930);
or U28415 (N_28415,N_27689,N_27531);
or U28416 (N_28416,N_27895,N_27584);
or U28417 (N_28417,N_27582,N_27937);
nand U28418 (N_28418,N_27707,N_27758);
xnor U28419 (N_28419,N_27781,N_27562);
nand U28420 (N_28420,N_27768,N_27749);
nand U28421 (N_28421,N_27653,N_27771);
or U28422 (N_28422,N_27774,N_27620);
and U28423 (N_28423,N_27702,N_27728);
nor U28424 (N_28424,N_27712,N_27756);
xnor U28425 (N_28425,N_27724,N_27633);
xnor U28426 (N_28426,N_27980,N_27897);
nor U28427 (N_28427,N_27893,N_27532);
and U28428 (N_28428,N_27828,N_27571);
nand U28429 (N_28429,N_27820,N_27679);
nor U28430 (N_28430,N_27650,N_27965);
xor U28431 (N_28431,N_27753,N_27851);
xor U28432 (N_28432,N_27769,N_27613);
xor U28433 (N_28433,N_27771,N_27701);
and U28434 (N_28434,N_27995,N_27865);
and U28435 (N_28435,N_27579,N_27768);
nand U28436 (N_28436,N_27691,N_27618);
and U28437 (N_28437,N_27834,N_27737);
and U28438 (N_28438,N_27789,N_27874);
and U28439 (N_28439,N_27803,N_27822);
nand U28440 (N_28440,N_27666,N_27962);
nor U28441 (N_28441,N_27736,N_27597);
nor U28442 (N_28442,N_27538,N_27870);
nand U28443 (N_28443,N_27763,N_27951);
nand U28444 (N_28444,N_27892,N_27734);
or U28445 (N_28445,N_27780,N_27731);
nor U28446 (N_28446,N_27621,N_27996);
and U28447 (N_28447,N_27616,N_27500);
nand U28448 (N_28448,N_27706,N_27844);
nand U28449 (N_28449,N_27727,N_27896);
nand U28450 (N_28450,N_27704,N_27554);
nor U28451 (N_28451,N_27704,N_27912);
xor U28452 (N_28452,N_27565,N_27910);
and U28453 (N_28453,N_27976,N_27786);
and U28454 (N_28454,N_27976,N_27587);
or U28455 (N_28455,N_27725,N_27801);
nand U28456 (N_28456,N_27812,N_27769);
nand U28457 (N_28457,N_27978,N_27585);
xor U28458 (N_28458,N_27739,N_27782);
or U28459 (N_28459,N_27642,N_27925);
nor U28460 (N_28460,N_27995,N_27968);
and U28461 (N_28461,N_27896,N_27904);
and U28462 (N_28462,N_27612,N_27555);
nand U28463 (N_28463,N_27740,N_27985);
nor U28464 (N_28464,N_27834,N_27782);
or U28465 (N_28465,N_27681,N_27691);
or U28466 (N_28466,N_27751,N_27982);
xnor U28467 (N_28467,N_27939,N_27873);
nand U28468 (N_28468,N_27580,N_27722);
nand U28469 (N_28469,N_27724,N_27735);
and U28470 (N_28470,N_27684,N_27620);
and U28471 (N_28471,N_27868,N_27791);
and U28472 (N_28472,N_27973,N_27813);
nor U28473 (N_28473,N_27849,N_27517);
nand U28474 (N_28474,N_27749,N_27696);
and U28475 (N_28475,N_27967,N_27942);
xor U28476 (N_28476,N_27802,N_27710);
nor U28477 (N_28477,N_27713,N_27837);
nor U28478 (N_28478,N_27945,N_27606);
xnor U28479 (N_28479,N_27929,N_27781);
nor U28480 (N_28480,N_27996,N_27500);
nand U28481 (N_28481,N_27863,N_27947);
and U28482 (N_28482,N_27999,N_27887);
and U28483 (N_28483,N_27885,N_27804);
or U28484 (N_28484,N_27647,N_27619);
xnor U28485 (N_28485,N_27971,N_27601);
or U28486 (N_28486,N_27826,N_27700);
nor U28487 (N_28487,N_27995,N_27503);
and U28488 (N_28488,N_27604,N_27697);
and U28489 (N_28489,N_27922,N_27688);
and U28490 (N_28490,N_27776,N_27535);
nor U28491 (N_28491,N_27765,N_27529);
and U28492 (N_28492,N_27509,N_27596);
xnor U28493 (N_28493,N_27996,N_27727);
nand U28494 (N_28494,N_27626,N_27552);
or U28495 (N_28495,N_27923,N_27715);
and U28496 (N_28496,N_27721,N_27665);
and U28497 (N_28497,N_27714,N_27744);
nand U28498 (N_28498,N_27960,N_27752);
and U28499 (N_28499,N_27777,N_27757);
xor U28500 (N_28500,N_28183,N_28210);
or U28501 (N_28501,N_28296,N_28464);
nor U28502 (N_28502,N_28345,N_28188);
xnor U28503 (N_28503,N_28440,N_28385);
nand U28504 (N_28504,N_28224,N_28186);
or U28505 (N_28505,N_28301,N_28145);
nor U28506 (N_28506,N_28014,N_28216);
nand U28507 (N_28507,N_28257,N_28326);
nand U28508 (N_28508,N_28007,N_28297);
nand U28509 (N_28509,N_28212,N_28499);
nand U28510 (N_28510,N_28276,N_28380);
or U28511 (N_28511,N_28189,N_28341);
nor U28512 (N_28512,N_28452,N_28338);
and U28513 (N_28513,N_28286,N_28194);
or U28514 (N_28514,N_28050,N_28364);
xor U28515 (N_28515,N_28316,N_28308);
nand U28516 (N_28516,N_28492,N_28233);
xnor U28517 (N_28517,N_28202,N_28156);
xnor U28518 (N_28518,N_28336,N_28391);
or U28519 (N_28519,N_28366,N_28182);
xnor U28520 (N_28520,N_28038,N_28491);
nor U28521 (N_28521,N_28018,N_28070);
and U28522 (N_28522,N_28221,N_28496);
nor U28523 (N_28523,N_28283,N_28135);
or U28524 (N_28524,N_28414,N_28150);
and U28525 (N_28525,N_28196,N_28284);
nor U28526 (N_28526,N_28035,N_28352);
or U28527 (N_28527,N_28081,N_28350);
and U28528 (N_28528,N_28054,N_28359);
nor U28529 (N_28529,N_28244,N_28343);
nor U28530 (N_28530,N_28164,N_28402);
and U28531 (N_28531,N_28108,N_28449);
nand U28532 (N_28532,N_28096,N_28044);
nand U28533 (N_28533,N_28084,N_28234);
nor U28534 (N_28534,N_28229,N_28117);
nand U28535 (N_28535,N_28079,N_28238);
nand U28536 (N_28536,N_28262,N_28255);
nand U28537 (N_28537,N_28066,N_28430);
and U28538 (N_28538,N_28217,N_28242);
xnor U28539 (N_28539,N_28024,N_28268);
nor U28540 (N_28540,N_28421,N_28002);
nand U28541 (N_28541,N_28494,N_28140);
or U28542 (N_28542,N_28057,N_28322);
xor U28543 (N_28543,N_28372,N_28171);
xnor U28544 (N_28544,N_28314,N_28407);
xor U28545 (N_28545,N_28434,N_28395);
or U28546 (N_28546,N_28468,N_28132);
and U28547 (N_28547,N_28142,N_28363);
and U28548 (N_28548,N_28305,N_28176);
and U28549 (N_28549,N_28017,N_28278);
xor U28550 (N_28550,N_28065,N_28049);
or U28551 (N_28551,N_28497,N_28046);
nor U28552 (N_28552,N_28149,N_28329);
or U28553 (N_28553,N_28428,N_28272);
or U28554 (N_28554,N_28040,N_28162);
xnor U28555 (N_28555,N_28377,N_28028);
nor U28556 (N_28556,N_28113,N_28174);
or U28557 (N_28557,N_28173,N_28201);
nor U28558 (N_28558,N_28073,N_28495);
xnor U28559 (N_28559,N_28409,N_28119);
nand U28560 (N_28560,N_28000,N_28125);
and U28561 (N_28561,N_28444,N_28203);
nand U28562 (N_28562,N_28193,N_28138);
or U28563 (N_28563,N_28413,N_28399);
nor U28564 (N_28564,N_28292,N_28127);
or U28565 (N_28565,N_28454,N_28223);
nor U28566 (N_28566,N_28141,N_28478);
nor U28567 (N_28567,N_28462,N_28102);
nor U28568 (N_28568,N_28170,N_28417);
or U28569 (N_28569,N_28342,N_28036);
xnor U28570 (N_28570,N_28195,N_28172);
nor U28571 (N_28571,N_28410,N_28348);
xor U28572 (N_28572,N_28277,N_28091);
nand U28573 (N_28573,N_28376,N_28146);
or U28574 (N_28574,N_28327,N_28041);
and U28575 (N_28575,N_28072,N_28431);
xor U28576 (N_28576,N_28163,N_28154);
and U28577 (N_28577,N_28360,N_28116);
nand U28578 (N_28578,N_28412,N_28351);
and U28579 (N_28579,N_28005,N_28300);
xnor U28580 (N_28580,N_28472,N_28441);
xor U28581 (N_28581,N_28482,N_28228);
xor U28582 (N_28582,N_28453,N_28393);
nor U28583 (N_28583,N_28064,N_28103);
nand U28584 (N_28584,N_28047,N_28282);
or U28585 (N_28585,N_28367,N_28248);
and U28586 (N_28586,N_28307,N_28168);
xor U28587 (N_28587,N_28205,N_28115);
and U28588 (N_28588,N_28129,N_28226);
xor U28589 (N_28589,N_28382,N_28012);
nand U28590 (N_28590,N_28298,N_28089);
and U28591 (N_28591,N_28134,N_28006);
and U28592 (N_28592,N_28427,N_28490);
or U28593 (N_28593,N_28076,N_28158);
xor U28594 (N_28594,N_28467,N_28152);
xor U28595 (N_28595,N_28355,N_28093);
nor U28596 (N_28596,N_28092,N_28261);
or U28597 (N_28597,N_28153,N_28107);
xor U28598 (N_28598,N_28267,N_28473);
or U28599 (N_28599,N_28251,N_28375);
or U28600 (N_28600,N_28269,N_28347);
xnor U28601 (N_28601,N_28397,N_28181);
nand U28602 (N_28602,N_28151,N_28404);
nor U28603 (N_28603,N_28423,N_28015);
xor U28604 (N_28604,N_28445,N_28361);
nor U28605 (N_28605,N_28324,N_28220);
or U28606 (N_28606,N_28253,N_28239);
and U28607 (N_28607,N_28470,N_28287);
nor U28608 (N_28608,N_28204,N_28457);
xnor U28609 (N_28609,N_28439,N_28143);
and U28610 (N_28610,N_28240,N_28087);
nand U28611 (N_28611,N_28334,N_28225);
xnor U28612 (N_28612,N_28099,N_28333);
xnor U28613 (N_28613,N_28003,N_28312);
nand U28614 (N_28614,N_28398,N_28048);
and U28615 (N_28615,N_28001,N_28022);
xor U28616 (N_28616,N_28386,N_28206);
and U28617 (N_28617,N_28455,N_28450);
nor U28618 (N_28618,N_28023,N_28053);
nor U28619 (N_28619,N_28458,N_28249);
or U28620 (N_28620,N_28388,N_28461);
nand U28621 (N_28621,N_28344,N_28227);
nor U28622 (N_28622,N_28291,N_28285);
and U28623 (N_28623,N_28281,N_28365);
or U28624 (N_28624,N_28483,N_28237);
and U28625 (N_28625,N_28088,N_28418);
and U28626 (N_28626,N_28354,N_28241);
or U28627 (N_28627,N_28466,N_28020);
and U28628 (N_28628,N_28067,N_28130);
and U28629 (N_28629,N_28406,N_28459);
nand U28630 (N_28630,N_28485,N_28318);
nor U28631 (N_28631,N_28469,N_28369);
and U28632 (N_28632,N_28396,N_28325);
or U28633 (N_28633,N_28498,N_28136);
and U28634 (N_28634,N_28021,N_28447);
and U28635 (N_28635,N_28471,N_28144);
nand U28636 (N_28636,N_28110,N_28254);
xor U28637 (N_28637,N_28013,N_28159);
and U28638 (N_28638,N_28480,N_28484);
or U28639 (N_28639,N_28207,N_28069);
xor U28640 (N_28640,N_28438,N_28009);
nand U28641 (N_28641,N_28190,N_28463);
nor U28642 (N_28642,N_28311,N_28169);
and U28643 (N_28643,N_28199,N_28200);
and U28644 (N_28644,N_28362,N_28394);
nor U28645 (N_28645,N_28105,N_28120);
nor U28646 (N_28646,N_28346,N_28258);
and U28647 (N_28647,N_28303,N_28451);
nand U28648 (N_28648,N_28299,N_28051);
nor U28649 (N_28649,N_28401,N_28353);
nor U28650 (N_28650,N_28264,N_28403);
xor U28651 (N_28651,N_28294,N_28033);
or U28652 (N_28652,N_28062,N_28486);
nor U28653 (N_28653,N_28232,N_28045);
nand U28654 (N_28654,N_28415,N_28160);
xor U28655 (N_28655,N_28074,N_28263);
xor U28656 (N_28656,N_28019,N_28106);
xor U28657 (N_28657,N_28139,N_28068);
xnor U28658 (N_28658,N_28295,N_28208);
nor U28659 (N_28659,N_28456,N_28101);
xnor U28660 (N_28660,N_28289,N_28097);
nor U28661 (N_28661,N_28493,N_28071);
xnor U28662 (N_28662,N_28392,N_28211);
and U28663 (N_28663,N_28331,N_28443);
or U28664 (N_28664,N_28155,N_28167);
and U28665 (N_28665,N_28250,N_28357);
nor U28666 (N_28666,N_28420,N_28077);
nor U28667 (N_28667,N_28187,N_28271);
xnor U28668 (N_28668,N_28236,N_28477);
nand U28669 (N_28669,N_28063,N_28209);
or U28670 (N_28670,N_28037,N_28039);
or U28671 (N_28671,N_28309,N_28320);
nor U28672 (N_28672,N_28059,N_28266);
and U28673 (N_28673,N_28137,N_28061);
nand U28674 (N_28674,N_28315,N_28387);
nand U28675 (N_28675,N_28374,N_28436);
xor U28676 (N_28676,N_28060,N_28270);
xnor U28677 (N_28677,N_28222,N_28008);
nand U28678 (N_28678,N_28476,N_28411);
xnor U28679 (N_28679,N_28288,N_28198);
or U28680 (N_28680,N_28133,N_28029);
nand U28681 (N_28681,N_28128,N_28104);
nand U28682 (N_28682,N_28381,N_28384);
nand U28683 (N_28683,N_28191,N_28100);
xor U28684 (N_28684,N_28058,N_28321);
or U28685 (N_28685,N_28379,N_28306);
nor U28686 (N_28686,N_28340,N_28405);
nor U28687 (N_28687,N_28313,N_28373);
or U28688 (N_28688,N_28435,N_28165);
or U28689 (N_28689,N_28370,N_28052);
and U28690 (N_28690,N_28056,N_28214);
or U28691 (N_28691,N_28332,N_28112);
xor U28692 (N_28692,N_28042,N_28004);
xnor U28693 (N_28693,N_28330,N_28437);
nand U28694 (N_28694,N_28323,N_28184);
or U28695 (N_28695,N_28218,N_28358);
nand U28696 (N_28696,N_28319,N_28368);
xnor U28697 (N_28697,N_28126,N_28460);
and U28698 (N_28698,N_28157,N_28031);
or U28699 (N_28699,N_28465,N_28197);
and U28700 (N_28700,N_28030,N_28481);
and U28701 (N_28701,N_28147,N_28349);
and U28702 (N_28702,N_28082,N_28078);
nor U28703 (N_28703,N_28419,N_28025);
and U28704 (N_28704,N_28090,N_28247);
and U28705 (N_28705,N_28335,N_28043);
or U28706 (N_28706,N_28246,N_28274);
nand U28707 (N_28707,N_28474,N_28339);
xnor U28708 (N_28708,N_28487,N_28055);
xor U28709 (N_28709,N_28083,N_28273);
nor U28710 (N_28710,N_28433,N_28293);
and U28711 (N_28711,N_28175,N_28026);
xnor U28712 (N_28712,N_28098,N_28429);
and U28713 (N_28713,N_28383,N_28243);
or U28714 (N_28714,N_28400,N_28075);
xor U28715 (N_28715,N_28011,N_28489);
nand U28716 (N_28716,N_28034,N_28279);
nor U28717 (N_28717,N_28275,N_28448);
nor U28718 (N_28718,N_28118,N_28389);
nand U28719 (N_28719,N_28179,N_28177);
xnor U28720 (N_28720,N_28425,N_28085);
xnor U28721 (N_28721,N_28131,N_28416);
nand U28722 (N_28722,N_28192,N_28231);
xor U28723 (N_28723,N_28280,N_28094);
nor U28724 (N_28724,N_28027,N_28185);
nor U28725 (N_28725,N_28032,N_28252);
xnor U28726 (N_28726,N_28260,N_28290);
nand U28727 (N_28727,N_28446,N_28180);
or U28728 (N_28728,N_28219,N_28086);
nand U28729 (N_28729,N_28356,N_28442);
or U28730 (N_28730,N_28337,N_28328);
xnor U28731 (N_28731,N_28488,N_28095);
and U28732 (N_28732,N_28310,N_28121);
and U28733 (N_28733,N_28124,N_28213);
and U28734 (N_28734,N_28148,N_28426);
xnor U28735 (N_28735,N_28245,N_28215);
xnor U28736 (N_28736,N_28230,N_28123);
nand U28737 (N_28737,N_28371,N_28408);
and U28738 (N_28738,N_28111,N_28161);
xor U28739 (N_28739,N_28479,N_28390);
xor U28740 (N_28740,N_28016,N_28304);
nand U28741 (N_28741,N_28259,N_28109);
xnor U28742 (N_28742,N_28432,N_28122);
nor U28743 (N_28743,N_28302,N_28378);
xor U28744 (N_28744,N_28422,N_28317);
and U28745 (N_28745,N_28080,N_28010);
nor U28746 (N_28746,N_28114,N_28235);
nand U28747 (N_28747,N_28424,N_28256);
nor U28748 (N_28748,N_28475,N_28265);
nand U28749 (N_28749,N_28166,N_28178);
and U28750 (N_28750,N_28373,N_28009);
or U28751 (N_28751,N_28004,N_28444);
nand U28752 (N_28752,N_28478,N_28246);
or U28753 (N_28753,N_28033,N_28348);
nor U28754 (N_28754,N_28208,N_28364);
nand U28755 (N_28755,N_28453,N_28016);
nand U28756 (N_28756,N_28337,N_28090);
nor U28757 (N_28757,N_28166,N_28389);
nand U28758 (N_28758,N_28478,N_28064);
xnor U28759 (N_28759,N_28376,N_28057);
nor U28760 (N_28760,N_28465,N_28030);
xor U28761 (N_28761,N_28252,N_28143);
or U28762 (N_28762,N_28165,N_28077);
xnor U28763 (N_28763,N_28266,N_28413);
xor U28764 (N_28764,N_28138,N_28162);
xor U28765 (N_28765,N_28139,N_28069);
nand U28766 (N_28766,N_28488,N_28055);
or U28767 (N_28767,N_28356,N_28270);
and U28768 (N_28768,N_28035,N_28055);
nand U28769 (N_28769,N_28154,N_28465);
xnor U28770 (N_28770,N_28022,N_28330);
nor U28771 (N_28771,N_28013,N_28328);
nand U28772 (N_28772,N_28286,N_28349);
xnor U28773 (N_28773,N_28311,N_28003);
or U28774 (N_28774,N_28244,N_28470);
xnor U28775 (N_28775,N_28229,N_28373);
or U28776 (N_28776,N_28020,N_28284);
nand U28777 (N_28777,N_28283,N_28390);
nor U28778 (N_28778,N_28438,N_28288);
nor U28779 (N_28779,N_28037,N_28256);
xor U28780 (N_28780,N_28224,N_28256);
nor U28781 (N_28781,N_28070,N_28481);
xnor U28782 (N_28782,N_28033,N_28323);
nand U28783 (N_28783,N_28415,N_28261);
nor U28784 (N_28784,N_28157,N_28449);
and U28785 (N_28785,N_28043,N_28435);
xor U28786 (N_28786,N_28290,N_28114);
xor U28787 (N_28787,N_28438,N_28094);
nor U28788 (N_28788,N_28040,N_28331);
and U28789 (N_28789,N_28388,N_28268);
xor U28790 (N_28790,N_28484,N_28363);
or U28791 (N_28791,N_28087,N_28456);
nand U28792 (N_28792,N_28355,N_28216);
and U28793 (N_28793,N_28124,N_28069);
nor U28794 (N_28794,N_28303,N_28264);
nor U28795 (N_28795,N_28115,N_28297);
xnor U28796 (N_28796,N_28141,N_28325);
and U28797 (N_28797,N_28164,N_28068);
nand U28798 (N_28798,N_28050,N_28104);
or U28799 (N_28799,N_28351,N_28490);
or U28800 (N_28800,N_28068,N_28315);
or U28801 (N_28801,N_28396,N_28286);
or U28802 (N_28802,N_28491,N_28452);
nand U28803 (N_28803,N_28431,N_28135);
nand U28804 (N_28804,N_28298,N_28286);
xnor U28805 (N_28805,N_28090,N_28172);
nor U28806 (N_28806,N_28120,N_28371);
xnor U28807 (N_28807,N_28181,N_28354);
nand U28808 (N_28808,N_28187,N_28407);
nand U28809 (N_28809,N_28055,N_28454);
and U28810 (N_28810,N_28482,N_28045);
and U28811 (N_28811,N_28153,N_28328);
nand U28812 (N_28812,N_28096,N_28032);
and U28813 (N_28813,N_28364,N_28163);
nor U28814 (N_28814,N_28391,N_28289);
xor U28815 (N_28815,N_28277,N_28292);
and U28816 (N_28816,N_28433,N_28439);
nand U28817 (N_28817,N_28351,N_28372);
nor U28818 (N_28818,N_28185,N_28046);
xor U28819 (N_28819,N_28466,N_28416);
or U28820 (N_28820,N_28207,N_28429);
xor U28821 (N_28821,N_28389,N_28427);
xnor U28822 (N_28822,N_28388,N_28170);
nand U28823 (N_28823,N_28038,N_28228);
and U28824 (N_28824,N_28389,N_28200);
nand U28825 (N_28825,N_28480,N_28250);
nor U28826 (N_28826,N_28084,N_28118);
nor U28827 (N_28827,N_28293,N_28146);
xnor U28828 (N_28828,N_28258,N_28073);
nor U28829 (N_28829,N_28254,N_28377);
or U28830 (N_28830,N_28469,N_28312);
nor U28831 (N_28831,N_28355,N_28343);
nor U28832 (N_28832,N_28388,N_28113);
and U28833 (N_28833,N_28233,N_28141);
or U28834 (N_28834,N_28212,N_28289);
nand U28835 (N_28835,N_28455,N_28494);
nor U28836 (N_28836,N_28141,N_28032);
nor U28837 (N_28837,N_28415,N_28200);
xor U28838 (N_28838,N_28394,N_28299);
nand U28839 (N_28839,N_28332,N_28196);
and U28840 (N_28840,N_28034,N_28365);
nand U28841 (N_28841,N_28278,N_28153);
and U28842 (N_28842,N_28487,N_28213);
nand U28843 (N_28843,N_28035,N_28373);
nor U28844 (N_28844,N_28167,N_28083);
nor U28845 (N_28845,N_28269,N_28105);
and U28846 (N_28846,N_28071,N_28436);
nor U28847 (N_28847,N_28470,N_28418);
or U28848 (N_28848,N_28233,N_28290);
nor U28849 (N_28849,N_28040,N_28489);
xor U28850 (N_28850,N_28128,N_28246);
nor U28851 (N_28851,N_28484,N_28211);
nor U28852 (N_28852,N_28056,N_28179);
nand U28853 (N_28853,N_28279,N_28291);
and U28854 (N_28854,N_28007,N_28424);
xor U28855 (N_28855,N_28472,N_28156);
xor U28856 (N_28856,N_28166,N_28068);
or U28857 (N_28857,N_28044,N_28015);
xnor U28858 (N_28858,N_28266,N_28112);
and U28859 (N_28859,N_28362,N_28349);
nor U28860 (N_28860,N_28364,N_28009);
nand U28861 (N_28861,N_28108,N_28494);
nor U28862 (N_28862,N_28187,N_28362);
nor U28863 (N_28863,N_28472,N_28019);
and U28864 (N_28864,N_28081,N_28287);
and U28865 (N_28865,N_28154,N_28051);
and U28866 (N_28866,N_28030,N_28427);
xor U28867 (N_28867,N_28440,N_28007);
or U28868 (N_28868,N_28232,N_28252);
xor U28869 (N_28869,N_28237,N_28291);
or U28870 (N_28870,N_28187,N_28019);
nor U28871 (N_28871,N_28469,N_28004);
or U28872 (N_28872,N_28218,N_28348);
and U28873 (N_28873,N_28300,N_28344);
xnor U28874 (N_28874,N_28184,N_28338);
or U28875 (N_28875,N_28329,N_28230);
xor U28876 (N_28876,N_28355,N_28248);
or U28877 (N_28877,N_28129,N_28062);
or U28878 (N_28878,N_28066,N_28456);
xor U28879 (N_28879,N_28330,N_28372);
xnor U28880 (N_28880,N_28122,N_28130);
and U28881 (N_28881,N_28117,N_28373);
or U28882 (N_28882,N_28220,N_28185);
and U28883 (N_28883,N_28230,N_28270);
nor U28884 (N_28884,N_28467,N_28130);
nand U28885 (N_28885,N_28196,N_28353);
nor U28886 (N_28886,N_28403,N_28297);
nor U28887 (N_28887,N_28445,N_28442);
xnor U28888 (N_28888,N_28281,N_28435);
xnor U28889 (N_28889,N_28011,N_28098);
or U28890 (N_28890,N_28094,N_28257);
or U28891 (N_28891,N_28077,N_28324);
and U28892 (N_28892,N_28469,N_28097);
xor U28893 (N_28893,N_28094,N_28090);
nor U28894 (N_28894,N_28458,N_28325);
nand U28895 (N_28895,N_28048,N_28365);
xnor U28896 (N_28896,N_28415,N_28074);
and U28897 (N_28897,N_28455,N_28354);
and U28898 (N_28898,N_28332,N_28026);
or U28899 (N_28899,N_28358,N_28243);
nor U28900 (N_28900,N_28376,N_28270);
nor U28901 (N_28901,N_28320,N_28242);
nor U28902 (N_28902,N_28388,N_28265);
nor U28903 (N_28903,N_28176,N_28105);
and U28904 (N_28904,N_28211,N_28483);
xor U28905 (N_28905,N_28405,N_28062);
and U28906 (N_28906,N_28106,N_28288);
nor U28907 (N_28907,N_28010,N_28049);
and U28908 (N_28908,N_28288,N_28234);
or U28909 (N_28909,N_28351,N_28093);
and U28910 (N_28910,N_28203,N_28248);
xor U28911 (N_28911,N_28287,N_28023);
and U28912 (N_28912,N_28040,N_28175);
nor U28913 (N_28913,N_28285,N_28222);
xor U28914 (N_28914,N_28442,N_28009);
nor U28915 (N_28915,N_28003,N_28036);
or U28916 (N_28916,N_28491,N_28460);
nand U28917 (N_28917,N_28284,N_28390);
or U28918 (N_28918,N_28199,N_28394);
xor U28919 (N_28919,N_28435,N_28188);
or U28920 (N_28920,N_28044,N_28118);
or U28921 (N_28921,N_28185,N_28349);
nand U28922 (N_28922,N_28490,N_28474);
nand U28923 (N_28923,N_28072,N_28101);
nand U28924 (N_28924,N_28047,N_28186);
and U28925 (N_28925,N_28028,N_28429);
and U28926 (N_28926,N_28420,N_28428);
and U28927 (N_28927,N_28384,N_28001);
and U28928 (N_28928,N_28104,N_28066);
or U28929 (N_28929,N_28486,N_28481);
nor U28930 (N_28930,N_28372,N_28326);
and U28931 (N_28931,N_28032,N_28178);
nor U28932 (N_28932,N_28198,N_28458);
and U28933 (N_28933,N_28139,N_28315);
or U28934 (N_28934,N_28127,N_28198);
nand U28935 (N_28935,N_28496,N_28432);
nand U28936 (N_28936,N_28148,N_28408);
xnor U28937 (N_28937,N_28106,N_28370);
and U28938 (N_28938,N_28488,N_28271);
nand U28939 (N_28939,N_28221,N_28289);
nand U28940 (N_28940,N_28414,N_28374);
or U28941 (N_28941,N_28029,N_28447);
xnor U28942 (N_28942,N_28113,N_28427);
or U28943 (N_28943,N_28495,N_28026);
or U28944 (N_28944,N_28220,N_28482);
xnor U28945 (N_28945,N_28218,N_28314);
or U28946 (N_28946,N_28116,N_28417);
nor U28947 (N_28947,N_28173,N_28224);
nor U28948 (N_28948,N_28124,N_28374);
nor U28949 (N_28949,N_28150,N_28368);
xor U28950 (N_28950,N_28271,N_28176);
and U28951 (N_28951,N_28414,N_28070);
and U28952 (N_28952,N_28266,N_28348);
nand U28953 (N_28953,N_28237,N_28019);
xnor U28954 (N_28954,N_28249,N_28086);
xnor U28955 (N_28955,N_28327,N_28260);
xor U28956 (N_28956,N_28393,N_28058);
nor U28957 (N_28957,N_28050,N_28149);
nor U28958 (N_28958,N_28412,N_28373);
or U28959 (N_28959,N_28234,N_28463);
xnor U28960 (N_28960,N_28044,N_28363);
and U28961 (N_28961,N_28226,N_28090);
and U28962 (N_28962,N_28196,N_28248);
and U28963 (N_28963,N_28350,N_28296);
xnor U28964 (N_28964,N_28307,N_28157);
or U28965 (N_28965,N_28107,N_28345);
nand U28966 (N_28966,N_28378,N_28390);
nor U28967 (N_28967,N_28328,N_28449);
xnor U28968 (N_28968,N_28077,N_28102);
nor U28969 (N_28969,N_28324,N_28391);
nand U28970 (N_28970,N_28148,N_28498);
or U28971 (N_28971,N_28031,N_28210);
nand U28972 (N_28972,N_28026,N_28424);
nand U28973 (N_28973,N_28110,N_28434);
and U28974 (N_28974,N_28398,N_28373);
nand U28975 (N_28975,N_28223,N_28192);
or U28976 (N_28976,N_28298,N_28359);
or U28977 (N_28977,N_28490,N_28060);
or U28978 (N_28978,N_28149,N_28117);
nor U28979 (N_28979,N_28196,N_28445);
and U28980 (N_28980,N_28280,N_28076);
or U28981 (N_28981,N_28097,N_28201);
or U28982 (N_28982,N_28020,N_28109);
nor U28983 (N_28983,N_28386,N_28407);
nand U28984 (N_28984,N_28212,N_28016);
and U28985 (N_28985,N_28068,N_28423);
and U28986 (N_28986,N_28497,N_28187);
nor U28987 (N_28987,N_28308,N_28459);
or U28988 (N_28988,N_28361,N_28421);
or U28989 (N_28989,N_28028,N_28375);
xnor U28990 (N_28990,N_28219,N_28194);
nor U28991 (N_28991,N_28023,N_28251);
nor U28992 (N_28992,N_28438,N_28103);
or U28993 (N_28993,N_28319,N_28493);
xnor U28994 (N_28994,N_28380,N_28146);
xnor U28995 (N_28995,N_28239,N_28160);
or U28996 (N_28996,N_28106,N_28462);
nor U28997 (N_28997,N_28482,N_28195);
nand U28998 (N_28998,N_28156,N_28358);
nand U28999 (N_28999,N_28254,N_28326);
and U29000 (N_29000,N_28557,N_28598);
nor U29001 (N_29001,N_28657,N_28514);
nand U29002 (N_29002,N_28510,N_28946);
nor U29003 (N_29003,N_28783,N_28823);
nand U29004 (N_29004,N_28794,N_28778);
xor U29005 (N_29005,N_28679,N_28831);
or U29006 (N_29006,N_28918,N_28885);
xnor U29007 (N_29007,N_28872,N_28743);
nor U29008 (N_29008,N_28636,N_28525);
nand U29009 (N_29009,N_28972,N_28907);
and U29010 (N_29010,N_28930,N_28655);
nand U29011 (N_29011,N_28995,N_28681);
nor U29012 (N_29012,N_28543,N_28713);
or U29013 (N_29013,N_28888,N_28711);
and U29014 (N_29014,N_28825,N_28998);
nand U29015 (N_29015,N_28773,N_28982);
nand U29016 (N_29016,N_28996,N_28620);
nand U29017 (N_29017,N_28715,N_28921);
nor U29018 (N_29018,N_28537,N_28853);
xnor U29019 (N_29019,N_28666,N_28746);
and U29020 (N_29020,N_28606,N_28754);
nand U29021 (N_29021,N_28965,N_28989);
nand U29022 (N_29022,N_28803,N_28765);
xnor U29023 (N_29023,N_28928,N_28667);
or U29024 (N_29024,N_28532,N_28534);
nand U29025 (N_29025,N_28821,N_28665);
xor U29026 (N_29026,N_28818,N_28864);
or U29027 (N_29027,N_28599,N_28707);
or U29028 (N_29028,N_28889,N_28772);
or U29029 (N_29029,N_28755,N_28670);
and U29030 (N_29030,N_28978,N_28986);
xnor U29031 (N_29031,N_28857,N_28571);
nand U29032 (N_29032,N_28844,N_28637);
nor U29033 (N_29033,N_28917,N_28662);
xor U29034 (N_29034,N_28682,N_28518);
or U29035 (N_29035,N_28870,N_28920);
or U29036 (N_29036,N_28816,N_28767);
nor U29037 (N_29037,N_28668,N_28869);
nor U29038 (N_29038,N_28898,N_28852);
nor U29039 (N_29039,N_28621,N_28674);
nand U29040 (N_29040,N_28550,N_28649);
and U29041 (N_29041,N_28939,N_28517);
or U29042 (N_29042,N_28584,N_28660);
and U29043 (N_29043,N_28762,N_28953);
and U29044 (N_29044,N_28776,N_28908);
xnor U29045 (N_29045,N_28728,N_28923);
nor U29046 (N_29046,N_28785,N_28507);
or U29047 (N_29047,N_28614,N_28568);
nand U29048 (N_29048,N_28651,N_28752);
and U29049 (N_29049,N_28603,N_28867);
xnor U29050 (N_29050,N_28904,N_28952);
or U29051 (N_29051,N_28847,N_28905);
and U29052 (N_29052,N_28860,N_28969);
xor U29053 (N_29053,N_28763,N_28868);
xor U29054 (N_29054,N_28798,N_28533);
xor U29055 (N_29055,N_28902,N_28795);
nor U29056 (N_29056,N_28569,N_28766);
xnor U29057 (N_29057,N_28784,N_28997);
and U29058 (N_29058,N_28677,N_28935);
and U29059 (N_29059,N_28782,N_28994);
nand U29060 (N_29060,N_28663,N_28516);
and U29061 (N_29061,N_28744,N_28940);
nand U29062 (N_29062,N_28694,N_28845);
xnor U29063 (N_29063,N_28900,N_28971);
nor U29064 (N_29064,N_28504,N_28683);
or U29065 (N_29065,N_28894,N_28709);
and U29066 (N_29066,N_28886,N_28600);
nand U29067 (N_29067,N_28704,N_28642);
xnor U29068 (N_29068,N_28501,N_28944);
and U29069 (N_29069,N_28559,N_28535);
and U29070 (N_29070,N_28645,N_28572);
nor U29071 (N_29071,N_28881,N_28549);
nand U29072 (N_29072,N_28725,N_28560);
xnor U29073 (N_29073,N_28701,N_28976);
and U29074 (N_29074,N_28901,N_28801);
nand U29075 (N_29075,N_28546,N_28689);
and U29076 (N_29076,N_28984,N_28903);
or U29077 (N_29077,N_28839,N_28574);
xor U29078 (N_29078,N_28884,N_28714);
xor U29079 (N_29079,N_28576,N_28523);
or U29080 (N_29080,N_28695,N_28836);
nor U29081 (N_29081,N_28826,N_28723);
nor U29082 (N_29082,N_28720,N_28628);
nand U29083 (N_29083,N_28545,N_28608);
or U29084 (N_29084,N_28999,N_28760);
nor U29085 (N_29085,N_28640,N_28583);
or U29086 (N_29086,N_28915,N_28506);
or U29087 (N_29087,N_28873,N_28697);
nand U29088 (N_29088,N_28502,N_28876);
nor U29089 (N_29089,N_28749,N_28722);
nor U29090 (N_29090,N_28968,N_28779);
nand U29091 (N_29091,N_28856,N_28592);
nor U29092 (N_29092,N_28974,N_28615);
xnor U29093 (N_29093,N_28815,N_28698);
nor U29094 (N_29094,N_28896,N_28964);
nor U29095 (N_29095,N_28623,N_28893);
nand U29096 (N_29096,N_28676,N_28751);
xnor U29097 (N_29097,N_28808,N_28846);
xor U29098 (N_29098,N_28612,N_28954);
nand U29099 (N_29099,N_28786,N_28519);
nand U29100 (N_29100,N_28792,N_28675);
or U29101 (N_29101,N_28759,N_28602);
and U29102 (N_29102,N_28883,N_28947);
nor U29103 (N_29103,N_28661,N_28540);
nand U29104 (N_29104,N_28813,N_28764);
or U29105 (N_29105,N_28820,N_28756);
or U29106 (N_29106,N_28804,N_28977);
nor U29107 (N_29107,N_28522,N_28937);
nand U29108 (N_29108,N_28956,N_28585);
or U29109 (N_29109,N_28841,N_28833);
or U29110 (N_29110,N_28521,N_28959);
or U29111 (N_29111,N_28787,N_28696);
nand U29112 (N_29112,N_28929,N_28919);
nor U29113 (N_29113,N_28828,N_28635);
and U29114 (N_29114,N_28992,N_28838);
xnor U29115 (N_29115,N_28578,N_28768);
nand U29116 (N_29116,N_28544,N_28793);
xnor U29117 (N_29117,N_28541,N_28684);
nor U29118 (N_29118,N_28987,N_28938);
nand U29119 (N_29119,N_28955,N_28513);
and U29120 (N_29120,N_28737,N_28575);
and U29121 (N_29121,N_28664,N_28879);
or U29122 (N_29122,N_28730,N_28593);
nand U29123 (N_29123,N_28729,N_28669);
nand U29124 (N_29124,N_28653,N_28530);
or U29125 (N_29125,N_28652,N_28678);
nor U29126 (N_29126,N_28973,N_28891);
xor U29127 (N_29127,N_28747,N_28587);
and U29128 (N_29128,N_28970,N_28866);
and U29129 (N_29129,N_28950,N_28622);
xnor U29130 (N_29130,N_28611,N_28877);
or U29131 (N_29131,N_28916,N_28805);
nand U29132 (N_29132,N_28563,N_28734);
or U29133 (N_29133,N_28790,N_28837);
xnor U29134 (N_29134,N_28648,N_28753);
and U29135 (N_29135,N_28840,N_28871);
and U29136 (N_29136,N_28774,N_28862);
xnor U29137 (N_29137,N_28547,N_28948);
or U29138 (N_29138,N_28692,N_28577);
and U29139 (N_29139,N_28738,N_28817);
and U29140 (N_29140,N_28634,N_28735);
or U29141 (N_29141,N_28878,N_28980);
nor U29142 (N_29142,N_28913,N_28671);
xor U29143 (N_29143,N_28581,N_28748);
xnor U29144 (N_29144,N_28539,N_28595);
and U29145 (N_29145,N_28761,N_28579);
nand U29146 (N_29146,N_28702,N_28797);
and U29147 (N_29147,N_28966,N_28536);
nor U29148 (N_29148,N_28941,N_28654);
nand U29149 (N_29149,N_28512,N_28520);
and U29150 (N_29150,N_28693,N_28528);
xor U29151 (N_29151,N_28960,N_28633);
or U29152 (N_29152,N_28629,N_28604);
xor U29153 (N_29153,N_28552,N_28607);
xor U29154 (N_29154,N_28850,N_28858);
or U29155 (N_29155,N_28957,N_28887);
nor U29156 (N_29156,N_28658,N_28788);
or U29157 (N_29157,N_28961,N_28807);
and U29158 (N_29158,N_28931,N_28863);
nand U29159 (N_29159,N_28527,N_28899);
or U29160 (N_29160,N_28851,N_28700);
nor U29161 (N_29161,N_28712,N_28812);
nand U29162 (N_29162,N_28742,N_28570);
nor U29163 (N_29163,N_28553,N_28609);
and U29164 (N_29164,N_28601,N_28508);
nand U29165 (N_29165,N_28538,N_28822);
or U29166 (N_29166,N_28529,N_28835);
or U29167 (N_29167,N_28686,N_28558);
and U29168 (N_29168,N_28796,N_28945);
and U29169 (N_29169,N_28848,N_28926);
nand U29170 (N_29170,N_28769,N_28710);
or U29171 (N_29171,N_28705,N_28906);
and U29172 (N_29172,N_28596,N_28699);
nand U29173 (N_29173,N_28582,N_28802);
nor U29174 (N_29174,N_28912,N_28988);
or U29175 (N_29175,N_28627,N_28827);
xnor U29176 (N_29176,N_28975,N_28925);
nor U29177 (N_29177,N_28731,N_28909);
nand U29178 (N_29178,N_28829,N_28580);
xor U29179 (N_29179,N_28511,N_28911);
xor U29180 (N_29180,N_28616,N_28687);
nor U29181 (N_29181,N_28922,N_28799);
or U29182 (N_29182,N_28554,N_28777);
nand U29183 (N_29183,N_28509,N_28810);
nand U29184 (N_29184,N_28605,N_28566);
nand U29185 (N_29185,N_28610,N_28875);
xor U29186 (N_29186,N_28983,N_28854);
or U29187 (N_29187,N_28650,N_28613);
nor U29188 (N_29188,N_28500,N_28617);
or U29189 (N_29189,N_28949,N_28562);
or U29190 (N_29190,N_28727,N_28526);
nand U29191 (N_29191,N_28505,N_28890);
nand U29192 (N_29192,N_28515,N_28910);
or U29193 (N_29193,N_28811,N_28586);
and U29194 (N_29194,N_28936,N_28619);
and U29195 (N_29195,N_28726,N_28745);
nand U29196 (N_29196,N_28685,N_28990);
nand U29197 (N_29197,N_28688,N_28943);
and U29198 (N_29198,N_28565,N_28809);
nor U29199 (N_29199,N_28741,N_28632);
nor U29200 (N_29200,N_28646,N_28724);
nor U29201 (N_29201,N_28591,N_28985);
and U29202 (N_29202,N_28732,N_28934);
and U29203 (N_29203,N_28631,N_28641);
or U29204 (N_29204,N_28895,N_28830);
or U29205 (N_29205,N_28639,N_28962);
xor U29206 (N_29206,N_28800,N_28740);
nand U29207 (N_29207,N_28716,N_28897);
nand U29208 (N_29208,N_28865,N_28806);
xnor U29209 (N_29209,N_28981,N_28880);
or U29210 (N_29210,N_28556,N_28503);
and U29211 (N_29211,N_28771,N_28861);
or U29212 (N_29212,N_28542,N_28524);
nand U29213 (N_29213,N_28832,N_28624);
xnor U29214 (N_29214,N_28991,N_28757);
and U29215 (N_29215,N_28551,N_28736);
nor U29216 (N_29216,N_28672,N_28892);
or U29217 (N_29217,N_28564,N_28680);
and U29218 (N_29218,N_28958,N_28643);
or U29219 (N_29219,N_28589,N_28842);
nor U29220 (N_29220,N_28882,N_28750);
and U29221 (N_29221,N_28791,N_28567);
nor U29222 (N_29222,N_28717,N_28758);
nor U29223 (N_29223,N_28561,N_28555);
xnor U29224 (N_29224,N_28588,N_28708);
nand U29225 (N_29225,N_28718,N_28690);
xnor U29226 (N_29226,N_28780,N_28594);
nor U29227 (N_29227,N_28967,N_28659);
nor U29228 (N_29228,N_28656,N_28819);
xor U29229 (N_29229,N_28932,N_28775);
nor U29230 (N_29230,N_28859,N_28781);
or U29231 (N_29231,N_28625,N_28590);
xnor U29232 (N_29232,N_28703,N_28573);
nand U29233 (N_29233,N_28963,N_28933);
and U29234 (N_29234,N_28706,N_28721);
xnor U29235 (N_29235,N_28874,N_28647);
and U29236 (N_29236,N_28673,N_28942);
xor U29237 (N_29237,N_28597,N_28739);
xnor U29238 (N_29238,N_28630,N_28733);
xor U29239 (N_29239,N_28834,N_28644);
or U29240 (N_29240,N_28993,N_28814);
xnor U29241 (N_29241,N_28548,N_28824);
nor U29242 (N_29242,N_28924,N_28843);
or U29243 (N_29243,N_28914,N_28849);
or U29244 (N_29244,N_28638,N_28789);
or U29245 (N_29245,N_28531,N_28770);
xor U29246 (N_29246,N_28927,N_28951);
and U29247 (N_29247,N_28719,N_28691);
and U29248 (N_29248,N_28618,N_28626);
nor U29249 (N_29249,N_28855,N_28979);
nand U29250 (N_29250,N_28764,N_28789);
nor U29251 (N_29251,N_28796,N_28805);
nand U29252 (N_29252,N_28660,N_28757);
or U29253 (N_29253,N_28635,N_28576);
and U29254 (N_29254,N_28822,N_28806);
nand U29255 (N_29255,N_28511,N_28936);
nor U29256 (N_29256,N_28651,N_28554);
and U29257 (N_29257,N_28817,N_28679);
xor U29258 (N_29258,N_28811,N_28605);
nor U29259 (N_29259,N_28760,N_28871);
and U29260 (N_29260,N_28793,N_28954);
xnor U29261 (N_29261,N_28708,N_28615);
nor U29262 (N_29262,N_28889,N_28942);
and U29263 (N_29263,N_28793,N_28779);
xnor U29264 (N_29264,N_28883,N_28815);
nand U29265 (N_29265,N_28999,N_28626);
or U29266 (N_29266,N_28896,N_28935);
nor U29267 (N_29267,N_28624,N_28917);
xnor U29268 (N_29268,N_28508,N_28972);
and U29269 (N_29269,N_28571,N_28834);
nor U29270 (N_29270,N_28755,N_28861);
or U29271 (N_29271,N_28831,N_28958);
nor U29272 (N_29272,N_28820,N_28605);
nand U29273 (N_29273,N_28913,N_28731);
xor U29274 (N_29274,N_28687,N_28544);
and U29275 (N_29275,N_28621,N_28850);
xnor U29276 (N_29276,N_28858,N_28581);
nand U29277 (N_29277,N_28676,N_28900);
xor U29278 (N_29278,N_28543,N_28516);
nor U29279 (N_29279,N_28598,N_28531);
nand U29280 (N_29280,N_28612,N_28515);
xor U29281 (N_29281,N_28663,N_28910);
and U29282 (N_29282,N_28710,N_28582);
and U29283 (N_29283,N_28903,N_28894);
or U29284 (N_29284,N_28701,N_28849);
and U29285 (N_29285,N_28624,N_28642);
xnor U29286 (N_29286,N_28898,N_28811);
nor U29287 (N_29287,N_28690,N_28630);
xor U29288 (N_29288,N_28625,N_28860);
xor U29289 (N_29289,N_28933,N_28846);
nand U29290 (N_29290,N_28988,N_28821);
nand U29291 (N_29291,N_28574,N_28671);
and U29292 (N_29292,N_28574,N_28797);
xnor U29293 (N_29293,N_28906,N_28833);
or U29294 (N_29294,N_28574,N_28577);
and U29295 (N_29295,N_28925,N_28747);
nand U29296 (N_29296,N_28792,N_28597);
or U29297 (N_29297,N_28529,N_28566);
xnor U29298 (N_29298,N_28686,N_28799);
or U29299 (N_29299,N_28653,N_28857);
and U29300 (N_29300,N_28865,N_28810);
xor U29301 (N_29301,N_28896,N_28627);
nor U29302 (N_29302,N_28541,N_28822);
or U29303 (N_29303,N_28693,N_28916);
nand U29304 (N_29304,N_28954,N_28558);
xnor U29305 (N_29305,N_28866,N_28963);
and U29306 (N_29306,N_28729,N_28709);
nor U29307 (N_29307,N_28561,N_28775);
and U29308 (N_29308,N_28518,N_28921);
nand U29309 (N_29309,N_28623,N_28843);
nor U29310 (N_29310,N_28684,N_28794);
xnor U29311 (N_29311,N_28826,N_28714);
and U29312 (N_29312,N_28532,N_28556);
xnor U29313 (N_29313,N_28843,N_28791);
or U29314 (N_29314,N_28971,N_28611);
nor U29315 (N_29315,N_28533,N_28967);
or U29316 (N_29316,N_28971,N_28712);
nand U29317 (N_29317,N_28887,N_28903);
or U29318 (N_29318,N_28825,N_28755);
nand U29319 (N_29319,N_28504,N_28655);
or U29320 (N_29320,N_28954,N_28876);
xor U29321 (N_29321,N_28798,N_28600);
or U29322 (N_29322,N_28846,N_28656);
xnor U29323 (N_29323,N_28555,N_28919);
or U29324 (N_29324,N_28991,N_28640);
xor U29325 (N_29325,N_28971,N_28636);
or U29326 (N_29326,N_28821,N_28687);
nor U29327 (N_29327,N_28947,N_28597);
or U29328 (N_29328,N_28841,N_28888);
xnor U29329 (N_29329,N_28958,N_28542);
nor U29330 (N_29330,N_28851,N_28921);
nand U29331 (N_29331,N_28880,N_28787);
or U29332 (N_29332,N_28912,N_28915);
nand U29333 (N_29333,N_28852,N_28543);
nand U29334 (N_29334,N_28740,N_28997);
or U29335 (N_29335,N_28608,N_28705);
and U29336 (N_29336,N_28734,N_28772);
and U29337 (N_29337,N_28783,N_28949);
nand U29338 (N_29338,N_28741,N_28506);
nand U29339 (N_29339,N_28661,N_28684);
xor U29340 (N_29340,N_28845,N_28973);
and U29341 (N_29341,N_28677,N_28920);
nor U29342 (N_29342,N_28571,N_28671);
nand U29343 (N_29343,N_28586,N_28643);
and U29344 (N_29344,N_28772,N_28963);
or U29345 (N_29345,N_28506,N_28881);
nor U29346 (N_29346,N_28921,N_28880);
and U29347 (N_29347,N_28606,N_28972);
nor U29348 (N_29348,N_28605,N_28805);
and U29349 (N_29349,N_28503,N_28957);
xor U29350 (N_29350,N_28582,N_28792);
or U29351 (N_29351,N_28940,N_28572);
nor U29352 (N_29352,N_28540,N_28708);
and U29353 (N_29353,N_28632,N_28619);
xnor U29354 (N_29354,N_28978,N_28681);
xnor U29355 (N_29355,N_28571,N_28508);
nand U29356 (N_29356,N_28877,N_28608);
nor U29357 (N_29357,N_28883,N_28702);
nor U29358 (N_29358,N_28994,N_28891);
or U29359 (N_29359,N_28966,N_28676);
and U29360 (N_29360,N_28992,N_28965);
nor U29361 (N_29361,N_28505,N_28881);
nor U29362 (N_29362,N_28886,N_28988);
and U29363 (N_29363,N_28702,N_28568);
xor U29364 (N_29364,N_28795,N_28693);
xor U29365 (N_29365,N_28533,N_28864);
nand U29366 (N_29366,N_28535,N_28711);
xnor U29367 (N_29367,N_28591,N_28865);
and U29368 (N_29368,N_28506,N_28667);
nand U29369 (N_29369,N_28934,N_28746);
nand U29370 (N_29370,N_28743,N_28876);
nor U29371 (N_29371,N_28752,N_28655);
nor U29372 (N_29372,N_28539,N_28772);
xor U29373 (N_29373,N_28640,N_28736);
nand U29374 (N_29374,N_28956,N_28686);
xnor U29375 (N_29375,N_28529,N_28628);
and U29376 (N_29376,N_28702,N_28937);
nor U29377 (N_29377,N_28934,N_28602);
nor U29378 (N_29378,N_28875,N_28790);
nor U29379 (N_29379,N_28776,N_28780);
nand U29380 (N_29380,N_28813,N_28649);
nor U29381 (N_29381,N_28648,N_28626);
and U29382 (N_29382,N_28971,N_28679);
nand U29383 (N_29383,N_28775,N_28844);
nand U29384 (N_29384,N_28605,N_28980);
nand U29385 (N_29385,N_28512,N_28985);
xnor U29386 (N_29386,N_28888,N_28600);
xor U29387 (N_29387,N_28626,N_28712);
nor U29388 (N_29388,N_28885,N_28941);
nand U29389 (N_29389,N_28571,N_28649);
and U29390 (N_29390,N_28800,N_28568);
nand U29391 (N_29391,N_28974,N_28945);
xor U29392 (N_29392,N_28960,N_28611);
nand U29393 (N_29393,N_28993,N_28827);
nor U29394 (N_29394,N_28619,N_28510);
nor U29395 (N_29395,N_28744,N_28811);
nand U29396 (N_29396,N_28565,N_28615);
nor U29397 (N_29397,N_28833,N_28580);
xnor U29398 (N_29398,N_28831,N_28696);
nor U29399 (N_29399,N_28687,N_28971);
nor U29400 (N_29400,N_28691,N_28508);
and U29401 (N_29401,N_28743,N_28735);
and U29402 (N_29402,N_28551,N_28912);
or U29403 (N_29403,N_28965,N_28948);
nor U29404 (N_29404,N_28641,N_28917);
xnor U29405 (N_29405,N_28503,N_28958);
xor U29406 (N_29406,N_28543,N_28790);
and U29407 (N_29407,N_28688,N_28752);
nand U29408 (N_29408,N_28809,N_28625);
nand U29409 (N_29409,N_28792,N_28846);
and U29410 (N_29410,N_28624,N_28933);
or U29411 (N_29411,N_28504,N_28868);
or U29412 (N_29412,N_28591,N_28589);
nand U29413 (N_29413,N_28815,N_28732);
or U29414 (N_29414,N_28732,N_28942);
nand U29415 (N_29415,N_28580,N_28534);
or U29416 (N_29416,N_28754,N_28509);
nor U29417 (N_29417,N_28686,N_28899);
nor U29418 (N_29418,N_28915,N_28754);
nor U29419 (N_29419,N_28711,N_28966);
nand U29420 (N_29420,N_28534,N_28941);
nand U29421 (N_29421,N_28768,N_28566);
nand U29422 (N_29422,N_28935,N_28841);
or U29423 (N_29423,N_28778,N_28960);
nand U29424 (N_29424,N_28906,N_28838);
or U29425 (N_29425,N_28508,N_28827);
nand U29426 (N_29426,N_28859,N_28780);
and U29427 (N_29427,N_28689,N_28968);
and U29428 (N_29428,N_28612,N_28756);
and U29429 (N_29429,N_28536,N_28999);
xor U29430 (N_29430,N_28783,N_28977);
xnor U29431 (N_29431,N_28698,N_28572);
or U29432 (N_29432,N_28878,N_28756);
nand U29433 (N_29433,N_28855,N_28936);
nor U29434 (N_29434,N_28879,N_28773);
nand U29435 (N_29435,N_28651,N_28577);
nand U29436 (N_29436,N_28737,N_28626);
or U29437 (N_29437,N_28617,N_28937);
xnor U29438 (N_29438,N_28950,N_28892);
or U29439 (N_29439,N_28553,N_28746);
nor U29440 (N_29440,N_28564,N_28698);
xnor U29441 (N_29441,N_28922,N_28831);
and U29442 (N_29442,N_28513,N_28782);
or U29443 (N_29443,N_28523,N_28789);
nand U29444 (N_29444,N_28656,N_28581);
nor U29445 (N_29445,N_28610,N_28791);
and U29446 (N_29446,N_28913,N_28708);
nand U29447 (N_29447,N_28800,N_28570);
xor U29448 (N_29448,N_28588,N_28668);
nand U29449 (N_29449,N_28513,N_28615);
nand U29450 (N_29450,N_28839,N_28659);
or U29451 (N_29451,N_28500,N_28765);
or U29452 (N_29452,N_28586,N_28510);
nor U29453 (N_29453,N_28729,N_28523);
xor U29454 (N_29454,N_28528,N_28633);
nor U29455 (N_29455,N_28593,N_28637);
and U29456 (N_29456,N_28605,N_28537);
nor U29457 (N_29457,N_28885,N_28780);
nand U29458 (N_29458,N_28934,N_28864);
xor U29459 (N_29459,N_28876,N_28723);
nand U29460 (N_29460,N_28539,N_28564);
and U29461 (N_29461,N_28834,N_28941);
nand U29462 (N_29462,N_28718,N_28924);
and U29463 (N_29463,N_28763,N_28825);
nor U29464 (N_29464,N_28888,N_28881);
nor U29465 (N_29465,N_28730,N_28920);
nand U29466 (N_29466,N_28979,N_28659);
or U29467 (N_29467,N_28899,N_28935);
nor U29468 (N_29468,N_28699,N_28542);
and U29469 (N_29469,N_28825,N_28871);
xor U29470 (N_29470,N_28543,N_28824);
nand U29471 (N_29471,N_28737,N_28578);
and U29472 (N_29472,N_28806,N_28625);
and U29473 (N_29473,N_28690,N_28657);
xor U29474 (N_29474,N_28620,N_28733);
or U29475 (N_29475,N_28622,N_28640);
nor U29476 (N_29476,N_28980,N_28915);
xor U29477 (N_29477,N_28973,N_28970);
nor U29478 (N_29478,N_28674,N_28623);
xnor U29479 (N_29479,N_28834,N_28725);
nand U29480 (N_29480,N_28943,N_28603);
and U29481 (N_29481,N_28751,N_28510);
and U29482 (N_29482,N_28606,N_28503);
or U29483 (N_29483,N_28544,N_28825);
nor U29484 (N_29484,N_28721,N_28990);
or U29485 (N_29485,N_28865,N_28748);
or U29486 (N_29486,N_28797,N_28956);
nand U29487 (N_29487,N_28869,N_28831);
nand U29488 (N_29488,N_28621,N_28889);
nand U29489 (N_29489,N_28621,N_28816);
xnor U29490 (N_29490,N_28921,N_28819);
xnor U29491 (N_29491,N_28749,N_28719);
and U29492 (N_29492,N_28548,N_28909);
and U29493 (N_29493,N_28810,N_28961);
and U29494 (N_29494,N_28881,N_28719);
and U29495 (N_29495,N_28594,N_28977);
or U29496 (N_29496,N_28705,N_28798);
nor U29497 (N_29497,N_28543,N_28561);
nand U29498 (N_29498,N_28853,N_28614);
nor U29499 (N_29499,N_28720,N_28565);
or U29500 (N_29500,N_29333,N_29279);
or U29501 (N_29501,N_29434,N_29470);
nand U29502 (N_29502,N_29008,N_29144);
xnor U29503 (N_29503,N_29000,N_29399);
or U29504 (N_29504,N_29360,N_29440);
xor U29505 (N_29505,N_29115,N_29067);
or U29506 (N_29506,N_29337,N_29283);
nor U29507 (N_29507,N_29353,N_29327);
nand U29508 (N_29508,N_29347,N_29173);
nor U29509 (N_29509,N_29082,N_29230);
nor U29510 (N_29510,N_29373,N_29338);
and U29511 (N_29511,N_29299,N_29296);
xnor U29512 (N_29512,N_29081,N_29344);
and U29513 (N_29513,N_29411,N_29492);
or U29514 (N_29514,N_29107,N_29392);
nand U29515 (N_29515,N_29346,N_29228);
xnor U29516 (N_29516,N_29331,N_29354);
and U29517 (N_29517,N_29127,N_29112);
xor U29518 (N_29518,N_29118,N_29076);
or U29519 (N_29519,N_29059,N_29223);
nor U29520 (N_29520,N_29456,N_29010);
nand U29521 (N_29521,N_29086,N_29121);
nand U29522 (N_29522,N_29015,N_29182);
nor U29523 (N_29523,N_29336,N_29320);
xnor U29524 (N_29524,N_29050,N_29164);
and U29525 (N_29525,N_29464,N_29437);
nor U29526 (N_29526,N_29404,N_29397);
or U29527 (N_29527,N_29140,N_29487);
or U29528 (N_29528,N_29055,N_29060);
or U29529 (N_29529,N_29466,N_29237);
and U29530 (N_29530,N_29039,N_29023);
and U29531 (N_29531,N_29251,N_29341);
xnor U29532 (N_29532,N_29161,N_29450);
nand U29533 (N_29533,N_29350,N_29137);
nand U29534 (N_29534,N_29190,N_29018);
or U29535 (N_29535,N_29097,N_29271);
nor U29536 (N_29536,N_29210,N_29222);
nand U29537 (N_29537,N_29075,N_29020);
xor U29538 (N_29538,N_29458,N_29229);
nand U29539 (N_29539,N_29294,N_29049);
and U29540 (N_29540,N_29195,N_29461);
and U29541 (N_29541,N_29430,N_29024);
nand U29542 (N_29542,N_29415,N_29034);
xnor U29543 (N_29543,N_29252,N_29138);
nor U29544 (N_29544,N_29315,N_29048);
and U29545 (N_29545,N_29258,N_29349);
or U29546 (N_29546,N_29145,N_29386);
xnor U29547 (N_29547,N_29358,N_29162);
nand U29548 (N_29548,N_29212,N_29125);
nand U29549 (N_29549,N_29382,N_29045);
nand U29550 (N_29550,N_29043,N_29316);
nand U29551 (N_29551,N_29484,N_29168);
xor U29552 (N_29552,N_29239,N_29468);
or U29553 (N_29553,N_29088,N_29499);
or U29554 (N_29554,N_29051,N_29384);
or U29555 (N_29555,N_29197,N_29135);
nand U29556 (N_29556,N_29038,N_29165);
nor U29557 (N_29557,N_29106,N_29019);
or U29558 (N_29558,N_29486,N_29143);
and U29559 (N_29559,N_29136,N_29198);
nor U29560 (N_29560,N_29236,N_29268);
and U29561 (N_29561,N_29416,N_29069);
xnor U29562 (N_29562,N_29080,N_29249);
nand U29563 (N_29563,N_29167,N_29184);
and U29564 (N_29564,N_29203,N_29063);
or U29565 (N_29565,N_29479,N_29278);
or U29566 (N_29566,N_29232,N_29070);
nand U29567 (N_29567,N_29231,N_29455);
and U29568 (N_29568,N_29058,N_29100);
xnor U29569 (N_29569,N_29032,N_29359);
nor U29570 (N_29570,N_29412,N_29089);
or U29571 (N_29571,N_29166,N_29219);
nor U29572 (N_29572,N_29340,N_29066);
nor U29573 (N_29573,N_29016,N_29240);
nor U29574 (N_29574,N_29157,N_29451);
nand U29575 (N_29575,N_29262,N_29409);
nor U29576 (N_29576,N_29188,N_29351);
or U29577 (N_29577,N_29323,N_29227);
or U29578 (N_29578,N_29348,N_29357);
xor U29579 (N_29579,N_29273,N_29319);
and U29580 (N_29580,N_29445,N_29491);
or U29581 (N_29581,N_29403,N_29079);
xor U29582 (N_29582,N_29306,N_29009);
or U29583 (N_29583,N_29269,N_29037);
nand U29584 (N_29584,N_29095,N_29194);
or U29585 (N_29585,N_29110,N_29021);
nor U29586 (N_29586,N_29224,N_29208);
nor U29587 (N_29587,N_29318,N_29093);
and U29588 (N_29588,N_29493,N_29314);
nand U29589 (N_29589,N_29036,N_29092);
nand U29590 (N_29590,N_29290,N_29098);
or U29591 (N_29591,N_29234,N_29207);
and U29592 (N_29592,N_29003,N_29176);
nand U29593 (N_29593,N_29419,N_29281);
or U29594 (N_29594,N_29396,N_29426);
nand U29595 (N_29595,N_29496,N_29463);
and U29596 (N_29596,N_29465,N_29431);
nand U29597 (N_29597,N_29180,N_29295);
nor U29598 (N_29598,N_29356,N_29413);
or U29599 (N_29599,N_29376,N_29477);
xnor U29600 (N_29600,N_29142,N_29117);
nor U29601 (N_29601,N_29233,N_29033);
nand U29602 (N_29602,N_29425,N_29343);
and U29603 (N_29603,N_29339,N_29150);
nand U29604 (N_29604,N_29196,N_29119);
xnor U29605 (N_29605,N_29122,N_29245);
xnor U29606 (N_29606,N_29213,N_29047);
and U29607 (N_29607,N_29374,N_29146);
nand U29608 (N_29608,N_29361,N_29061);
xor U29609 (N_29609,N_29124,N_29427);
and U29610 (N_29610,N_29334,N_29056);
nor U29611 (N_29611,N_29453,N_29375);
xor U29612 (N_29612,N_29191,N_29389);
nand U29613 (N_29613,N_29482,N_29292);
or U29614 (N_29614,N_29495,N_29209);
or U29615 (N_29615,N_29474,N_29387);
and U29616 (N_29616,N_29498,N_29275);
nor U29617 (N_29617,N_29276,N_29104);
xnor U29618 (N_29618,N_29041,N_29446);
or U29619 (N_29619,N_29134,N_29305);
nor U29620 (N_29620,N_29368,N_29235);
nor U29621 (N_29621,N_29307,N_29154);
nand U29622 (N_29622,N_29454,N_29225);
or U29623 (N_29623,N_29129,N_29291);
nand U29624 (N_29624,N_29027,N_29408);
and U29625 (N_29625,N_29324,N_29226);
xor U29626 (N_29626,N_29149,N_29469);
or U29627 (N_29627,N_29052,N_29418);
nor U29628 (N_29628,N_29062,N_29332);
and U29629 (N_29629,N_29270,N_29345);
xnor U29630 (N_29630,N_29172,N_29030);
and U29631 (N_29631,N_29179,N_29366);
nand U29632 (N_29632,N_29090,N_29029);
nor U29633 (N_29633,N_29309,N_29256);
nor U29634 (N_29634,N_29028,N_29113);
nand U29635 (N_29635,N_29116,N_29204);
and U29636 (N_29636,N_29417,N_29467);
nor U29637 (N_29637,N_29057,N_29201);
nor U29638 (N_29638,N_29065,N_29111);
nand U29639 (N_29639,N_29071,N_29485);
xor U29640 (N_29640,N_29311,N_29211);
or U29641 (N_29641,N_29308,N_29429);
nand U29642 (N_29642,N_29402,N_29302);
nand U29643 (N_29643,N_29202,N_29388);
nor U29644 (N_29644,N_29293,N_29253);
xor U29645 (N_29645,N_29178,N_29126);
nor U29646 (N_29646,N_29013,N_29254);
nand U29647 (N_29647,N_29014,N_29006);
nor U29648 (N_29648,N_29329,N_29420);
or U29649 (N_29649,N_29170,N_29216);
nand U29650 (N_29650,N_29459,N_29321);
nor U29651 (N_29651,N_29310,N_29200);
nor U29652 (N_29652,N_29432,N_29390);
nand U29653 (N_29653,N_29159,N_29289);
or U29654 (N_29654,N_29365,N_29266);
nand U29655 (N_29655,N_29328,N_29087);
nor U29656 (N_29656,N_29449,N_29246);
nand U29657 (N_29657,N_29217,N_29114);
or U29658 (N_29658,N_29109,N_29395);
and U29659 (N_29659,N_29448,N_29322);
and U29660 (N_29660,N_29263,N_29105);
nor U29661 (N_29661,N_29439,N_29367);
nand U29662 (N_29662,N_29285,N_29436);
or U29663 (N_29663,N_29181,N_29096);
xor U29664 (N_29664,N_29193,N_29185);
nor U29665 (N_29665,N_29460,N_29379);
nand U29666 (N_29666,N_29005,N_29101);
and U29667 (N_29667,N_29447,N_29264);
or U29668 (N_29668,N_29152,N_29383);
xnor U29669 (N_29669,N_29011,N_29335);
xnor U29670 (N_29670,N_29192,N_29280);
or U29671 (N_29671,N_29001,N_29241);
and U29672 (N_29672,N_29085,N_29133);
or U29673 (N_29673,N_29481,N_29099);
xnor U29674 (N_29674,N_29094,N_29444);
nand U29675 (N_29675,N_29288,N_29364);
nand U29676 (N_29676,N_29186,N_29483);
nand U29677 (N_29677,N_29406,N_29068);
xnor U29678 (N_29678,N_29132,N_29401);
and U29679 (N_29679,N_29205,N_29083);
and U29680 (N_29680,N_29298,N_29489);
nand U29681 (N_29681,N_29371,N_29177);
xnor U29682 (N_29682,N_29073,N_29064);
xnor U29683 (N_29683,N_29480,N_29171);
nand U29684 (N_29684,N_29035,N_29274);
or U29685 (N_29685,N_29091,N_29398);
and U29686 (N_29686,N_29442,N_29490);
nor U29687 (N_29687,N_29370,N_29473);
xor U29688 (N_29688,N_29244,N_29218);
xor U29689 (N_29689,N_29151,N_29300);
and U29690 (N_29690,N_29072,N_29153);
or U29691 (N_29691,N_29312,N_29247);
and U29692 (N_29692,N_29031,N_29287);
nand U29693 (N_29693,N_29054,N_29243);
xnor U29694 (N_29694,N_29025,N_29433);
or U29695 (N_29695,N_29488,N_29206);
and U29696 (N_29696,N_29255,N_29123);
nor U29697 (N_29697,N_29272,N_29163);
xnor U29698 (N_29698,N_29317,N_29261);
and U29699 (N_29699,N_29120,N_29325);
or U29700 (N_29700,N_29257,N_29297);
nor U29701 (N_29701,N_29372,N_29304);
nand U29702 (N_29702,N_29183,N_29260);
or U29703 (N_29703,N_29326,N_29084);
nand U29704 (N_29704,N_29284,N_29221);
xor U29705 (N_29705,N_29475,N_29017);
nor U29706 (N_29706,N_29022,N_29303);
xor U29707 (N_29707,N_29053,N_29405);
and U29708 (N_29708,N_29128,N_29002);
nand U29709 (N_29709,N_29435,N_29378);
and U29710 (N_29710,N_29074,N_29497);
nand U29711 (N_29711,N_29199,N_29410);
and U29712 (N_29712,N_29385,N_29301);
xor U29713 (N_29713,N_29393,N_29160);
xnor U29714 (N_29714,N_29220,N_29369);
or U29715 (N_29715,N_29286,N_29428);
or U29716 (N_29716,N_29250,N_29423);
and U29717 (N_29717,N_29248,N_29342);
nor U29718 (N_29718,N_29044,N_29380);
nor U29719 (N_29719,N_29141,N_29130);
xor U29720 (N_29720,N_29238,N_29478);
nor U29721 (N_29721,N_29147,N_29363);
xor U29722 (N_29722,N_29155,N_29352);
xor U29723 (N_29723,N_29494,N_29169);
nor U29724 (N_29724,N_29441,N_29452);
nor U29725 (N_29725,N_29422,N_29004);
nor U29726 (N_29726,N_29443,N_29215);
and U29727 (N_29727,N_29046,N_29077);
nand U29728 (N_29728,N_29242,N_29313);
nand U29729 (N_29729,N_29391,N_29026);
or U29730 (N_29730,N_29421,N_29189);
nand U29731 (N_29731,N_29394,N_29148);
xor U29732 (N_29732,N_29174,N_29040);
or U29733 (N_29733,N_29078,N_29265);
nand U29734 (N_29734,N_29330,N_29012);
and U29735 (N_29735,N_29438,N_29007);
xor U29736 (N_29736,N_29472,N_29377);
nand U29737 (N_29737,N_29103,N_29259);
or U29738 (N_29738,N_29400,N_29414);
or U29739 (N_29739,N_29102,N_29424);
and U29740 (N_29740,N_29108,N_29381);
xor U29741 (N_29741,N_29158,N_29476);
nand U29742 (N_29742,N_29131,N_29042);
and U29743 (N_29743,N_29139,N_29462);
nand U29744 (N_29744,N_29187,N_29355);
nor U29745 (N_29745,N_29457,N_29175);
and U29746 (N_29746,N_29277,N_29471);
nor U29747 (N_29747,N_29156,N_29214);
nand U29748 (N_29748,N_29362,N_29282);
nor U29749 (N_29749,N_29407,N_29267);
nand U29750 (N_29750,N_29355,N_29122);
nor U29751 (N_29751,N_29142,N_29029);
nand U29752 (N_29752,N_29044,N_29131);
and U29753 (N_29753,N_29350,N_29424);
and U29754 (N_29754,N_29473,N_29475);
or U29755 (N_29755,N_29323,N_29101);
xnor U29756 (N_29756,N_29400,N_29107);
nor U29757 (N_29757,N_29379,N_29244);
or U29758 (N_29758,N_29366,N_29269);
and U29759 (N_29759,N_29296,N_29417);
xnor U29760 (N_29760,N_29497,N_29250);
and U29761 (N_29761,N_29473,N_29229);
nand U29762 (N_29762,N_29058,N_29048);
and U29763 (N_29763,N_29202,N_29143);
nor U29764 (N_29764,N_29220,N_29269);
nor U29765 (N_29765,N_29067,N_29037);
nor U29766 (N_29766,N_29128,N_29216);
nor U29767 (N_29767,N_29004,N_29488);
nor U29768 (N_29768,N_29384,N_29451);
xnor U29769 (N_29769,N_29234,N_29490);
nand U29770 (N_29770,N_29180,N_29181);
xnor U29771 (N_29771,N_29348,N_29125);
and U29772 (N_29772,N_29234,N_29208);
and U29773 (N_29773,N_29162,N_29428);
and U29774 (N_29774,N_29041,N_29173);
xor U29775 (N_29775,N_29016,N_29267);
xnor U29776 (N_29776,N_29183,N_29253);
or U29777 (N_29777,N_29020,N_29127);
or U29778 (N_29778,N_29403,N_29437);
xnor U29779 (N_29779,N_29400,N_29202);
or U29780 (N_29780,N_29301,N_29295);
nor U29781 (N_29781,N_29267,N_29450);
nand U29782 (N_29782,N_29040,N_29299);
nor U29783 (N_29783,N_29458,N_29196);
nand U29784 (N_29784,N_29037,N_29327);
xnor U29785 (N_29785,N_29105,N_29223);
nand U29786 (N_29786,N_29243,N_29171);
or U29787 (N_29787,N_29389,N_29051);
nor U29788 (N_29788,N_29309,N_29325);
and U29789 (N_29789,N_29172,N_29056);
xor U29790 (N_29790,N_29243,N_29058);
or U29791 (N_29791,N_29130,N_29335);
xnor U29792 (N_29792,N_29215,N_29471);
nand U29793 (N_29793,N_29358,N_29213);
and U29794 (N_29794,N_29153,N_29014);
and U29795 (N_29795,N_29299,N_29149);
and U29796 (N_29796,N_29489,N_29175);
nand U29797 (N_29797,N_29387,N_29199);
or U29798 (N_29798,N_29085,N_29105);
or U29799 (N_29799,N_29056,N_29083);
xor U29800 (N_29800,N_29436,N_29152);
xnor U29801 (N_29801,N_29231,N_29453);
nor U29802 (N_29802,N_29168,N_29311);
nor U29803 (N_29803,N_29265,N_29282);
nor U29804 (N_29804,N_29119,N_29438);
nor U29805 (N_29805,N_29463,N_29266);
xor U29806 (N_29806,N_29397,N_29125);
or U29807 (N_29807,N_29113,N_29001);
and U29808 (N_29808,N_29426,N_29187);
nand U29809 (N_29809,N_29285,N_29489);
xnor U29810 (N_29810,N_29156,N_29074);
or U29811 (N_29811,N_29410,N_29451);
nor U29812 (N_29812,N_29195,N_29363);
nor U29813 (N_29813,N_29042,N_29488);
xnor U29814 (N_29814,N_29133,N_29363);
nor U29815 (N_29815,N_29087,N_29019);
xor U29816 (N_29816,N_29425,N_29479);
nor U29817 (N_29817,N_29039,N_29468);
and U29818 (N_29818,N_29280,N_29463);
nor U29819 (N_29819,N_29114,N_29488);
xor U29820 (N_29820,N_29131,N_29182);
xnor U29821 (N_29821,N_29090,N_29436);
xor U29822 (N_29822,N_29370,N_29397);
and U29823 (N_29823,N_29089,N_29414);
or U29824 (N_29824,N_29119,N_29344);
and U29825 (N_29825,N_29156,N_29269);
nand U29826 (N_29826,N_29369,N_29066);
xnor U29827 (N_29827,N_29213,N_29110);
or U29828 (N_29828,N_29078,N_29217);
nand U29829 (N_29829,N_29072,N_29460);
and U29830 (N_29830,N_29219,N_29483);
or U29831 (N_29831,N_29285,N_29018);
xor U29832 (N_29832,N_29073,N_29185);
or U29833 (N_29833,N_29292,N_29425);
xor U29834 (N_29834,N_29388,N_29441);
and U29835 (N_29835,N_29360,N_29110);
or U29836 (N_29836,N_29312,N_29422);
nand U29837 (N_29837,N_29292,N_29117);
xor U29838 (N_29838,N_29239,N_29424);
nand U29839 (N_29839,N_29412,N_29260);
xnor U29840 (N_29840,N_29324,N_29380);
and U29841 (N_29841,N_29433,N_29395);
and U29842 (N_29842,N_29366,N_29486);
or U29843 (N_29843,N_29008,N_29146);
nor U29844 (N_29844,N_29243,N_29343);
or U29845 (N_29845,N_29207,N_29494);
or U29846 (N_29846,N_29224,N_29099);
xor U29847 (N_29847,N_29044,N_29425);
or U29848 (N_29848,N_29453,N_29205);
nand U29849 (N_29849,N_29234,N_29107);
or U29850 (N_29850,N_29310,N_29479);
and U29851 (N_29851,N_29287,N_29414);
and U29852 (N_29852,N_29049,N_29146);
and U29853 (N_29853,N_29058,N_29163);
nand U29854 (N_29854,N_29062,N_29492);
nand U29855 (N_29855,N_29245,N_29020);
and U29856 (N_29856,N_29041,N_29015);
nand U29857 (N_29857,N_29479,N_29056);
nand U29858 (N_29858,N_29408,N_29165);
or U29859 (N_29859,N_29146,N_29251);
xor U29860 (N_29860,N_29076,N_29091);
and U29861 (N_29861,N_29357,N_29458);
and U29862 (N_29862,N_29138,N_29288);
nor U29863 (N_29863,N_29148,N_29109);
xor U29864 (N_29864,N_29139,N_29271);
or U29865 (N_29865,N_29025,N_29443);
xnor U29866 (N_29866,N_29138,N_29060);
xnor U29867 (N_29867,N_29225,N_29257);
nand U29868 (N_29868,N_29262,N_29001);
or U29869 (N_29869,N_29266,N_29166);
xnor U29870 (N_29870,N_29372,N_29296);
nand U29871 (N_29871,N_29342,N_29090);
and U29872 (N_29872,N_29053,N_29227);
and U29873 (N_29873,N_29136,N_29230);
or U29874 (N_29874,N_29290,N_29046);
xnor U29875 (N_29875,N_29319,N_29349);
nand U29876 (N_29876,N_29319,N_29080);
nand U29877 (N_29877,N_29308,N_29022);
or U29878 (N_29878,N_29335,N_29418);
nor U29879 (N_29879,N_29461,N_29077);
and U29880 (N_29880,N_29315,N_29285);
nor U29881 (N_29881,N_29452,N_29120);
nand U29882 (N_29882,N_29164,N_29165);
and U29883 (N_29883,N_29057,N_29298);
xor U29884 (N_29884,N_29423,N_29147);
nor U29885 (N_29885,N_29283,N_29486);
nand U29886 (N_29886,N_29353,N_29014);
nor U29887 (N_29887,N_29271,N_29122);
nand U29888 (N_29888,N_29016,N_29343);
or U29889 (N_29889,N_29062,N_29123);
nand U29890 (N_29890,N_29158,N_29077);
or U29891 (N_29891,N_29374,N_29452);
or U29892 (N_29892,N_29319,N_29270);
nand U29893 (N_29893,N_29430,N_29100);
or U29894 (N_29894,N_29314,N_29116);
or U29895 (N_29895,N_29423,N_29021);
or U29896 (N_29896,N_29410,N_29416);
xor U29897 (N_29897,N_29003,N_29080);
or U29898 (N_29898,N_29148,N_29128);
nand U29899 (N_29899,N_29275,N_29397);
xnor U29900 (N_29900,N_29425,N_29478);
and U29901 (N_29901,N_29357,N_29370);
xnor U29902 (N_29902,N_29232,N_29119);
xor U29903 (N_29903,N_29432,N_29371);
nor U29904 (N_29904,N_29063,N_29409);
nand U29905 (N_29905,N_29495,N_29282);
and U29906 (N_29906,N_29166,N_29347);
xor U29907 (N_29907,N_29233,N_29462);
or U29908 (N_29908,N_29215,N_29420);
nand U29909 (N_29909,N_29044,N_29426);
nor U29910 (N_29910,N_29459,N_29238);
nand U29911 (N_29911,N_29221,N_29288);
nor U29912 (N_29912,N_29174,N_29486);
xor U29913 (N_29913,N_29239,N_29442);
nand U29914 (N_29914,N_29406,N_29200);
nand U29915 (N_29915,N_29292,N_29064);
nand U29916 (N_29916,N_29102,N_29311);
xnor U29917 (N_29917,N_29471,N_29128);
and U29918 (N_29918,N_29192,N_29255);
and U29919 (N_29919,N_29079,N_29050);
xnor U29920 (N_29920,N_29430,N_29477);
or U29921 (N_29921,N_29304,N_29225);
nand U29922 (N_29922,N_29386,N_29388);
xnor U29923 (N_29923,N_29372,N_29053);
and U29924 (N_29924,N_29153,N_29047);
and U29925 (N_29925,N_29397,N_29055);
nand U29926 (N_29926,N_29071,N_29372);
and U29927 (N_29927,N_29384,N_29495);
nor U29928 (N_29928,N_29082,N_29430);
nand U29929 (N_29929,N_29113,N_29213);
xor U29930 (N_29930,N_29196,N_29075);
and U29931 (N_29931,N_29302,N_29275);
and U29932 (N_29932,N_29395,N_29042);
nand U29933 (N_29933,N_29402,N_29004);
or U29934 (N_29934,N_29430,N_29461);
nand U29935 (N_29935,N_29422,N_29216);
xor U29936 (N_29936,N_29188,N_29075);
nor U29937 (N_29937,N_29066,N_29464);
nand U29938 (N_29938,N_29240,N_29391);
nand U29939 (N_29939,N_29024,N_29255);
nor U29940 (N_29940,N_29068,N_29186);
and U29941 (N_29941,N_29440,N_29342);
and U29942 (N_29942,N_29482,N_29314);
or U29943 (N_29943,N_29405,N_29016);
or U29944 (N_29944,N_29080,N_29322);
xnor U29945 (N_29945,N_29105,N_29402);
nor U29946 (N_29946,N_29422,N_29325);
xnor U29947 (N_29947,N_29342,N_29296);
or U29948 (N_29948,N_29126,N_29094);
nor U29949 (N_29949,N_29354,N_29021);
and U29950 (N_29950,N_29329,N_29383);
or U29951 (N_29951,N_29260,N_29464);
or U29952 (N_29952,N_29041,N_29433);
or U29953 (N_29953,N_29052,N_29401);
or U29954 (N_29954,N_29061,N_29146);
and U29955 (N_29955,N_29072,N_29442);
nor U29956 (N_29956,N_29462,N_29386);
nand U29957 (N_29957,N_29389,N_29086);
or U29958 (N_29958,N_29083,N_29250);
or U29959 (N_29959,N_29051,N_29030);
nand U29960 (N_29960,N_29090,N_29018);
nand U29961 (N_29961,N_29267,N_29105);
xor U29962 (N_29962,N_29019,N_29027);
or U29963 (N_29963,N_29399,N_29050);
and U29964 (N_29964,N_29214,N_29099);
and U29965 (N_29965,N_29163,N_29498);
nor U29966 (N_29966,N_29439,N_29330);
xor U29967 (N_29967,N_29448,N_29435);
and U29968 (N_29968,N_29062,N_29079);
xor U29969 (N_29969,N_29464,N_29309);
or U29970 (N_29970,N_29484,N_29313);
or U29971 (N_29971,N_29077,N_29006);
and U29972 (N_29972,N_29469,N_29432);
or U29973 (N_29973,N_29009,N_29196);
nand U29974 (N_29974,N_29341,N_29202);
and U29975 (N_29975,N_29376,N_29400);
nor U29976 (N_29976,N_29423,N_29448);
nand U29977 (N_29977,N_29361,N_29496);
nor U29978 (N_29978,N_29121,N_29295);
xor U29979 (N_29979,N_29278,N_29404);
xnor U29980 (N_29980,N_29335,N_29394);
or U29981 (N_29981,N_29087,N_29290);
nor U29982 (N_29982,N_29064,N_29201);
xnor U29983 (N_29983,N_29247,N_29107);
nand U29984 (N_29984,N_29187,N_29106);
or U29985 (N_29985,N_29126,N_29377);
and U29986 (N_29986,N_29351,N_29158);
nor U29987 (N_29987,N_29327,N_29428);
and U29988 (N_29988,N_29081,N_29111);
nor U29989 (N_29989,N_29092,N_29379);
nand U29990 (N_29990,N_29139,N_29167);
xor U29991 (N_29991,N_29418,N_29285);
or U29992 (N_29992,N_29224,N_29461);
xnor U29993 (N_29993,N_29459,N_29495);
and U29994 (N_29994,N_29486,N_29375);
nor U29995 (N_29995,N_29153,N_29302);
xor U29996 (N_29996,N_29196,N_29310);
nor U29997 (N_29997,N_29490,N_29039);
nand U29998 (N_29998,N_29090,N_29291);
nand U29999 (N_29999,N_29016,N_29373);
and UO_0 (O_0,N_29710,N_29924);
xor UO_1 (O_1,N_29984,N_29927);
and UO_2 (O_2,N_29776,N_29723);
nand UO_3 (O_3,N_29964,N_29649);
xnor UO_4 (O_4,N_29840,N_29731);
or UO_5 (O_5,N_29683,N_29711);
nor UO_6 (O_6,N_29559,N_29989);
or UO_7 (O_7,N_29629,N_29586);
and UO_8 (O_8,N_29846,N_29635);
nor UO_9 (O_9,N_29952,N_29859);
nand UO_10 (O_10,N_29739,N_29783);
xnor UO_11 (O_11,N_29521,N_29729);
xnor UO_12 (O_12,N_29779,N_29724);
nand UO_13 (O_13,N_29614,N_29680);
or UO_14 (O_14,N_29882,N_29975);
nor UO_15 (O_15,N_29827,N_29722);
xor UO_16 (O_16,N_29906,N_29808);
nand UO_17 (O_17,N_29583,N_29895);
or UO_18 (O_18,N_29805,N_29616);
nor UO_19 (O_19,N_29738,N_29575);
xor UO_20 (O_20,N_29702,N_29932);
or UO_21 (O_21,N_29581,N_29834);
nand UO_22 (O_22,N_29589,N_29830);
nand UO_23 (O_23,N_29662,N_29936);
and UO_24 (O_24,N_29844,N_29871);
xnor UO_25 (O_25,N_29945,N_29909);
or UO_26 (O_26,N_29647,N_29637);
xor UO_27 (O_27,N_29878,N_29623);
or UO_28 (O_28,N_29593,N_29555);
and UO_29 (O_29,N_29822,N_29853);
nor UO_30 (O_30,N_29770,N_29917);
xor UO_31 (O_31,N_29860,N_29737);
nor UO_32 (O_32,N_29991,N_29780);
nand UO_33 (O_33,N_29801,N_29526);
nor UO_34 (O_34,N_29619,N_29606);
or UO_35 (O_35,N_29698,N_29762);
nand UO_36 (O_36,N_29661,N_29784);
nand UO_37 (O_37,N_29501,N_29990);
or UO_38 (O_38,N_29654,N_29807);
and UO_39 (O_39,N_29818,N_29733);
or UO_40 (O_40,N_29931,N_29512);
or UO_41 (O_41,N_29605,N_29778);
and UO_42 (O_42,N_29685,N_29826);
nor UO_43 (O_43,N_29595,N_29673);
and UO_44 (O_44,N_29796,N_29572);
or UO_45 (O_45,N_29771,N_29811);
nor UO_46 (O_46,N_29716,N_29672);
and UO_47 (O_47,N_29536,N_29767);
xnor UO_48 (O_48,N_29633,N_29751);
nand UO_49 (O_49,N_29634,N_29865);
or UO_50 (O_50,N_29684,N_29790);
nor UO_51 (O_51,N_29901,N_29929);
and UO_52 (O_52,N_29546,N_29838);
nand UO_53 (O_53,N_29788,N_29873);
nor UO_54 (O_54,N_29877,N_29653);
xnor UO_55 (O_55,N_29824,N_29884);
or UO_56 (O_56,N_29506,N_29785);
nor UO_57 (O_57,N_29735,N_29502);
or UO_58 (O_58,N_29695,N_29626);
nor UO_59 (O_59,N_29837,N_29617);
xor UO_60 (O_60,N_29576,N_29571);
and UO_61 (O_61,N_29786,N_29912);
nor UO_62 (O_62,N_29919,N_29957);
xor UO_63 (O_63,N_29675,N_29507);
and UO_64 (O_64,N_29930,N_29892);
and UO_65 (O_65,N_29823,N_29750);
nand UO_66 (O_66,N_29959,N_29712);
nor UO_67 (O_67,N_29797,N_29569);
nor UO_68 (O_68,N_29718,N_29773);
and UO_69 (O_69,N_29696,N_29627);
and UO_70 (O_70,N_29632,N_29867);
or UO_71 (O_71,N_29851,N_29579);
nand UO_72 (O_72,N_29578,N_29941);
and UO_73 (O_73,N_29652,N_29803);
xor UO_74 (O_74,N_29821,N_29791);
and UO_75 (O_75,N_29999,N_29510);
nor UO_76 (O_76,N_29624,N_29709);
and UO_77 (O_77,N_29728,N_29833);
xnor UO_78 (O_78,N_29670,N_29641);
or UO_79 (O_79,N_29925,N_29886);
and UO_80 (O_80,N_29518,N_29721);
xnor UO_81 (O_81,N_29688,N_29839);
nor UO_82 (O_82,N_29643,N_29962);
xor UO_83 (O_83,N_29676,N_29782);
and UO_84 (O_84,N_29757,N_29525);
nand UO_85 (O_85,N_29793,N_29667);
nor UO_86 (O_86,N_29631,N_29544);
nor UO_87 (O_87,N_29677,N_29642);
xnor UO_88 (O_88,N_29538,N_29923);
xor UO_89 (O_89,N_29529,N_29868);
and UO_90 (O_90,N_29855,N_29814);
nand UO_91 (O_91,N_29939,N_29727);
nor UO_92 (O_92,N_29749,N_29800);
xnor UO_93 (O_93,N_29610,N_29553);
xnor UO_94 (O_94,N_29541,N_29713);
nor UO_95 (O_95,N_29556,N_29996);
nor UO_96 (O_96,N_29597,N_29831);
and UO_97 (O_97,N_29956,N_29948);
xnor UO_98 (O_98,N_29520,N_29516);
or UO_99 (O_99,N_29903,N_29899);
nand UO_100 (O_100,N_29781,N_29994);
nor UO_101 (O_101,N_29655,N_29955);
nor UO_102 (O_102,N_29706,N_29812);
xnor UO_103 (O_103,N_29875,N_29752);
nor UO_104 (O_104,N_29674,N_29947);
xnor UO_105 (O_105,N_29935,N_29567);
nor UO_106 (O_106,N_29763,N_29740);
and UO_107 (O_107,N_29787,N_29732);
nor UO_108 (O_108,N_29756,N_29777);
or UO_109 (O_109,N_29598,N_29792);
and UO_110 (O_110,N_29986,N_29527);
xor UO_111 (O_111,N_29967,N_29568);
or UO_112 (O_112,N_29715,N_29974);
or UO_113 (O_113,N_29864,N_29644);
or UO_114 (O_114,N_29705,N_29726);
nor UO_115 (O_115,N_29973,N_29842);
nand UO_116 (O_116,N_29646,N_29584);
xor UO_117 (O_117,N_29717,N_29650);
nand UO_118 (O_118,N_29651,N_29671);
xor UO_119 (O_119,N_29622,N_29630);
nand UO_120 (O_120,N_29745,N_29640);
or UO_121 (O_121,N_29806,N_29534);
xor UO_122 (O_122,N_29772,N_29754);
xnor UO_123 (O_123,N_29628,N_29703);
or UO_124 (O_124,N_29841,N_29609);
nand UO_125 (O_125,N_29523,N_29983);
nor UO_126 (O_126,N_29938,N_29774);
nor UO_127 (O_127,N_29748,N_29596);
xnor UO_128 (O_128,N_29942,N_29928);
nand UO_129 (O_129,N_29816,N_29764);
nand UO_130 (O_130,N_29890,N_29580);
or UO_131 (O_131,N_29656,N_29563);
or UO_132 (O_132,N_29547,N_29940);
nor UO_133 (O_133,N_29730,N_29746);
nand UO_134 (O_134,N_29809,N_29590);
xor UO_135 (O_135,N_29588,N_29835);
and UO_136 (O_136,N_29550,N_29845);
and UO_137 (O_137,N_29829,N_29592);
xnor UO_138 (O_138,N_29560,N_29858);
xnor UO_139 (O_139,N_29561,N_29530);
nand UO_140 (O_140,N_29690,N_29539);
nand UO_141 (O_141,N_29982,N_29686);
nor UO_142 (O_142,N_29618,N_29564);
and UO_143 (O_143,N_29852,N_29665);
nor UO_144 (O_144,N_29922,N_29719);
or UO_145 (O_145,N_29620,N_29766);
nor UO_146 (O_146,N_29689,N_29638);
and UO_147 (O_147,N_29504,N_29992);
nor UO_148 (O_148,N_29532,N_29968);
nand UO_149 (O_149,N_29863,N_29625);
or UO_150 (O_150,N_29921,N_29613);
nor UO_151 (O_151,N_29548,N_29760);
or UO_152 (O_152,N_29997,N_29987);
xnor UO_153 (O_153,N_29993,N_29639);
nor UO_154 (O_154,N_29820,N_29798);
or UO_155 (O_155,N_29607,N_29519);
nand UO_156 (O_156,N_29802,N_29509);
xnor UO_157 (O_157,N_29615,N_29602);
nand UO_158 (O_158,N_29843,N_29914);
nor UO_159 (O_159,N_29599,N_29891);
or UO_160 (O_160,N_29954,N_29794);
or UO_161 (O_161,N_29761,N_29795);
nand UO_162 (O_162,N_29995,N_29699);
xnor UO_163 (O_163,N_29704,N_29552);
xor UO_164 (O_164,N_29894,N_29681);
or UO_165 (O_165,N_29513,N_29870);
xnor UO_166 (O_166,N_29604,N_29701);
or UO_167 (O_167,N_29988,N_29958);
xor UO_168 (O_168,N_29543,N_29979);
xnor UO_169 (O_169,N_29789,N_29668);
or UO_170 (O_170,N_29741,N_29562);
and UO_171 (O_171,N_29893,N_29692);
nor UO_172 (O_172,N_29765,N_29907);
nor UO_173 (O_173,N_29888,N_29687);
xnor UO_174 (O_174,N_29832,N_29946);
nand UO_175 (O_175,N_29889,N_29697);
and UO_176 (O_176,N_29966,N_29769);
or UO_177 (O_177,N_29856,N_29902);
xor UO_178 (O_178,N_29531,N_29514);
nor UO_179 (O_179,N_29700,N_29587);
nand UO_180 (O_180,N_29883,N_29522);
xor UO_181 (O_181,N_29679,N_29911);
nand UO_182 (O_182,N_29554,N_29933);
or UO_183 (O_183,N_29848,N_29528);
nor UO_184 (O_184,N_29904,N_29775);
or UO_185 (O_185,N_29658,N_29664);
nor UO_186 (O_186,N_29998,N_29603);
nor UO_187 (O_187,N_29913,N_29612);
xnor UO_188 (O_188,N_29537,N_29768);
nand UO_189 (O_189,N_29978,N_29657);
nand UO_190 (O_190,N_29582,N_29758);
xnor UO_191 (O_191,N_29885,N_29535);
nand UO_192 (O_192,N_29972,N_29574);
xor UO_193 (O_193,N_29850,N_29515);
xnor UO_194 (O_194,N_29645,N_29608);
xnor UO_195 (O_195,N_29743,N_29817);
xnor UO_196 (O_196,N_29573,N_29896);
or UO_197 (O_197,N_29815,N_29511);
xnor UO_198 (O_198,N_29934,N_29551);
or UO_199 (O_199,N_29611,N_29866);
xnor UO_200 (O_200,N_29950,N_29755);
nor UO_201 (O_201,N_29505,N_29804);
and UO_202 (O_202,N_29862,N_29985);
xnor UO_203 (O_203,N_29980,N_29854);
nor UO_204 (O_204,N_29881,N_29937);
or UO_205 (O_205,N_29874,N_29825);
nand UO_206 (O_206,N_29594,N_29545);
xnor UO_207 (O_207,N_29707,N_29747);
nand UO_208 (O_208,N_29542,N_29669);
nor UO_209 (O_209,N_29557,N_29857);
and UO_210 (O_210,N_29570,N_29900);
xnor UO_211 (O_211,N_29869,N_29678);
xnor UO_212 (O_212,N_29663,N_29971);
or UO_213 (O_213,N_29585,N_29915);
nand UO_214 (O_214,N_29648,N_29943);
nor UO_215 (O_215,N_29880,N_29836);
nand UO_216 (O_216,N_29819,N_29508);
nand UO_217 (O_217,N_29714,N_29524);
or UO_218 (O_218,N_29977,N_29799);
xor UO_219 (O_219,N_29759,N_29879);
or UO_220 (O_220,N_29636,N_29744);
nand UO_221 (O_221,N_29549,N_29736);
nand UO_222 (O_222,N_29566,N_29944);
and UO_223 (O_223,N_29887,N_29970);
nor UO_224 (O_224,N_29953,N_29905);
nor UO_225 (O_225,N_29708,N_29898);
xor UO_226 (O_226,N_29813,N_29600);
and UO_227 (O_227,N_29897,N_29565);
or UO_228 (O_228,N_29682,N_29533);
xor UO_229 (O_229,N_29861,N_29753);
nor UO_230 (O_230,N_29558,N_29910);
xor UO_231 (O_231,N_29949,N_29540);
and UO_232 (O_232,N_29969,N_29577);
nor UO_233 (O_233,N_29500,N_29965);
nand UO_234 (O_234,N_29847,N_29976);
or UO_235 (O_235,N_29963,N_29981);
or UO_236 (O_236,N_29916,N_29659);
nor UO_237 (O_237,N_29693,N_29725);
nor UO_238 (O_238,N_29926,N_29694);
nor UO_239 (O_239,N_29742,N_29621);
nand UO_240 (O_240,N_29720,N_29591);
or UO_241 (O_241,N_29908,N_29951);
nand UO_242 (O_242,N_29734,N_29517);
nor UO_243 (O_243,N_29660,N_29920);
nand UO_244 (O_244,N_29601,N_29691);
or UO_245 (O_245,N_29918,N_29503);
or UO_246 (O_246,N_29849,N_29872);
nor UO_247 (O_247,N_29876,N_29810);
xnor UO_248 (O_248,N_29666,N_29828);
or UO_249 (O_249,N_29961,N_29960);
xnor UO_250 (O_250,N_29823,N_29676);
xor UO_251 (O_251,N_29706,N_29589);
nor UO_252 (O_252,N_29857,N_29623);
and UO_253 (O_253,N_29695,N_29771);
nand UO_254 (O_254,N_29892,N_29855);
xor UO_255 (O_255,N_29732,N_29580);
and UO_256 (O_256,N_29565,N_29834);
or UO_257 (O_257,N_29805,N_29580);
nand UO_258 (O_258,N_29698,N_29666);
nand UO_259 (O_259,N_29865,N_29947);
or UO_260 (O_260,N_29679,N_29940);
xor UO_261 (O_261,N_29534,N_29678);
nor UO_262 (O_262,N_29990,N_29546);
nor UO_263 (O_263,N_29618,N_29552);
nand UO_264 (O_264,N_29717,N_29584);
or UO_265 (O_265,N_29540,N_29803);
or UO_266 (O_266,N_29592,N_29611);
nor UO_267 (O_267,N_29794,N_29873);
nor UO_268 (O_268,N_29849,N_29676);
xor UO_269 (O_269,N_29853,N_29568);
xnor UO_270 (O_270,N_29857,N_29794);
and UO_271 (O_271,N_29619,N_29654);
nand UO_272 (O_272,N_29883,N_29918);
and UO_273 (O_273,N_29696,N_29674);
nor UO_274 (O_274,N_29805,N_29786);
nor UO_275 (O_275,N_29890,N_29899);
nor UO_276 (O_276,N_29828,N_29870);
xor UO_277 (O_277,N_29522,N_29808);
xnor UO_278 (O_278,N_29745,N_29502);
nand UO_279 (O_279,N_29550,N_29831);
xnor UO_280 (O_280,N_29977,N_29830);
xor UO_281 (O_281,N_29956,N_29826);
and UO_282 (O_282,N_29895,N_29501);
xnor UO_283 (O_283,N_29858,N_29585);
xor UO_284 (O_284,N_29749,N_29984);
nor UO_285 (O_285,N_29754,N_29673);
xor UO_286 (O_286,N_29690,N_29815);
or UO_287 (O_287,N_29756,N_29911);
nor UO_288 (O_288,N_29616,N_29932);
or UO_289 (O_289,N_29544,N_29578);
and UO_290 (O_290,N_29961,N_29853);
and UO_291 (O_291,N_29830,N_29711);
or UO_292 (O_292,N_29799,N_29944);
or UO_293 (O_293,N_29949,N_29738);
nor UO_294 (O_294,N_29569,N_29964);
and UO_295 (O_295,N_29895,N_29635);
nand UO_296 (O_296,N_29750,N_29558);
nor UO_297 (O_297,N_29744,N_29515);
nand UO_298 (O_298,N_29684,N_29958);
xnor UO_299 (O_299,N_29980,N_29697);
xor UO_300 (O_300,N_29536,N_29835);
nor UO_301 (O_301,N_29883,N_29582);
nand UO_302 (O_302,N_29541,N_29573);
or UO_303 (O_303,N_29779,N_29684);
nor UO_304 (O_304,N_29521,N_29945);
nand UO_305 (O_305,N_29614,N_29938);
nor UO_306 (O_306,N_29670,N_29721);
xnor UO_307 (O_307,N_29931,N_29797);
or UO_308 (O_308,N_29770,N_29633);
and UO_309 (O_309,N_29538,N_29503);
xor UO_310 (O_310,N_29639,N_29749);
or UO_311 (O_311,N_29652,N_29710);
xnor UO_312 (O_312,N_29964,N_29552);
nor UO_313 (O_313,N_29723,N_29826);
nand UO_314 (O_314,N_29734,N_29870);
nand UO_315 (O_315,N_29671,N_29554);
or UO_316 (O_316,N_29721,N_29549);
nor UO_317 (O_317,N_29807,N_29972);
xor UO_318 (O_318,N_29725,N_29846);
and UO_319 (O_319,N_29520,N_29851);
nand UO_320 (O_320,N_29898,N_29884);
and UO_321 (O_321,N_29821,N_29786);
and UO_322 (O_322,N_29509,N_29667);
xor UO_323 (O_323,N_29929,N_29917);
or UO_324 (O_324,N_29640,N_29948);
xnor UO_325 (O_325,N_29527,N_29773);
nor UO_326 (O_326,N_29675,N_29607);
or UO_327 (O_327,N_29861,N_29549);
nor UO_328 (O_328,N_29816,N_29790);
nor UO_329 (O_329,N_29780,N_29622);
nor UO_330 (O_330,N_29800,N_29601);
and UO_331 (O_331,N_29793,N_29896);
xor UO_332 (O_332,N_29691,N_29686);
nand UO_333 (O_333,N_29838,N_29677);
or UO_334 (O_334,N_29805,N_29549);
xnor UO_335 (O_335,N_29678,N_29913);
xor UO_336 (O_336,N_29653,N_29921);
nand UO_337 (O_337,N_29957,N_29509);
xnor UO_338 (O_338,N_29502,N_29835);
or UO_339 (O_339,N_29585,N_29651);
nor UO_340 (O_340,N_29690,N_29610);
nor UO_341 (O_341,N_29863,N_29758);
nor UO_342 (O_342,N_29964,N_29846);
or UO_343 (O_343,N_29589,N_29935);
nand UO_344 (O_344,N_29585,N_29685);
and UO_345 (O_345,N_29819,N_29763);
or UO_346 (O_346,N_29725,N_29700);
nor UO_347 (O_347,N_29958,N_29903);
nor UO_348 (O_348,N_29629,N_29624);
xor UO_349 (O_349,N_29506,N_29537);
and UO_350 (O_350,N_29899,N_29615);
nor UO_351 (O_351,N_29637,N_29689);
and UO_352 (O_352,N_29957,N_29802);
nand UO_353 (O_353,N_29758,N_29759);
nand UO_354 (O_354,N_29894,N_29668);
or UO_355 (O_355,N_29694,N_29709);
xor UO_356 (O_356,N_29859,N_29766);
nand UO_357 (O_357,N_29733,N_29587);
nand UO_358 (O_358,N_29629,N_29758);
and UO_359 (O_359,N_29620,N_29517);
nand UO_360 (O_360,N_29736,N_29669);
nor UO_361 (O_361,N_29739,N_29789);
or UO_362 (O_362,N_29762,N_29924);
nor UO_363 (O_363,N_29983,N_29551);
nor UO_364 (O_364,N_29889,N_29931);
nand UO_365 (O_365,N_29623,N_29797);
or UO_366 (O_366,N_29907,N_29875);
xnor UO_367 (O_367,N_29671,N_29690);
nand UO_368 (O_368,N_29634,N_29684);
nor UO_369 (O_369,N_29504,N_29559);
nand UO_370 (O_370,N_29778,N_29884);
and UO_371 (O_371,N_29984,N_29529);
nor UO_372 (O_372,N_29944,N_29589);
xor UO_373 (O_373,N_29671,N_29739);
and UO_374 (O_374,N_29965,N_29539);
xor UO_375 (O_375,N_29993,N_29937);
nand UO_376 (O_376,N_29633,N_29956);
and UO_377 (O_377,N_29545,N_29956);
or UO_378 (O_378,N_29789,N_29817);
nor UO_379 (O_379,N_29996,N_29899);
nor UO_380 (O_380,N_29611,N_29610);
xor UO_381 (O_381,N_29669,N_29845);
and UO_382 (O_382,N_29660,N_29903);
nand UO_383 (O_383,N_29870,N_29671);
and UO_384 (O_384,N_29947,N_29573);
xnor UO_385 (O_385,N_29861,N_29777);
xor UO_386 (O_386,N_29727,N_29794);
nand UO_387 (O_387,N_29557,N_29839);
nand UO_388 (O_388,N_29998,N_29803);
or UO_389 (O_389,N_29537,N_29790);
nand UO_390 (O_390,N_29889,N_29686);
nor UO_391 (O_391,N_29936,N_29964);
and UO_392 (O_392,N_29510,N_29981);
nand UO_393 (O_393,N_29592,N_29848);
xnor UO_394 (O_394,N_29880,N_29778);
and UO_395 (O_395,N_29569,N_29813);
nor UO_396 (O_396,N_29647,N_29624);
or UO_397 (O_397,N_29860,N_29672);
xor UO_398 (O_398,N_29827,N_29769);
and UO_399 (O_399,N_29737,N_29987);
or UO_400 (O_400,N_29849,N_29522);
or UO_401 (O_401,N_29505,N_29585);
or UO_402 (O_402,N_29999,N_29992);
and UO_403 (O_403,N_29831,N_29626);
or UO_404 (O_404,N_29505,N_29930);
nand UO_405 (O_405,N_29769,N_29778);
nor UO_406 (O_406,N_29715,N_29643);
and UO_407 (O_407,N_29740,N_29538);
nor UO_408 (O_408,N_29932,N_29594);
nor UO_409 (O_409,N_29939,N_29721);
nor UO_410 (O_410,N_29695,N_29934);
and UO_411 (O_411,N_29884,N_29821);
nand UO_412 (O_412,N_29634,N_29999);
and UO_413 (O_413,N_29949,N_29862);
and UO_414 (O_414,N_29677,N_29656);
nand UO_415 (O_415,N_29811,N_29622);
xnor UO_416 (O_416,N_29748,N_29859);
xnor UO_417 (O_417,N_29507,N_29741);
nand UO_418 (O_418,N_29807,N_29939);
nor UO_419 (O_419,N_29593,N_29954);
nand UO_420 (O_420,N_29942,N_29986);
nand UO_421 (O_421,N_29668,N_29976);
nor UO_422 (O_422,N_29590,N_29540);
xnor UO_423 (O_423,N_29508,N_29595);
and UO_424 (O_424,N_29835,N_29811);
nand UO_425 (O_425,N_29548,N_29940);
nor UO_426 (O_426,N_29512,N_29817);
nand UO_427 (O_427,N_29969,N_29749);
nand UO_428 (O_428,N_29614,N_29993);
and UO_429 (O_429,N_29777,N_29746);
xnor UO_430 (O_430,N_29512,N_29624);
and UO_431 (O_431,N_29738,N_29652);
nand UO_432 (O_432,N_29914,N_29832);
and UO_433 (O_433,N_29572,N_29691);
or UO_434 (O_434,N_29766,N_29623);
nor UO_435 (O_435,N_29690,N_29850);
and UO_436 (O_436,N_29923,N_29578);
or UO_437 (O_437,N_29621,N_29773);
or UO_438 (O_438,N_29796,N_29709);
nand UO_439 (O_439,N_29907,N_29567);
nand UO_440 (O_440,N_29888,N_29732);
nand UO_441 (O_441,N_29919,N_29769);
and UO_442 (O_442,N_29670,N_29682);
or UO_443 (O_443,N_29834,N_29665);
nand UO_444 (O_444,N_29865,N_29826);
xor UO_445 (O_445,N_29855,N_29524);
nand UO_446 (O_446,N_29970,N_29873);
and UO_447 (O_447,N_29506,N_29894);
xnor UO_448 (O_448,N_29972,N_29718);
nand UO_449 (O_449,N_29963,N_29959);
or UO_450 (O_450,N_29883,N_29539);
xnor UO_451 (O_451,N_29521,N_29807);
or UO_452 (O_452,N_29524,N_29856);
nand UO_453 (O_453,N_29690,N_29523);
nor UO_454 (O_454,N_29722,N_29888);
nand UO_455 (O_455,N_29678,N_29543);
xor UO_456 (O_456,N_29879,N_29770);
or UO_457 (O_457,N_29687,N_29816);
nor UO_458 (O_458,N_29887,N_29739);
nand UO_459 (O_459,N_29536,N_29837);
nand UO_460 (O_460,N_29595,N_29913);
xnor UO_461 (O_461,N_29788,N_29712);
nand UO_462 (O_462,N_29846,N_29579);
xor UO_463 (O_463,N_29702,N_29549);
or UO_464 (O_464,N_29752,N_29822);
nand UO_465 (O_465,N_29786,N_29830);
and UO_466 (O_466,N_29639,N_29675);
nand UO_467 (O_467,N_29605,N_29918);
xnor UO_468 (O_468,N_29590,N_29971);
xnor UO_469 (O_469,N_29875,N_29570);
nor UO_470 (O_470,N_29772,N_29725);
nand UO_471 (O_471,N_29532,N_29805);
xnor UO_472 (O_472,N_29820,N_29583);
or UO_473 (O_473,N_29588,N_29599);
and UO_474 (O_474,N_29937,N_29818);
or UO_475 (O_475,N_29790,N_29854);
xor UO_476 (O_476,N_29873,N_29938);
xor UO_477 (O_477,N_29690,N_29691);
or UO_478 (O_478,N_29594,N_29884);
or UO_479 (O_479,N_29791,N_29942);
or UO_480 (O_480,N_29732,N_29716);
or UO_481 (O_481,N_29645,N_29577);
xnor UO_482 (O_482,N_29606,N_29841);
xor UO_483 (O_483,N_29716,N_29779);
or UO_484 (O_484,N_29722,N_29977);
nor UO_485 (O_485,N_29701,N_29579);
xor UO_486 (O_486,N_29712,N_29738);
or UO_487 (O_487,N_29508,N_29533);
or UO_488 (O_488,N_29812,N_29592);
nor UO_489 (O_489,N_29536,N_29515);
and UO_490 (O_490,N_29724,N_29843);
nand UO_491 (O_491,N_29640,N_29998);
or UO_492 (O_492,N_29975,N_29855);
nor UO_493 (O_493,N_29982,N_29902);
nand UO_494 (O_494,N_29719,N_29723);
nand UO_495 (O_495,N_29750,N_29610);
or UO_496 (O_496,N_29549,N_29525);
and UO_497 (O_497,N_29703,N_29849);
nand UO_498 (O_498,N_29819,N_29850);
and UO_499 (O_499,N_29878,N_29514);
xnor UO_500 (O_500,N_29699,N_29629);
xnor UO_501 (O_501,N_29800,N_29628);
nor UO_502 (O_502,N_29556,N_29642);
and UO_503 (O_503,N_29705,N_29681);
nor UO_504 (O_504,N_29835,N_29523);
xnor UO_505 (O_505,N_29998,N_29601);
nor UO_506 (O_506,N_29546,N_29769);
or UO_507 (O_507,N_29505,N_29793);
and UO_508 (O_508,N_29970,N_29852);
nand UO_509 (O_509,N_29699,N_29914);
nor UO_510 (O_510,N_29779,N_29683);
xnor UO_511 (O_511,N_29839,N_29931);
nor UO_512 (O_512,N_29721,N_29531);
or UO_513 (O_513,N_29953,N_29903);
nand UO_514 (O_514,N_29992,N_29547);
or UO_515 (O_515,N_29911,N_29814);
and UO_516 (O_516,N_29725,N_29902);
nand UO_517 (O_517,N_29969,N_29951);
nand UO_518 (O_518,N_29509,N_29674);
xor UO_519 (O_519,N_29757,N_29822);
or UO_520 (O_520,N_29912,N_29799);
nor UO_521 (O_521,N_29519,N_29989);
or UO_522 (O_522,N_29702,N_29914);
nor UO_523 (O_523,N_29642,N_29903);
nand UO_524 (O_524,N_29682,N_29901);
or UO_525 (O_525,N_29830,N_29594);
xor UO_526 (O_526,N_29849,N_29679);
nor UO_527 (O_527,N_29889,N_29681);
nand UO_528 (O_528,N_29545,N_29765);
xor UO_529 (O_529,N_29926,N_29891);
xor UO_530 (O_530,N_29879,N_29563);
and UO_531 (O_531,N_29726,N_29622);
nor UO_532 (O_532,N_29522,N_29788);
xor UO_533 (O_533,N_29763,N_29606);
or UO_534 (O_534,N_29949,N_29821);
nor UO_535 (O_535,N_29653,N_29523);
nor UO_536 (O_536,N_29760,N_29951);
xor UO_537 (O_537,N_29880,N_29916);
and UO_538 (O_538,N_29829,N_29767);
and UO_539 (O_539,N_29766,N_29511);
nor UO_540 (O_540,N_29694,N_29957);
and UO_541 (O_541,N_29738,N_29934);
or UO_542 (O_542,N_29931,N_29752);
nand UO_543 (O_543,N_29799,N_29928);
xnor UO_544 (O_544,N_29757,N_29714);
xnor UO_545 (O_545,N_29501,N_29526);
nor UO_546 (O_546,N_29619,N_29574);
nor UO_547 (O_547,N_29855,N_29616);
nand UO_548 (O_548,N_29632,N_29526);
nand UO_549 (O_549,N_29798,N_29695);
nor UO_550 (O_550,N_29920,N_29738);
or UO_551 (O_551,N_29777,N_29796);
or UO_552 (O_552,N_29820,N_29793);
nor UO_553 (O_553,N_29536,N_29836);
nor UO_554 (O_554,N_29837,N_29741);
nand UO_555 (O_555,N_29862,N_29680);
and UO_556 (O_556,N_29698,N_29884);
xor UO_557 (O_557,N_29795,N_29703);
or UO_558 (O_558,N_29968,N_29530);
nor UO_559 (O_559,N_29690,N_29806);
nand UO_560 (O_560,N_29736,N_29514);
nor UO_561 (O_561,N_29574,N_29586);
and UO_562 (O_562,N_29602,N_29612);
and UO_563 (O_563,N_29956,N_29728);
nor UO_564 (O_564,N_29908,N_29608);
xor UO_565 (O_565,N_29606,N_29762);
xor UO_566 (O_566,N_29509,N_29940);
nor UO_567 (O_567,N_29816,N_29838);
nor UO_568 (O_568,N_29542,N_29689);
or UO_569 (O_569,N_29661,N_29538);
nor UO_570 (O_570,N_29545,N_29708);
xor UO_571 (O_571,N_29953,N_29756);
nor UO_572 (O_572,N_29950,N_29737);
and UO_573 (O_573,N_29873,N_29811);
xor UO_574 (O_574,N_29803,N_29579);
nor UO_575 (O_575,N_29577,N_29732);
nand UO_576 (O_576,N_29549,N_29959);
or UO_577 (O_577,N_29987,N_29671);
nor UO_578 (O_578,N_29890,N_29772);
nor UO_579 (O_579,N_29607,N_29595);
or UO_580 (O_580,N_29839,N_29866);
or UO_581 (O_581,N_29617,N_29989);
and UO_582 (O_582,N_29924,N_29696);
nand UO_583 (O_583,N_29869,N_29727);
nor UO_584 (O_584,N_29544,N_29528);
nor UO_585 (O_585,N_29883,N_29923);
nand UO_586 (O_586,N_29592,N_29513);
and UO_587 (O_587,N_29972,N_29633);
xnor UO_588 (O_588,N_29801,N_29988);
nor UO_589 (O_589,N_29836,N_29819);
xnor UO_590 (O_590,N_29951,N_29692);
and UO_591 (O_591,N_29614,N_29894);
or UO_592 (O_592,N_29883,N_29773);
xnor UO_593 (O_593,N_29579,N_29575);
or UO_594 (O_594,N_29736,N_29656);
nor UO_595 (O_595,N_29704,N_29985);
and UO_596 (O_596,N_29876,N_29806);
nand UO_597 (O_597,N_29762,N_29568);
xnor UO_598 (O_598,N_29846,N_29734);
xnor UO_599 (O_599,N_29987,N_29609);
nor UO_600 (O_600,N_29881,N_29674);
or UO_601 (O_601,N_29994,N_29503);
xnor UO_602 (O_602,N_29844,N_29855);
and UO_603 (O_603,N_29650,N_29728);
nor UO_604 (O_604,N_29525,N_29697);
nand UO_605 (O_605,N_29986,N_29950);
xor UO_606 (O_606,N_29698,N_29785);
nor UO_607 (O_607,N_29920,N_29541);
nor UO_608 (O_608,N_29536,N_29949);
nand UO_609 (O_609,N_29703,N_29941);
nand UO_610 (O_610,N_29688,N_29700);
and UO_611 (O_611,N_29699,N_29916);
nand UO_612 (O_612,N_29894,N_29884);
or UO_613 (O_613,N_29798,N_29572);
nor UO_614 (O_614,N_29897,N_29806);
xnor UO_615 (O_615,N_29753,N_29806);
nand UO_616 (O_616,N_29816,N_29908);
or UO_617 (O_617,N_29876,N_29828);
and UO_618 (O_618,N_29555,N_29857);
or UO_619 (O_619,N_29766,N_29700);
nand UO_620 (O_620,N_29665,N_29980);
nor UO_621 (O_621,N_29706,N_29922);
xor UO_622 (O_622,N_29692,N_29571);
nand UO_623 (O_623,N_29643,N_29798);
nand UO_624 (O_624,N_29678,N_29879);
nor UO_625 (O_625,N_29858,N_29562);
xor UO_626 (O_626,N_29914,N_29776);
xnor UO_627 (O_627,N_29563,N_29751);
or UO_628 (O_628,N_29503,N_29936);
nor UO_629 (O_629,N_29522,N_29546);
nor UO_630 (O_630,N_29782,N_29789);
and UO_631 (O_631,N_29746,N_29818);
and UO_632 (O_632,N_29569,N_29960);
nor UO_633 (O_633,N_29850,N_29870);
and UO_634 (O_634,N_29872,N_29966);
and UO_635 (O_635,N_29808,N_29851);
and UO_636 (O_636,N_29840,N_29735);
or UO_637 (O_637,N_29578,N_29807);
nor UO_638 (O_638,N_29981,N_29655);
and UO_639 (O_639,N_29875,N_29586);
or UO_640 (O_640,N_29605,N_29644);
nor UO_641 (O_641,N_29793,N_29964);
xnor UO_642 (O_642,N_29525,N_29684);
nand UO_643 (O_643,N_29926,N_29602);
nand UO_644 (O_644,N_29727,N_29825);
nor UO_645 (O_645,N_29850,N_29987);
and UO_646 (O_646,N_29627,N_29554);
nor UO_647 (O_647,N_29978,N_29970);
nor UO_648 (O_648,N_29650,N_29878);
nand UO_649 (O_649,N_29832,N_29789);
xor UO_650 (O_650,N_29796,N_29693);
nand UO_651 (O_651,N_29621,N_29800);
nand UO_652 (O_652,N_29604,N_29664);
xor UO_653 (O_653,N_29953,N_29860);
xor UO_654 (O_654,N_29954,N_29576);
nor UO_655 (O_655,N_29659,N_29867);
xor UO_656 (O_656,N_29920,N_29649);
or UO_657 (O_657,N_29916,N_29858);
xor UO_658 (O_658,N_29876,N_29696);
nor UO_659 (O_659,N_29517,N_29880);
nand UO_660 (O_660,N_29913,N_29625);
xor UO_661 (O_661,N_29505,N_29964);
nand UO_662 (O_662,N_29729,N_29771);
nor UO_663 (O_663,N_29886,N_29502);
xor UO_664 (O_664,N_29982,N_29688);
nand UO_665 (O_665,N_29799,N_29573);
nand UO_666 (O_666,N_29557,N_29884);
nor UO_667 (O_667,N_29986,N_29620);
or UO_668 (O_668,N_29791,N_29716);
xnor UO_669 (O_669,N_29725,N_29949);
or UO_670 (O_670,N_29847,N_29740);
and UO_671 (O_671,N_29841,N_29842);
or UO_672 (O_672,N_29916,N_29751);
xnor UO_673 (O_673,N_29686,N_29822);
nand UO_674 (O_674,N_29873,N_29759);
and UO_675 (O_675,N_29812,N_29983);
and UO_676 (O_676,N_29831,N_29873);
xor UO_677 (O_677,N_29941,N_29877);
nor UO_678 (O_678,N_29708,N_29670);
and UO_679 (O_679,N_29554,N_29630);
or UO_680 (O_680,N_29823,N_29960);
nand UO_681 (O_681,N_29988,N_29841);
and UO_682 (O_682,N_29698,N_29592);
nor UO_683 (O_683,N_29590,N_29747);
or UO_684 (O_684,N_29511,N_29823);
and UO_685 (O_685,N_29625,N_29601);
or UO_686 (O_686,N_29566,N_29993);
nand UO_687 (O_687,N_29693,N_29985);
and UO_688 (O_688,N_29641,N_29723);
nand UO_689 (O_689,N_29753,N_29759);
xor UO_690 (O_690,N_29940,N_29999);
or UO_691 (O_691,N_29820,N_29738);
nand UO_692 (O_692,N_29551,N_29813);
nor UO_693 (O_693,N_29865,N_29836);
or UO_694 (O_694,N_29648,N_29998);
xor UO_695 (O_695,N_29992,N_29822);
and UO_696 (O_696,N_29926,N_29608);
xnor UO_697 (O_697,N_29681,N_29547);
and UO_698 (O_698,N_29954,N_29960);
nand UO_699 (O_699,N_29852,N_29684);
and UO_700 (O_700,N_29931,N_29965);
nand UO_701 (O_701,N_29991,N_29749);
nor UO_702 (O_702,N_29850,N_29895);
nand UO_703 (O_703,N_29505,N_29661);
and UO_704 (O_704,N_29800,N_29508);
nor UO_705 (O_705,N_29828,N_29604);
and UO_706 (O_706,N_29546,N_29642);
or UO_707 (O_707,N_29950,N_29744);
nor UO_708 (O_708,N_29722,N_29925);
and UO_709 (O_709,N_29514,N_29894);
xnor UO_710 (O_710,N_29916,N_29847);
or UO_711 (O_711,N_29600,N_29765);
nand UO_712 (O_712,N_29638,N_29865);
or UO_713 (O_713,N_29903,N_29921);
xor UO_714 (O_714,N_29632,N_29738);
and UO_715 (O_715,N_29784,N_29650);
nor UO_716 (O_716,N_29683,N_29733);
or UO_717 (O_717,N_29666,N_29944);
nor UO_718 (O_718,N_29619,N_29585);
or UO_719 (O_719,N_29678,N_29774);
nor UO_720 (O_720,N_29515,N_29942);
or UO_721 (O_721,N_29732,N_29749);
or UO_722 (O_722,N_29672,N_29617);
and UO_723 (O_723,N_29799,N_29623);
nand UO_724 (O_724,N_29913,N_29902);
nor UO_725 (O_725,N_29731,N_29898);
or UO_726 (O_726,N_29664,N_29921);
or UO_727 (O_727,N_29543,N_29916);
or UO_728 (O_728,N_29789,N_29988);
xor UO_729 (O_729,N_29913,N_29677);
or UO_730 (O_730,N_29964,N_29717);
or UO_731 (O_731,N_29936,N_29654);
nand UO_732 (O_732,N_29961,N_29539);
or UO_733 (O_733,N_29829,N_29921);
xnor UO_734 (O_734,N_29962,N_29794);
and UO_735 (O_735,N_29697,N_29822);
xnor UO_736 (O_736,N_29766,N_29817);
nand UO_737 (O_737,N_29862,N_29633);
xnor UO_738 (O_738,N_29648,N_29883);
or UO_739 (O_739,N_29805,N_29693);
or UO_740 (O_740,N_29962,N_29546);
xnor UO_741 (O_741,N_29789,N_29737);
xnor UO_742 (O_742,N_29681,N_29508);
nor UO_743 (O_743,N_29689,N_29727);
or UO_744 (O_744,N_29716,N_29594);
nor UO_745 (O_745,N_29687,N_29910);
nor UO_746 (O_746,N_29545,N_29650);
nand UO_747 (O_747,N_29694,N_29749);
and UO_748 (O_748,N_29944,N_29560);
or UO_749 (O_749,N_29976,N_29882);
or UO_750 (O_750,N_29997,N_29535);
nor UO_751 (O_751,N_29790,N_29754);
or UO_752 (O_752,N_29531,N_29708);
nand UO_753 (O_753,N_29800,N_29774);
nand UO_754 (O_754,N_29762,N_29566);
and UO_755 (O_755,N_29855,N_29700);
nor UO_756 (O_756,N_29934,N_29769);
and UO_757 (O_757,N_29565,N_29695);
nor UO_758 (O_758,N_29953,N_29508);
and UO_759 (O_759,N_29905,N_29691);
nand UO_760 (O_760,N_29842,N_29591);
nand UO_761 (O_761,N_29588,N_29773);
xnor UO_762 (O_762,N_29805,N_29883);
nand UO_763 (O_763,N_29590,N_29837);
or UO_764 (O_764,N_29983,N_29521);
xor UO_765 (O_765,N_29895,N_29707);
or UO_766 (O_766,N_29982,N_29907);
xor UO_767 (O_767,N_29598,N_29642);
or UO_768 (O_768,N_29644,N_29501);
and UO_769 (O_769,N_29637,N_29782);
or UO_770 (O_770,N_29889,N_29607);
or UO_771 (O_771,N_29547,N_29854);
nand UO_772 (O_772,N_29519,N_29880);
or UO_773 (O_773,N_29856,N_29935);
nor UO_774 (O_774,N_29784,N_29897);
nor UO_775 (O_775,N_29831,N_29536);
xor UO_776 (O_776,N_29730,N_29573);
or UO_777 (O_777,N_29885,N_29634);
and UO_778 (O_778,N_29924,N_29869);
nor UO_779 (O_779,N_29550,N_29681);
and UO_780 (O_780,N_29875,N_29727);
xnor UO_781 (O_781,N_29891,N_29909);
nand UO_782 (O_782,N_29624,N_29539);
nor UO_783 (O_783,N_29628,N_29742);
and UO_784 (O_784,N_29581,N_29867);
nor UO_785 (O_785,N_29559,N_29985);
xor UO_786 (O_786,N_29509,N_29859);
nand UO_787 (O_787,N_29565,N_29638);
nor UO_788 (O_788,N_29569,N_29752);
xor UO_789 (O_789,N_29552,N_29537);
nor UO_790 (O_790,N_29734,N_29947);
nand UO_791 (O_791,N_29940,N_29541);
nand UO_792 (O_792,N_29625,N_29652);
nand UO_793 (O_793,N_29933,N_29623);
nand UO_794 (O_794,N_29962,N_29721);
or UO_795 (O_795,N_29989,N_29901);
xnor UO_796 (O_796,N_29943,N_29703);
nor UO_797 (O_797,N_29806,N_29975);
and UO_798 (O_798,N_29724,N_29938);
xor UO_799 (O_799,N_29549,N_29941);
or UO_800 (O_800,N_29554,N_29535);
nand UO_801 (O_801,N_29988,N_29600);
nand UO_802 (O_802,N_29574,N_29550);
nor UO_803 (O_803,N_29716,N_29505);
nand UO_804 (O_804,N_29534,N_29923);
xor UO_805 (O_805,N_29516,N_29652);
nand UO_806 (O_806,N_29891,N_29617);
and UO_807 (O_807,N_29707,N_29740);
nor UO_808 (O_808,N_29554,N_29812);
and UO_809 (O_809,N_29882,N_29710);
and UO_810 (O_810,N_29725,N_29962);
nand UO_811 (O_811,N_29750,N_29759);
nand UO_812 (O_812,N_29859,N_29652);
and UO_813 (O_813,N_29591,N_29683);
nand UO_814 (O_814,N_29856,N_29580);
or UO_815 (O_815,N_29533,N_29575);
and UO_816 (O_816,N_29742,N_29537);
nand UO_817 (O_817,N_29587,N_29654);
xnor UO_818 (O_818,N_29777,N_29820);
xnor UO_819 (O_819,N_29629,N_29800);
nor UO_820 (O_820,N_29840,N_29687);
xor UO_821 (O_821,N_29504,N_29783);
nand UO_822 (O_822,N_29604,N_29698);
nand UO_823 (O_823,N_29918,N_29687);
or UO_824 (O_824,N_29854,N_29990);
nor UO_825 (O_825,N_29531,N_29625);
nand UO_826 (O_826,N_29643,N_29629);
nand UO_827 (O_827,N_29953,N_29598);
and UO_828 (O_828,N_29583,N_29624);
nor UO_829 (O_829,N_29544,N_29681);
xor UO_830 (O_830,N_29663,N_29968);
and UO_831 (O_831,N_29694,N_29941);
nand UO_832 (O_832,N_29525,N_29554);
and UO_833 (O_833,N_29786,N_29916);
or UO_834 (O_834,N_29871,N_29928);
nand UO_835 (O_835,N_29703,N_29887);
nand UO_836 (O_836,N_29691,N_29854);
nor UO_837 (O_837,N_29880,N_29769);
nand UO_838 (O_838,N_29993,N_29597);
or UO_839 (O_839,N_29735,N_29743);
or UO_840 (O_840,N_29770,N_29671);
xnor UO_841 (O_841,N_29624,N_29952);
nand UO_842 (O_842,N_29621,N_29971);
nand UO_843 (O_843,N_29542,N_29798);
or UO_844 (O_844,N_29955,N_29859);
xnor UO_845 (O_845,N_29900,N_29768);
nor UO_846 (O_846,N_29508,N_29752);
nand UO_847 (O_847,N_29830,N_29552);
nand UO_848 (O_848,N_29758,N_29938);
and UO_849 (O_849,N_29857,N_29655);
xor UO_850 (O_850,N_29599,N_29786);
xnor UO_851 (O_851,N_29992,N_29570);
nand UO_852 (O_852,N_29913,N_29690);
xnor UO_853 (O_853,N_29564,N_29663);
nand UO_854 (O_854,N_29590,N_29784);
and UO_855 (O_855,N_29941,N_29922);
nand UO_856 (O_856,N_29538,N_29771);
xor UO_857 (O_857,N_29707,N_29596);
xor UO_858 (O_858,N_29901,N_29515);
and UO_859 (O_859,N_29624,N_29701);
and UO_860 (O_860,N_29993,N_29853);
nand UO_861 (O_861,N_29884,N_29677);
and UO_862 (O_862,N_29723,N_29556);
xnor UO_863 (O_863,N_29640,N_29776);
or UO_864 (O_864,N_29685,N_29837);
and UO_865 (O_865,N_29595,N_29669);
or UO_866 (O_866,N_29612,N_29855);
and UO_867 (O_867,N_29746,N_29656);
nor UO_868 (O_868,N_29706,N_29791);
nand UO_869 (O_869,N_29883,N_29725);
nor UO_870 (O_870,N_29639,N_29641);
xor UO_871 (O_871,N_29952,N_29770);
and UO_872 (O_872,N_29935,N_29564);
nand UO_873 (O_873,N_29649,N_29582);
nor UO_874 (O_874,N_29800,N_29863);
xnor UO_875 (O_875,N_29716,N_29842);
and UO_876 (O_876,N_29639,N_29510);
and UO_877 (O_877,N_29866,N_29648);
and UO_878 (O_878,N_29611,N_29756);
or UO_879 (O_879,N_29654,N_29608);
nor UO_880 (O_880,N_29600,N_29803);
or UO_881 (O_881,N_29826,N_29958);
and UO_882 (O_882,N_29946,N_29680);
and UO_883 (O_883,N_29848,N_29644);
nand UO_884 (O_884,N_29645,N_29965);
and UO_885 (O_885,N_29921,N_29940);
xor UO_886 (O_886,N_29988,N_29821);
nor UO_887 (O_887,N_29767,N_29998);
nand UO_888 (O_888,N_29849,N_29862);
and UO_889 (O_889,N_29623,N_29740);
or UO_890 (O_890,N_29744,N_29543);
and UO_891 (O_891,N_29658,N_29536);
nand UO_892 (O_892,N_29556,N_29703);
nand UO_893 (O_893,N_29789,N_29972);
or UO_894 (O_894,N_29503,N_29931);
nor UO_895 (O_895,N_29999,N_29934);
xor UO_896 (O_896,N_29998,N_29577);
xnor UO_897 (O_897,N_29559,N_29874);
nand UO_898 (O_898,N_29735,N_29931);
xnor UO_899 (O_899,N_29751,N_29554);
or UO_900 (O_900,N_29886,N_29913);
nor UO_901 (O_901,N_29892,N_29917);
xnor UO_902 (O_902,N_29601,N_29955);
nand UO_903 (O_903,N_29513,N_29986);
and UO_904 (O_904,N_29838,N_29975);
nor UO_905 (O_905,N_29757,N_29686);
xor UO_906 (O_906,N_29654,N_29542);
or UO_907 (O_907,N_29631,N_29924);
nand UO_908 (O_908,N_29779,N_29972);
xnor UO_909 (O_909,N_29813,N_29676);
and UO_910 (O_910,N_29749,N_29850);
xor UO_911 (O_911,N_29519,N_29758);
and UO_912 (O_912,N_29565,N_29829);
xor UO_913 (O_913,N_29979,N_29691);
or UO_914 (O_914,N_29780,N_29828);
nor UO_915 (O_915,N_29864,N_29755);
xor UO_916 (O_916,N_29502,N_29647);
nor UO_917 (O_917,N_29519,N_29918);
nand UO_918 (O_918,N_29804,N_29570);
nor UO_919 (O_919,N_29974,N_29904);
or UO_920 (O_920,N_29600,N_29698);
or UO_921 (O_921,N_29580,N_29834);
nor UO_922 (O_922,N_29980,N_29724);
xor UO_923 (O_923,N_29690,N_29655);
and UO_924 (O_924,N_29959,N_29672);
or UO_925 (O_925,N_29804,N_29742);
xor UO_926 (O_926,N_29936,N_29740);
nand UO_927 (O_927,N_29848,N_29596);
nand UO_928 (O_928,N_29817,N_29846);
or UO_929 (O_929,N_29970,N_29889);
nand UO_930 (O_930,N_29759,N_29668);
nor UO_931 (O_931,N_29661,N_29958);
and UO_932 (O_932,N_29577,N_29957);
nor UO_933 (O_933,N_29901,N_29897);
nand UO_934 (O_934,N_29842,N_29932);
and UO_935 (O_935,N_29593,N_29835);
nor UO_936 (O_936,N_29670,N_29980);
nor UO_937 (O_937,N_29658,N_29682);
nor UO_938 (O_938,N_29822,N_29918);
nand UO_939 (O_939,N_29729,N_29954);
xor UO_940 (O_940,N_29929,N_29719);
or UO_941 (O_941,N_29684,N_29900);
xor UO_942 (O_942,N_29592,N_29912);
and UO_943 (O_943,N_29824,N_29866);
nand UO_944 (O_944,N_29576,N_29714);
nand UO_945 (O_945,N_29747,N_29715);
xor UO_946 (O_946,N_29830,N_29817);
xnor UO_947 (O_947,N_29793,N_29517);
nand UO_948 (O_948,N_29561,N_29542);
nor UO_949 (O_949,N_29730,N_29953);
or UO_950 (O_950,N_29644,N_29738);
and UO_951 (O_951,N_29925,N_29887);
nor UO_952 (O_952,N_29774,N_29601);
nor UO_953 (O_953,N_29550,N_29689);
nor UO_954 (O_954,N_29963,N_29791);
nor UO_955 (O_955,N_29533,N_29673);
nand UO_956 (O_956,N_29644,N_29959);
or UO_957 (O_957,N_29511,N_29542);
nor UO_958 (O_958,N_29710,N_29725);
nor UO_959 (O_959,N_29567,N_29830);
nand UO_960 (O_960,N_29765,N_29517);
or UO_961 (O_961,N_29513,N_29512);
and UO_962 (O_962,N_29823,N_29860);
xnor UO_963 (O_963,N_29816,N_29566);
and UO_964 (O_964,N_29801,N_29917);
nor UO_965 (O_965,N_29764,N_29814);
xor UO_966 (O_966,N_29888,N_29619);
nor UO_967 (O_967,N_29936,N_29858);
and UO_968 (O_968,N_29715,N_29717);
and UO_969 (O_969,N_29593,N_29822);
or UO_970 (O_970,N_29822,N_29756);
and UO_971 (O_971,N_29552,N_29798);
xor UO_972 (O_972,N_29928,N_29567);
or UO_973 (O_973,N_29581,N_29549);
xor UO_974 (O_974,N_29899,N_29978);
xnor UO_975 (O_975,N_29768,N_29523);
and UO_976 (O_976,N_29746,N_29838);
xor UO_977 (O_977,N_29531,N_29572);
or UO_978 (O_978,N_29933,N_29516);
and UO_979 (O_979,N_29908,N_29672);
or UO_980 (O_980,N_29710,N_29755);
or UO_981 (O_981,N_29532,N_29802);
nand UO_982 (O_982,N_29587,N_29799);
xor UO_983 (O_983,N_29648,N_29788);
and UO_984 (O_984,N_29892,N_29881);
or UO_985 (O_985,N_29910,N_29598);
and UO_986 (O_986,N_29852,N_29714);
xor UO_987 (O_987,N_29917,N_29946);
xor UO_988 (O_988,N_29573,N_29517);
xor UO_989 (O_989,N_29836,N_29856);
xnor UO_990 (O_990,N_29503,N_29972);
xnor UO_991 (O_991,N_29735,N_29676);
nand UO_992 (O_992,N_29937,N_29555);
nor UO_993 (O_993,N_29833,N_29564);
or UO_994 (O_994,N_29587,N_29839);
nand UO_995 (O_995,N_29819,N_29584);
and UO_996 (O_996,N_29693,N_29620);
xor UO_997 (O_997,N_29810,N_29723);
nor UO_998 (O_998,N_29535,N_29971);
xnor UO_999 (O_999,N_29786,N_29801);
xor UO_1000 (O_1000,N_29569,N_29656);
nor UO_1001 (O_1001,N_29573,N_29780);
xnor UO_1002 (O_1002,N_29579,N_29871);
nor UO_1003 (O_1003,N_29998,N_29817);
nand UO_1004 (O_1004,N_29975,N_29878);
xor UO_1005 (O_1005,N_29710,N_29949);
xnor UO_1006 (O_1006,N_29847,N_29811);
xnor UO_1007 (O_1007,N_29986,N_29679);
nor UO_1008 (O_1008,N_29922,N_29623);
or UO_1009 (O_1009,N_29652,N_29771);
nand UO_1010 (O_1010,N_29648,N_29799);
and UO_1011 (O_1011,N_29627,N_29762);
nand UO_1012 (O_1012,N_29649,N_29691);
or UO_1013 (O_1013,N_29866,N_29804);
or UO_1014 (O_1014,N_29797,N_29722);
nor UO_1015 (O_1015,N_29520,N_29519);
or UO_1016 (O_1016,N_29932,N_29914);
nand UO_1017 (O_1017,N_29501,N_29699);
xor UO_1018 (O_1018,N_29642,N_29723);
and UO_1019 (O_1019,N_29552,N_29784);
xor UO_1020 (O_1020,N_29983,N_29918);
nor UO_1021 (O_1021,N_29746,N_29501);
xnor UO_1022 (O_1022,N_29599,N_29969);
nand UO_1023 (O_1023,N_29653,N_29600);
nor UO_1024 (O_1024,N_29637,N_29882);
and UO_1025 (O_1025,N_29780,N_29673);
or UO_1026 (O_1026,N_29517,N_29947);
xnor UO_1027 (O_1027,N_29645,N_29969);
xnor UO_1028 (O_1028,N_29508,N_29757);
nor UO_1029 (O_1029,N_29630,N_29625);
xor UO_1030 (O_1030,N_29709,N_29920);
nor UO_1031 (O_1031,N_29850,N_29558);
nor UO_1032 (O_1032,N_29728,N_29517);
and UO_1033 (O_1033,N_29870,N_29781);
xnor UO_1034 (O_1034,N_29515,N_29944);
nand UO_1035 (O_1035,N_29755,N_29806);
and UO_1036 (O_1036,N_29653,N_29553);
xnor UO_1037 (O_1037,N_29798,N_29575);
nor UO_1038 (O_1038,N_29918,N_29557);
xor UO_1039 (O_1039,N_29586,N_29982);
nand UO_1040 (O_1040,N_29703,N_29748);
and UO_1041 (O_1041,N_29963,N_29525);
or UO_1042 (O_1042,N_29812,N_29681);
nand UO_1043 (O_1043,N_29624,N_29812);
nand UO_1044 (O_1044,N_29806,N_29554);
and UO_1045 (O_1045,N_29816,N_29746);
nor UO_1046 (O_1046,N_29604,N_29942);
nor UO_1047 (O_1047,N_29702,N_29887);
nand UO_1048 (O_1048,N_29738,N_29554);
nand UO_1049 (O_1049,N_29552,N_29608);
or UO_1050 (O_1050,N_29980,N_29520);
nor UO_1051 (O_1051,N_29909,N_29981);
nor UO_1052 (O_1052,N_29724,N_29729);
nor UO_1053 (O_1053,N_29890,N_29629);
nand UO_1054 (O_1054,N_29747,N_29664);
or UO_1055 (O_1055,N_29705,N_29523);
nand UO_1056 (O_1056,N_29763,N_29807);
or UO_1057 (O_1057,N_29650,N_29611);
nor UO_1058 (O_1058,N_29541,N_29574);
and UO_1059 (O_1059,N_29609,N_29506);
nor UO_1060 (O_1060,N_29735,N_29637);
nand UO_1061 (O_1061,N_29638,N_29972);
and UO_1062 (O_1062,N_29506,N_29955);
nand UO_1063 (O_1063,N_29623,N_29975);
nor UO_1064 (O_1064,N_29897,N_29520);
nor UO_1065 (O_1065,N_29767,N_29656);
or UO_1066 (O_1066,N_29990,N_29554);
nor UO_1067 (O_1067,N_29750,N_29562);
nor UO_1068 (O_1068,N_29816,N_29751);
or UO_1069 (O_1069,N_29897,N_29633);
and UO_1070 (O_1070,N_29930,N_29664);
or UO_1071 (O_1071,N_29807,N_29985);
xnor UO_1072 (O_1072,N_29562,N_29721);
xor UO_1073 (O_1073,N_29964,N_29577);
or UO_1074 (O_1074,N_29603,N_29909);
xor UO_1075 (O_1075,N_29956,N_29726);
or UO_1076 (O_1076,N_29727,N_29583);
or UO_1077 (O_1077,N_29812,N_29851);
xnor UO_1078 (O_1078,N_29568,N_29735);
nor UO_1079 (O_1079,N_29815,N_29961);
nor UO_1080 (O_1080,N_29714,N_29508);
xor UO_1081 (O_1081,N_29887,N_29769);
xor UO_1082 (O_1082,N_29700,N_29582);
nand UO_1083 (O_1083,N_29686,N_29887);
and UO_1084 (O_1084,N_29830,N_29839);
and UO_1085 (O_1085,N_29897,N_29600);
nor UO_1086 (O_1086,N_29930,N_29553);
and UO_1087 (O_1087,N_29530,N_29959);
nor UO_1088 (O_1088,N_29687,N_29622);
nand UO_1089 (O_1089,N_29887,N_29521);
nor UO_1090 (O_1090,N_29559,N_29924);
or UO_1091 (O_1091,N_29596,N_29500);
xnor UO_1092 (O_1092,N_29727,N_29570);
nand UO_1093 (O_1093,N_29604,N_29603);
or UO_1094 (O_1094,N_29667,N_29715);
nor UO_1095 (O_1095,N_29571,N_29951);
and UO_1096 (O_1096,N_29722,N_29781);
nor UO_1097 (O_1097,N_29676,N_29753);
nor UO_1098 (O_1098,N_29983,N_29815);
or UO_1099 (O_1099,N_29533,N_29513);
and UO_1100 (O_1100,N_29803,N_29722);
and UO_1101 (O_1101,N_29691,N_29689);
and UO_1102 (O_1102,N_29785,N_29553);
xor UO_1103 (O_1103,N_29966,N_29593);
and UO_1104 (O_1104,N_29760,N_29817);
and UO_1105 (O_1105,N_29564,N_29736);
nor UO_1106 (O_1106,N_29569,N_29634);
or UO_1107 (O_1107,N_29939,N_29524);
nor UO_1108 (O_1108,N_29997,N_29843);
nor UO_1109 (O_1109,N_29880,N_29553);
xnor UO_1110 (O_1110,N_29890,N_29881);
or UO_1111 (O_1111,N_29567,N_29568);
xor UO_1112 (O_1112,N_29598,N_29844);
and UO_1113 (O_1113,N_29893,N_29514);
or UO_1114 (O_1114,N_29719,N_29821);
nor UO_1115 (O_1115,N_29630,N_29972);
or UO_1116 (O_1116,N_29943,N_29960);
or UO_1117 (O_1117,N_29743,N_29971);
and UO_1118 (O_1118,N_29625,N_29968);
xor UO_1119 (O_1119,N_29858,N_29896);
and UO_1120 (O_1120,N_29912,N_29885);
xor UO_1121 (O_1121,N_29789,N_29941);
xnor UO_1122 (O_1122,N_29786,N_29842);
nand UO_1123 (O_1123,N_29957,N_29719);
nor UO_1124 (O_1124,N_29740,N_29640);
and UO_1125 (O_1125,N_29630,N_29698);
xor UO_1126 (O_1126,N_29726,N_29821);
nor UO_1127 (O_1127,N_29816,N_29555);
or UO_1128 (O_1128,N_29980,N_29718);
nor UO_1129 (O_1129,N_29932,N_29531);
and UO_1130 (O_1130,N_29506,N_29886);
xor UO_1131 (O_1131,N_29799,N_29667);
xnor UO_1132 (O_1132,N_29815,N_29939);
nand UO_1133 (O_1133,N_29886,N_29921);
nor UO_1134 (O_1134,N_29941,N_29622);
and UO_1135 (O_1135,N_29797,N_29862);
nor UO_1136 (O_1136,N_29849,N_29599);
nand UO_1137 (O_1137,N_29795,N_29562);
nand UO_1138 (O_1138,N_29826,N_29613);
and UO_1139 (O_1139,N_29580,N_29711);
or UO_1140 (O_1140,N_29748,N_29734);
xor UO_1141 (O_1141,N_29926,N_29607);
and UO_1142 (O_1142,N_29501,N_29747);
nand UO_1143 (O_1143,N_29714,N_29925);
nor UO_1144 (O_1144,N_29950,N_29507);
xor UO_1145 (O_1145,N_29928,N_29863);
xor UO_1146 (O_1146,N_29601,N_29681);
or UO_1147 (O_1147,N_29646,N_29828);
nand UO_1148 (O_1148,N_29761,N_29668);
and UO_1149 (O_1149,N_29648,N_29668);
nor UO_1150 (O_1150,N_29709,N_29924);
and UO_1151 (O_1151,N_29645,N_29872);
nand UO_1152 (O_1152,N_29921,N_29860);
nor UO_1153 (O_1153,N_29524,N_29687);
nor UO_1154 (O_1154,N_29827,N_29689);
nor UO_1155 (O_1155,N_29728,N_29678);
nor UO_1156 (O_1156,N_29584,N_29956);
nand UO_1157 (O_1157,N_29743,N_29830);
nor UO_1158 (O_1158,N_29785,N_29604);
nand UO_1159 (O_1159,N_29714,N_29680);
nor UO_1160 (O_1160,N_29714,N_29724);
or UO_1161 (O_1161,N_29673,N_29906);
or UO_1162 (O_1162,N_29872,N_29868);
or UO_1163 (O_1163,N_29605,N_29962);
and UO_1164 (O_1164,N_29811,N_29765);
and UO_1165 (O_1165,N_29893,N_29970);
and UO_1166 (O_1166,N_29745,N_29612);
xnor UO_1167 (O_1167,N_29560,N_29994);
or UO_1168 (O_1168,N_29588,N_29547);
xor UO_1169 (O_1169,N_29994,N_29778);
and UO_1170 (O_1170,N_29970,N_29936);
and UO_1171 (O_1171,N_29831,N_29770);
xnor UO_1172 (O_1172,N_29809,N_29872);
and UO_1173 (O_1173,N_29551,N_29766);
xnor UO_1174 (O_1174,N_29942,N_29792);
xnor UO_1175 (O_1175,N_29556,N_29549);
or UO_1176 (O_1176,N_29962,N_29964);
nand UO_1177 (O_1177,N_29564,N_29961);
nor UO_1178 (O_1178,N_29873,N_29630);
nor UO_1179 (O_1179,N_29613,N_29638);
or UO_1180 (O_1180,N_29895,N_29625);
nor UO_1181 (O_1181,N_29860,N_29863);
xnor UO_1182 (O_1182,N_29522,N_29512);
nor UO_1183 (O_1183,N_29612,N_29702);
nand UO_1184 (O_1184,N_29724,N_29691);
nand UO_1185 (O_1185,N_29720,N_29667);
or UO_1186 (O_1186,N_29694,N_29504);
nor UO_1187 (O_1187,N_29737,N_29585);
nor UO_1188 (O_1188,N_29881,N_29941);
nor UO_1189 (O_1189,N_29907,N_29832);
and UO_1190 (O_1190,N_29712,N_29943);
xnor UO_1191 (O_1191,N_29938,N_29989);
and UO_1192 (O_1192,N_29971,N_29832);
nand UO_1193 (O_1193,N_29729,N_29623);
nand UO_1194 (O_1194,N_29515,N_29694);
nand UO_1195 (O_1195,N_29575,N_29908);
or UO_1196 (O_1196,N_29628,N_29820);
or UO_1197 (O_1197,N_29587,N_29770);
or UO_1198 (O_1198,N_29572,N_29789);
or UO_1199 (O_1199,N_29692,N_29628);
or UO_1200 (O_1200,N_29842,N_29905);
xnor UO_1201 (O_1201,N_29943,N_29846);
nand UO_1202 (O_1202,N_29734,N_29737);
xor UO_1203 (O_1203,N_29761,N_29508);
nand UO_1204 (O_1204,N_29741,N_29629);
xor UO_1205 (O_1205,N_29715,N_29611);
or UO_1206 (O_1206,N_29872,N_29667);
nor UO_1207 (O_1207,N_29673,N_29599);
nand UO_1208 (O_1208,N_29896,N_29773);
or UO_1209 (O_1209,N_29952,N_29766);
nor UO_1210 (O_1210,N_29650,N_29637);
xor UO_1211 (O_1211,N_29741,N_29687);
and UO_1212 (O_1212,N_29624,N_29661);
nand UO_1213 (O_1213,N_29980,N_29944);
or UO_1214 (O_1214,N_29866,N_29984);
xor UO_1215 (O_1215,N_29806,N_29963);
xnor UO_1216 (O_1216,N_29674,N_29860);
xor UO_1217 (O_1217,N_29881,N_29846);
xor UO_1218 (O_1218,N_29934,N_29898);
nor UO_1219 (O_1219,N_29727,N_29774);
nand UO_1220 (O_1220,N_29842,N_29604);
xnor UO_1221 (O_1221,N_29817,N_29683);
xor UO_1222 (O_1222,N_29591,N_29749);
xor UO_1223 (O_1223,N_29756,N_29848);
or UO_1224 (O_1224,N_29673,N_29742);
nor UO_1225 (O_1225,N_29547,N_29713);
or UO_1226 (O_1226,N_29668,N_29658);
or UO_1227 (O_1227,N_29951,N_29876);
and UO_1228 (O_1228,N_29854,N_29817);
and UO_1229 (O_1229,N_29888,N_29539);
xnor UO_1230 (O_1230,N_29558,N_29848);
or UO_1231 (O_1231,N_29936,N_29928);
nor UO_1232 (O_1232,N_29818,N_29729);
nor UO_1233 (O_1233,N_29517,N_29943);
or UO_1234 (O_1234,N_29804,N_29895);
nand UO_1235 (O_1235,N_29727,N_29636);
nor UO_1236 (O_1236,N_29661,N_29788);
or UO_1237 (O_1237,N_29719,N_29897);
or UO_1238 (O_1238,N_29659,N_29673);
xnor UO_1239 (O_1239,N_29758,N_29539);
or UO_1240 (O_1240,N_29855,N_29789);
nand UO_1241 (O_1241,N_29749,N_29508);
nor UO_1242 (O_1242,N_29874,N_29668);
and UO_1243 (O_1243,N_29619,N_29556);
nor UO_1244 (O_1244,N_29971,N_29984);
xnor UO_1245 (O_1245,N_29617,N_29556);
nor UO_1246 (O_1246,N_29627,N_29950);
nor UO_1247 (O_1247,N_29837,N_29734);
or UO_1248 (O_1248,N_29801,N_29795);
xnor UO_1249 (O_1249,N_29845,N_29893);
nand UO_1250 (O_1250,N_29894,N_29704);
nor UO_1251 (O_1251,N_29589,N_29581);
xor UO_1252 (O_1252,N_29741,N_29910);
or UO_1253 (O_1253,N_29514,N_29843);
and UO_1254 (O_1254,N_29547,N_29699);
nand UO_1255 (O_1255,N_29713,N_29527);
nand UO_1256 (O_1256,N_29817,N_29571);
nor UO_1257 (O_1257,N_29628,N_29944);
or UO_1258 (O_1258,N_29754,N_29803);
or UO_1259 (O_1259,N_29567,N_29588);
or UO_1260 (O_1260,N_29817,N_29549);
and UO_1261 (O_1261,N_29550,N_29699);
or UO_1262 (O_1262,N_29958,N_29741);
nand UO_1263 (O_1263,N_29684,N_29991);
or UO_1264 (O_1264,N_29579,N_29896);
nor UO_1265 (O_1265,N_29560,N_29899);
or UO_1266 (O_1266,N_29745,N_29516);
nand UO_1267 (O_1267,N_29533,N_29839);
or UO_1268 (O_1268,N_29774,N_29540);
nor UO_1269 (O_1269,N_29520,N_29680);
and UO_1270 (O_1270,N_29666,N_29713);
xor UO_1271 (O_1271,N_29709,N_29570);
and UO_1272 (O_1272,N_29554,N_29919);
xor UO_1273 (O_1273,N_29876,N_29983);
xnor UO_1274 (O_1274,N_29633,N_29582);
nor UO_1275 (O_1275,N_29889,N_29988);
nand UO_1276 (O_1276,N_29512,N_29713);
nand UO_1277 (O_1277,N_29634,N_29527);
xor UO_1278 (O_1278,N_29745,N_29649);
or UO_1279 (O_1279,N_29645,N_29880);
or UO_1280 (O_1280,N_29601,N_29798);
nand UO_1281 (O_1281,N_29753,N_29859);
nand UO_1282 (O_1282,N_29738,N_29813);
xor UO_1283 (O_1283,N_29876,N_29687);
nor UO_1284 (O_1284,N_29618,N_29679);
and UO_1285 (O_1285,N_29972,N_29563);
xnor UO_1286 (O_1286,N_29796,N_29659);
nor UO_1287 (O_1287,N_29905,N_29720);
and UO_1288 (O_1288,N_29985,N_29960);
and UO_1289 (O_1289,N_29765,N_29850);
and UO_1290 (O_1290,N_29627,N_29834);
or UO_1291 (O_1291,N_29666,N_29926);
xnor UO_1292 (O_1292,N_29622,N_29501);
or UO_1293 (O_1293,N_29635,N_29929);
nor UO_1294 (O_1294,N_29988,N_29543);
or UO_1295 (O_1295,N_29902,N_29547);
nor UO_1296 (O_1296,N_29540,N_29634);
nor UO_1297 (O_1297,N_29582,N_29659);
xnor UO_1298 (O_1298,N_29959,N_29755);
nor UO_1299 (O_1299,N_29779,N_29746);
xnor UO_1300 (O_1300,N_29846,N_29835);
xnor UO_1301 (O_1301,N_29507,N_29536);
and UO_1302 (O_1302,N_29934,N_29674);
and UO_1303 (O_1303,N_29532,N_29547);
or UO_1304 (O_1304,N_29708,N_29691);
xnor UO_1305 (O_1305,N_29694,N_29866);
or UO_1306 (O_1306,N_29616,N_29770);
xnor UO_1307 (O_1307,N_29913,N_29848);
xor UO_1308 (O_1308,N_29760,N_29829);
or UO_1309 (O_1309,N_29824,N_29541);
xor UO_1310 (O_1310,N_29964,N_29517);
and UO_1311 (O_1311,N_29603,N_29829);
or UO_1312 (O_1312,N_29513,N_29809);
xnor UO_1313 (O_1313,N_29509,N_29853);
and UO_1314 (O_1314,N_29712,N_29559);
nand UO_1315 (O_1315,N_29776,N_29754);
nand UO_1316 (O_1316,N_29946,N_29741);
xor UO_1317 (O_1317,N_29817,N_29874);
and UO_1318 (O_1318,N_29559,N_29676);
or UO_1319 (O_1319,N_29869,N_29713);
nand UO_1320 (O_1320,N_29727,N_29759);
nor UO_1321 (O_1321,N_29532,N_29887);
and UO_1322 (O_1322,N_29710,N_29546);
nor UO_1323 (O_1323,N_29785,N_29697);
xor UO_1324 (O_1324,N_29692,N_29903);
and UO_1325 (O_1325,N_29591,N_29934);
nor UO_1326 (O_1326,N_29616,N_29650);
nor UO_1327 (O_1327,N_29515,N_29905);
nor UO_1328 (O_1328,N_29886,N_29796);
or UO_1329 (O_1329,N_29822,N_29894);
nand UO_1330 (O_1330,N_29996,N_29768);
nor UO_1331 (O_1331,N_29870,N_29528);
or UO_1332 (O_1332,N_29785,N_29731);
nor UO_1333 (O_1333,N_29864,N_29965);
and UO_1334 (O_1334,N_29508,N_29642);
xnor UO_1335 (O_1335,N_29831,N_29996);
nor UO_1336 (O_1336,N_29688,N_29699);
xor UO_1337 (O_1337,N_29644,N_29593);
nand UO_1338 (O_1338,N_29519,N_29589);
xor UO_1339 (O_1339,N_29664,N_29571);
and UO_1340 (O_1340,N_29890,N_29839);
and UO_1341 (O_1341,N_29543,N_29944);
nand UO_1342 (O_1342,N_29520,N_29568);
nor UO_1343 (O_1343,N_29796,N_29878);
or UO_1344 (O_1344,N_29665,N_29740);
nor UO_1345 (O_1345,N_29557,N_29561);
xor UO_1346 (O_1346,N_29624,N_29646);
and UO_1347 (O_1347,N_29826,N_29721);
nor UO_1348 (O_1348,N_29845,N_29668);
and UO_1349 (O_1349,N_29547,N_29745);
xor UO_1350 (O_1350,N_29679,N_29613);
xor UO_1351 (O_1351,N_29775,N_29570);
and UO_1352 (O_1352,N_29997,N_29663);
nand UO_1353 (O_1353,N_29939,N_29521);
nor UO_1354 (O_1354,N_29593,N_29674);
xor UO_1355 (O_1355,N_29876,N_29843);
nor UO_1356 (O_1356,N_29567,N_29923);
xor UO_1357 (O_1357,N_29947,N_29609);
nand UO_1358 (O_1358,N_29850,N_29893);
nand UO_1359 (O_1359,N_29824,N_29583);
or UO_1360 (O_1360,N_29557,N_29519);
nor UO_1361 (O_1361,N_29686,N_29518);
and UO_1362 (O_1362,N_29932,N_29533);
or UO_1363 (O_1363,N_29837,N_29922);
xor UO_1364 (O_1364,N_29588,N_29648);
nor UO_1365 (O_1365,N_29977,N_29981);
nand UO_1366 (O_1366,N_29938,N_29812);
or UO_1367 (O_1367,N_29749,N_29976);
nand UO_1368 (O_1368,N_29910,N_29915);
nand UO_1369 (O_1369,N_29847,N_29591);
nor UO_1370 (O_1370,N_29545,N_29998);
or UO_1371 (O_1371,N_29910,N_29706);
or UO_1372 (O_1372,N_29501,N_29606);
and UO_1373 (O_1373,N_29541,N_29936);
and UO_1374 (O_1374,N_29864,N_29565);
xor UO_1375 (O_1375,N_29951,N_29546);
nand UO_1376 (O_1376,N_29582,N_29964);
nand UO_1377 (O_1377,N_29784,N_29800);
and UO_1378 (O_1378,N_29635,N_29646);
xor UO_1379 (O_1379,N_29542,N_29813);
nand UO_1380 (O_1380,N_29541,N_29736);
and UO_1381 (O_1381,N_29756,N_29875);
nor UO_1382 (O_1382,N_29769,N_29605);
xnor UO_1383 (O_1383,N_29978,N_29792);
and UO_1384 (O_1384,N_29975,N_29835);
nand UO_1385 (O_1385,N_29744,N_29943);
xor UO_1386 (O_1386,N_29917,N_29836);
or UO_1387 (O_1387,N_29629,N_29529);
nor UO_1388 (O_1388,N_29725,N_29923);
nor UO_1389 (O_1389,N_29930,N_29550);
xor UO_1390 (O_1390,N_29737,N_29630);
nand UO_1391 (O_1391,N_29926,N_29598);
and UO_1392 (O_1392,N_29967,N_29954);
nor UO_1393 (O_1393,N_29928,N_29685);
and UO_1394 (O_1394,N_29784,N_29848);
or UO_1395 (O_1395,N_29759,N_29528);
and UO_1396 (O_1396,N_29740,N_29872);
and UO_1397 (O_1397,N_29707,N_29770);
xnor UO_1398 (O_1398,N_29909,N_29946);
and UO_1399 (O_1399,N_29827,N_29877);
and UO_1400 (O_1400,N_29709,N_29697);
nand UO_1401 (O_1401,N_29768,N_29890);
or UO_1402 (O_1402,N_29934,N_29852);
nand UO_1403 (O_1403,N_29720,N_29569);
and UO_1404 (O_1404,N_29838,N_29907);
xnor UO_1405 (O_1405,N_29708,N_29528);
and UO_1406 (O_1406,N_29640,N_29827);
or UO_1407 (O_1407,N_29703,N_29594);
and UO_1408 (O_1408,N_29593,N_29847);
or UO_1409 (O_1409,N_29999,N_29504);
and UO_1410 (O_1410,N_29757,N_29731);
or UO_1411 (O_1411,N_29852,N_29965);
xor UO_1412 (O_1412,N_29634,N_29642);
xnor UO_1413 (O_1413,N_29714,N_29616);
and UO_1414 (O_1414,N_29816,N_29998);
nor UO_1415 (O_1415,N_29609,N_29597);
nor UO_1416 (O_1416,N_29957,N_29822);
and UO_1417 (O_1417,N_29548,N_29931);
xnor UO_1418 (O_1418,N_29600,N_29681);
nand UO_1419 (O_1419,N_29606,N_29972);
nor UO_1420 (O_1420,N_29604,N_29522);
xor UO_1421 (O_1421,N_29772,N_29971);
and UO_1422 (O_1422,N_29553,N_29537);
and UO_1423 (O_1423,N_29562,N_29963);
and UO_1424 (O_1424,N_29632,N_29531);
nor UO_1425 (O_1425,N_29634,N_29973);
or UO_1426 (O_1426,N_29821,N_29752);
nand UO_1427 (O_1427,N_29953,N_29716);
nor UO_1428 (O_1428,N_29781,N_29566);
or UO_1429 (O_1429,N_29672,N_29802);
and UO_1430 (O_1430,N_29784,N_29508);
and UO_1431 (O_1431,N_29958,N_29601);
and UO_1432 (O_1432,N_29989,N_29993);
xnor UO_1433 (O_1433,N_29916,N_29899);
xor UO_1434 (O_1434,N_29926,N_29739);
xnor UO_1435 (O_1435,N_29717,N_29629);
and UO_1436 (O_1436,N_29631,N_29753);
and UO_1437 (O_1437,N_29657,N_29628);
nand UO_1438 (O_1438,N_29521,N_29824);
or UO_1439 (O_1439,N_29923,N_29811);
nor UO_1440 (O_1440,N_29738,N_29890);
or UO_1441 (O_1441,N_29810,N_29666);
nand UO_1442 (O_1442,N_29835,N_29863);
or UO_1443 (O_1443,N_29534,N_29770);
and UO_1444 (O_1444,N_29684,N_29600);
and UO_1445 (O_1445,N_29547,N_29536);
nand UO_1446 (O_1446,N_29618,N_29788);
xor UO_1447 (O_1447,N_29988,N_29859);
nand UO_1448 (O_1448,N_29770,N_29840);
and UO_1449 (O_1449,N_29539,N_29535);
nor UO_1450 (O_1450,N_29628,N_29756);
nor UO_1451 (O_1451,N_29610,N_29635);
nor UO_1452 (O_1452,N_29714,N_29664);
nand UO_1453 (O_1453,N_29672,N_29845);
or UO_1454 (O_1454,N_29559,N_29952);
nor UO_1455 (O_1455,N_29713,N_29578);
or UO_1456 (O_1456,N_29619,N_29715);
xnor UO_1457 (O_1457,N_29585,N_29795);
and UO_1458 (O_1458,N_29840,N_29695);
nand UO_1459 (O_1459,N_29620,N_29652);
nor UO_1460 (O_1460,N_29786,N_29695);
or UO_1461 (O_1461,N_29845,N_29927);
nor UO_1462 (O_1462,N_29939,N_29633);
and UO_1463 (O_1463,N_29930,N_29992);
nor UO_1464 (O_1464,N_29793,N_29562);
xor UO_1465 (O_1465,N_29611,N_29674);
and UO_1466 (O_1466,N_29750,N_29928);
and UO_1467 (O_1467,N_29610,N_29891);
and UO_1468 (O_1468,N_29550,N_29834);
xor UO_1469 (O_1469,N_29861,N_29996);
xor UO_1470 (O_1470,N_29541,N_29562);
or UO_1471 (O_1471,N_29542,N_29627);
xor UO_1472 (O_1472,N_29771,N_29594);
xnor UO_1473 (O_1473,N_29841,N_29875);
nand UO_1474 (O_1474,N_29536,N_29610);
or UO_1475 (O_1475,N_29916,N_29574);
xnor UO_1476 (O_1476,N_29589,N_29882);
nor UO_1477 (O_1477,N_29738,N_29843);
and UO_1478 (O_1478,N_29944,N_29698);
or UO_1479 (O_1479,N_29638,N_29607);
xor UO_1480 (O_1480,N_29821,N_29886);
nand UO_1481 (O_1481,N_29537,N_29697);
and UO_1482 (O_1482,N_29613,N_29931);
nand UO_1483 (O_1483,N_29889,N_29962);
xor UO_1484 (O_1484,N_29573,N_29848);
or UO_1485 (O_1485,N_29721,N_29508);
and UO_1486 (O_1486,N_29609,N_29804);
and UO_1487 (O_1487,N_29860,N_29788);
xor UO_1488 (O_1488,N_29539,N_29995);
nor UO_1489 (O_1489,N_29926,N_29677);
and UO_1490 (O_1490,N_29673,N_29713);
and UO_1491 (O_1491,N_29761,N_29811);
and UO_1492 (O_1492,N_29561,N_29882);
nor UO_1493 (O_1493,N_29741,N_29969);
xor UO_1494 (O_1494,N_29501,N_29560);
nand UO_1495 (O_1495,N_29780,N_29611);
xor UO_1496 (O_1496,N_29930,N_29590);
nand UO_1497 (O_1497,N_29751,N_29718);
xor UO_1498 (O_1498,N_29720,N_29594);
nand UO_1499 (O_1499,N_29872,N_29970);
nand UO_1500 (O_1500,N_29905,N_29707);
xnor UO_1501 (O_1501,N_29603,N_29632);
xnor UO_1502 (O_1502,N_29647,N_29795);
xnor UO_1503 (O_1503,N_29638,N_29789);
xnor UO_1504 (O_1504,N_29534,N_29953);
nor UO_1505 (O_1505,N_29668,N_29904);
nor UO_1506 (O_1506,N_29667,N_29542);
nand UO_1507 (O_1507,N_29716,N_29541);
nor UO_1508 (O_1508,N_29809,N_29913);
nor UO_1509 (O_1509,N_29552,N_29739);
xnor UO_1510 (O_1510,N_29980,N_29838);
and UO_1511 (O_1511,N_29571,N_29699);
or UO_1512 (O_1512,N_29638,N_29552);
nand UO_1513 (O_1513,N_29931,N_29649);
xor UO_1514 (O_1514,N_29789,N_29905);
nand UO_1515 (O_1515,N_29832,N_29864);
nor UO_1516 (O_1516,N_29560,N_29630);
nor UO_1517 (O_1517,N_29875,N_29910);
xor UO_1518 (O_1518,N_29663,N_29788);
and UO_1519 (O_1519,N_29794,N_29892);
nand UO_1520 (O_1520,N_29989,N_29772);
nor UO_1521 (O_1521,N_29891,N_29984);
and UO_1522 (O_1522,N_29602,N_29756);
nor UO_1523 (O_1523,N_29661,N_29531);
and UO_1524 (O_1524,N_29682,N_29690);
nor UO_1525 (O_1525,N_29994,N_29760);
nor UO_1526 (O_1526,N_29573,N_29963);
nor UO_1527 (O_1527,N_29528,N_29763);
nor UO_1528 (O_1528,N_29819,N_29597);
nor UO_1529 (O_1529,N_29779,N_29785);
xor UO_1530 (O_1530,N_29974,N_29717);
and UO_1531 (O_1531,N_29690,N_29961);
nand UO_1532 (O_1532,N_29901,N_29621);
nand UO_1533 (O_1533,N_29769,N_29817);
nand UO_1534 (O_1534,N_29594,N_29782);
and UO_1535 (O_1535,N_29740,N_29889);
and UO_1536 (O_1536,N_29591,N_29997);
xor UO_1537 (O_1537,N_29952,N_29578);
xnor UO_1538 (O_1538,N_29996,N_29612);
and UO_1539 (O_1539,N_29904,N_29945);
and UO_1540 (O_1540,N_29748,N_29549);
and UO_1541 (O_1541,N_29827,N_29797);
nor UO_1542 (O_1542,N_29627,N_29925);
and UO_1543 (O_1543,N_29831,N_29624);
nand UO_1544 (O_1544,N_29875,N_29660);
and UO_1545 (O_1545,N_29671,N_29542);
nand UO_1546 (O_1546,N_29831,N_29503);
and UO_1547 (O_1547,N_29631,N_29599);
nand UO_1548 (O_1548,N_29921,N_29821);
and UO_1549 (O_1549,N_29904,N_29606);
and UO_1550 (O_1550,N_29957,N_29826);
or UO_1551 (O_1551,N_29651,N_29655);
nor UO_1552 (O_1552,N_29843,N_29546);
and UO_1553 (O_1553,N_29868,N_29823);
xor UO_1554 (O_1554,N_29700,N_29612);
or UO_1555 (O_1555,N_29918,N_29706);
nand UO_1556 (O_1556,N_29654,N_29930);
nor UO_1557 (O_1557,N_29560,N_29589);
and UO_1558 (O_1558,N_29927,N_29866);
or UO_1559 (O_1559,N_29815,N_29749);
nand UO_1560 (O_1560,N_29619,N_29675);
or UO_1561 (O_1561,N_29571,N_29620);
nor UO_1562 (O_1562,N_29743,N_29663);
xnor UO_1563 (O_1563,N_29933,N_29964);
xor UO_1564 (O_1564,N_29511,N_29671);
nand UO_1565 (O_1565,N_29717,N_29528);
and UO_1566 (O_1566,N_29982,N_29753);
and UO_1567 (O_1567,N_29595,N_29745);
xnor UO_1568 (O_1568,N_29558,N_29987);
xor UO_1569 (O_1569,N_29979,N_29556);
or UO_1570 (O_1570,N_29813,N_29845);
and UO_1571 (O_1571,N_29579,N_29807);
nor UO_1572 (O_1572,N_29555,N_29592);
or UO_1573 (O_1573,N_29736,N_29851);
and UO_1574 (O_1574,N_29902,N_29806);
and UO_1575 (O_1575,N_29798,N_29761);
xnor UO_1576 (O_1576,N_29876,N_29894);
xnor UO_1577 (O_1577,N_29676,N_29652);
or UO_1578 (O_1578,N_29590,N_29620);
nor UO_1579 (O_1579,N_29781,N_29504);
nor UO_1580 (O_1580,N_29610,N_29971);
and UO_1581 (O_1581,N_29944,N_29906);
nand UO_1582 (O_1582,N_29767,N_29932);
xnor UO_1583 (O_1583,N_29773,N_29577);
or UO_1584 (O_1584,N_29872,N_29844);
and UO_1585 (O_1585,N_29723,N_29541);
nor UO_1586 (O_1586,N_29629,N_29862);
xnor UO_1587 (O_1587,N_29904,N_29509);
and UO_1588 (O_1588,N_29725,N_29946);
xnor UO_1589 (O_1589,N_29782,N_29902);
nor UO_1590 (O_1590,N_29831,N_29556);
nand UO_1591 (O_1591,N_29520,N_29515);
or UO_1592 (O_1592,N_29515,N_29620);
nand UO_1593 (O_1593,N_29674,N_29505);
xor UO_1594 (O_1594,N_29798,N_29814);
xnor UO_1595 (O_1595,N_29879,N_29606);
nor UO_1596 (O_1596,N_29751,N_29778);
and UO_1597 (O_1597,N_29795,N_29868);
and UO_1598 (O_1598,N_29500,N_29914);
or UO_1599 (O_1599,N_29847,N_29790);
nand UO_1600 (O_1600,N_29894,N_29546);
or UO_1601 (O_1601,N_29987,N_29800);
nand UO_1602 (O_1602,N_29907,N_29761);
xor UO_1603 (O_1603,N_29873,N_29898);
nor UO_1604 (O_1604,N_29705,N_29895);
or UO_1605 (O_1605,N_29678,N_29823);
and UO_1606 (O_1606,N_29940,N_29970);
and UO_1607 (O_1607,N_29847,N_29547);
nor UO_1608 (O_1608,N_29666,N_29900);
xnor UO_1609 (O_1609,N_29896,N_29886);
xnor UO_1610 (O_1610,N_29898,N_29700);
or UO_1611 (O_1611,N_29940,N_29976);
xor UO_1612 (O_1612,N_29859,N_29986);
nand UO_1613 (O_1613,N_29911,N_29660);
or UO_1614 (O_1614,N_29920,N_29856);
xnor UO_1615 (O_1615,N_29510,N_29805);
and UO_1616 (O_1616,N_29687,N_29683);
nor UO_1617 (O_1617,N_29639,N_29809);
xor UO_1618 (O_1618,N_29695,N_29750);
and UO_1619 (O_1619,N_29567,N_29947);
or UO_1620 (O_1620,N_29964,N_29800);
and UO_1621 (O_1621,N_29657,N_29961);
xnor UO_1622 (O_1622,N_29797,N_29668);
and UO_1623 (O_1623,N_29883,N_29683);
nand UO_1624 (O_1624,N_29874,N_29623);
nor UO_1625 (O_1625,N_29872,N_29804);
nand UO_1626 (O_1626,N_29957,N_29995);
or UO_1627 (O_1627,N_29977,N_29740);
nand UO_1628 (O_1628,N_29867,N_29953);
xnor UO_1629 (O_1629,N_29937,N_29514);
or UO_1630 (O_1630,N_29826,N_29959);
or UO_1631 (O_1631,N_29841,N_29517);
nor UO_1632 (O_1632,N_29695,N_29831);
or UO_1633 (O_1633,N_29884,N_29875);
nor UO_1634 (O_1634,N_29731,N_29744);
or UO_1635 (O_1635,N_29683,N_29519);
xnor UO_1636 (O_1636,N_29732,N_29545);
or UO_1637 (O_1637,N_29729,N_29859);
or UO_1638 (O_1638,N_29823,N_29684);
or UO_1639 (O_1639,N_29580,N_29994);
nand UO_1640 (O_1640,N_29601,N_29924);
nor UO_1641 (O_1641,N_29936,N_29902);
xor UO_1642 (O_1642,N_29735,N_29595);
xor UO_1643 (O_1643,N_29925,N_29883);
and UO_1644 (O_1644,N_29656,N_29701);
xnor UO_1645 (O_1645,N_29769,N_29745);
nand UO_1646 (O_1646,N_29650,N_29974);
nor UO_1647 (O_1647,N_29684,N_29868);
and UO_1648 (O_1648,N_29775,N_29785);
nor UO_1649 (O_1649,N_29983,N_29923);
and UO_1650 (O_1650,N_29556,N_29684);
nand UO_1651 (O_1651,N_29710,N_29806);
nor UO_1652 (O_1652,N_29810,N_29714);
nor UO_1653 (O_1653,N_29693,N_29978);
xnor UO_1654 (O_1654,N_29598,N_29917);
nor UO_1655 (O_1655,N_29809,N_29977);
nand UO_1656 (O_1656,N_29992,N_29503);
xor UO_1657 (O_1657,N_29703,N_29854);
xor UO_1658 (O_1658,N_29938,N_29534);
xnor UO_1659 (O_1659,N_29950,N_29931);
nand UO_1660 (O_1660,N_29611,N_29749);
and UO_1661 (O_1661,N_29697,N_29844);
nand UO_1662 (O_1662,N_29945,N_29885);
xor UO_1663 (O_1663,N_29970,N_29510);
or UO_1664 (O_1664,N_29713,N_29569);
and UO_1665 (O_1665,N_29636,N_29658);
nand UO_1666 (O_1666,N_29633,N_29573);
nand UO_1667 (O_1667,N_29623,N_29724);
nor UO_1668 (O_1668,N_29817,N_29664);
nor UO_1669 (O_1669,N_29505,N_29737);
or UO_1670 (O_1670,N_29530,N_29743);
xnor UO_1671 (O_1671,N_29995,N_29929);
or UO_1672 (O_1672,N_29723,N_29686);
nand UO_1673 (O_1673,N_29813,N_29790);
and UO_1674 (O_1674,N_29847,N_29957);
or UO_1675 (O_1675,N_29997,N_29628);
and UO_1676 (O_1676,N_29852,N_29963);
nor UO_1677 (O_1677,N_29796,N_29707);
xor UO_1678 (O_1678,N_29740,N_29825);
and UO_1679 (O_1679,N_29835,N_29562);
nor UO_1680 (O_1680,N_29573,N_29651);
nor UO_1681 (O_1681,N_29823,N_29966);
xor UO_1682 (O_1682,N_29573,N_29817);
or UO_1683 (O_1683,N_29529,N_29563);
and UO_1684 (O_1684,N_29532,N_29610);
or UO_1685 (O_1685,N_29914,N_29924);
or UO_1686 (O_1686,N_29623,N_29569);
nor UO_1687 (O_1687,N_29717,N_29728);
and UO_1688 (O_1688,N_29801,N_29877);
nor UO_1689 (O_1689,N_29619,N_29980);
xnor UO_1690 (O_1690,N_29557,N_29872);
and UO_1691 (O_1691,N_29810,N_29766);
xor UO_1692 (O_1692,N_29966,N_29679);
nand UO_1693 (O_1693,N_29676,N_29748);
xnor UO_1694 (O_1694,N_29548,N_29511);
xor UO_1695 (O_1695,N_29630,N_29940);
and UO_1696 (O_1696,N_29804,N_29779);
nor UO_1697 (O_1697,N_29640,N_29943);
xnor UO_1698 (O_1698,N_29570,N_29620);
nand UO_1699 (O_1699,N_29892,N_29508);
nand UO_1700 (O_1700,N_29711,N_29770);
nor UO_1701 (O_1701,N_29899,N_29554);
and UO_1702 (O_1702,N_29556,N_29536);
nand UO_1703 (O_1703,N_29517,N_29873);
xor UO_1704 (O_1704,N_29661,N_29877);
nand UO_1705 (O_1705,N_29731,N_29948);
xnor UO_1706 (O_1706,N_29567,N_29964);
xor UO_1707 (O_1707,N_29882,N_29780);
xor UO_1708 (O_1708,N_29546,N_29620);
or UO_1709 (O_1709,N_29713,N_29687);
xnor UO_1710 (O_1710,N_29777,N_29753);
nand UO_1711 (O_1711,N_29722,N_29881);
and UO_1712 (O_1712,N_29812,N_29546);
xnor UO_1713 (O_1713,N_29823,N_29669);
xnor UO_1714 (O_1714,N_29607,N_29714);
or UO_1715 (O_1715,N_29992,N_29770);
and UO_1716 (O_1716,N_29507,N_29945);
and UO_1717 (O_1717,N_29746,N_29712);
nand UO_1718 (O_1718,N_29517,N_29872);
nand UO_1719 (O_1719,N_29885,N_29933);
nand UO_1720 (O_1720,N_29630,N_29929);
xnor UO_1721 (O_1721,N_29702,N_29850);
nand UO_1722 (O_1722,N_29706,N_29513);
or UO_1723 (O_1723,N_29537,N_29899);
xnor UO_1724 (O_1724,N_29629,N_29607);
nand UO_1725 (O_1725,N_29686,N_29977);
nand UO_1726 (O_1726,N_29624,N_29879);
xor UO_1727 (O_1727,N_29621,N_29730);
and UO_1728 (O_1728,N_29529,N_29615);
and UO_1729 (O_1729,N_29567,N_29689);
xnor UO_1730 (O_1730,N_29724,N_29841);
and UO_1731 (O_1731,N_29555,N_29877);
xor UO_1732 (O_1732,N_29902,N_29912);
xor UO_1733 (O_1733,N_29766,N_29530);
xor UO_1734 (O_1734,N_29884,N_29805);
xnor UO_1735 (O_1735,N_29587,N_29735);
xnor UO_1736 (O_1736,N_29881,N_29837);
or UO_1737 (O_1737,N_29952,N_29553);
or UO_1738 (O_1738,N_29648,N_29680);
nand UO_1739 (O_1739,N_29604,N_29663);
nor UO_1740 (O_1740,N_29880,N_29738);
xor UO_1741 (O_1741,N_29667,N_29619);
nor UO_1742 (O_1742,N_29737,N_29607);
and UO_1743 (O_1743,N_29683,N_29726);
nor UO_1744 (O_1744,N_29862,N_29997);
or UO_1745 (O_1745,N_29933,N_29579);
or UO_1746 (O_1746,N_29803,N_29933);
or UO_1747 (O_1747,N_29675,N_29569);
nand UO_1748 (O_1748,N_29964,N_29730);
xor UO_1749 (O_1749,N_29768,N_29749);
or UO_1750 (O_1750,N_29697,N_29507);
nor UO_1751 (O_1751,N_29995,N_29848);
nor UO_1752 (O_1752,N_29566,N_29913);
nor UO_1753 (O_1753,N_29754,N_29973);
nor UO_1754 (O_1754,N_29579,N_29662);
or UO_1755 (O_1755,N_29678,N_29872);
or UO_1756 (O_1756,N_29935,N_29695);
nor UO_1757 (O_1757,N_29780,N_29661);
nor UO_1758 (O_1758,N_29509,N_29916);
nand UO_1759 (O_1759,N_29602,N_29763);
nor UO_1760 (O_1760,N_29944,N_29529);
nor UO_1761 (O_1761,N_29571,N_29842);
or UO_1762 (O_1762,N_29552,N_29991);
nor UO_1763 (O_1763,N_29642,N_29801);
and UO_1764 (O_1764,N_29908,N_29564);
and UO_1765 (O_1765,N_29876,N_29626);
nand UO_1766 (O_1766,N_29615,N_29826);
xor UO_1767 (O_1767,N_29920,N_29936);
nand UO_1768 (O_1768,N_29878,N_29656);
xor UO_1769 (O_1769,N_29738,N_29685);
nand UO_1770 (O_1770,N_29994,N_29765);
and UO_1771 (O_1771,N_29693,N_29626);
xnor UO_1772 (O_1772,N_29996,N_29671);
nand UO_1773 (O_1773,N_29919,N_29737);
or UO_1774 (O_1774,N_29589,N_29998);
nor UO_1775 (O_1775,N_29585,N_29656);
nand UO_1776 (O_1776,N_29685,N_29693);
xor UO_1777 (O_1777,N_29602,N_29643);
nor UO_1778 (O_1778,N_29753,N_29590);
nor UO_1779 (O_1779,N_29734,N_29756);
nand UO_1780 (O_1780,N_29671,N_29763);
or UO_1781 (O_1781,N_29782,N_29504);
xnor UO_1782 (O_1782,N_29798,N_29859);
and UO_1783 (O_1783,N_29774,N_29973);
xnor UO_1784 (O_1784,N_29561,N_29866);
xor UO_1785 (O_1785,N_29576,N_29749);
nand UO_1786 (O_1786,N_29506,N_29991);
xnor UO_1787 (O_1787,N_29556,N_29559);
nand UO_1788 (O_1788,N_29615,N_29556);
xnor UO_1789 (O_1789,N_29881,N_29592);
or UO_1790 (O_1790,N_29727,N_29694);
and UO_1791 (O_1791,N_29892,N_29581);
xnor UO_1792 (O_1792,N_29856,N_29843);
xor UO_1793 (O_1793,N_29612,N_29728);
nor UO_1794 (O_1794,N_29986,N_29888);
or UO_1795 (O_1795,N_29779,N_29561);
xnor UO_1796 (O_1796,N_29751,N_29888);
and UO_1797 (O_1797,N_29909,N_29721);
xor UO_1798 (O_1798,N_29907,N_29888);
nor UO_1799 (O_1799,N_29506,N_29517);
or UO_1800 (O_1800,N_29596,N_29602);
nor UO_1801 (O_1801,N_29992,N_29572);
and UO_1802 (O_1802,N_29798,N_29555);
nor UO_1803 (O_1803,N_29552,N_29942);
nor UO_1804 (O_1804,N_29874,N_29596);
or UO_1805 (O_1805,N_29502,N_29547);
and UO_1806 (O_1806,N_29967,N_29684);
nand UO_1807 (O_1807,N_29968,N_29567);
nand UO_1808 (O_1808,N_29881,N_29767);
or UO_1809 (O_1809,N_29921,N_29811);
nand UO_1810 (O_1810,N_29764,N_29540);
xor UO_1811 (O_1811,N_29845,N_29555);
nand UO_1812 (O_1812,N_29957,N_29740);
and UO_1813 (O_1813,N_29672,N_29668);
or UO_1814 (O_1814,N_29705,N_29524);
and UO_1815 (O_1815,N_29874,N_29750);
nor UO_1816 (O_1816,N_29915,N_29925);
or UO_1817 (O_1817,N_29590,N_29776);
nand UO_1818 (O_1818,N_29789,N_29564);
xor UO_1819 (O_1819,N_29576,N_29734);
nor UO_1820 (O_1820,N_29587,N_29990);
or UO_1821 (O_1821,N_29787,N_29783);
and UO_1822 (O_1822,N_29610,N_29588);
or UO_1823 (O_1823,N_29730,N_29813);
or UO_1824 (O_1824,N_29919,N_29922);
nor UO_1825 (O_1825,N_29922,N_29778);
nand UO_1826 (O_1826,N_29711,N_29848);
nand UO_1827 (O_1827,N_29932,N_29843);
or UO_1828 (O_1828,N_29787,N_29980);
nor UO_1829 (O_1829,N_29886,N_29999);
nand UO_1830 (O_1830,N_29862,N_29908);
or UO_1831 (O_1831,N_29533,N_29550);
and UO_1832 (O_1832,N_29567,N_29569);
nor UO_1833 (O_1833,N_29680,N_29721);
or UO_1834 (O_1834,N_29775,N_29947);
or UO_1835 (O_1835,N_29751,N_29689);
xor UO_1836 (O_1836,N_29549,N_29994);
nor UO_1837 (O_1837,N_29792,N_29802);
xnor UO_1838 (O_1838,N_29644,N_29651);
nor UO_1839 (O_1839,N_29864,N_29886);
nand UO_1840 (O_1840,N_29968,N_29908);
nor UO_1841 (O_1841,N_29653,N_29948);
nand UO_1842 (O_1842,N_29803,N_29505);
nor UO_1843 (O_1843,N_29707,N_29592);
or UO_1844 (O_1844,N_29828,N_29532);
or UO_1845 (O_1845,N_29810,N_29572);
nor UO_1846 (O_1846,N_29819,N_29815);
nor UO_1847 (O_1847,N_29949,N_29627);
xor UO_1848 (O_1848,N_29595,N_29950);
xnor UO_1849 (O_1849,N_29636,N_29812);
nand UO_1850 (O_1850,N_29527,N_29685);
nand UO_1851 (O_1851,N_29742,N_29917);
and UO_1852 (O_1852,N_29974,N_29695);
xnor UO_1853 (O_1853,N_29512,N_29922);
nor UO_1854 (O_1854,N_29948,N_29755);
nand UO_1855 (O_1855,N_29956,N_29985);
and UO_1856 (O_1856,N_29621,N_29628);
xnor UO_1857 (O_1857,N_29567,N_29990);
and UO_1858 (O_1858,N_29530,N_29704);
or UO_1859 (O_1859,N_29637,N_29850);
xnor UO_1860 (O_1860,N_29643,N_29721);
nor UO_1861 (O_1861,N_29616,N_29677);
nand UO_1862 (O_1862,N_29917,N_29833);
nand UO_1863 (O_1863,N_29726,N_29698);
xor UO_1864 (O_1864,N_29772,N_29683);
nor UO_1865 (O_1865,N_29816,N_29878);
nand UO_1866 (O_1866,N_29702,N_29778);
nand UO_1867 (O_1867,N_29796,N_29596);
nor UO_1868 (O_1868,N_29808,N_29743);
nor UO_1869 (O_1869,N_29834,N_29839);
and UO_1870 (O_1870,N_29741,N_29959);
or UO_1871 (O_1871,N_29687,N_29989);
nor UO_1872 (O_1872,N_29603,N_29528);
nand UO_1873 (O_1873,N_29550,N_29774);
xnor UO_1874 (O_1874,N_29938,N_29771);
nand UO_1875 (O_1875,N_29959,N_29690);
or UO_1876 (O_1876,N_29634,N_29800);
nor UO_1877 (O_1877,N_29961,N_29919);
and UO_1878 (O_1878,N_29594,N_29934);
and UO_1879 (O_1879,N_29779,N_29992);
nand UO_1880 (O_1880,N_29715,N_29914);
and UO_1881 (O_1881,N_29566,N_29865);
nor UO_1882 (O_1882,N_29791,N_29569);
or UO_1883 (O_1883,N_29741,N_29575);
xnor UO_1884 (O_1884,N_29738,N_29851);
xor UO_1885 (O_1885,N_29925,N_29776);
xnor UO_1886 (O_1886,N_29793,N_29528);
and UO_1887 (O_1887,N_29545,N_29887);
nand UO_1888 (O_1888,N_29943,N_29948);
xor UO_1889 (O_1889,N_29886,N_29932);
nand UO_1890 (O_1890,N_29943,N_29586);
or UO_1891 (O_1891,N_29815,N_29509);
nor UO_1892 (O_1892,N_29536,N_29503);
xnor UO_1893 (O_1893,N_29713,N_29709);
or UO_1894 (O_1894,N_29995,N_29899);
and UO_1895 (O_1895,N_29890,N_29885);
nand UO_1896 (O_1896,N_29585,N_29925);
nand UO_1897 (O_1897,N_29559,N_29585);
xor UO_1898 (O_1898,N_29566,N_29727);
and UO_1899 (O_1899,N_29659,N_29815);
nand UO_1900 (O_1900,N_29530,N_29908);
nor UO_1901 (O_1901,N_29826,N_29925);
or UO_1902 (O_1902,N_29785,N_29819);
nor UO_1903 (O_1903,N_29565,N_29802);
nor UO_1904 (O_1904,N_29695,N_29984);
or UO_1905 (O_1905,N_29718,N_29782);
nand UO_1906 (O_1906,N_29747,N_29702);
xnor UO_1907 (O_1907,N_29976,N_29820);
xor UO_1908 (O_1908,N_29885,N_29733);
or UO_1909 (O_1909,N_29530,N_29758);
xor UO_1910 (O_1910,N_29591,N_29985);
nand UO_1911 (O_1911,N_29965,N_29563);
nor UO_1912 (O_1912,N_29566,N_29879);
and UO_1913 (O_1913,N_29883,N_29814);
nor UO_1914 (O_1914,N_29714,N_29676);
xnor UO_1915 (O_1915,N_29531,N_29666);
and UO_1916 (O_1916,N_29868,N_29738);
or UO_1917 (O_1917,N_29699,N_29826);
nor UO_1918 (O_1918,N_29506,N_29617);
nand UO_1919 (O_1919,N_29527,N_29644);
nand UO_1920 (O_1920,N_29658,N_29654);
or UO_1921 (O_1921,N_29739,N_29651);
nor UO_1922 (O_1922,N_29975,N_29786);
xor UO_1923 (O_1923,N_29958,N_29501);
or UO_1924 (O_1924,N_29728,N_29548);
nor UO_1925 (O_1925,N_29727,N_29608);
nor UO_1926 (O_1926,N_29967,N_29989);
nand UO_1927 (O_1927,N_29828,N_29995);
nand UO_1928 (O_1928,N_29703,N_29820);
nor UO_1929 (O_1929,N_29823,N_29794);
xor UO_1930 (O_1930,N_29857,N_29759);
or UO_1931 (O_1931,N_29716,N_29553);
or UO_1932 (O_1932,N_29512,N_29537);
or UO_1933 (O_1933,N_29709,N_29724);
xor UO_1934 (O_1934,N_29687,N_29537);
nor UO_1935 (O_1935,N_29955,N_29616);
nand UO_1936 (O_1936,N_29562,N_29540);
xor UO_1937 (O_1937,N_29632,N_29904);
nand UO_1938 (O_1938,N_29677,N_29756);
nand UO_1939 (O_1939,N_29861,N_29521);
nand UO_1940 (O_1940,N_29561,N_29878);
or UO_1941 (O_1941,N_29900,N_29774);
nor UO_1942 (O_1942,N_29692,N_29838);
xor UO_1943 (O_1943,N_29875,N_29788);
nor UO_1944 (O_1944,N_29802,N_29971);
xnor UO_1945 (O_1945,N_29968,N_29550);
or UO_1946 (O_1946,N_29564,N_29750);
and UO_1947 (O_1947,N_29782,N_29575);
or UO_1948 (O_1948,N_29560,N_29685);
xor UO_1949 (O_1949,N_29681,N_29946);
nand UO_1950 (O_1950,N_29718,N_29905);
or UO_1951 (O_1951,N_29740,N_29820);
and UO_1952 (O_1952,N_29822,N_29522);
or UO_1953 (O_1953,N_29585,N_29772);
and UO_1954 (O_1954,N_29599,N_29674);
or UO_1955 (O_1955,N_29936,N_29527);
and UO_1956 (O_1956,N_29513,N_29738);
xnor UO_1957 (O_1957,N_29611,N_29576);
xor UO_1958 (O_1958,N_29881,N_29954);
nand UO_1959 (O_1959,N_29934,N_29726);
or UO_1960 (O_1960,N_29825,N_29590);
nor UO_1961 (O_1961,N_29977,N_29927);
nand UO_1962 (O_1962,N_29916,N_29933);
or UO_1963 (O_1963,N_29831,N_29951);
and UO_1964 (O_1964,N_29771,N_29707);
xor UO_1965 (O_1965,N_29889,N_29906);
xnor UO_1966 (O_1966,N_29841,N_29865);
nor UO_1967 (O_1967,N_29643,N_29537);
nand UO_1968 (O_1968,N_29762,N_29611);
and UO_1969 (O_1969,N_29741,N_29875);
xnor UO_1970 (O_1970,N_29833,N_29633);
or UO_1971 (O_1971,N_29646,N_29827);
nor UO_1972 (O_1972,N_29929,N_29846);
or UO_1973 (O_1973,N_29955,N_29633);
and UO_1974 (O_1974,N_29923,N_29604);
or UO_1975 (O_1975,N_29950,N_29695);
or UO_1976 (O_1976,N_29784,N_29806);
or UO_1977 (O_1977,N_29796,N_29726);
and UO_1978 (O_1978,N_29587,N_29793);
and UO_1979 (O_1979,N_29563,N_29606);
and UO_1980 (O_1980,N_29899,N_29667);
or UO_1981 (O_1981,N_29645,N_29747);
nand UO_1982 (O_1982,N_29783,N_29748);
and UO_1983 (O_1983,N_29957,N_29508);
or UO_1984 (O_1984,N_29877,N_29519);
nor UO_1985 (O_1985,N_29710,N_29886);
xnor UO_1986 (O_1986,N_29646,N_29568);
nor UO_1987 (O_1987,N_29950,N_29913);
nand UO_1988 (O_1988,N_29879,N_29500);
or UO_1989 (O_1989,N_29748,N_29852);
xor UO_1990 (O_1990,N_29538,N_29624);
or UO_1991 (O_1991,N_29546,N_29840);
and UO_1992 (O_1992,N_29840,N_29559);
nand UO_1993 (O_1993,N_29554,N_29676);
nor UO_1994 (O_1994,N_29758,N_29708);
nand UO_1995 (O_1995,N_29651,N_29858);
nand UO_1996 (O_1996,N_29694,N_29970);
or UO_1997 (O_1997,N_29697,N_29796);
xor UO_1998 (O_1998,N_29639,N_29862);
xor UO_1999 (O_1999,N_29652,N_29818);
or UO_2000 (O_2000,N_29638,N_29919);
and UO_2001 (O_2001,N_29521,N_29586);
and UO_2002 (O_2002,N_29820,N_29936);
and UO_2003 (O_2003,N_29690,N_29697);
nor UO_2004 (O_2004,N_29966,N_29524);
xor UO_2005 (O_2005,N_29595,N_29988);
xnor UO_2006 (O_2006,N_29727,N_29843);
and UO_2007 (O_2007,N_29983,N_29911);
xor UO_2008 (O_2008,N_29917,N_29807);
or UO_2009 (O_2009,N_29702,N_29972);
nor UO_2010 (O_2010,N_29869,N_29561);
nor UO_2011 (O_2011,N_29793,N_29866);
nor UO_2012 (O_2012,N_29932,N_29772);
nand UO_2013 (O_2013,N_29596,N_29587);
xor UO_2014 (O_2014,N_29620,N_29810);
and UO_2015 (O_2015,N_29626,N_29945);
nand UO_2016 (O_2016,N_29827,N_29699);
nand UO_2017 (O_2017,N_29585,N_29804);
xor UO_2018 (O_2018,N_29787,N_29726);
xor UO_2019 (O_2019,N_29787,N_29596);
and UO_2020 (O_2020,N_29994,N_29874);
xor UO_2021 (O_2021,N_29500,N_29622);
xnor UO_2022 (O_2022,N_29521,N_29773);
nor UO_2023 (O_2023,N_29791,N_29688);
nor UO_2024 (O_2024,N_29888,N_29876);
or UO_2025 (O_2025,N_29745,N_29871);
nor UO_2026 (O_2026,N_29993,N_29817);
nand UO_2027 (O_2027,N_29946,N_29925);
nand UO_2028 (O_2028,N_29940,N_29655);
xnor UO_2029 (O_2029,N_29675,N_29604);
or UO_2030 (O_2030,N_29852,N_29946);
xnor UO_2031 (O_2031,N_29692,N_29890);
and UO_2032 (O_2032,N_29532,N_29980);
xnor UO_2033 (O_2033,N_29682,N_29798);
xor UO_2034 (O_2034,N_29641,N_29614);
nand UO_2035 (O_2035,N_29603,N_29694);
xor UO_2036 (O_2036,N_29555,N_29921);
nand UO_2037 (O_2037,N_29785,N_29890);
or UO_2038 (O_2038,N_29695,N_29875);
nand UO_2039 (O_2039,N_29721,N_29568);
nand UO_2040 (O_2040,N_29523,N_29940);
nor UO_2041 (O_2041,N_29907,N_29545);
nand UO_2042 (O_2042,N_29981,N_29716);
nand UO_2043 (O_2043,N_29664,N_29951);
or UO_2044 (O_2044,N_29861,N_29759);
and UO_2045 (O_2045,N_29598,N_29692);
nand UO_2046 (O_2046,N_29765,N_29931);
nor UO_2047 (O_2047,N_29587,N_29562);
or UO_2048 (O_2048,N_29699,N_29503);
nor UO_2049 (O_2049,N_29805,N_29610);
nand UO_2050 (O_2050,N_29631,N_29795);
or UO_2051 (O_2051,N_29811,N_29799);
nor UO_2052 (O_2052,N_29941,N_29771);
and UO_2053 (O_2053,N_29599,N_29606);
and UO_2054 (O_2054,N_29667,N_29612);
or UO_2055 (O_2055,N_29831,N_29872);
and UO_2056 (O_2056,N_29934,N_29560);
nand UO_2057 (O_2057,N_29711,N_29635);
or UO_2058 (O_2058,N_29972,N_29765);
or UO_2059 (O_2059,N_29666,N_29747);
and UO_2060 (O_2060,N_29546,N_29848);
xor UO_2061 (O_2061,N_29756,N_29580);
xnor UO_2062 (O_2062,N_29757,N_29887);
nor UO_2063 (O_2063,N_29676,N_29964);
or UO_2064 (O_2064,N_29582,N_29600);
or UO_2065 (O_2065,N_29568,N_29654);
and UO_2066 (O_2066,N_29686,N_29566);
and UO_2067 (O_2067,N_29690,N_29954);
xor UO_2068 (O_2068,N_29865,N_29927);
or UO_2069 (O_2069,N_29519,N_29575);
xnor UO_2070 (O_2070,N_29842,N_29692);
nor UO_2071 (O_2071,N_29563,N_29862);
nand UO_2072 (O_2072,N_29717,N_29935);
nand UO_2073 (O_2073,N_29887,N_29753);
xor UO_2074 (O_2074,N_29957,N_29661);
nor UO_2075 (O_2075,N_29656,N_29848);
nand UO_2076 (O_2076,N_29957,N_29518);
and UO_2077 (O_2077,N_29909,N_29547);
nand UO_2078 (O_2078,N_29818,N_29738);
nor UO_2079 (O_2079,N_29702,N_29783);
nand UO_2080 (O_2080,N_29901,N_29592);
and UO_2081 (O_2081,N_29678,N_29808);
nand UO_2082 (O_2082,N_29924,N_29796);
nand UO_2083 (O_2083,N_29790,N_29857);
and UO_2084 (O_2084,N_29833,N_29980);
or UO_2085 (O_2085,N_29787,N_29824);
nand UO_2086 (O_2086,N_29646,N_29518);
or UO_2087 (O_2087,N_29539,N_29984);
or UO_2088 (O_2088,N_29958,N_29515);
or UO_2089 (O_2089,N_29502,N_29689);
nor UO_2090 (O_2090,N_29778,N_29663);
or UO_2091 (O_2091,N_29893,N_29889);
nor UO_2092 (O_2092,N_29523,N_29979);
nand UO_2093 (O_2093,N_29520,N_29662);
nand UO_2094 (O_2094,N_29566,N_29968);
nor UO_2095 (O_2095,N_29715,N_29999);
and UO_2096 (O_2096,N_29635,N_29952);
xnor UO_2097 (O_2097,N_29945,N_29791);
and UO_2098 (O_2098,N_29626,N_29904);
xnor UO_2099 (O_2099,N_29622,N_29844);
and UO_2100 (O_2100,N_29571,N_29980);
xor UO_2101 (O_2101,N_29991,N_29529);
and UO_2102 (O_2102,N_29552,N_29650);
or UO_2103 (O_2103,N_29527,N_29505);
nor UO_2104 (O_2104,N_29688,N_29826);
nand UO_2105 (O_2105,N_29784,N_29602);
and UO_2106 (O_2106,N_29992,N_29717);
and UO_2107 (O_2107,N_29973,N_29751);
or UO_2108 (O_2108,N_29610,N_29821);
or UO_2109 (O_2109,N_29870,N_29962);
nand UO_2110 (O_2110,N_29835,N_29608);
and UO_2111 (O_2111,N_29574,N_29628);
nand UO_2112 (O_2112,N_29809,N_29888);
nand UO_2113 (O_2113,N_29794,N_29697);
xnor UO_2114 (O_2114,N_29883,N_29559);
or UO_2115 (O_2115,N_29829,N_29602);
nor UO_2116 (O_2116,N_29882,N_29621);
or UO_2117 (O_2117,N_29839,N_29654);
xnor UO_2118 (O_2118,N_29827,N_29919);
nand UO_2119 (O_2119,N_29632,N_29594);
xor UO_2120 (O_2120,N_29889,N_29907);
and UO_2121 (O_2121,N_29970,N_29915);
nor UO_2122 (O_2122,N_29737,N_29664);
nand UO_2123 (O_2123,N_29737,N_29739);
nand UO_2124 (O_2124,N_29964,N_29651);
or UO_2125 (O_2125,N_29907,N_29655);
and UO_2126 (O_2126,N_29909,N_29962);
and UO_2127 (O_2127,N_29574,N_29985);
nand UO_2128 (O_2128,N_29701,N_29503);
and UO_2129 (O_2129,N_29674,N_29561);
nor UO_2130 (O_2130,N_29830,N_29774);
nor UO_2131 (O_2131,N_29890,N_29852);
nor UO_2132 (O_2132,N_29595,N_29873);
or UO_2133 (O_2133,N_29844,N_29763);
or UO_2134 (O_2134,N_29912,N_29824);
and UO_2135 (O_2135,N_29999,N_29626);
and UO_2136 (O_2136,N_29741,N_29732);
nand UO_2137 (O_2137,N_29711,N_29532);
nor UO_2138 (O_2138,N_29552,N_29894);
and UO_2139 (O_2139,N_29782,N_29518);
xnor UO_2140 (O_2140,N_29944,N_29957);
and UO_2141 (O_2141,N_29711,N_29703);
and UO_2142 (O_2142,N_29840,N_29885);
nor UO_2143 (O_2143,N_29899,N_29650);
and UO_2144 (O_2144,N_29587,N_29559);
or UO_2145 (O_2145,N_29900,N_29565);
and UO_2146 (O_2146,N_29811,N_29688);
xor UO_2147 (O_2147,N_29813,N_29570);
and UO_2148 (O_2148,N_29533,N_29812);
xor UO_2149 (O_2149,N_29870,N_29559);
xor UO_2150 (O_2150,N_29746,N_29696);
and UO_2151 (O_2151,N_29984,N_29570);
nor UO_2152 (O_2152,N_29549,N_29623);
nor UO_2153 (O_2153,N_29698,N_29782);
nand UO_2154 (O_2154,N_29644,N_29777);
nand UO_2155 (O_2155,N_29739,N_29793);
xnor UO_2156 (O_2156,N_29861,N_29799);
nor UO_2157 (O_2157,N_29642,N_29554);
or UO_2158 (O_2158,N_29612,N_29682);
or UO_2159 (O_2159,N_29914,N_29773);
xor UO_2160 (O_2160,N_29764,N_29554);
nand UO_2161 (O_2161,N_29875,N_29517);
nor UO_2162 (O_2162,N_29645,N_29802);
nor UO_2163 (O_2163,N_29957,N_29506);
xnor UO_2164 (O_2164,N_29879,N_29546);
xnor UO_2165 (O_2165,N_29598,N_29696);
and UO_2166 (O_2166,N_29816,N_29509);
nor UO_2167 (O_2167,N_29762,N_29948);
nor UO_2168 (O_2168,N_29746,N_29507);
nor UO_2169 (O_2169,N_29626,N_29833);
or UO_2170 (O_2170,N_29616,N_29995);
xor UO_2171 (O_2171,N_29906,N_29724);
nor UO_2172 (O_2172,N_29868,N_29780);
nand UO_2173 (O_2173,N_29579,N_29746);
nor UO_2174 (O_2174,N_29910,N_29840);
nor UO_2175 (O_2175,N_29871,N_29524);
or UO_2176 (O_2176,N_29721,N_29811);
and UO_2177 (O_2177,N_29744,N_29968);
and UO_2178 (O_2178,N_29943,N_29835);
and UO_2179 (O_2179,N_29801,N_29566);
nor UO_2180 (O_2180,N_29563,N_29790);
nand UO_2181 (O_2181,N_29874,N_29626);
xor UO_2182 (O_2182,N_29921,N_29744);
nand UO_2183 (O_2183,N_29718,N_29655);
nand UO_2184 (O_2184,N_29984,N_29569);
nand UO_2185 (O_2185,N_29936,N_29759);
or UO_2186 (O_2186,N_29862,N_29824);
nor UO_2187 (O_2187,N_29692,N_29831);
nor UO_2188 (O_2188,N_29953,N_29714);
or UO_2189 (O_2189,N_29598,N_29720);
xor UO_2190 (O_2190,N_29649,N_29594);
and UO_2191 (O_2191,N_29764,N_29629);
and UO_2192 (O_2192,N_29959,N_29649);
nand UO_2193 (O_2193,N_29833,N_29961);
and UO_2194 (O_2194,N_29678,N_29783);
or UO_2195 (O_2195,N_29858,N_29509);
or UO_2196 (O_2196,N_29882,N_29958);
or UO_2197 (O_2197,N_29915,N_29708);
or UO_2198 (O_2198,N_29851,N_29541);
or UO_2199 (O_2199,N_29552,N_29933);
nor UO_2200 (O_2200,N_29635,N_29997);
nand UO_2201 (O_2201,N_29510,N_29524);
or UO_2202 (O_2202,N_29677,N_29880);
nor UO_2203 (O_2203,N_29691,N_29648);
xor UO_2204 (O_2204,N_29797,N_29905);
and UO_2205 (O_2205,N_29548,N_29969);
nand UO_2206 (O_2206,N_29952,N_29863);
xnor UO_2207 (O_2207,N_29937,N_29621);
or UO_2208 (O_2208,N_29658,N_29638);
or UO_2209 (O_2209,N_29523,N_29550);
nor UO_2210 (O_2210,N_29710,N_29981);
and UO_2211 (O_2211,N_29542,N_29724);
xor UO_2212 (O_2212,N_29649,N_29838);
or UO_2213 (O_2213,N_29646,N_29532);
or UO_2214 (O_2214,N_29943,N_29794);
and UO_2215 (O_2215,N_29958,N_29891);
and UO_2216 (O_2216,N_29524,N_29777);
and UO_2217 (O_2217,N_29973,N_29544);
and UO_2218 (O_2218,N_29558,N_29532);
and UO_2219 (O_2219,N_29984,N_29917);
nand UO_2220 (O_2220,N_29944,N_29748);
nor UO_2221 (O_2221,N_29975,N_29771);
and UO_2222 (O_2222,N_29803,N_29918);
nand UO_2223 (O_2223,N_29709,N_29916);
or UO_2224 (O_2224,N_29956,N_29756);
nor UO_2225 (O_2225,N_29842,N_29513);
and UO_2226 (O_2226,N_29794,N_29804);
nor UO_2227 (O_2227,N_29698,N_29602);
and UO_2228 (O_2228,N_29793,N_29655);
and UO_2229 (O_2229,N_29586,N_29541);
xnor UO_2230 (O_2230,N_29845,N_29675);
and UO_2231 (O_2231,N_29723,N_29709);
xor UO_2232 (O_2232,N_29955,N_29954);
and UO_2233 (O_2233,N_29851,N_29728);
nand UO_2234 (O_2234,N_29922,N_29986);
or UO_2235 (O_2235,N_29848,N_29795);
nor UO_2236 (O_2236,N_29580,N_29928);
and UO_2237 (O_2237,N_29908,N_29821);
xnor UO_2238 (O_2238,N_29994,N_29796);
xor UO_2239 (O_2239,N_29980,N_29819);
nor UO_2240 (O_2240,N_29951,N_29608);
or UO_2241 (O_2241,N_29845,N_29627);
nand UO_2242 (O_2242,N_29740,N_29962);
xnor UO_2243 (O_2243,N_29641,N_29746);
and UO_2244 (O_2244,N_29515,N_29767);
and UO_2245 (O_2245,N_29849,N_29831);
xnor UO_2246 (O_2246,N_29748,N_29526);
and UO_2247 (O_2247,N_29922,N_29790);
nand UO_2248 (O_2248,N_29860,N_29692);
and UO_2249 (O_2249,N_29959,N_29928);
nor UO_2250 (O_2250,N_29886,N_29861);
nand UO_2251 (O_2251,N_29553,N_29751);
nand UO_2252 (O_2252,N_29756,N_29988);
nor UO_2253 (O_2253,N_29904,N_29546);
xnor UO_2254 (O_2254,N_29983,N_29532);
nand UO_2255 (O_2255,N_29512,N_29569);
or UO_2256 (O_2256,N_29921,N_29518);
nor UO_2257 (O_2257,N_29987,N_29985);
or UO_2258 (O_2258,N_29532,N_29801);
nor UO_2259 (O_2259,N_29982,N_29874);
and UO_2260 (O_2260,N_29624,N_29749);
and UO_2261 (O_2261,N_29569,N_29712);
and UO_2262 (O_2262,N_29986,N_29612);
nand UO_2263 (O_2263,N_29527,N_29677);
xor UO_2264 (O_2264,N_29854,N_29572);
nor UO_2265 (O_2265,N_29661,N_29736);
nand UO_2266 (O_2266,N_29724,N_29910);
xnor UO_2267 (O_2267,N_29651,N_29619);
nor UO_2268 (O_2268,N_29834,N_29620);
and UO_2269 (O_2269,N_29502,N_29900);
and UO_2270 (O_2270,N_29527,N_29668);
nor UO_2271 (O_2271,N_29568,N_29839);
xor UO_2272 (O_2272,N_29823,N_29521);
nand UO_2273 (O_2273,N_29922,N_29676);
nand UO_2274 (O_2274,N_29637,N_29723);
xnor UO_2275 (O_2275,N_29856,N_29979);
and UO_2276 (O_2276,N_29961,N_29583);
or UO_2277 (O_2277,N_29985,N_29858);
or UO_2278 (O_2278,N_29549,N_29652);
nor UO_2279 (O_2279,N_29686,N_29879);
nand UO_2280 (O_2280,N_29514,N_29698);
nor UO_2281 (O_2281,N_29561,N_29991);
xnor UO_2282 (O_2282,N_29780,N_29753);
and UO_2283 (O_2283,N_29619,N_29530);
and UO_2284 (O_2284,N_29999,N_29643);
and UO_2285 (O_2285,N_29662,N_29843);
and UO_2286 (O_2286,N_29615,N_29886);
and UO_2287 (O_2287,N_29822,N_29813);
and UO_2288 (O_2288,N_29731,N_29694);
and UO_2289 (O_2289,N_29580,N_29501);
nor UO_2290 (O_2290,N_29957,N_29504);
nor UO_2291 (O_2291,N_29855,N_29564);
nor UO_2292 (O_2292,N_29766,N_29862);
xor UO_2293 (O_2293,N_29733,N_29581);
nor UO_2294 (O_2294,N_29623,N_29895);
nand UO_2295 (O_2295,N_29710,N_29644);
xor UO_2296 (O_2296,N_29570,N_29906);
or UO_2297 (O_2297,N_29690,N_29925);
nor UO_2298 (O_2298,N_29638,N_29679);
and UO_2299 (O_2299,N_29925,N_29741);
or UO_2300 (O_2300,N_29966,N_29668);
nor UO_2301 (O_2301,N_29944,N_29976);
nor UO_2302 (O_2302,N_29899,N_29552);
xor UO_2303 (O_2303,N_29725,N_29910);
or UO_2304 (O_2304,N_29632,N_29957);
nand UO_2305 (O_2305,N_29715,N_29817);
and UO_2306 (O_2306,N_29758,N_29678);
or UO_2307 (O_2307,N_29517,N_29585);
or UO_2308 (O_2308,N_29660,N_29661);
nand UO_2309 (O_2309,N_29822,N_29572);
and UO_2310 (O_2310,N_29727,N_29932);
nor UO_2311 (O_2311,N_29756,N_29675);
or UO_2312 (O_2312,N_29552,N_29921);
and UO_2313 (O_2313,N_29525,N_29646);
nor UO_2314 (O_2314,N_29719,N_29778);
or UO_2315 (O_2315,N_29966,N_29582);
nor UO_2316 (O_2316,N_29511,N_29727);
nand UO_2317 (O_2317,N_29947,N_29895);
or UO_2318 (O_2318,N_29985,N_29854);
nand UO_2319 (O_2319,N_29728,N_29785);
nand UO_2320 (O_2320,N_29661,N_29707);
and UO_2321 (O_2321,N_29739,N_29837);
xor UO_2322 (O_2322,N_29713,N_29516);
nor UO_2323 (O_2323,N_29753,N_29979);
xnor UO_2324 (O_2324,N_29952,N_29515);
nor UO_2325 (O_2325,N_29508,N_29795);
or UO_2326 (O_2326,N_29551,N_29571);
or UO_2327 (O_2327,N_29515,N_29935);
nor UO_2328 (O_2328,N_29868,N_29674);
or UO_2329 (O_2329,N_29915,N_29596);
xnor UO_2330 (O_2330,N_29800,N_29804);
or UO_2331 (O_2331,N_29722,N_29964);
nor UO_2332 (O_2332,N_29900,N_29627);
nor UO_2333 (O_2333,N_29892,N_29860);
xor UO_2334 (O_2334,N_29710,N_29787);
nand UO_2335 (O_2335,N_29743,N_29631);
or UO_2336 (O_2336,N_29727,N_29505);
xor UO_2337 (O_2337,N_29571,N_29908);
nand UO_2338 (O_2338,N_29577,N_29896);
or UO_2339 (O_2339,N_29603,N_29995);
or UO_2340 (O_2340,N_29657,N_29771);
xnor UO_2341 (O_2341,N_29896,N_29964);
nand UO_2342 (O_2342,N_29912,N_29977);
nand UO_2343 (O_2343,N_29600,N_29527);
nor UO_2344 (O_2344,N_29685,N_29715);
nand UO_2345 (O_2345,N_29827,N_29724);
xnor UO_2346 (O_2346,N_29924,N_29562);
xor UO_2347 (O_2347,N_29849,N_29788);
nand UO_2348 (O_2348,N_29704,N_29988);
nand UO_2349 (O_2349,N_29962,N_29701);
nand UO_2350 (O_2350,N_29913,N_29880);
xnor UO_2351 (O_2351,N_29722,N_29562);
or UO_2352 (O_2352,N_29580,N_29960);
xnor UO_2353 (O_2353,N_29941,N_29957);
nor UO_2354 (O_2354,N_29796,N_29648);
or UO_2355 (O_2355,N_29536,N_29770);
nor UO_2356 (O_2356,N_29787,N_29825);
and UO_2357 (O_2357,N_29543,N_29608);
or UO_2358 (O_2358,N_29633,N_29711);
nor UO_2359 (O_2359,N_29836,N_29918);
nor UO_2360 (O_2360,N_29900,N_29839);
or UO_2361 (O_2361,N_29661,N_29940);
nand UO_2362 (O_2362,N_29930,N_29622);
nand UO_2363 (O_2363,N_29968,N_29549);
xor UO_2364 (O_2364,N_29949,N_29694);
or UO_2365 (O_2365,N_29581,N_29511);
xnor UO_2366 (O_2366,N_29921,N_29618);
and UO_2367 (O_2367,N_29833,N_29596);
and UO_2368 (O_2368,N_29678,N_29593);
nor UO_2369 (O_2369,N_29744,N_29615);
nand UO_2370 (O_2370,N_29728,N_29749);
xor UO_2371 (O_2371,N_29521,N_29719);
nand UO_2372 (O_2372,N_29981,N_29647);
and UO_2373 (O_2373,N_29949,N_29990);
nor UO_2374 (O_2374,N_29820,N_29926);
xnor UO_2375 (O_2375,N_29952,N_29735);
and UO_2376 (O_2376,N_29927,N_29712);
xor UO_2377 (O_2377,N_29900,N_29729);
or UO_2378 (O_2378,N_29961,N_29603);
or UO_2379 (O_2379,N_29990,N_29964);
xor UO_2380 (O_2380,N_29742,N_29957);
nand UO_2381 (O_2381,N_29588,N_29540);
xor UO_2382 (O_2382,N_29657,N_29998);
or UO_2383 (O_2383,N_29579,N_29612);
xor UO_2384 (O_2384,N_29552,N_29888);
nand UO_2385 (O_2385,N_29712,N_29711);
nand UO_2386 (O_2386,N_29873,N_29767);
nand UO_2387 (O_2387,N_29574,N_29806);
nor UO_2388 (O_2388,N_29751,N_29984);
or UO_2389 (O_2389,N_29826,N_29727);
nor UO_2390 (O_2390,N_29648,N_29649);
xnor UO_2391 (O_2391,N_29673,N_29781);
or UO_2392 (O_2392,N_29621,N_29702);
xnor UO_2393 (O_2393,N_29719,N_29532);
nor UO_2394 (O_2394,N_29667,N_29648);
nor UO_2395 (O_2395,N_29685,N_29831);
and UO_2396 (O_2396,N_29715,N_29874);
xor UO_2397 (O_2397,N_29755,N_29854);
nor UO_2398 (O_2398,N_29667,N_29626);
and UO_2399 (O_2399,N_29834,N_29993);
and UO_2400 (O_2400,N_29856,N_29570);
nor UO_2401 (O_2401,N_29546,N_29633);
xor UO_2402 (O_2402,N_29783,N_29809);
or UO_2403 (O_2403,N_29584,N_29795);
and UO_2404 (O_2404,N_29760,N_29721);
and UO_2405 (O_2405,N_29641,N_29652);
or UO_2406 (O_2406,N_29942,N_29685);
and UO_2407 (O_2407,N_29945,N_29532);
xnor UO_2408 (O_2408,N_29915,N_29626);
or UO_2409 (O_2409,N_29854,N_29776);
nor UO_2410 (O_2410,N_29616,N_29877);
or UO_2411 (O_2411,N_29717,N_29746);
nor UO_2412 (O_2412,N_29912,N_29791);
nor UO_2413 (O_2413,N_29748,N_29798);
xnor UO_2414 (O_2414,N_29517,N_29889);
and UO_2415 (O_2415,N_29774,N_29559);
nor UO_2416 (O_2416,N_29505,N_29698);
nand UO_2417 (O_2417,N_29614,N_29610);
or UO_2418 (O_2418,N_29718,N_29624);
or UO_2419 (O_2419,N_29761,N_29683);
or UO_2420 (O_2420,N_29958,N_29769);
and UO_2421 (O_2421,N_29837,N_29703);
xor UO_2422 (O_2422,N_29800,N_29844);
xnor UO_2423 (O_2423,N_29947,N_29800);
nor UO_2424 (O_2424,N_29812,N_29630);
xnor UO_2425 (O_2425,N_29916,N_29937);
nand UO_2426 (O_2426,N_29883,N_29896);
xnor UO_2427 (O_2427,N_29886,N_29664);
nor UO_2428 (O_2428,N_29504,N_29630);
or UO_2429 (O_2429,N_29645,N_29729);
xnor UO_2430 (O_2430,N_29659,N_29992);
or UO_2431 (O_2431,N_29571,N_29693);
or UO_2432 (O_2432,N_29981,N_29727);
or UO_2433 (O_2433,N_29771,N_29770);
xor UO_2434 (O_2434,N_29604,N_29936);
nand UO_2435 (O_2435,N_29877,N_29972);
xnor UO_2436 (O_2436,N_29948,N_29711);
and UO_2437 (O_2437,N_29720,N_29921);
and UO_2438 (O_2438,N_29990,N_29609);
xor UO_2439 (O_2439,N_29611,N_29533);
nand UO_2440 (O_2440,N_29548,N_29522);
or UO_2441 (O_2441,N_29526,N_29500);
or UO_2442 (O_2442,N_29836,N_29726);
nor UO_2443 (O_2443,N_29678,N_29719);
or UO_2444 (O_2444,N_29556,N_29905);
or UO_2445 (O_2445,N_29839,N_29818);
and UO_2446 (O_2446,N_29875,N_29633);
and UO_2447 (O_2447,N_29800,N_29670);
or UO_2448 (O_2448,N_29656,N_29995);
nand UO_2449 (O_2449,N_29599,N_29761);
nand UO_2450 (O_2450,N_29877,N_29758);
and UO_2451 (O_2451,N_29741,N_29546);
nand UO_2452 (O_2452,N_29835,N_29613);
and UO_2453 (O_2453,N_29990,N_29717);
nor UO_2454 (O_2454,N_29604,N_29687);
or UO_2455 (O_2455,N_29852,N_29581);
xor UO_2456 (O_2456,N_29628,N_29931);
nor UO_2457 (O_2457,N_29724,N_29769);
nor UO_2458 (O_2458,N_29925,N_29944);
and UO_2459 (O_2459,N_29546,N_29985);
nand UO_2460 (O_2460,N_29782,N_29856);
xnor UO_2461 (O_2461,N_29781,N_29862);
nor UO_2462 (O_2462,N_29936,N_29912);
xor UO_2463 (O_2463,N_29753,N_29911);
and UO_2464 (O_2464,N_29911,N_29873);
nand UO_2465 (O_2465,N_29775,N_29817);
and UO_2466 (O_2466,N_29695,N_29673);
xnor UO_2467 (O_2467,N_29825,N_29582);
and UO_2468 (O_2468,N_29861,N_29942);
nor UO_2469 (O_2469,N_29802,N_29958);
and UO_2470 (O_2470,N_29916,N_29531);
nand UO_2471 (O_2471,N_29512,N_29872);
xnor UO_2472 (O_2472,N_29704,N_29706);
nor UO_2473 (O_2473,N_29759,N_29959);
and UO_2474 (O_2474,N_29864,N_29812);
and UO_2475 (O_2475,N_29605,N_29796);
and UO_2476 (O_2476,N_29704,N_29628);
nand UO_2477 (O_2477,N_29918,N_29987);
and UO_2478 (O_2478,N_29851,N_29768);
nor UO_2479 (O_2479,N_29960,N_29511);
and UO_2480 (O_2480,N_29594,N_29630);
nor UO_2481 (O_2481,N_29762,N_29764);
nand UO_2482 (O_2482,N_29750,N_29931);
nand UO_2483 (O_2483,N_29754,N_29763);
and UO_2484 (O_2484,N_29579,N_29688);
xnor UO_2485 (O_2485,N_29875,N_29700);
xor UO_2486 (O_2486,N_29572,N_29701);
xor UO_2487 (O_2487,N_29858,N_29724);
nand UO_2488 (O_2488,N_29653,N_29988);
xor UO_2489 (O_2489,N_29537,N_29592);
nor UO_2490 (O_2490,N_29790,N_29965);
xnor UO_2491 (O_2491,N_29721,N_29888);
and UO_2492 (O_2492,N_29514,N_29502);
nand UO_2493 (O_2493,N_29616,N_29929);
and UO_2494 (O_2494,N_29947,N_29759);
xnor UO_2495 (O_2495,N_29647,N_29599);
nand UO_2496 (O_2496,N_29829,N_29686);
xnor UO_2497 (O_2497,N_29741,N_29517);
or UO_2498 (O_2498,N_29794,N_29896);
or UO_2499 (O_2499,N_29505,N_29965);
and UO_2500 (O_2500,N_29718,N_29951);
or UO_2501 (O_2501,N_29788,N_29948);
and UO_2502 (O_2502,N_29612,N_29863);
xnor UO_2503 (O_2503,N_29544,N_29598);
and UO_2504 (O_2504,N_29874,N_29902);
nor UO_2505 (O_2505,N_29919,N_29875);
nand UO_2506 (O_2506,N_29804,N_29820);
or UO_2507 (O_2507,N_29602,N_29603);
or UO_2508 (O_2508,N_29686,N_29685);
xor UO_2509 (O_2509,N_29625,N_29569);
nand UO_2510 (O_2510,N_29634,N_29568);
xnor UO_2511 (O_2511,N_29735,N_29772);
nand UO_2512 (O_2512,N_29538,N_29972);
nand UO_2513 (O_2513,N_29951,N_29795);
nor UO_2514 (O_2514,N_29561,N_29597);
or UO_2515 (O_2515,N_29673,N_29913);
or UO_2516 (O_2516,N_29780,N_29748);
and UO_2517 (O_2517,N_29572,N_29987);
and UO_2518 (O_2518,N_29721,N_29718);
nand UO_2519 (O_2519,N_29770,N_29847);
and UO_2520 (O_2520,N_29961,N_29517);
xor UO_2521 (O_2521,N_29988,N_29829);
xor UO_2522 (O_2522,N_29881,N_29532);
or UO_2523 (O_2523,N_29654,N_29737);
and UO_2524 (O_2524,N_29727,N_29895);
nor UO_2525 (O_2525,N_29730,N_29981);
and UO_2526 (O_2526,N_29839,N_29736);
nand UO_2527 (O_2527,N_29748,N_29533);
or UO_2528 (O_2528,N_29790,N_29993);
or UO_2529 (O_2529,N_29870,N_29570);
or UO_2530 (O_2530,N_29560,N_29970);
nor UO_2531 (O_2531,N_29769,N_29505);
xor UO_2532 (O_2532,N_29660,N_29789);
or UO_2533 (O_2533,N_29602,N_29640);
and UO_2534 (O_2534,N_29955,N_29878);
or UO_2535 (O_2535,N_29732,N_29658);
and UO_2536 (O_2536,N_29584,N_29594);
or UO_2537 (O_2537,N_29771,N_29747);
or UO_2538 (O_2538,N_29920,N_29727);
or UO_2539 (O_2539,N_29844,N_29550);
nand UO_2540 (O_2540,N_29900,N_29688);
or UO_2541 (O_2541,N_29972,N_29796);
nand UO_2542 (O_2542,N_29549,N_29683);
or UO_2543 (O_2543,N_29856,N_29696);
and UO_2544 (O_2544,N_29668,N_29705);
or UO_2545 (O_2545,N_29657,N_29675);
nor UO_2546 (O_2546,N_29532,N_29939);
or UO_2547 (O_2547,N_29696,N_29785);
or UO_2548 (O_2548,N_29756,N_29806);
or UO_2549 (O_2549,N_29854,N_29509);
and UO_2550 (O_2550,N_29597,N_29610);
nand UO_2551 (O_2551,N_29676,N_29707);
or UO_2552 (O_2552,N_29816,N_29715);
xnor UO_2553 (O_2553,N_29581,N_29531);
nand UO_2554 (O_2554,N_29690,N_29955);
and UO_2555 (O_2555,N_29822,N_29568);
and UO_2556 (O_2556,N_29764,N_29667);
nor UO_2557 (O_2557,N_29791,N_29737);
nand UO_2558 (O_2558,N_29527,N_29643);
or UO_2559 (O_2559,N_29513,N_29565);
nand UO_2560 (O_2560,N_29834,N_29886);
nand UO_2561 (O_2561,N_29796,N_29724);
nor UO_2562 (O_2562,N_29609,N_29580);
and UO_2563 (O_2563,N_29640,N_29652);
nor UO_2564 (O_2564,N_29992,N_29556);
xor UO_2565 (O_2565,N_29775,N_29820);
xor UO_2566 (O_2566,N_29751,N_29589);
nand UO_2567 (O_2567,N_29947,N_29705);
or UO_2568 (O_2568,N_29741,N_29902);
nor UO_2569 (O_2569,N_29682,N_29527);
nand UO_2570 (O_2570,N_29521,N_29503);
xnor UO_2571 (O_2571,N_29720,N_29888);
nor UO_2572 (O_2572,N_29678,N_29744);
xnor UO_2573 (O_2573,N_29987,N_29560);
nor UO_2574 (O_2574,N_29946,N_29864);
xor UO_2575 (O_2575,N_29887,N_29844);
and UO_2576 (O_2576,N_29505,N_29647);
nand UO_2577 (O_2577,N_29733,N_29509);
and UO_2578 (O_2578,N_29691,N_29531);
xnor UO_2579 (O_2579,N_29851,N_29676);
xnor UO_2580 (O_2580,N_29785,N_29888);
nand UO_2581 (O_2581,N_29631,N_29949);
and UO_2582 (O_2582,N_29511,N_29624);
or UO_2583 (O_2583,N_29553,N_29615);
xnor UO_2584 (O_2584,N_29775,N_29583);
or UO_2585 (O_2585,N_29609,N_29867);
xnor UO_2586 (O_2586,N_29682,N_29940);
xor UO_2587 (O_2587,N_29554,N_29552);
and UO_2588 (O_2588,N_29943,N_29731);
or UO_2589 (O_2589,N_29503,N_29832);
nand UO_2590 (O_2590,N_29806,N_29904);
or UO_2591 (O_2591,N_29642,N_29705);
and UO_2592 (O_2592,N_29825,N_29717);
and UO_2593 (O_2593,N_29807,N_29905);
nor UO_2594 (O_2594,N_29949,N_29868);
or UO_2595 (O_2595,N_29711,N_29907);
nand UO_2596 (O_2596,N_29981,N_29964);
xnor UO_2597 (O_2597,N_29524,N_29815);
and UO_2598 (O_2598,N_29900,N_29537);
nand UO_2599 (O_2599,N_29961,N_29596);
and UO_2600 (O_2600,N_29769,N_29644);
nand UO_2601 (O_2601,N_29609,N_29870);
and UO_2602 (O_2602,N_29849,N_29656);
and UO_2603 (O_2603,N_29761,N_29764);
or UO_2604 (O_2604,N_29860,N_29651);
nor UO_2605 (O_2605,N_29939,N_29666);
or UO_2606 (O_2606,N_29822,N_29681);
nor UO_2607 (O_2607,N_29602,N_29574);
or UO_2608 (O_2608,N_29984,N_29932);
and UO_2609 (O_2609,N_29622,N_29910);
xnor UO_2610 (O_2610,N_29625,N_29894);
nand UO_2611 (O_2611,N_29862,N_29933);
xnor UO_2612 (O_2612,N_29590,N_29932);
and UO_2613 (O_2613,N_29674,N_29775);
xor UO_2614 (O_2614,N_29871,N_29858);
or UO_2615 (O_2615,N_29945,N_29989);
nor UO_2616 (O_2616,N_29931,N_29591);
xnor UO_2617 (O_2617,N_29846,N_29516);
xnor UO_2618 (O_2618,N_29677,N_29621);
and UO_2619 (O_2619,N_29654,N_29806);
xor UO_2620 (O_2620,N_29658,N_29831);
and UO_2621 (O_2621,N_29502,N_29876);
nor UO_2622 (O_2622,N_29933,N_29622);
nand UO_2623 (O_2623,N_29866,N_29533);
nand UO_2624 (O_2624,N_29523,N_29884);
and UO_2625 (O_2625,N_29776,N_29563);
nand UO_2626 (O_2626,N_29756,N_29717);
nand UO_2627 (O_2627,N_29938,N_29701);
nand UO_2628 (O_2628,N_29830,N_29620);
nand UO_2629 (O_2629,N_29724,N_29770);
or UO_2630 (O_2630,N_29633,N_29784);
or UO_2631 (O_2631,N_29726,N_29754);
xor UO_2632 (O_2632,N_29672,N_29611);
or UO_2633 (O_2633,N_29639,N_29863);
or UO_2634 (O_2634,N_29982,N_29861);
nand UO_2635 (O_2635,N_29899,N_29607);
and UO_2636 (O_2636,N_29767,N_29752);
nor UO_2637 (O_2637,N_29674,N_29671);
or UO_2638 (O_2638,N_29760,N_29832);
and UO_2639 (O_2639,N_29656,N_29886);
nor UO_2640 (O_2640,N_29831,N_29893);
and UO_2641 (O_2641,N_29765,N_29701);
or UO_2642 (O_2642,N_29564,N_29887);
xor UO_2643 (O_2643,N_29525,N_29685);
nor UO_2644 (O_2644,N_29898,N_29941);
xnor UO_2645 (O_2645,N_29695,N_29710);
xnor UO_2646 (O_2646,N_29548,N_29632);
nand UO_2647 (O_2647,N_29865,N_29777);
and UO_2648 (O_2648,N_29861,N_29654);
and UO_2649 (O_2649,N_29624,N_29735);
or UO_2650 (O_2650,N_29566,N_29967);
and UO_2651 (O_2651,N_29827,N_29954);
or UO_2652 (O_2652,N_29605,N_29552);
nor UO_2653 (O_2653,N_29875,N_29959);
xor UO_2654 (O_2654,N_29867,N_29668);
nor UO_2655 (O_2655,N_29836,N_29556);
and UO_2656 (O_2656,N_29599,N_29508);
nor UO_2657 (O_2657,N_29880,N_29817);
nand UO_2658 (O_2658,N_29927,N_29781);
or UO_2659 (O_2659,N_29748,N_29583);
xnor UO_2660 (O_2660,N_29560,N_29575);
and UO_2661 (O_2661,N_29590,N_29866);
xor UO_2662 (O_2662,N_29990,N_29732);
xnor UO_2663 (O_2663,N_29975,N_29951);
xor UO_2664 (O_2664,N_29920,N_29747);
nor UO_2665 (O_2665,N_29966,N_29877);
or UO_2666 (O_2666,N_29819,N_29812);
and UO_2667 (O_2667,N_29634,N_29868);
nor UO_2668 (O_2668,N_29908,N_29558);
xnor UO_2669 (O_2669,N_29709,N_29574);
xnor UO_2670 (O_2670,N_29601,N_29704);
and UO_2671 (O_2671,N_29560,N_29716);
or UO_2672 (O_2672,N_29541,N_29718);
or UO_2673 (O_2673,N_29923,N_29642);
nand UO_2674 (O_2674,N_29621,N_29604);
or UO_2675 (O_2675,N_29874,N_29876);
or UO_2676 (O_2676,N_29521,N_29842);
xor UO_2677 (O_2677,N_29545,N_29666);
xor UO_2678 (O_2678,N_29648,N_29531);
nand UO_2679 (O_2679,N_29554,N_29974);
or UO_2680 (O_2680,N_29742,N_29744);
nor UO_2681 (O_2681,N_29708,N_29765);
xor UO_2682 (O_2682,N_29777,N_29850);
xnor UO_2683 (O_2683,N_29837,N_29706);
and UO_2684 (O_2684,N_29795,N_29544);
nor UO_2685 (O_2685,N_29882,N_29911);
or UO_2686 (O_2686,N_29733,N_29560);
or UO_2687 (O_2687,N_29841,N_29666);
or UO_2688 (O_2688,N_29803,N_29947);
nand UO_2689 (O_2689,N_29734,N_29633);
and UO_2690 (O_2690,N_29631,N_29620);
xor UO_2691 (O_2691,N_29684,N_29725);
nor UO_2692 (O_2692,N_29986,N_29960);
and UO_2693 (O_2693,N_29749,N_29951);
xnor UO_2694 (O_2694,N_29760,N_29999);
nand UO_2695 (O_2695,N_29690,N_29726);
or UO_2696 (O_2696,N_29823,N_29539);
nand UO_2697 (O_2697,N_29661,N_29888);
nand UO_2698 (O_2698,N_29921,N_29500);
nand UO_2699 (O_2699,N_29778,N_29582);
nand UO_2700 (O_2700,N_29748,N_29541);
nor UO_2701 (O_2701,N_29852,N_29593);
nor UO_2702 (O_2702,N_29519,N_29518);
xnor UO_2703 (O_2703,N_29944,N_29687);
nand UO_2704 (O_2704,N_29915,N_29923);
xor UO_2705 (O_2705,N_29715,N_29791);
and UO_2706 (O_2706,N_29727,N_29948);
or UO_2707 (O_2707,N_29870,N_29721);
and UO_2708 (O_2708,N_29517,N_29998);
nor UO_2709 (O_2709,N_29998,N_29886);
or UO_2710 (O_2710,N_29746,N_29654);
or UO_2711 (O_2711,N_29702,N_29525);
and UO_2712 (O_2712,N_29504,N_29681);
nand UO_2713 (O_2713,N_29595,N_29784);
and UO_2714 (O_2714,N_29917,N_29689);
nor UO_2715 (O_2715,N_29687,N_29565);
nand UO_2716 (O_2716,N_29903,N_29580);
xnor UO_2717 (O_2717,N_29986,N_29845);
xnor UO_2718 (O_2718,N_29523,N_29584);
and UO_2719 (O_2719,N_29852,N_29899);
xor UO_2720 (O_2720,N_29889,N_29610);
and UO_2721 (O_2721,N_29991,N_29590);
or UO_2722 (O_2722,N_29683,N_29813);
nand UO_2723 (O_2723,N_29655,N_29770);
nand UO_2724 (O_2724,N_29567,N_29911);
nor UO_2725 (O_2725,N_29811,N_29603);
nor UO_2726 (O_2726,N_29791,N_29526);
xor UO_2727 (O_2727,N_29738,N_29546);
nand UO_2728 (O_2728,N_29746,N_29597);
nand UO_2729 (O_2729,N_29981,N_29677);
xor UO_2730 (O_2730,N_29777,N_29765);
nor UO_2731 (O_2731,N_29683,N_29561);
xor UO_2732 (O_2732,N_29627,N_29929);
nand UO_2733 (O_2733,N_29830,N_29695);
nor UO_2734 (O_2734,N_29784,N_29733);
xnor UO_2735 (O_2735,N_29625,N_29802);
xnor UO_2736 (O_2736,N_29913,N_29915);
nor UO_2737 (O_2737,N_29888,N_29504);
xor UO_2738 (O_2738,N_29650,N_29729);
nor UO_2739 (O_2739,N_29904,N_29548);
nand UO_2740 (O_2740,N_29697,N_29589);
or UO_2741 (O_2741,N_29504,N_29894);
xnor UO_2742 (O_2742,N_29809,N_29880);
nor UO_2743 (O_2743,N_29601,N_29513);
nand UO_2744 (O_2744,N_29890,N_29853);
nor UO_2745 (O_2745,N_29981,N_29969);
nand UO_2746 (O_2746,N_29980,N_29912);
nand UO_2747 (O_2747,N_29904,N_29909);
or UO_2748 (O_2748,N_29822,N_29570);
nand UO_2749 (O_2749,N_29799,N_29873);
xnor UO_2750 (O_2750,N_29787,N_29599);
or UO_2751 (O_2751,N_29704,N_29582);
xnor UO_2752 (O_2752,N_29621,N_29854);
nand UO_2753 (O_2753,N_29762,N_29607);
xnor UO_2754 (O_2754,N_29935,N_29927);
xor UO_2755 (O_2755,N_29522,N_29782);
or UO_2756 (O_2756,N_29855,N_29743);
and UO_2757 (O_2757,N_29908,N_29976);
or UO_2758 (O_2758,N_29681,N_29799);
nor UO_2759 (O_2759,N_29535,N_29684);
nand UO_2760 (O_2760,N_29848,N_29777);
and UO_2761 (O_2761,N_29675,N_29668);
xnor UO_2762 (O_2762,N_29708,N_29788);
nor UO_2763 (O_2763,N_29863,N_29573);
nor UO_2764 (O_2764,N_29864,N_29668);
and UO_2765 (O_2765,N_29927,N_29664);
nand UO_2766 (O_2766,N_29688,N_29979);
nand UO_2767 (O_2767,N_29907,N_29857);
nand UO_2768 (O_2768,N_29795,N_29965);
xnor UO_2769 (O_2769,N_29566,N_29712);
or UO_2770 (O_2770,N_29855,N_29505);
nor UO_2771 (O_2771,N_29940,N_29508);
and UO_2772 (O_2772,N_29809,N_29832);
nand UO_2773 (O_2773,N_29963,N_29572);
or UO_2774 (O_2774,N_29935,N_29886);
nand UO_2775 (O_2775,N_29640,N_29687);
nand UO_2776 (O_2776,N_29790,N_29860);
and UO_2777 (O_2777,N_29958,N_29698);
and UO_2778 (O_2778,N_29538,N_29633);
nand UO_2779 (O_2779,N_29902,N_29567);
nand UO_2780 (O_2780,N_29747,N_29794);
xor UO_2781 (O_2781,N_29698,N_29763);
or UO_2782 (O_2782,N_29634,N_29629);
and UO_2783 (O_2783,N_29615,N_29599);
or UO_2784 (O_2784,N_29968,N_29603);
nor UO_2785 (O_2785,N_29945,N_29826);
nand UO_2786 (O_2786,N_29819,N_29921);
or UO_2787 (O_2787,N_29537,N_29563);
nand UO_2788 (O_2788,N_29973,N_29951);
nand UO_2789 (O_2789,N_29835,N_29847);
or UO_2790 (O_2790,N_29869,N_29560);
and UO_2791 (O_2791,N_29742,N_29548);
xor UO_2792 (O_2792,N_29835,N_29795);
or UO_2793 (O_2793,N_29722,N_29721);
xnor UO_2794 (O_2794,N_29571,N_29633);
nor UO_2795 (O_2795,N_29892,N_29791);
nor UO_2796 (O_2796,N_29776,N_29802);
nand UO_2797 (O_2797,N_29544,N_29789);
and UO_2798 (O_2798,N_29855,N_29574);
nor UO_2799 (O_2799,N_29832,N_29925);
or UO_2800 (O_2800,N_29655,N_29521);
or UO_2801 (O_2801,N_29740,N_29635);
nand UO_2802 (O_2802,N_29737,N_29992);
or UO_2803 (O_2803,N_29860,N_29817);
and UO_2804 (O_2804,N_29705,N_29928);
nand UO_2805 (O_2805,N_29859,N_29662);
and UO_2806 (O_2806,N_29674,N_29903);
xnor UO_2807 (O_2807,N_29866,N_29701);
or UO_2808 (O_2808,N_29688,N_29697);
nor UO_2809 (O_2809,N_29903,N_29890);
nand UO_2810 (O_2810,N_29792,N_29658);
and UO_2811 (O_2811,N_29692,N_29635);
and UO_2812 (O_2812,N_29529,N_29969);
nand UO_2813 (O_2813,N_29654,N_29804);
nand UO_2814 (O_2814,N_29527,N_29877);
nand UO_2815 (O_2815,N_29636,N_29890);
nand UO_2816 (O_2816,N_29590,N_29595);
xnor UO_2817 (O_2817,N_29956,N_29731);
nor UO_2818 (O_2818,N_29624,N_29957);
and UO_2819 (O_2819,N_29533,N_29921);
nor UO_2820 (O_2820,N_29996,N_29983);
or UO_2821 (O_2821,N_29830,N_29797);
or UO_2822 (O_2822,N_29693,N_29690);
nand UO_2823 (O_2823,N_29706,N_29644);
xnor UO_2824 (O_2824,N_29560,N_29666);
nand UO_2825 (O_2825,N_29691,N_29974);
and UO_2826 (O_2826,N_29699,N_29968);
xor UO_2827 (O_2827,N_29817,N_29904);
nor UO_2828 (O_2828,N_29640,N_29503);
and UO_2829 (O_2829,N_29801,N_29717);
nand UO_2830 (O_2830,N_29657,N_29552);
nor UO_2831 (O_2831,N_29592,N_29834);
nor UO_2832 (O_2832,N_29526,N_29974);
or UO_2833 (O_2833,N_29658,N_29894);
nor UO_2834 (O_2834,N_29933,N_29902);
and UO_2835 (O_2835,N_29911,N_29730);
nand UO_2836 (O_2836,N_29824,N_29570);
nor UO_2837 (O_2837,N_29574,N_29617);
nand UO_2838 (O_2838,N_29609,N_29938);
nand UO_2839 (O_2839,N_29949,N_29542);
nor UO_2840 (O_2840,N_29839,N_29509);
xnor UO_2841 (O_2841,N_29928,N_29855);
nand UO_2842 (O_2842,N_29965,N_29688);
or UO_2843 (O_2843,N_29660,N_29714);
nand UO_2844 (O_2844,N_29695,N_29641);
nand UO_2845 (O_2845,N_29602,N_29646);
xor UO_2846 (O_2846,N_29777,N_29623);
and UO_2847 (O_2847,N_29657,N_29603);
nand UO_2848 (O_2848,N_29642,N_29905);
or UO_2849 (O_2849,N_29669,N_29680);
xnor UO_2850 (O_2850,N_29598,N_29566);
nor UO_2851 (O_2851,N_29704,N_29810);
and UO_2852 (O_2852,N_29813,N_29618);
and UO_2853 (O_2853,N_29935,N_29591);
nor UO_2854 (O_2854,N_29554,N_29861);
or UO_2855 (O_2855,N_29969,N_29905);
or UO_2856 (O_2856,N_29663,N_29793);
or UO_2857 (O_2857,N_29629,N_29808);
or UO_2858 (O_2858,N_29715,N_29597);
and UO_2859 (O_2859,N_29964,N_29969);
and UO_2860 (O_2860,N_29682,N_29644);
or UO_2861 (O_2861,N_29503,N_29746);
and UO_2862 (O_2862,N_29708,N_29771);
and UO_2863 (O_2863,N_29838,N_29535);
and UO_2864 (O_2864,N_29844,N_29979);
nand UO_2865 (O_2865,N_29694,N_29676);
xor UO_2866 (O_2866,N_29523,N_29746);
xor UO_2867 (O_2867,N_29664,N_29754);
xnor UO_2868 (O_2868,N_29881,N_29682);
nor UO_2869 (O_2869,N_29936,N_29580);
nand UO_2870 (O_2870,N_29957,N_29929);
and UO_2871 (O_2871,N_29522,N_29777);
nor UO_2872 (O_2872,N_29505,N_29898);
xor UO_2873 (O_2873,N_29999,N_29822);
nand UO_2874 (O_2874,N_29696,N_29872);
nor UO_2875 (O_2875,N_29971,N_29765);
nor UO_2876 (O_2876,N_29548,N_29574);
nand UO_2877 (O_2877,N_29713,N_29556);
nor UO_2878 (O_2878,N_29888,N_29973);
nor UO_2879 (O_2879,N_29761,N_29884);
nor UO_2880 (O_2880,N_29837,N_29986);
nor UO_2881 (O_2881,N_29900,N_29973);
xnor UO_2882 (O_2882,N_29613,N_29985);
nor UO_2883 (O_2883,N_29923,N_29545);
or UO_2884 (O_2884,N_29597,N_29575);
or UO_2885 (O_2885,N_29670,N_29811);
or UO_2886 (O_2886,N_29906,N_29876);
nand UO_2887 (O_2887,N_29898,N_29815);
xor UO_2888 (O_2888,N_29782,N_29943);
and UO_2889 (O_2889,N_29950,N_29949);
and UO_2890 (O_2890,N_29971,N_29741);
nor UO_2891 (O_2891,N_29906,N_29932);
nand UO_2892 (O_2892,N_29621,N_29582);
and UO_2893 (O_2893,N_29798,N_29890);
xor UO_2894 (O_2894,N_29592,N_29943);
nand UO_2895 (O_2895,N_29601,N_29509);
and UO_2896 (O_2896,N_29770,N_29686);
xor UO_2897 (O_2897,N_29776,N_29562);
xor UO_2898 (O_2898,N_29716,N_29513);
nand UO_2899 (O_2899,N_29615,N_29516);
nor UO_2900 (O_2900,N_29630,N_29600);
and UO_2901 (O_2901,N_29835,N_29650);
or UO_2902 (O_2902,N_29709,N_29787);
xnor UO_2903 (O_2903,N_29625,N_29542);
xor UO_2904 (O_2904,N_29553,N_29992);
nor UO_2905 (O_2905,N_29725,N_29617);
and UO_2906 (O_2906,N_29887,N_29674);
and UO_2907 (O_2907,N_29583,N_29508);
nor UO_2908 (O_2908,N_29721,N_29817);
xor UO_2909 (O_2909,N_29536,N_29983);
nand UO_2910 (O_2910,N_29765,N_29949);
or UO_2911 (O_2911,N_29667,N_29802);
nand UO_2912 (O_2912,N_29906,N_29870);
xor UO_2913 (O_2913,N_29621,N_29553);
and UO_2914 (O_2914,N_29944,N_29935);
nor UO_2915 (O_2915,N_29587,N_29964);
xnor UO_2916 (O_2916,N_29595,N_29655);
nand UO_2917 (O_2917,N_29577,N_29951);
xor UO_2918 (O_2918,N_29813,N_29656);
nor UO_2919 (O_2919,N_29786,N_29658);
or UO_2920 (O_2920,N_29944,N_29565);
or UO_2921 (O_2921,N_29518,N_29725);
or UO_2922 (O_2922,N_29883,N_29510);
xor UO_2923 (O_2923,N_29653,N_29581);
nand UO_2924 (O_2924,N_29577,N_29649);
nor UO_2925 (O_2925,N_29802,N_29646);
nand UO_2926 (O_2926,N_29559,N_29832);
nand UO_2927 (O_2927,N_29607,N_29873);
nor UO_2928 (O_2928,N_29875,N_29621);
and UO_2929 (O_2929,N_29968,N_29606);
nor UO_2930 (O_2930,N_29574,N_29799);
nand UO_2931 (O_2931,N_29530,N_29878);
nor UO_2932 (O_2932,N_29672,N_29658);
nand UO_2933 (O_2933,N_29665,N_29660);
and UO_2934 (O_2934,N_29948,N_29959);
and UO_2935 (O_2935,N_29643,N_29768);
nor UO_2936 (O_2936,N_29638,N_29705);
nor UO_2937 (O_2937,N_29521,N_29818);
or UO_2938 (O_2938,N_29701,N_29622);
nor UO_2939 (O_2939,N_29706,N_29765);
nand UO_2940 (O_2940,N_29956,N_29547);
nand UO_2941 (O_2941,N_29761,N_29546);
nor UO_2942 (O_2942,N_29617,N_29775);
nand UO_2943 (O_2943,N_29506,N_29835);
nand UO_2944 (O_2944,N_29846,N_29755);
xor UO_2945 (O_2945,N_29730,N_29857);
or UO_2946 (O_2946,N_29776,N_29886);
xor UO_2947 (O_2947,N_29758,N_29511);
nand UO_2948 (O_2948,N_29624,N_29955);
xor UO_2949 (O_2949,N_29502,N_29945);
nor UO_2950 (O_2950,N_29634,N_29605);
and UO_2951 (O_2951,N_29846,N_29664);
xor UO_2952 (O_2952,N_29615,N_29860);
nor UO_2953 (O_2953,N_29693,N_29686);
and UO_2954 (O_2954,N_29643,N_29720);
nand UO_2955 (O_2955,N_29836,N_29835);
nor UO_2956 (O_2956,N_29923,N_29503);
xor UO_2957 (O_2957,N_29839,N_29763);
nor UO_2958 (O_2958,N_29586,N_29624);
xor UO_2959 (O_2959,N_29500,N_29857);
xor UO_2960 (O_2960,N_29987,N_29993);
nand UO_2961 (O_2961,N_29509,N_29549);
nand UO_2962 (O_2962,N_29699,N_29920);
xor UO_2963 (O_2963,N_29988,N_29675);
and UO_2964 (O_2964,N_29684,N_29627);
and UO_2965 (O_2965,N_29966,N_29775);
or UO_2966 (O_2966,N_29882,N_29826);
or UO_2967 (O_2967,N_29563,N_29599);
nor UO_2968 (O_2968,N_29875,N_29909);
or UO_2969 (O_2969,N_29604,N_29918);
and UO_2970 (O_2970,N_29684,N_29792);
nor UO_2971 (O_2971,N_29657,N_29568);
and UO_2972 (O_2972,N_29710,N_29604);
nand UO_2973 (O_2973,N_29629,N_29893);
nor UO_2974 (O_2974,N_29621,N_29786);
nor UO_2975 (O_2975,N_29636,N_29641);
xnor UO_2976 (O_2976,N_29932,N_29516);
or UO_2977 (O_2977,N_29594,N_29707);
xor UO_2978 (O_2978,N_29722,N_29999);
nor UO_2979 (O_2979,N_29772,N_29705);
nor UO_2980 (O_2980,N_29545,N_29958);
or UO_2981 (O_2981,N_29685,N_29702);
or UO_2982 (O_2982,N_29773,N_29906);
nand UO_2983 (O_2983,N_29804,N_29591);
nor UO_2984 (O_2984,N_29795,N_29815);
and UO_2985 (O_2985,N_29586,N_29818);
and UO_2986 (O_2986,N_29523,N_29737);
xnor UO_2987 (O_2987,N_29812,N_29898);
nand UO_2988 (O_2988,N_29953,N_29672);
nor UO_2989 (O_2989,N_29859,N_29512);
nand UO_2990 (O_2990,N_29872,N_29846);
nand UO_2991 (O_2991,N_29715,N_29694);
and UO_2992 (O_2992,N_29636,N_29967);
xor UO_2993 (O_2993,N_29526,N_29649);
nand UO_2994 (O_2994,N_29892,N_29885);
and UO_2995 (O_2995,N_29835,N_29639);
xnor UO_2996 (O_2996,N_29662,N_29676);
nand UO_2997 (O_2997,N_29967,N_29735);
or UO_2998 (O_2998,N_29539,N_29826);
nor UO_2999 (O_2999,N_29922,N_29839);
or UO_3000 (O_3000,N_29873,N_29847);
or UO_3001 (O_3001,N_29789,N_29532);
xnor UO_3002 (O_3002,N_29653,N_29509);
nand UO_3003 (O_3003,N_29739,N_29645);
xnor UO_3004 (O_3004,N_29506,N_29539);
or UO_3005 (O_3005,N_29848,N_29845);
xnor UO_3006 (O_3006,N_29647,N_29651);
and UO_3007 (O_3007,N_29646,N_29830);
nor UO_3008 (O_3008,N_29835,N_29708);
nand UO_3009 (O_3009,N_29744,N_29982);
or UO_3010 (O_3010,N_29693,N_29544);
and UO_3011 (O_3011,N_29827,N_29774);
or UO_3012 (O_3012,N_29514,N_29603);
nor UO_3013 (O_3013,N_29518,N_29784);
nand UO_3014 (O_3014,N_29838,N_29734);
nor UO_3015 (O_3015,N_29709,N_29522);
xor UO_3016 (O_3016,N_29832,N_29563);
nor UO_3017 (O_3017,N_29954,N_29890);
nand UO_3018 (O_3018,N_29933,N_29861);
nand UO_3019 (O_3019,N_29884,N_29895);
nor UO_3020 (O_3020,N_29930,N_29905);
nor UO_3021 (O_3021,N_29997,N_29516);
nor UO_3022 (O_3022,N_29673,N_29627);
and UO_3023 (O_3023,N_29567,N_29779);
xor UO_3024 (O_3024,N_29784,N_29709);
xor UO_3025 (O_3025,N_29633,N_29685);
and UO_3026 (O_3026,N_29663,N_29826);
xnor UO_3027 (O_3027,N_29789,N_29850);
or UO_3028 (O_3028,N_29821,N_29549);
or UO_3029 (O_3029,N_29528,N_29899);
or UO_3030 (O_3030,N_29708,N_29868);
nand UO_3031 (O_3031,N_29885,N_29729);
nand UO_3032 (O_3032,N_29987,N_29594);
or UO_3033 (O_3033,N_29703,N_29956);
nor UO_3034 (O_3034,N_29786,N_29525);
and UO_3035 (O_3035,N_29974,N_29828);
nor UO_3036 (O_3036,N_29837,N_29992);
xnor UO_3037 (O_3037,N_29506,N_29776);
and UO_3038 (O_3038,N_29580,N_29871);
or UO_3039 (O_3039,N_29930,N_29802);
nand UO_3040 (O_3040,N_29704,N_29514);
nand UO_3041 (O_3041,N_29970,N_29993);
nor UO_3042 (O_3042,N_29970,N_29744);
or UO_3043 (O_3043,N_29682,N_29834);
nand UO_3044 (O_3044,N_29775,N_29645);
and UO_3045 (O_3045,N_29787,N_29687);
and UO_3046 (O_3046,N_29572,N_29834);
or UO_3047 (O_3047,N_29671,N_29896);
or UO_3048 (O_3048,N_29716,N_29675);
xor UO_3049 (O_3049,N_29757,N_29756);
nor UO_3050 (O_3050,N_29899,N_29734);
or UO_3051 (O_3051,N_29840,N_29590);
nor UO_3052 (O_3052,N_29817,N_29805);
nand UO_3053 (O_3053,N_29574,N_29545);
nand UO_3054 (O_3054,N_29617,N_29942);
xnor UO_3055 (O_3055,N_29761,N_29994);
or UO_3056 (O_3056,N_29993,N_29873);
or UO_3057 (O_3057,N_29513,N_29895);
nor UO_3058 (O_3058,N_29535,N_29721);
nand UO_3059 (O_3059,N_29581,N_29540);
xnor UO_3060 (O_3060,N_29713,N_29870);
or UO_3061 (O_3061,N_29620,N_29553);
and UO_3062 (O_3062,N_29977,N_29802);
xnor UO_3063 (O_3063,N_29911,N_29580);
and UO_3064 (O_3064,N_29651,N_29524);
and UO_3065 (O_3065,N_29999,N_29995);
nand UO_3066 (O_3066,N_29946,N_29765);
nor UO_3067 (O_3067,N_29889,N_29713);
and UO_3068 (O_3068,N_29648,N_29817);
and UO_3069 (O_3069,N_29820,N_29829);
or UO_3070 (O_3070,N_29755,N_29902);
or UO_3071 (O_3071,N_29820,N_29508);
and UO_3072 (O_3072,N_29991,N_29899);
nand UO_3073 (O_3073,N_29777,N_29946);
nor UO_3074 (O_3074,N_29789,N_29756);
and UO_3075 (O_3075,N_29865,N_29676);
nor UO_3076 (O_3076,N_29962,N_29544);
xor UO_3077 (O_3077,N_29675,N_29856);
and UO_3078 (O_3078,N_29767,N_29754);
nand UO_3079 (O_3079,N_29825,N_29905);
nor UO_3080 (O_3080,N_29836,N_29864);
or UO_3081 (O_3081,N_29953,N_29996);
or UO_3082 (O_3082,N_29679,N_29672);
nor UO_3083 (O_3083,N_29519,N_29884);
or UO_3084 (O_3084,N_29649,N_29576);
nand UO_3085 (O_3085,N_29739,N_29546);
and UO_3086 (O_3086,N_29879,N_29778);
and UO_3087 (O_3087,N_29591,N_29635);
or UO_3088 (O_3088,N_29826,N_29999);
nand UO_3089 (O_3089,N_29774,N_29878);
and UO_3090 (O_3090,N_29949,N_29902);
nor UO_3091 (O_3091,N_29779,N_29524);
xnor UO_3092 (O_3092,N_29953,N_29617);
nand UO_3093 (O_3093,N_29671,N_29803);
nand UO_3094 (O_3094,N_29748,N_29945);
and UO_3095 (O_3095,N_29959,N_29506);
and UO_3096 (O_3096,N_29604,N_29689);
nor UO_3097 (O_3097,N_29739,N_29771);
xor UO_3098 (O_3098,N_29768,N_29849);
and UO_3099 (O_3099,N_29860,N_29846);
xor UO_3100 (O_3100,N_29619,N_29941);
and UO_3101 (O_3101,N_29767,N_29867);
or UO_3102 (O_3102,N_29676,N_29593);
nor UO_3103 (O_3103,N_29802,N_29818);
nor UO_3104 (O_3104,N_29548,N_29630);
nand UO_3105 (O_3105,N_29538,N_29587);
nand UO_3106 (O_3106,N_29926,N_29652);
or UO_3107 (O_3107,N_29753,N_29956);
or UO_3108 (O_3108,N_29983,N_29614);
or UO_3109 (O_3109,N_29598,N_29580);
nor UO_3110 (O_3110,N_29617,N_29796);
or UO_3111 (O_3111,N_29897,N_29561);
nand UO_3112 (O_3112,N_29604,N_29950);
and UO_3113 (O_3113,N_29510,N_29836);
or UO_3114 (O_3114,N_29984,N_29764);
or UO_3115 (O_3115,N_29588,N_29679);
xnor UO_3116 (O_3116,N_29754,N_29925);
and UO_3117 (O_3117,N_29742,N_29597);
or UO_3118 (O_3118,N_29626,N_29650);
nor UO_3119 (O_3119,N_29795,N_29749);
or UO_3120 (O_3120,N_29617,N_29804);
xor UO_3121 (O_3121,N_29632,N_29931);
or UO_3122 (O_3122,N_29633,N_29950);
nor UO_3123 (O_3123,N_29830,N_29569);
nor UO_3124 (O_3124,N_29578,N_29888);
xnor UO_3125 (O_3125,N_29943,N_29999);
nor UO_3126 (O_3126,N_29551,N_29802);
nor UO_3127 (O_3127,N_29824,N_29605);
xnor UO_3128 (O_3128,N_29633,N_29541);
nor UO_3129 (O_3129,N_29908,N_29550);
nor UO_3130 (O_3130,N_29621,N_29515);
nand UO_3131 (O_3131,N_29980,N_29781);
xor UO_3132 (O_3132,N_29536,N_29677);
nand UO_3133 (O_3133,N_29996,N_29533);
nor UO_3134 (O_3134,N_29732,N_29641);
nor UO_3135 (O_3135,N_29657,N_29892);
xnor UO_3136 (O_3136,N_29771,N_29750);
xor UO_3137 (O_3137,N_29752,N_29561);
xor UO_3138 (O_3138,N_29587,N_29719);
nor UO_3139 (O_3139,N_29827,N_29831);
nor UO_3140 (O_3140,N_29984,N_29556);
nor UO_3141 (O_3141,N_29579,N_29939);
nand UO_3142 (O_3142,N_29916,N_29825);
xor UO_3143 (O_3143,N_29515,N_29603);
xnor UO_3144 (O_3144,N_29631,N_29704);
xnor UO_3145 (O_3145,N_29586,N_29559);
xor UO_3146 (O_3146,N_29506,N_29581);
nand UO_3147 (O_3147,N_29592,N_29736);
or UO_3148 (O_3148,N_29571,N_29613);
or UO_3149 (O_3149,N_29729,N_29911);
and UO_3150 (O_3150,N_29824,N_29779);
or UO_3151 (O_3151,N_29532,N_29734);
nand UO_3152 (O_3152,N_29868,N_29899);
or UO_3153 (O_3153,N_29760,N_29953);
xor UO_3154 (O_3154,N_29593,N_29774);
xnor UO_3155 (O_3155,N_29664,N_29655);
and UO_3156 (O_3156,N_29554,N_29593);
nor UO_3157 (O_3157,N_29704,N_29834);
and UO_3158 (O_3158,N_29714,N_29546);
nor UO_3159 (O_3159,N_29563,N_29755);
or UO_3160 (O_3160,N_29619,N_29723);
or UO_3161 (O_3161,N_29666,N_29542);
nor UO_3162 (O_3162,N_29589,N_29646);
nand UO_3163 (O_3163,N_29636,N_29587);
nor UO_3164 (O_3164,N_29850,N_29521);
xnor UO_3165 (O_3165,N_29829,N_29561);
or UO_3166 (O_3166,N_29890,N_29787);
nand UO_3167 (O_3167,N_29552,N_29622);
or UO_3168 (O_3168,N_29923,N_29816);
and UO_3169 (O_3169,N_29902,N_29960);
xnor UO_3170 (O_3170,N_29671,N_29751);
xnor UO_3171 (O_3171,N_29969,N_29658);
nand UO_3172 (O_3172,N_29749,N_29664);
nor UO_3173 (O_3173,N_29677,N_29661);
nor UO_3174 (O_3174,N_29561,N_29673);
or UO_3175 (O_3175,N_29762,N_29734);
or UO_3176 (O_3176,N_29895,N_29700);
nand UO_3177 (O_3177,N_29766,N_29637);
xnor UO_3178 (O_3178,N_29675,N_29959);
nand UO_3179 (O_3179,N_29933,N_29641);
xor UO_3180 (O_3180,N_29878,N_29935);
nor UO_3181 (O_3181,N_29853,N_29578);
or UO_3182 (O_3182,N_29968,N_29770);
xnor UO_3183 (O_3183,N_29723,N_29825);
or UO_3184 (O_3184,N_29504,N_29912);
nand UO_3185 (O_3185,N_29649,N_29937);
nor UO_3186 (O_3186,N_29982,N_29721);
xnor UO_3187 (O_3187,N_29755,N_29662);
or UO_3188 (O_3188,N_29641,N_29501);
and UO_3189 (O_3189,N_29826,N_29913);
nand UO_3190 (O_3190,N_29632,N_29866);
xnor UO_3191 (O_3191,N_29666,N_29503);
or UO_3192 (O_3192,N_29794,N_29967);
or UO_3193 (O_3193,N_29883,N_29643);
xnor UO_3194 (O_3194,N_29870,N_29951);
xnor UO_3195 (O_3195,N_29839,N_29867);
and UO_3196 (O_3196,N_29697,N_29926);
and UO_3197 (O_3197,N_29736,N_29843);
or UO_3198 (O_3198,N_29647,N_29898);
nand UO_3199 (O_3199,N_29775,N_29789);
xnor UO_3200 (O_3200,N_29992,N_29546);
and UO_3201 (O_3201,N_29658,N_29992);
and UO_3202 (O_3202,N_29941,N_29572);
nand UO_3203 (O_3203,N_29889,N_29701);
nand UO_3204 (O_3204,N_29700,N_29701);
nor UO_3205 (O_3205,N_29855,N_29838);
nor UO_3206 (O_3206,N_29563,N_29981);
and UO_3207 (O_3207,N_29680,N_29949);
and UO_3208 (O_3208,N_29563,N_29803);
nor UO_3209 (O_3209,N_29639,N_29677);
and UO_3210 (O_3210,N_29600,N_29736);
or UO_3211 (O_3211,N_29504,N_29537);
xor UO_3212 (O_3212,N_29785,N_29631);
nand UO_3213 (O_3213,N_29601,N_29912);
and UO_3214 (O_3214,N_29736,N_29774);
and UO_3215 (O_3215,N_29838,N_29755);
xnor UO_3216 (O_3216,N_29779,N_29773);
xor UO_3217 (O_3217,N_29773,N_29897);
and UO_3218 (O_3218,N_29532,N_29876);
and UO_3219 (O_3219,N_29881,N_29649);
or UO_3220 (O_3220,N_29518,N_29778);
nand UO_3221 (O_3221,N_29741,N_29654);
or UO_3222 (O_3222,N_29891,N_29914);
and UO_3223 (O_3223,N_29929,N_29855);
nand UO_3224 (O_3224,N_29741,N_29725);
nand UO_3225 (O_3225,N_29535,N_29792);
or UO_3226 (O_3226,N_29501,N_29864);
or UO_3227 (O_3227,N_29826,N_29626);
or UO_3228 (O_3228,N_29638,N_29596);
or UO_3229 (O_3229,N_29797,N_29815);
xor UO_3230 (O_3230,N_29739,N_29767);
or UO_3231 (O_3231,N_29636,N_29920);
or UO_3232 (O_3232,N_29709,N_29710);
and UO_3233 (O_3233,N_29881,N_29893);
nor UO_3234 (O_3234,N_29989,N_29800);
xor UO_3235 (O_3235,N_29965,N_29597);
and UO_3236 (O_3236,N_29637,N_29636);
and UO_3237 (O_3237,N_29874,N_29726);
xnor UO_3238 (O_3238,N_29633,N_29926);
nor UO_3239 (O_3239,N_29791,N_29792);
nor UO_3240 (O_3240,N_29598,N_29829);
or UO_3241 (O_3241,N_29571,N_29728);
nand UO_3242 (O_3242,N_29764,N_29610);
nor UO_3243 (O_3243,N_29758,N_29779);
nand UO_3244 (O_3244,N_29642,N_29842);
nor UO_3245 (O_3245,N_29563,N_29847);
and UO_3246 (O_3246,N_29542,N_29772);
nand UO_3247 (O_3247,N_29881,N_29578);
and UO_3248 (O_3248,N_29782,N_29819);
and UO_3249 (O_3249,N_29919,N_29873);
nand UO_3250 (O_3250,N_29791,N_29845);
or UO_3251 (O_3251,N_29500,N_29502);
nor UO_3252 (O_3252,N_29605,N_29883);
or UO_3253 (O_3253,N_29927,N_29513);
nor UO_3254 (O_3254,N_29552,N_29574);
nor UO_3255 (O_3255,N_29588,N_29898);
xor UO_3256 (O_3256,N_29814,N_29695);
nor UO_3257 (O_3257,N_29524,N_29528);
xnor UO_3258 (O_3258,N_29974,N_29769);
nor UO_3259 (O_3259,N_29656,N_29958);
or UO_3260 (O_3260,N_29532,N_29520);
xor UO_3261 (O_3261,N_29731,N_29852);
nand UO_3262 (O_3262,N_29651,N_29894);
xnor UO_3263 (O_3263,N_29559,N_29684);
xnor UO_3264 (O_3264,N_29781,N_29691);
and UO_3265 (O_3265,N_29953,N_29769);
xor UO_3266 (O_3266,N_29687,N_29533);
and UO_3267 (O_3267,N_29704,N_29993);
nand UO_3268 (O_3268,N_29932,N_29622);
nor UO_3269 (O_3269,N_29980,N_29975);
nand UO_3270 (O_3270,N_29781,N_29979);
or UO_3271 (O_3271,N_29995,N_29847);
nand UO_3272 (O_3272,N_29670,N_29569);
nor UO_3273 (O_3273,N_29751,N_29630);
xor UO_3274 (O_3274,N_29894,N_29984);
nand UO_3275 (O_3275,N_29631,N_29791);
nand UO_3276 (O_3276,N_29941,N_29626);
nor UO_3277 (O_3277,N_29806,N_29731);
or UO_3278 (O_3278,N_29892,N_29944);
nand UO_3279 (O_3279,N_29633,N_29602);
nand UO_3280 (O_3280,N_29615,N_29619);
xnor UO_3281 (O_3281,N_29605,N_29601);
nor UO_3282 (O_3282,N_29707,N_29983);
and UO_3283 (O_3283,N_29968,N_29812);
nor UO_3284 (O_3284,N_29549,N_29815);
nand UO_3285 (O_3285,N_29787,N_29949);
nand UO_3286 (O_3286,N_29821,N_29984);
xor UO_3287 (O_3287,N_29682,N_29550);
nand UO_3288 (O_3288,N_29998,N_29585);
or UO_3289 (O_3289,N_29702,N_29631);
and UO_3290 (O_3290,N_29930,N_29706);
nand UO_3291 (O_3291,N_29673,N_29516);
xor UO_3292 (O_3292,N_29818,N_29749);
nand UO_3293 (O_3293,N_29725,N_29507);
or UO_3294 (O_3294,N_29726,N_29760);
nand UO_3295 (O_3295,N_29907,N_29862);
or UO_3296 (O_3296,N_29725,N_29919);
xnor UO_3297 (O_3297,N_29511,N_29791);
xor UO_3298 (O_3298,N_29639,N_29752);
and UO_3299 (O_3299,N_29802,N_29554);
and UO_3300 (O_3300,N_29707,N_29884);
nand UO_3301 (O_3301,N_29971,N_29896);
nor UO_3302 (O_3302,N_29756,N_29536);
nand UO_3303 (O_3303,N_29937,N_29783);
xor UO_3304 (O_3304,N_29827,N_29653);
and UO_3305 (O_3305,N_29951,N_29558);
xor UO_3306 (O_3306,N_29835,N_29762);
and UO_3307 (O_3307,N_29956,N_29679);
xor UO_3308 (O_3308,N_29559,N_29549);
xor UO_3309 (O_3309,N_29602,N_29729);
and UO_3310 (O_3310,N_29649,N_29827);
or UO_3311 (O_3311,N_29769,N_29945);
nand UO_3312 (O_3312,N_29667,N_29732);
xor UO_3313 (O_3313,N_29860,N_29890);
nor UO_3314 (O_3314,N_29576,N_29636);
xor UO_3315 (O_3315,N_29813,N_29610);
nand UO_3316 (O_3316,N_29525,N_29810);
and UO_3317 (O_3317,N_29784,N_29828);
or UO_3318 (O_3318,N_29516,N_29558);
or UO_3319 (O_3319,N_29783,N_29501);
and UO_3320 (O_3320,N_29535,N_29564);
and UO_3321 (O_3321,N_29571,N_29780);
and UO_3322 (O_3322,N_29509,N_29719);
and UO_3323 (O_3323,N_29835,N_29591);
nor UO_3324 (O_3324,N_29583,N_29767);
nor UO_3325 (O_3325,N_29800,N_29520);
nor UO_3326 (O_3326,N_29870,N_29984);
or UO_3327 (O_3327,N_29691,N_29826);
or UO_3328 (O_3328,N_29607,N_29650);
xnor UO_3329 (O_3329,N_29685,N_29798);
and UO_3330 (O_3330,N_29696,N_29556);
xor UO_3331 (O_3331,N_29590,N_29628);
nor UO_3332 (O_3332,N_29821,N_29940);
nor UO_3333 (O_3333,N_29791,N_29886);
xnor UO_3334 (O_3334,N_29953,N_29888);
nand UO_3335 (O_3335,N_29724,N_29926);
and UO_3336 (O_3336,N_29681,N_29505);
or UO_3337 (O_3337,N_29526,N_29582);
nand UO_3338 (O_3338,N_29798,N_29636);
nor UO_3339 (O_3339,N_29990,N_29892);
and UO_3340 (O_3340,N_29525,N_29713);
or UO_3341 (O_3341,N_29842,N_29626);
or UO_3342 (O_3342,N_29742,N_29726);
xnor UO_3343 (O_3343,N_29528,N_29580);
nor UO_3344 (O_3344,N_29963,N_29697);
or UO_3345 (O_3345,N_29545,N_29554);
and UO_3346 (O_3346,N_29779,N_29551);
or UO_3347 (O_3347,N_29642,N_29662);
nor UO_3348 (O_3348,N_29695,N_29633);
nor UO_3349 (O_3349,N_29763,N_29944);
or UO_3350 (O_3350,N_29951,N_29729);
xor UO_3351 (O_3351,N_29871,N_29877);
nand UO_3352 (O_3352,N_29900,N_29763);
xor UO_3353 (O_3353,N_29583,N_29995);
nand UO_3354 (O_3354,N_29564,N_29959);
nand UO_3355 (O_3355,N_29776,N_29749);
nand UO_3356 (O_3356,N_29534,N_29721);
or UO_3357 (O_3357,N_29696,N_29564);
and UO_3358 (O_3358,N_29751,N_29883);
nor UO_3359 (O_3359,N_29908,N_29698);
nand UO_3360 (O_3360,N_29688,N_29560);
nor UO_3361 (O_3361,N_29584,N_29987);
and UO_3362 (O_3362,N_29637,N_29847);
xnor UO_3363 (O_3363,N_29839,N_29903);
or UO_3364 (O_3364,N_29781,N_29942);
or UO_3365 (O_3365,N_29816,N_29653);
and UO_3366 (O_3366,N_29762,N_29858);
and UO_3367 (O_3367,N_29866,N_29662);
nor UO_3368 (O_3368,N_29816,N_29777);
nand UO_3369 (O_3369,N_29678,N_29503);
and UO_3370 (O_3370,N_29843,N_29529);
and UO_3371 (O_3371,N_29701,N_29990);
and UO_3372 (O_3372,N_29690,N_29865);
and UO_3373 (O_3373,N_29764,N_29693);
xor UO_3374 (O_3374,N_29583,N_29584);
or UO_3375 (O_3375,N_29868,N_29589);
nor UO_3376 (O_3376,N_29781,N_29941);
xor UO_3377 (O_3377,N_29549,N_29808);
nand UO_3378 (O_3378,N_29508,N_29660);
or UO_3379 (O_3379,N_29518,N_29880);
xnor UO_3380 (O_3380,N_29715,N_29813);
xnor UO_3381 (O_3381,N_29992,N_29771);
or UO_3382 (O_3382,N_29633,N_29696);
xnor UO_3383 (O_3383,N_29604,N_29796);
nor UO_3384 (O_3384,N_29665,N_29805);
or UO_3385 (O_3385,N_29764,N_29791);
nand UO_3386 (O_3386,N_29998,N_29707);
and UO_3387 (O_3387,N_29596,N_29916);
xor UO_3388 (O_3388,N_29578,N_29747);
or UO_3389 (O_3389,N_29799,N_29773);
nand UO_3390 (O_3390,N_29562,N_29778);
and UO_3391 (O_3391,N_29762,N_29928);
nand UO_3392 (O_3392,N_29809,N_29753);
nor UO_3393 (O_3393,N_29709,N_29691);
nand UO_3394 (O_3394,N_29915,N_29957);
or UO_3395 (O_3395,N_29782,N_29919);
nand UO_3396 (O_3396,N_29820,N_29622);
nand UO_3397 (O_3397,N_29925,N_29549);
nand UO_3398 (O_3398,N_29676,N_29861);
or UO_3399 (O_3399,N_29556,N_29506);
xnor UO_3400 (O_3400,N_29822,N_29977);
and UO_3401 (O_3401,N_29912,N_29542);
and UO_3402 (O_3402,N_29849,N_29519);
xnor UO_3403 (O_3403,N_29627,N_29656);
nand UO_3404 (O_3404,N_29746,N_29860);
nor UO_3405 (O_3405,N_29910,N_29960);
nand UO_3406 (O_3406,N_29881,N_29598);
xnor UO_3407 (O_3407,N_29627,N_29807);
or UO_3408 (O_3408,N_29866,N_29745);
and UO_3409 (O_3409,N_29518,N_29575);
and UO_3410 (O_3410,N_29757,N_29905);
and UO_3411 (O_3411,N_29751,N_29896);
nor UO_3412 (O_3412,N_29608,N_29507);
or UO_3413 (O_3413,N_29569,N_29974);
nor UO_3414 (O_3414,N_29529,N_29507);
or UO_3415 (O_3415,N_29961,N_29601);
nor UO_3416 (O_3416,N_29979,N_29718);
and UO_3417 (O_3417,N_29795,N_29877);
nand UO_3418 (O_3418,N_29876,N_29974);
xor UO_3419 (O_3419,N_29758,N_29627);
nor UO_3420 (O_3420,N_29597,N_29887);
or UO_3421 (O_3421,N_29990,N_29509);
and UO_3422 (O_3422,N_29682,N_29568);
and UO_3423 (O_3423,N_29846,N_29661);
nand UO_3424 (O_3424,N_29922,N_29785);
xor UO_3425 (O_3425,N_29650,N_29856);
or UO_3426 (O_3426,N_29674,N_29991);
and UO_3427 (O_3427,N_29680,N_29988);
nand UO_3428 (O_3428,N_29672,N_29528);
nor UO_3429 (O_3429,N_29858,N_29884);
nand UO_3430 (O_3430,N_29548,N_29874);
or UO_3431 (O_3431,N_29856,N_29682);
and UO_3432 (O_3432,N_29639,N_29635);
or UO_3433 (O_3433,N_29821,N_29683);
or UO_3434 (O_3434,N_29624,N_29906);
nor UO_3435 (O_3435,N_29642,N_29762);
or UO_3436 (O_3436,N_29674,N_29511);
and UO_3437 (O_3437,N_29731,N_29959);
and UO_3438 (O_3438,N_29756,N_29903);
and UO_3439 (O_3439,N_29624,N_29738);
or UO_3440 (O_3440,N_29663,N_29552);
or UO_3441 (O_3441,N_29968,N_29974);
nand UO_3442 (O_3442,N_29512,N_29863);
or UO_3443 (O_3443,N_29688,N_29879);
or UO_3444 (O_3444,N_29686,N_29543);
nor UO_3445 (O_3445,N_29977,N_29854);
nor UO_3446 (O_3446,N_29758,N_29919);
nor UO_3447 (O_3447,N_29716,N_29625);
nand UO_3448 (O_3448,N_29845,N_29648);
or UO_3449 (O_3449,N_29734,N_29614);
nand UO_3450 (O_3450,N_29831,N_29834);
xnor UO_3451 (O_3451,N_29740,N_29556);
nand UO_3452 (O_3452,N_29597,N_29820);
xor UO_3453 (O_3453,N_29837,N_29580);
xnor UO_3454 (O_3454,N_29653,N_29726);
xor UO_3455 (O_3455,N_29535,N_29970);
nand UO_3456 (O_3456,N_29722,N_29603);
or UO_3457 (O_3457,N_29898,N_29621);
nand UO_3458 (O_3458,N_29772,N_29745);
xor UO_3459 (O_3459,N_29843,N_29891);
nand UO_3460 (O_3460,N_29554,N_29661);
nand UO_3461 (O_3461,N_29936,N_29531);
nand UO_3462 (O_3462,N_29505,N_29649);
nor UO_3463 (O_3463,N_29894,N_29592);
nand UO_3464 (O_3464,N_29617,N_29851);
nor UO_3465 (O_3465,N_29810,N_29755);
nand UO_3466 (O_3466,N_29602,N_29588);
nand UO_3467 (O_3467,N_29626,N_29970);
and UO_3468 (O_3468,N_29706,N_29795);
xnor UO_3469 (O_3469,N_29872,N_29855);
xnor UO_3470 (O_3470,N_29588,N_29823);
nor UO_3471 (O_3471,N_29682,N_29747);
xor UO_3472 (O_3472,N_29650,N_29657);
nor UO_3473 (O_3473,N_29653,N_29907);
xnor UO_3474 (O_3474,N_29868,N_29957);
nand UO_3475 (O_3475,N_29572,N_29770);
nor UO_3476 (O_3476,N_29551,N_29957);
or UO_3477 (O_3477,N_29987,N_29972);
xor UO_3478 (O_3478,N_29668,N_29871);
xnor UO_3479 (O_3479,N_29560,N_29637);
nor UO_3480 (O_3480,N_29839,N_29675);
or UO_3481 (O_3481,N_29818,N_29721);
or UO_3482 (O_3482,N_29577,N_29825);
nand UO_3483 (O_3483,N_29726,N_29851);
nand UO_3484 (O_3484,N_29809,N_29547);
nor UO_3485 (O_3485,N_29909,N_29855);
xor UO_3486 (O_3486,N_29505,N_29555);
nor UO_3487 (O_3487,N_29618,N_29684);
and UO_3488 (O_3488,N_29703,N_29575);
nor UO_3489 (O_3489,N_29943,N_29803);
and UO_3490 (O_3490,N_29791,N_29628);
and UO_3491 (O_3491,N_29534,N_29894);
nand UO_3492 (O_3492,N_29875,N_29515);
nor UO_3493 (O_3493,N_29618,N_29888);
nor UO_3494 (O_3494,N_29558,N_29925);
or UO_3495 (O_3495,N_29873,N_29672);
or UO_3496 (O_3496,N_29680,N_29997);
nand UO_3497 (O_3497,N_29840,N_29588);
nand UO_3498 (O_3498,N_29806,N_29877);
nor UO_3499 (O_3499,N_29946,N_29610);
endmodule