module basic_500_3000_500_15_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_309,In_387);
nor U1 (N_1,In_201,In_446);
or U2 (N_2,In_110,In_37);
xnor U3 (N_3,In_415,In_278);
nand U4 (N_4,In_329,In_475);
and U5 (N_5,In_60,In_109);
or U6 (N_6,In_254,In_346);
nand U7 (N_7,In_372,In_455);
xor U8 (N_8,In_351,In_232);
xor U9 (N_9,In_331,In_29);
xor U10 (N_10,In_177,In_236);
and U11 (N_11,In_404,In_179);
or U12 (N_12,In_343,In_382);
xor U13 (N_13,In_27,In_389);
xor U14 (N_14,In_456,In_216);
nor U15 (N_15,In_134,In_35);
nor U16 (N_16,In_116,In_454);
and U17 (N_17,In_198,In_125);
or U18 (N_18,In_374,In_299);
xor U19 (N_19,In_25,In_368);
and U20 (N_20,In_132,In_195);
xor U21 (N_21,In_225,In_405);
nand U22 (N_22,In_439,In_99);
xor U23 (N_23,In_321,In_154);
or U24 (N_24,In_170,In_428);
and U25 (N_25,In_396,In_365);
nand U26 (N_26,In_265,In_214);
or U27 (N_27,In_70,In_104);
nor U28 (N_28,In_465,In_2);
nand U29 (N_29,In_87,In_360);
nand U30 (N_30,In_267,In_74);
xnor U31 (N_31,In_234,In_102);
or U32 (N_32,In_129,In_275);
xor U33 (N_33,In_75,In_85);
nand U34 (N_34,In_491,In_196);
nand U35 (N_35,In_332,In_478);
nor U36 (N_36,In_51,In_176);
nor U37 (N_37,In_274,In_369);
and U38 (N_38,In_357,In_143);
or U39 (N_39,In_48,In_14);
nor U40 (N_40,In_121,In_130);
and U41 (N_41,In_440,In_392);
xnor U42 (N_42,In_305,In_127);
nand U43 (N_43,In_342,In_341);
or U44 (N_44,In_24,In_150);
and U45 (N_45,In_221,In_126);
nand U46 (N_46,In_311,In_431);
or U47 (N_47,In_292,In_97);
or U48 (N_48,In_249,In_119);
or U49 (N_49,In_304,In_194);
xnor U50 (N_50,In_349,In_277);
nand U51 (N_51,In_107,In_412);
nand U52 (N_52,In_448,In_94);
or U53 (N_53,In_61,In_33);
xnor U54 (N_54,In_21,In_380);
or U55 (N_55,In_339,In_282);
xnor U56 (N_56,In_203,In_247);
or U57 (N_57,In_135,In_86);
and U58 (N_58,In_231,In_89);
nand U59 (N_59,In_316,In_464);
or U60 (N_60,In_229,In_312);
xor U61 (N_61,In_65,In_363);
and U62 (N_62,In_113,In_18);
xnor U63 (N_63,In_178,In_174);
or U64 (N_64,In_444,In_62);
and U65 (N_65,In_451,In_480);
nor U66 (N_66,In_41,In_139);
and U67 (N_67,In_11,In_463);
xnor U68 (N_68,In_34,In_373);
xnor U69 (N_69,In_257,In_435);
and U70 (N_70,In_199,In_106);
nor U71 (N_71,In_297,In_430);
nand U72 (N_72,In_181,In_59);
and U73 (N_73,In_447,In_419);
or U74 (N_74,In_418,In_36);
xnor U75 (N_75,In_204,In_111);
or U76 (N_76,In_58,In_192);
or U77 (N_77,In_128,In_17);
xnor U78 (N_78,In_337,In_398);
nand U79 (N_79,In_457,In_131);
xnor U80 (N_80,In_492,In_461);
nand U81 (N_81,In_393,In_407);
and U82 (N_82,In_361,In_416);
nor U83 (N_83,In_52,In_384);
or U84 (N_84,In_397,In_133);
xnor U85 (N_85,In_210,In_490);
nor U86 (N_86,In_100,In_146);
and U87 (N_87,In_251,In_426);
and U88 (N_88,In_244,In_468);
nand U89 (N_89,In_445,In_255);
xnor U90 (N_90,In_4,In_161);
nor U91 (N_91,In_458,In_471);
nor U92 (N_92,In_84,In_486);
and U93 (N_93,In_413,In_103);
xnor U94 (N_94,In_497,In_166);
xnor U95 (N_95,In_91,In_200);
xor U96 (N_96,In_487,In_302);
or U97 (N_97,In_0,In_264);
xnor U98 (N_98,In_43,In_6);
xnor U99 (N_99,In_144,In_235);
nand U100 (N_100,In_273,In_239);
or U101 (N_101,In_64,In_326);
and U102 (N_102,In_50,In_452);
or U103 (N_103,In_420,In_317);
and U104 (N_104,In_148,In_423);
xnor U105 (N_105,In_485,In_336);
nand U106 (N_106,In_72,In_472);
nor U107 (N_107,In_180,In_163);
nor U108 (N_108,In_69,In_40);
or U109 (N_109,In_173,In_172);
nor U110 (N_110,In_95,In_145);
and U111 (N_111,In_46,In_303);
nor U112 (N_112,In_429,In_295);
nand U113 (N_113,In_286,In_375);
and U114 (N_114,In_352,In_307);
xor U115 (N_115,In_39,In_425);
xnor U116 (N_116,In_290,In_226);
and U117 (N_117,In_324,In_66);
and U118 (N_118,In_269,In_390);
or U119 (N_119,In_340,In_259);
nand U120 (N_120,In_151,In_45);
nand U121 (N_121,In_386,In_495);
xnor U122 (N_122,In_344,In_322);
xnor U123 (N_123,In_301,In_358);
nor U124 (N_124,In_80,In_142);
xnor U125 (N_125,In_88,In_12);
nand U126 (N_126,In_314,In_28);
nand U127 (N_127,In_206,In_421);
or U128 (N_128,In_83,In_207);
or U129 (N_129,In_400,In_320);
nor U130 (N_130,In_245,In_289);
or U131 (N_131,In_489,In_15);
nor U132 (N_132,In_399,In_325);
and U133 (N_133,In_153,In_479);
nor U134 (N_134,In_496,In_186);
nor U135 (N_135,In_473,In_138);
xor U136 (N_136,In_484,In_188);
nand U137 (N_137,In_197,In_175);
nand U138 (N_138,In_350,In_476);
nor U139 (N_139,In_162,In_68);
nand U140 (N_140,In_22,In_168);
and U141 (N_141,In_474,In_8);
nor U142 (N_142,In_183,In_93);
or U143 (N_143,In_152,In_228);
or U144 (N_144,In_268,In_248);
and U145 (N_145,In_262,In_345);
nand U146 (N_146,In_417,In_354);
or U147 (N_147,In_137,In_370);
nand U148 (N_148,In_258,In_120);
nand U149 (N_149,In_184,In_403);
and U150 (N_150,In_434,In_44);
xor U151 (N_151,In_298,In_79);
xnor U152 (N_152,In_433,In_217);
nand U153 (N_153,In_124,In_218);
nor U154 (N_154,In_371,In_73);
or U155 (N_155,In_157,In_283);
nand U156 (N_156,In_466,In_334);
xnor U157 (N_157,In_13,In_300);
or U158 (N_158,In_438,In_294);
and U159 (N_159,In_315,In_205);
xnor U160 (N_160,In_424,In_185);
or U161 (N_161,In_394,In_285);
or U162 (N_162,In_243,In_385);
or U163 (N_163,In_92,In_366);
nand U164 (N_164,In_499,In_155);
and U165 (N_165,In_388,In_356);
nand U166 (N_166,In_171,In_237);
nor U167 (N_167,In_391,In_488);
xnor U168 (N_168,In_401,In_77);
or U169 (N_169,In_459,In_383);
nor U170 (N_170,In_253,In_67);
nor U171 (N_171,In_213,In_19);
and U172 (N_172,In_9,In_31);
and U173 (N_173,In_240,In_140);
and U174 (N_174,In_323,In_427);
nor U175 (N_175,In_462,In_402);
xnor U176 (N_176,In_256,In_112);
or U177 (N_177,In_165,In_441);
nand U178 (N_178,In_63,In_147);
nand U179 (N_179,In_76,In_81);
or U180 (N_180,In_212,In_190);
nor U181 (N_181,In_362,In_182);
nor U182 (N_182,In_310,In_313);
and U183 (N_183,In_115,In_20);
or U184 (N_184,In_260,In_449);
and U185 (N_185,In_364,In_261);
nor U186 (N_186,In_348,In_101);
nand U187 (N_187,In_319,In_280);
nand U188 (N_188,In_381,In_54);
nor U189 (N_189,In_498,In_284);
or U190 (N_190,In_276,In_90);
nand U191 (N_191,In_470,In_271);
and U192 (N_192,In_494,In_223);
xnor U193 (N_193,In_98,In_202);
and U194 (N_194,In_26,In_30);
and U195 (N_195,In_327,In_266);
xor U196 (N_196,In_159,In_436);
and U197 (N_197,In_414,In_122);
xnor U198 (N_198,In_7,In_469);
nand U199 (N_199,In_270,In_306);
nor U200 (N_200,In_246,In_211);
xnor U201 (N_201,N_36,N_24);
nand U202 (N_202,N_17,N_55);
and U203 (N_203,N_125,In_49);
xnor U204 (N_204,In_411,N_74);
and U205 (N_205,N_44,N_185);
nor U206 (N_206,N_188,N_15);
and U207 (N_207,N_97,In_395);
nor U208 (N_208,N_41,N_169);
xor U209 (N_209,In_32,In_1);
and U210 (N_210,N_143,In_408);
nand U211 (N_211,N_162,In_296);
xor U212 (N_212,In_208,N_4);
nand U213 (N_213,N_56,In_118);
and U214 (N_214,In_355,In_482);
nor U215 (N_215,N_49,N_95);
xnor U216 (N_216,N_141,N_147);
and U217 (N_217,N_152,In_38);
nor U218 (N_218,N_106,N_8);
xor U219 (N_219,N_187,In_330);
xnor U220 (N_220,N_75,In_141);
nand U221 (N_221,N_117,N_170);
nor U222 (N_222,N_87,N_83);
xnor U223 (N_223,N_21,In_432);
nand U224 (N_224,N_22,N_151);
nor U225 (N_225,In_238,In_10);
xor U226 (N_226,N_149,In_224);
nand U227 (N_227,N_67,N_119);
and U228 (N_228,N_127,N_25);
nor U229 (N_229,In_227,N_157);
or U230 (N_230,In_376,N_70);
nor U231 (N_231,N_72,N_91);
nand U232 (N_232,In_291,In_483);
nand U233 (N_233,In_279,N_103);
xor U234 (N_234,N_62,In_82);
or U235 (N_235,N_9,N_68);
and U236 (N_236,In_47,N_28);
or U237 (N_237,N_148,N_175);
nor U238 (N_238,N_66,In_56);
and U239 (N_239,N_124,In_149);
xor U240 (N_240,N_166,N_34);
or U241 (N_241,In_338,In_193);
and U242 (N_242,N_191,In_233);
nor U243 (N_243,N_42,In_3);
xor U244 (N_244,In_123,In_117);
or U245 (N_245,N_113,In_281);
and U246 (N_246,In_164,N_190);
and U247 (N_247,In_460,In_450);
nor U248 (N_248,N_105,In_189);
nor U249 (N_249,N_111,N_77);
nor U250 (N_250,In_55,N_108);
and U251 (N_251,N_81,In_42);
nand U252 (N_252,N_2,N_13);
nor U253 (N_253,N_153,N_14);
xor U254 (N_254,In_191,N_135);
and U255 (N_255,N_159,N_23);
nor U256 (N_256,N_154,N_1);
or U257 (N_257,N_73,In_169);
nor U258 (N_258,N_19,N_7);
or U259 (N_259,N_30,In_263);
nand U260 (N_260,N_189,In_220);
nor U261 (N_261,N_5,N_100);
or U262 (N_262,In_481,In_328);
xnor U263 (N_263,In_367,In_287);
xnor U264 (N_264,N_161,In_406);
and U265 (N_265,N_51,N_12);
and U266 (N_266,N_122,N_82);
and U267 (N_267,N_0,In_187);
nor U268 (N_268,N_94,In_250);
nor U269 (N_269,N_120,In_160);
nor U270 (N_270,In_57,In_272);
or U271 (N_271,N_184,N_35);
nand U272 (N_272,N_88,N_144);
nand U273 (N_273,N_61,N_172);
xor U274 (N_274,N_6,N_54);
xnor U275 (N_275,N_59,N_78);
and U276 (N_276,N_58,N_195);
xor U277 (N_277,N_114,N_27);
and U278 (N_278,N_193,N_43);
or U279 (N_279,N_137,N_96);
or U280 (N_280,N_116,In_308);
and U281 (N_281,In_96,In_437);
xor U282 (N_282,N_40,In_230);
xnor U283 (N_283,N_174,N_198);
nor U284 (N_284,N_89,N_145);
and U285 (N_285,N_121,N_65);
xor U286 (N_286,N_128,N_32);
nand U287 (N_287,N_3,In_78);
and U288 (N_288,N_92,N_53);
nand U289 (N_289,N_176,N_26);
and U290 (N_290,N_150,N_156);
or U291 (N_291,N_52,N_38);
and U292 (N_292,N_183,N_186);
nor U293 (N_293,N_133,N_134);
or U294 (N_294,N_178,N_197);
or U295 (N_295,N_93,N_192);
nand U296 (N_296,In_333,In_347);
or U297 (N_297,N_194,N_131);
xor U298 (N_298,N_139,In_288);
or U299 (N_299,N_29,N_196);
nand U300 (N_300,N_37,N_199);
and U301 (N_301,In_467,In_219);
and U302 (N_302,N_146,N_181);
nor U303 (N_303,N_142,N_84);
or U304 (N_304,In_377,N_71);
xor U305 (N_305,In_453,N_101);
and U306 (N_306,In_493,In_108);
nand U307 (N_307,N_140,In_53);
and U308 (N_308,In_71,N_138);
or U309 (N_309,N_57,N_79);
or U310 (N_310,N_46,N_39);
nor U311 (N_311,In_252,In_5);
xnor U312 (N_312,N_130,In_442);
or U313 (N_313,In_215,N_20);
xor U314 (N_314,N_136,N_104);
or U315 (N_315,N_80,In_353);
xor U316 (N_316,N_112,In_158);
nand U317 (N_317,In_241,In_242);
nand U318 (N_318,In_114,N_171);
or U319 (N_319,N_33,N_45);
nor U320 (N_320,In_156,In_422);
or U321 (N_321,In_335,N_18);
xor U322 (N_322,In_136,N_64);
xnor U323 (N_323,In_105,N_177);
and U324 (N_324,In_222,In_477);
xnor U325 (N_325,N_98,In_409);
xnor U326 (N_326,In_443,In_378);
xor U327 (N_327,N_102,N_164);
nand U328 (N_328,N_182,In_167);
nand U329 (N_329,N_86,In_16);
nand U330 (N_330,N_165,In_359);
nand U331 (N_331,In_209,N_69);
nor U332 (N_332,N_168,N_180);
nand U333 (N_333,N_76,N_173);
xor U334 (N_334,N_129,N_10);
or U335 (N_335,N_16,N_48);
or U336 (N_336,N_179,N_31);
or U337 (N_337,N_132,N_123);
xnor U338 (N_338,N_11,N_109);
and U339 (N_339,In_410,N_110);
nand U340 (N_340,N_85,N_63);
nor U341 (N_341,In_379,N_115);
nor U342 (N_342,N_155,N_167);
and U343 (N_343,N_160,N_99);
nand U344 (N_344,N_90,In_23);
or U345 (N_345,N_50,N_158);
and U346 (N_346,N_126,N_47);
and U347 (N_347,N_118,N_107);
nand U348 (N_348,In_318,N_163);
and U349 (N_349,In_293,N_60);
nor U350 (N_350,In_219,N_131);
or U351 (N_351,N_97,N_115);
and U352 (N_352,In_23,N_115);
or U353 (N_353,N_49,In_330);
xor U354 (N_354,N_121,N_159);
and U355 (N_355,In_55,N_81);
nor U356 (N_356,N_149,N_5);
xor U357 (N_357,N_96,N_10);
or U358 (N_358,In_149,N_123);
nor U359 (N_359,In_53,N_69);
nor U360 (N_360,N_0,N_111);
and U361 (N_361,N_92,N_100);
and U362 (N_362,In_10,N_109);
xor U363 (N_363,N_3,In_238);
nand U364 (N_364,N_14,N_9);
or U365 (N_365,In_411,N_163);
nand U366 (N_366,In_411,N_33);
nor U367 (N_367,In_409,In_437);
nand U368 (N_368,N_160,N_148);
nand U369 (N_369,N_155,In_108);
nor U370 (N_370,N_44,N_191);
and U371 (N_371,N_181,N_176);
nor U372 (N_372,N_92,N_167);
nor U373 (N_373,N_98,In_3);
or U374 (N_374,In_82,In_410);
and U375 (N_375,In_450,N_2);
nor U376 (N_376,N_94,N_3);
and U377 (N_377,N_45,N_129);
and U378 (N_378,N_69,N_12);
or U379 (N_379,N_74,In_56);
nor U380 (N_380,N_51,N_76);
nor U381 (N_381,In_193,N_121);
or U382 (N_382,N_29,In_16);
nor U383 (N_383,N_61,N_164);
and U384 (N_384,N_192,N_29);
and U385 (N_385,In_187,N_189);
nor U386 (N_386,N_142,In_211);
or U387 (N_387,N_74,N_97);
xnor U388 (N_388,In_437,N_91);
xnor U389 (N_389,N_61,In_105);
or U390 (N_390,In_32,N_33);
or U391 (N_391,In_318,N_157);
xor U392 (N_392,N_198,N_50);
xor U393 (N_393,N_182,In_187);
nor U394 (N_394,N_0,In_296);
and U395 (N_395,N_65,In_359);
and U396 (N_396,N_42,In_227);
nand U397 (N_397,In_252,N_78);
nor U398 (N_398,N_161,N_82);
nand U399 (N_399,In_105,N_141);
xnor U400 (N_400,N_280,N_242);
xor U401 (N_401,N_363,N_246);
xor U402 (N_402,N_353,N_385);
nand U403 (N_403,N_360,N_228);
or U404 (N_404,N_296,N_319);
nor U405 (N_405,N_239,N_315);
or U406 (N_406,N_376,N_369);
or U407 (N_407,N_210,N_271);
nand U408 (N_408,N_278,N_313);
nand U409 (N_409,N_295,N_336);
or U410 (N_410,N_279,N_331);
or U411 (N_411,N_343,N_221);
nand U412 (N_412,N_260,N_229);
nor U413 (N_413,N_332,N_371);
nand U414 (N_414,N_291,N_316);
or U415 (N_415,N_232,N_300);
nor U416 (N_416,N_350,N_390);
and U417 (N_417,N_344,N_352);
nand U418 (N_418,N_354,N_285);
nand U419 (N_419,N_374,N_327);
xnor U420 (N_420,N_357,N_202);
or U421 (N_421,N_233,N_310);
xor U422 (N_422,N_306,N_224);
or U423 (N_423,N_388,N_397);
or U424 (N_424,N_366,N_234);
nand U425 (N_425,N_253,N_265);
or U426 (N_426,N_240,N_267);
nor U427 (N_427,N_255,N_348);
and U428 (N_428,N_220,N_378);
and U429 (N_429,N_261,N_399);
xor U430 (N_430,N_322,N_257);
nand U431 (N_431,N_303,N_200);
or U432 (N_432,N_236,N_201);
nor U433 (N_433,N_218,N_335);
xor U434 (N_434,N_324,N_274);
nand U435 (N_435,N_245,N_283);
nand U436 (N_436,N_387,N_273);
nand U437 (N_437,N_297,N_386);
nor U438 (N_438,N_365,N_225);
xor U439 (N_439,N_321,N_393);
or U440 (N_440,N_219,N_275);
or U441 (N_441,N_308,N_312);
nor U442 (N_442,N_241,N_395);
and U443 (N_443,N_337,N_311);
nand U444 (N_444,N_268,N_284);
nand U445 (N_445,N_290,N_345);
and U446 (N_446,N_329,N_282);
nor U447 (N_447,N_288,N_227);
xnor U448 (N_448,N_341,N_398);
xor U449 (N_449,N_252,N_272);
nor U450 (N_450,N_379,N_359);
nand U451 (N_451,N_207,N_342);
and U452 (N_452,N_269,N_286);
xor U453 (N_453,N_320,N_307);
nor U454 (N_454,N_334,N_368);
nor U455 (N_455,N_209,N_380);
xnor U456 (N_456,N_340,N_264);
and U457 (N_457,N_262,N_301);
or U458 (N_458,N_223,N_333);
nand U459 (N_459,N_214,N_205);
or U460 (N_460,N_249,N_394);
nor U461 (N_461,N_304,N_277);
nand U462 (N_462,N_356,N_248);
nor U463 (N_463,N_254,N_287);
nand U464 (N_464,N_384,N_361);
nor U465 (N_465,N_381,N_293);
nand U466 (N_466,N_317,N_247);
and U467 (N_467,N_230,N_302);
and U468 (N_468,N_203,N_314);
and U469 (N_469,N_256,N_211);
nand U470 (N_470,N_222,N_270);
nand U471 (N_471,N_367,N_305);
nand U472 (N_472,N_237,N_281);
and U473 (N_473,N_251,N_358);
or U474 (N_474,N_382,N_318);
nor U475 (N_475,N_309,N_235);
nand U476 (N_476,N_391,N_266);
or U477 (N_477,N_392,N_289);
and U478 (N_478,N_243,N_294);
xor U479 (N_479,N_346,N_217);
nand U480 (N_480,N_373,N_347);
and U481 (N_481,N_326,N_226);
nand U482 (N_482,N_396,N_259);
and U483 (N_483,N_276,N_215);
nand U484 (N_484,N_238,N_355);
xor U485 (N_485,N_377,N_299);
xnor U486 (N_486,N_328,N_330);
and U487 (N_487,N_364,N_213);
nand U488 (N_488,N_339,N_349);
nand U489 (N_489,N_208,N_204);
xor U490 (N_490,N_212,N_375);
nand U491 (N_491,N_351,N_362);
and U492 (N_492,N_370,N_389);
xnor U493 (N_493,N_206,N_298);
xnor U494 (N_494,N_325,N_323);
or U495 (N_495,N_231,N_258);
or U496 (N_496,N_263,N_383);
xnor U497 (N_497,N_372,N_250);
nor U498 (N_498,N_292,N_338);
and U499 (N_499,N_244,N_216);
nor U500 (N_500,N_293,N_310);
and U501 (N_501,N_263,N_308);
or U502 (N_502,N_355,N_398);
nand U503 (N_503,N_258,N_396);
nand U504 (N_504,N_377,N_311);
xor U505 (N_505,N_332,N_333);
nand U506 (N_506,N_274,N_320);
or U507 (N_507,N_391,N_230);
or U508 (N_508,N_200,N_395);
nor U509 (N_509,N_372,N_203);
and U510 (N_510,N_397,N_255);
xnor U511 (N_511,N_273,N_377);
or U512 (N_512,N_363,N_280);
and U513 (N_513,N_224,N_285);
nor U514 (N_514,N_261,N_219);
or U515 (N_515,N_350,N_244);
xor U516 (N_516,N_298,N_304);
nor U517 (N_517,N_312,N_280);
xor U518 (N_518,N_254,N_381);
xnor U519 (N_519,N_279,N_377);
and U520 (N_520,N_371,N_357);
or U521 (N_521,N_273,N_370);
xnor U522 (N_522,N_327,N_246);
and U523 (N_523,N_292,N_265);
or U524 (N_524,N_259,N_215);
nor U525 (N_525,N_317,N_248);
nand U526 (N_526,N_337,N_289);
nand U527 (N_527,N_366,N_233);
nand U528 (N_528,N_207,N_251);
nand U529 (N_529,N_355,N_345);
or U530 (N_530,N_364,N_325);
nand U531 (N_531,N_278,N_357);
nor U532 (N_532,N_326,N_237);
and U533 (N_533,N_380,N_245);
or U534 (N_534,N_251,N_298);
nand U535 (N_535,N_258,N_288);
and U536 (N_536,N_254,N_322);
or U537 (N_537,N_313,N_277);
xor U538 (N_538,N_220,N_365);
xor U539 (N_539,N_234,N_287);
or U540 (N_540,N_350,N_299);
nor U541 (N_541,N_370,N_303);
xnor U542 (N_542,N_329,N_398);
or U543 (N_543,N_265,N_218);
nand U544 (N_544,N_222,N_293);
and U545 (N_545,N_392,N_388);
xnor U546 (N_546,N_259,N_384);
and U547 (N_547,N_249,N_381);
nand U548 (N_548,N_286,N_299);
xnor U549 (N_549,N_348,N_221);
nand U550 (N_550,N_270,N_290);
nand U551 (N_551,N_390,N_202);
xor U552 (N_552,N_281,N_322);
or U553 (N_553,N_366,N_206);
nand U554 (N_554,N_357,N_232);
nand U555 (N_555,N_264,N_339);
nor U556 (N_556,N_253,N_205);
or U557 (N_557,N_277,N_324);
xnor U558 (N_558,N_393,N_244);
nor U559 (N_559,N_285,N_206);
xor U560 (N_560,N_399,N_201);
xor U561 (N_561,N_213,N_371);
nand U562 (N_562,N_253,N_395);
xnor U563 (N_563,N_305,N_318);
xor U564 (N_564,N_376,N_218);
xnor U565 (N_565,N_393,N_224);
xor U566 (N_566,N_302,N_266);
or U567 (N_567,N_273,N_227);
or U568 (N_568,N_312,N_316);
nand U569 (N_569,N_274,N_215);
xor U570 (N_570,N_363,N_381);
xnor U571 (N_571,N_284,N_228);
xor U572 (N_572,N_271,N_288);
or U573 (N_573,N_396,N_374);
or U574 (N_574,N_373,N_389);
nand U575 (N_575,N_275,N_259);
or U576 (N_576,N_357,N_230);
or U577 (N_577,N_251,N_341);
nor U578 (N_578,N_321,N_240);
xor U579 (N_579,N_393,N_243);
or U580 (N_580,N_326,N_219);
xnor U581 (N_581,N_299,N_276);
xor U582 (N_582,N_222,N_291);
or U583 (N_583,N_342,N_270);
or U584 (N_584,N_254,N_259);
and U585 (N_585,N_321,N_265);
nand U586 (N_586,N_305,N_329);
or U587 (N_587,N_263,N_236);
nor U588 (N_588,N_322,N_248);
nand U589 (N_589,N_294,N_235);
xor U590 (N_590,N_340,N_250);
nor U591 (N_591,N_346,N_225);
nor U592 (N_592,N_285,N_244);
and U593 (N_593,N_334,N_365);
xnor U594 (N_594,N_229,N_338);
xor U595 (N_595,N_200,N_309);
and U596 (N_596,N_282,N_261);
and U597 (N_597,N_327,N_208);
nor U598 (N_598,N_240,N_348);
nand U599 (N_599,N_357,N_264);
nor U600 (N_600,N_535,N_560);
nand U601 (N_601,N_492,N_568);
xnor U602 (N_602,N_542,N_454);
nor U603 (N_603,N_462,N_520);
or U604 (N_604,N_427,N_569);
and U605 (N_605,N_475,N_436);
nor U606 (N_606,N_419,N_460);
nor U607 (N_607,N_512,N_582);
nand U608 (N_608,N_485,N_437);
or U609 (N_609,N_575,N_450);
or U610 (N_610,N_482,N_537);
or U611 (N_611,N_589,N_412);
nor U612 (N_612,N_544,N_457);
nand U613 (N_613,N_581,N_596);
xnor U614 (N_614,N_456,N_578);
xor U615 (N_615,N_556,N_525);
or U616 (N_616,N_442,N_477);
xnor U617 (N_617,N_481,N_528);
nor U618 (N_618,N_496,N_583);
nor U619 (N_619,N_425,N_409);
xnor U620 (N_620,N_504,N_444);
xor U621 (N_621,N_598,N_593);
nor U622 (N_622,N_577,N_490);
xnor U623 (N_623,N_500,N_495);
nand U624 (N_624,N_432,N_426);
nand U625 (N_625,N_558,N_452);
and U626 (N_626,N_552,N_403);
and U627 (N_627,N_584,N_549);
nand U628 (N_628,N_592,N_562);
and U629 (N_629,N_458,N_428);
nand U630 (N_630,N_449,N_588);
xor U631 (N_631,N_599,N_546);
xor U632 (N_632,N_423,N_540);
nand U633 (N_633,N_410,N_503);
and U634 (N_634,N_561,N_463);
nand U635 (N_635,N_406,N_587);
nand U636 (N_636,N_564,N_418);
xor U637 (N_637,N_572,N_590);
and U638 (N_638,N_545,N_483);
or U639 (N_639,N_422,N_438);
nand U640 (N_640,N_515,N_506);
nand U641 (N_641,N_470,N_411);
or U642 (N_642,N_529,N_484);
nor U643 (N_643,N_447,N_404);
or U644 (N_644,N_448,N_479);
xor U645 (N_645,N_571,N_510);
nand U646 (N_646,N_513,N_408);
or U647 (N_647,N_517,N_420);
or U648 (N_648,N_459,N_526);
nand U649 (N_649,N_467,N_471);
or U650 (N_650,N_402,N_440);
nand U651 (N_651,N_521,N_469);
and U652 (N_652,N_509,N_430);
nand U653 (N_653,N_541,N_416);
or U654 (N_654,N_468,N_434);
and U655 (N_655,N_579,N_480);
xor U656 (N_656,N_439,N_514);
nor U657 (N_657,N_565,N_415);
and U658 (N_658,N_405,N_421);
nand U659 (N_659,N_555,N_538);
xor U660 (N_660,N_511,N_497);
and U661 (N_661,N_400,N_414);
xor U662 (N_662,N_488,N_570);
and U663 (N_663,N_566,N_473);
nor U664 (N_664,N_554,N_543);
and U665 (N_665,N_465,N_435);
or U666 (N_666,N_519,N_474);
and U667 (N_667,N_585,N_586);
nor U668 (N_668,N_595,N_516);
and U669 (N_669,N_498,N_464);
nor U670 (N_670,N_573,N_550);
xor U671 (N_671,N_576,N_597);
nor U672 (N_672,N_413,N_445);
nand U673 (N_673,N_505,N_494);
and U674 (N_674,N_489,N_431);
nor U675 (N_675,N_441,N_524);
or U676 (N_676,N_594,N_493);
nor U677 (N_677,N_446,N_534);
xnor U678 (N_678,N_508,N_522);
or U679 (N_679,N_417,N_523);
xor U680 (N_680,N_502,N_472);
and U681 (N_681,N_407,N_518);
or U682 (N_682,N_557,N_547);
nor U683 (N_683,N_461,N_527);
or U684 (N_684,N_539,N_499);
nand U685 (N_685,N_491,N_401);
nand U686 (N_686,N_487,N_533);
xnor U687 (N_687,N_574,N_429);
or U688 (N_688,N_531,N_563);
nor U689 (N_689,N_553,N_536);
nand U690 (N_690,N_424,N_453);
xnor U691 (N_691,N_443,N_478);
nor U692 (N_692,N_551,N_486);
or U693 (N_693,N_433,N_580);
or U694 (N_694,N_466,N_451);
nand U695 (N_695,N_567,N_476);
nand U696 (N_696,N_532,N_507);
or U697 (N_697,N_548,N_591);
nand U698 (N_698,N_559,N_530);
and U699 (N_699,N_501,N_455);
nand U700 (N_700,N_516,N_513);
and U701 (N_701,N_412,N_517);
nand U702 (N_702,N_556,N_580);
nand U703 (N_703,N_428,N_575);
or U704 (N_704,N_463,N_426);
nand U705 (N_705,N_577,N_468);
nor U706 (N_706,N_587,N_569);
and U707 (N_707,N_420,N_575);
or U708 (N_708,N_462,N_424);
nor U709 (N_709,N_587,N_422);
xor U710 (N_710,N_416,N_574);
nor U711 (N_711,N_569,N_432);
or U712 (N_712,N_587,N_586);
nor U713 (N_713,N_419,N_453);
nand U714 (N_714,N_412,N_575);
nor U715 (N_715,N_403,N_585);
or U716 (N_716,N_446,N_566);
or U717 (N_717,N_576,N_475);
or U718 (N_718,N_578,N_598);
nand U719 (N_719,N_419,N_521);
nand U720 (N_720,N_585,N_432);
and U721 (N_721,N_575,N_580);
nand U722 (N_722,N_408,N_583);
nor U723 (N_723,N_539,N_594);
xor U724 (N_724,N_530,N_507);
xor U725 (N_725,N_530,N_442);
nand U726 (N_726,N_408,N_431);
or U727 (N_727,N_458,N_518);
or U728 (N_728,N_422,N_543);
nand U729 (N_729,N_428,N_410);
nand U730 (N_730,N_560,N_524);
xor U731 (N_731,N_449,N_445);
nor U732 (N_732,N_499,N_425);
nor U733 (N_733,N_489,N_444);
nor U734 (N_734,N_463,N_576);
or U735 (N_735,N_439,N_512);
nand U736 (N_736,N_403,N_589);
or U737 (N_737,N_515,N_554);
and U738 (N_738,N_453,N_560);
or U739 (N_739,N_502,N_435);
xnor U740 (N_740,N_429,N_472);
xnor U741 (N_741,N_500,N_467);
or U742 (N_742,N_474,N_475);
xor U743 (N_743,N_501,N_402);
or U744 (N_744,N_528,N_521);
and U745 (N_745,N_455,N_419);
xnor U746 (N_746,N_570,N_532);
xor U747 (N_747,N_561,N_479);
and U748 (N_748,N_531,N_451);
or U749 (N_749,N_446,N_544);
and U750 (N_750,N_442,N_544);
or U751 (N_751,N_464,N_470);
or U752 (N_752,N_447,N_463);
nor U753 (N_753,N_505,N_497);
or U754 (N_754,N_583,N_487);
or U755 (N_755,N_451,N_526);
xnor U756 (N_756,N_433,N_447);
or U757 (N_757,N_489,N_582);
nand U758 (N_758,N_480,N_468);
nor U759 (N_759,N_426,N_524);
and U760 (N_760,N_536,N_517);
nand U761 (N_761,N_584,N_456);
nand U762 (N_762,N_417,N_538);
xnor U763 (N_763,N_582,N_590);
and U764 (N_764,N_498,N_591);
or U765 (N_765,N_421,N_484);
xnor U766 (N_766,N_527,N_446);
nand U767 (N_767,N_449,N_434);
and U768 (N_768,N_545,N_476);
or U769 (N_769,N_595,N_480);
or U770 (N_770,N_598,N_513);
and U771 (N_771,N_496,N_480);
or U772 (N_772,N_590,N_433);
xnor U773 (N_773,N_553,N_451);
nor U774 (N_774,N_499,N_545);
xnor U775 (N_775,N_512,N_436);
or U776 (N_776,N_551,N_589);
nor U777 (N_777,N_433,N_430);
or U778 (N_778,N_575,N_534);
nor U779 (N_779,N_512,N_584);
nand U780 (N_780,N_438,N_536);
and U781 (N_781,N_401,N_405);
or U782 (N_782,N_439,N_560);
or U783 (N_783,N_577,N_497);
and U784 (N_784,N_430,N_412);
nand U785 (N_785,N_426,N_405);
and U786 (N_786,N_402,N_493);
or U787 (N_787,N_568,N_497);
and U788 (N_788,N_496,N_527);
and U789 (N_789,N_570,N_420);
or U790 (N_790,N_431,N_517);
xnor U791 (N_791,N_444,N_583);
and U792 (N_792,N_554,N_561);
and U793 (N_793,N_551,N_431);
nand U794 (N_794,N_525,N_567);
nor U795 (N_795,N_471,N_521);
and U796 (N_796,N_502,N_560);
nand U797 (N_797,N_574,N_424);
and U798 (N_798,N_403,N_509);
xnor U799 (N_799,N_438,N_552);
nand U800 (N_800,N_791,N_732);
and U801 (N_801,N_676,N_753);
xnor U802 (N_802,N_746,N_778);
xnor U803 (N_803,N_694,N_772);
and U804 (N_804,N_667,N_610);
and U805 (N_805,N_755,N_630);
or U806 (N_806,N_699,N_708);
nand U807 (N_807,N_724,N_602);
xor U808 (N_808,N_726,N_795);
and U809 (N_809,N_693,N_767);
and U810 (N_810,N_617,N_671);
or U811 (N_811,N_731,N_689);
xor U812 (N_812,N_710,N_759);
nor U813 (N_813,N_733,N_611);
nand U814 (N_814,N_612,N_656);
nand U815 (N_815,N_715,N_714);
nand U816 (N_816,N_628,N_793);
nand U817 (N_817,N_758,N_763);
nand U818 (N_818,N_723,N_616);
nor U819 (N_819,N_734,N_675);
and U820 (N_820,N_635,N_697);
or U821 (N_821,N_701,N_727);
and U822 (N_822,N_608,N_662);
and U823 (N_823,N_797,N_738);
xnor U824 (N_824,N_629,N_752);
xor U825 (N_825,N_606,N_601);
or U826 (N_826,N_653,N_679);
or U827 (N_827,N_775,N_650);
nor U828 (N_828,N_777,N_786);
nand U829 (N_829,N_771,N_631);
nand U830 (N_830,N_741,N_687);
nand U831 (N_831,N_640,N_622);
nor U832 (N_832,N_773,N_742);
or U833 (N_833,N_678,N_692);
nor U834 (N_834,N_737,N_688);
or U835 (N_835,N_750,N_729);
or U836 (N_836,N_661,N_794);
xor U837 (N_837,N_613,N_695);
nand U838 (N_838,N_717,N_761);
xor U839 (N_839,N_757,N_637);
nand U840 (N_840,N_636,N_633);
or U841 (N_841,N_747,N_624);
nor U842 (N_842,N_706,N_762);
xor U843 (N_843,N_685,N_625);
nand U844 (N_844,N_647,N_626);
and U845 (N_845,N_751,N_618);
nor U846 (N_846,N_691,N_720);
nand U847 (N_847,N_649,N_658);
nand U848 (N_848,N_765,N_621);
nand U849 (N_849,N_743,N_638);
and U850 (N_850,N_620,N_632);
nor U851 (N_851,N_668,N_686);
xnor U852 (N_852,N_645,N_604);
nand U853 (N_853,N_756,N_799);
and U854 (N_854,N_718,N_739);
or U855 (N_855,N_615,N_768);
and U856 (N_856,N_677,N_779);
and U857 (N_857,N_744,N_785);
nor U858 (N_858,N_764,N_627);
nand U859 (N_859,N_774,N_722);
xnor U860 (N_860,N_787,N_790);
or U861 (N_861,N_725,N_760);
nand U862 (N_862,N_745,N_769);
nor U863 (N_863,N_670,N_709);
or U864 (N_864,N_711,N_700);
nand U865 (N_865,N_784,N_639);
xnor U866 (N_866,N_748,N_607);
or U867 (N_867,N_707,N_614);
and U868 (N_868,N_643,N_703);
and U869 (N_869,N_754,N_672);
xor U870 (N_870,N_713,N_735);
nor U871 (N_871,N_644,N_776);
and U872 (N_872,N_641,N_654);
xor U873 (N_873,N_704,N_659);
or U874 (N_874,N_736,N_719);
and U875 (N_875,N_796,N_634);
or U876 (N_876,N_766,N_721);
nor U877 (N_877,N_792,N_783);
xnor U878 (N_878,N_646,N_674);
and U879 (N_879,N_690,N_663);
and U880 (N_880,N_666,N_680);
nor U881 (N_881,N_696,N_664);
and U882 (N_882,N_728,N_652);
nor U883 (N_883,N_605,N_673);
nand U884 (N_884,N_788,N_609);
xor U885 (N_885,N_623,N_603);
xnor U886 (N_886,N_698,N_780);
and U887 (N_887,N_665,N_684);
and U888 (N_888,N_657,N_782);
nand U889 (N_889,N_619,N_682);
nand U890 (N_890,N_770,N_798);
nor U891 (N_891,N_681,N_600);
xnor U892 (N_892,N_712,N_789);
nor U893 (N_893,N_730,N_749);
or U894 (N_894,N_716,N_660);
xnor U895 (N_895,N_648,N_683);
or U896 (N_896,N_702,N_655);
or U897 (N_897,N_669,N_642);
or U898 (N_898,N_740,N_651);
or U899 (N_899,N_705,N_781);
or U900 (N_900,N_715,N_613);
and U901 (N_901,N_791,N_661);
nor U902 (N_902,N_654,N_684);
or U903 (N_903,N_744,N_601);
or U904 (N_904,N_658,N_698);
xor U905 (N_905,N_674,N_797);
and U906 (N_906,N_678,N_771);
or U907 (N_907,N_631,N_719);
xor U908 (N_908,N_636,N_776);
or U909 (N_909,N_666,N_660);
nor U910 (N_910,N_757,N_693);
or U911 (N_911,N_746,N_668);
and U912 (N_912,N_665,N_766);
and U913 (N_913,N_709,N_762);
and U914 (N_914,N_623,N_718);
nand U915 (N_915,N_777,N_646);
nand U916 (N_916,N_716,N_772);
and U917 (N_917,N_739,N_607);
and U918 (N_918,N_781,N_732);
nor U919 (N_919,N_741,N_783);
or U920 (N_920,N_736,N_777);
nand U921 (N_921,N_631,N_786);
nand U922 (N_922,N_798,N_690);
xor U923 (N_923,N_610,N_618);
nand U924 (N_924,N_662,N_630);
nand U925 (N_925,N_796,N_765);
nand U926 (N_926,N_691,N_642);
xor U927 (N_927,N_644,N_715);
and U928 (N_928,N_642,N_730);
and U929 (N_929,N_765,N_674);
or U930 (N_930,N_682,N_784);
xor U931 (N_931,N_664,N_767);
or U932 (N_932,N_737,N_785);
and U933 (N_933,N_609,N_688);
or U934 (N_934,N_757,N_796);
or U935 (N_935,N_636,N_755);
nor U936 (N_936,N_775,N_643);
or U937 (N_937,N_766,N_645);
and U938 (N_938,N_746,N_628);
nand U939 (N_939,N_606,N_713);
nor U940 (N_940,N_644,N_732);
and U941 (N_941,N_601,N_763);
and U942 (N_942,N_606,N_723);
and U943 (N_943,N_769,N_739);
or U944 (N_944,N_687,N_635);
and U945 (N_945,N_609,N_762);
nand U946 (N_946,N_602,N_662);
or U947 (N_947,N_662,N_660);
xnor U948 (N_948,N_689,N_755);
nor U949 (N_949,N_660,N_663);
and U950 (N_950,N_653,N_638);
nand U951 (N_951,N_707,N_633);
nand U952 (N_952,N_604,N_689);
nor U953 (N_953,N_700,N_663);
xor U954 (N_954,N_648,N_791);
xor U955 (N_955,N_794,N_730);
or U956 (N_956,N_765,N_706);
xor U957 (N_957,N_662,N_658);
or U958 (N_958,N_636,N_747);
xor U959 (N_959,N_772,N_636);
xnor U960 (N_960,N_639,N_692);
nand U961 (N_961,N_763,N_760);
xnor U962 (N_962,N_629,N_667);
or U963 (N_963,N_605,N_786);
xor U964 (N_964,N_782,N_730);
or U965 (N_965,N_768,N_776);
or U966 (N_966,N_764,N_610);
and U967 (N_967,N_677,N_717);
and U968 (N_968,N_669,N_790);
and U969 (N_969,N_692,N_721);
or U970 (N_970,N_627,N_739);
and U971 (N_971,N_674,N_666);
and U972 (N_972,N_786,N_699);
nor U973 (N_973,N_642,N_769);
nand U974 (N_974,N_655,N_794);
nand U975 (N_975,N_757,N_751);
or U976 (N_976,N_779,N_722);
xor U977 (N_977,N_711,N_642);
and U978 (N_978,N_716,N_722);
nor U979 (N_979,N_628,N_606);
nor U980 (N_980,N_624,N_725);
nor U981 (N_981,N_745,N_710);
nor U982 (N_982,N_761,N_721);
nor U983 (N_983,N_690,N_697);
or U984 (N_984,N_695,N_601);
or U985 (N_985,N_741,N_600);
nor U986 (N_986,N_749,N_791);
nor U987 (N_987,N_611,N_646);
nor U988 (N_988,N_647,N_750);
or U989 (N_989,N_605,N_781);
nand U990 (N_990,N_753,N_707);
xor U991 (N_991,N_731,N_718);
xor U992 (N_992,N_678,N_795);
nor U993 (N_993,N_700,N_626);
and U994 (N_994,N_744,N_787);
nand U995 (N_995,N_728,N_671);
or U996 (N_996,N_698,N_774);
nand U997 (N_997,N_767,N_614);
xor U998 (N_998,N_796,N_624);
and U999 (N_999,N_658,N_746);
xor U1000 (N_1000,N_901,N_944);
xnor U1001 (N_1001,N_829,N_823);
nand U1002 (N_1002,N_894,N_980);
or U1003 (N_1003,N_983,N_819);
nand U1004 (N_1004,N_938,N_943);
nand U1005 (N_1005,N_878,N_916);
and U1006 (N_1006,N_842,N_923);
xor U1007 (N_1007,N_886,N_979);
nand U1008 (N_1008,N_847,N_942);
nand U1009 (N_1009,N_826,N_871);
and U1010 (N_1010,N_991,N_985);
and U1011 (N_1011,N_876,N_987);
nand U1012 (N_1012,N_899,N_904);
and U1013 (N_1013,N_990,N_867);
and U1014 (N_1014,N_900,N_828);
nand U1015 (N_1015,N_844,N_925);
nand U1016 (N_1016,N_947,N_814);
and U1017 (N_1017,N_855,N_965);
and U1018 (N_1018,N_888,N_946);
xor U1019 (N_1019,N_984,N_885);
and U1020 (N_1020,N_841,N_920);
xor U1021 (N_1021,N_875,N_800);
nand U1022 (N_1022,N_997,N_910);
xnor U1023 (N_1023,N_845,N_858);
xor U1024 (N_1024,N_902,N_941);
nor U1025 (N_1025,N_807,N_939);
nand U1026 (N_1026,N_884,N_966);
or U1027 (N_1027,N_957,N_958);
nand U1028 (N_1028,N_811,N_852);
nor U1029 (N_1029,N_860,N_869);
and U1030 (N_1030,N_940,N_896);
and U1031 (N_1031,N_935,N_952);
nor U1032 (N_1032,N_851,N_948);
xnor U1033 (N_1033,N_830,N_827);
xor U1034 (N_1034,N_953,N_812);
xnor U1035 (N_1035,N_839,N_908);
nand U1036 (N_1036,N_934,N_959);
nor U1037 (N_1037,N_868,N_950);
or U1038 (N_1038,N_872,N_915);
or U1039 (N_1039,N_955,N_808);
or U1040 (N_1040,N_994,N_913);
nor U1041 (N_1041,N_992,N_967);
nand U1042 (N_1042,N_893,N_975);
nor U1043 (N_1043,N_835,N_949);
and U1044 (N_1044,N_898,N_846);
xor U1045 (N_1045,N_906,N_929);
or U1046 (N_1046,N_854,N_971);
or U1047 (N_1047,N_870,N_936);
xnor U1048 (N_1048,N_905,N_882);
xnor U1049 (N_1049,N_801,N_804);
nor U1050 (N_1050,N_861,N_810);
or U1051 (N_1051,N_856,N_805);
nor U1052 (N_1052,N_892,N_977);
nor U1053 (N_1053,N_931,N_877);
or U1054 (N_1054,N_866,N_933);
xor U1055 (N_1055,N_802,N_821);
xor U1056 (N_1056,N_982,N_956);
or U1057 (N_1057,N_837,N_998);
nor U1058 (N_1058,N_817,N_917);
xnor U1059 (N_1059,N_895,N_849);
nor U1060 (N_1060,N_918,N_838);
and U1061 (N_1061,N_961,N_962);
or U1062 (N_1062,N_822,N_924);
or U1063 (N_1063,N_907,N_927);
and U1064 (N_1064,N_824,N_909);
and U1065 (N_1065,N_889,N_865);
nor U1066 (N_1066,N_996,N_825);
xnor U1067 (N_1067,N_863,N_848);
nor U1068 (N_1068,N_930,N_969);
and U1069 (N_1069,N_932,N_883);
nand U1070 (N_1070,N_911,N_981);
nor U1071 (N_1071,N_989,N_970);
xor U1072 (N_1072,N_926,N_862);
and U1073 (N_1073,N_857,N_963);
nor U1074 (N_1074,N_874,N_903);
or U1075 (N_1075,N_937,N_813);
nand U1076 (N_1076,N_864,N_880);
and U1077 (N_1077,N_978,N_836);
and U1078 (N_1078,N_891,N_974);
and U1079 (N_1079,N_831,N_954);
nand U1080 (N_1080,N_832,N_993);
xor U1081 (N_1081,N_890,N_815);
nand U1082 (N_1082,N_853,N_964);
nor U1083 (N_1083,N_818,N_897);
and U1084 (N_1084,N_945,N_973);
nand U1085 (N_1085,N_879,N_976);
or U1086 (N_1086,N_887,N_986);
nor U1087 (N_1087,N_951,N_921);
nor U1088 (N_1088,N_843,N_919);
and U1089 (N_1089,N_999,N_914);
nand U1090 (N_1090,N_928,N_995);
nor U1091 (N_1091,N_922,N_820);
and U1092 (N_1092,N_833,N_803);
nor U1093 (N_1093,N_873,N_912);
xor U1094 (N_1094,N_988,N_850);
or U1095 (N_1095,N_816,N_840);
nand U1096 (N_1096,N_809,N_859);
nand U1097 (N_1097,N_806,N_972);
nor U1098 (N_1098,N_960,N_834);
nand U1099 (N_1099,N_881,N_968);
nand U1100 (N_1100,N_813,N_994);
and U1101 (N_1101,N_854,N_896);
xnor U1102 (N_1102,N_868,N_969);
and U1103 (N_1103,N_905,N_988);
nor U1104 (N_1104,N_972,N_832);
xnor U1105 (N_1105,N_810,N_912);
and U1106 (N_1106,N_923,N_936);
xnor U1107 (N_1107,N_976,N_818);
xor U1108 (N_1108,N_928,N_831);
nand U1109 (N_1109,N_918,N_886);
or U1110 (N_1110,N_820,N_842);
nor U1111 (N_1111,N_902,N_961);
xor U1112 (N_1112,N_909,N_991);
nor U1113 (N_1113,N_877,N_938);
and U1114 (N_1114,N_870,N_996);
xor U1115 (N_1115,N_830,N_985);
and U1116 (N_1116,N_801,N_829);
xor U1117 (N_1117,N_894,N_914);
nand U1118 (N_1118,N_866,N_896);
nand U1119 (N_1119,N_827,N_912);
or U1120 (N_1120,N_971,N_906);
nor U1121 (N_1121,N_995,N_911);
nand U1122 (N_1122,N_817,N_955);
nand U1123 (N_1123,N_807,N_952);
and U1124 (N_1124,N_879,N_885);
nand U1125 (N_1125,N_824,N_801);
and U1126 (N_1126,N_947,N_895);
and U1127 (N_1127,N_894,N_919);
nor U1128 (N_1128,N_957,N_998);
and U1129 (N_1129,N_965,N_871);
nor U1130 (N_1130,N_911,N_953);
and U1131 (N_1131,N_868,N_819);
nand U1132 (N_1132,N_853,N_953);
and U1133 (N_1133,N_992,N_928);
or U1134 (N_1134,N_929,N_948);
or U1135 (N_1135,N_933,N_829);
nand U1136 (N_1136,N_936,N_913);
xnor U1137 (N_1137,N_975,N_963);
and U1138 (N_1138,N_855,N_906);
or U1139 (N_1139,N_905,N_817);
or U1140 (N_1140,N_996,N_844);
nand U1141 (N_1141,N_996,N_946);
nand U1142 (N_1142,N_867,N_858);
nand U1143 (N_1143,N_838,N_860);
nand U1144 (N_1144,N_890,N_936);
nor U1145 (N_1145,N_924,N_904);
xnor U1146 (N_1146,N_903,N_965);
nand U1147 (N_1147,N_927,N_862);
xor U1148 (N_1148,N_949,N_908);
xor U1149 (N_1149,N_963,N_972);
nor U1150 (N_1150,N_833,N_809);
xnor U1151 (N_1151,N_814,N_929);
nor U1152 (N_1152,N_908,N_848);
and U1153 (N_1153,N_936,N_924);
and U1154 (N_1154,N_805,N_874);
nand U1155 (N_1155,N_954,N_917);
and U1156 (N_1156,N_890,N_946);
or U1157 (N_1157,N_938,N_958);
nor U1158 (N_1158,N_845,N_895);
or U1159 (N_1159,N_938,N_927);
nor U1160 (N_1160,N_828,N_891);
and U1161 (N_1161,N_957,N_829);
or U1162 (N_1162,N_829,N_834);
and U1163 (N_1163,N_801,N_916);
and U1164 (N_1164,N_906,N_988);
nor U1165 (N_1165,N_933,N_957);
or U1166 (N_1166,N_907,N_854);
xnor U1167 (N_1167,N_906,N_859);
and U1168 (N_1168,N_879,N_914);
nand U1169 (N_1169,N_802,N_866);
nor U1170 (N_1170,N_841,N_842);
and U1171 (N_1171,N_891,N_880);
or U1172 (N_1172,N_828,N_896);
xor U1173 (N_1173,N_985,N_874);
nand U1174 (N_1174,N_823,N_806);
xnor U1175 (N_1175,N_988,N_954);
xor U1176 (N_1176,N_816,N_830);
nor U1177 (N_1177,N_802,N_874);
and U1178 (N_1178,N_964,N_971);
and U1179 (N_1179,N_843,N_846);
nor U1180 (N_1180,N_981,N_995);
nor U1181 (N_1181,N_986,N_930);
or U1182 (N_1182,N_918,N_807);
xor U1183 (N_1183,N_850,N_956);
nor U1184 (N_1184,N_980,N_925);
nand U1185 (N_1185,N_837,N_888);
and U1186 (N_1186,N_844,N_853);
or U1187 (N_1187,N_824,N_914);
or U1188 (N_1188,N_805,N_931);
nand U1189 (N_1189,N_995,N_945);
or U1190 (N_1190,N_842,N_984);
nand U1191 (N_1191,N_807,N_933);
nand U1192 (N_1192,N_831,N_842);
nand U1193 (N_1193,N_953,N_963);
xor U1194 (N_1194,N_923,N_905);
and U1195 (N_1195,N_837,N_928);
nor U1196 (N_1196,N_974,N_940);
nand U1197 (N_1197,N_819,N_891);
nand U1198 (N_1198,N_911,N_970);
or U1199 (N_1199,N_826,N_901);
xor U1200 (N_1200,N_1083,N_1148);
and U1201 (N_1201,N_1048,N_1017);
or U1202 (N_1202,N_1137,N_1061);
nor U1203 (N_1203,N_1098,N_1093);
or U1204 (N_1204,N_1167,N_1043);
xnor U1205 (N_1205,N_1127,N_1195);
nand U1206 (N_1206,N_1159,N_1006);
nor U1207 (N_1207,N_1193,N_1084);
xor U1208 (N_1208,N_1199,N_1066);
nor U1209 (N_1209,N_1038,N_1042);
nor U1210 (N_1210,N_1179,N_1082);
xor U1211 (N_1211,N_1001,N_1138);
nand U1212 (N_1212,N_1015,N_1079);
xor U1213 (N_1213,N_1026,N_1142);
nor U1214 (N_1214,N_1172,N_1099);
nand U1215 (N_1215,N_1040,N_1152);
or U1216 (N_1216,N_1019,N_1034);
and U1217 (N_1217,N_1182,N_1056);
xor U1218 (N_1218,N_1149,N_1071);
and U1219 (N_1219,N_1030,N_1129);
and U1220 (N_1220,N_1090,N_1065);
xnor U1221 (N_1221,N_1198,N_1119);
xnor U1222 (N_1222,N_1134,N_1155);
xor U1223 (N_1223,N_1097,N_1100);
and U1224 (N_1224,N_1184,N_1028);
nor U1225 (N_1225,N_1140,N_1116);
nand U1226 (N_1226,N_1133,N_1053);
or U1227 (N_1227,N_1151,N_1005);
xnor U1228 (N_1228,N_1135,N_1191);
xnor U1229 (N_1229,N_1096,N_1032);
xnor U1230 (N_1230,N_1020,N_1077);
nor U1231 (N_1231,N_1076,N_1080);
nor U1232 (N_1232,N_1009,N_1130);
nand U1233 (N_1233,N_1037,N_1108);
nand U1234 (N_1234,N_1059,N_1021);
nor U1235 (N_1235,N_1062,N_1194);
and U1236 (N_1236,N_1163,N_1041);
or U1237 (N_1237,N_1132,N_1058);
and U1238 (N_1238,N_1075,N_1057);
xor U1239 (N_1239,N_1143,N_1124);
or U1240 (N_1240,N_1016,N_1117);
and U1241 (N_1241,N_1039,N_1007);
and U1242 (N_1242,N_1035,N_1012);
nor U1243 (N_1243,N_1175,N_1153);
or U1244 (N_1244,N_1081,N_1114);
nand U1245 (N_1245,N_1121,N_1031);
or U1246 (N_1246,N_1085,N_1089);
and U1247 (N_1247,N_1045,N_1050);
nand U1248 (N_1248,N_1046,N_1189);
nor U1249 (N_1249,N_1073,N_1122);
nor U1250 (N_1250,N_1010,N_1144);
nand U1251 (N_1251,N_1023,N_1154);
xnor U1252 (N_1252,N_1025,N_1111);
nor U1253 (N_1253,N_1173,N_1150);
nor U1254 (N_1254,N_1139,N_1044);
nand U1255 (N_1255,N_1180,N_1051);
or U1256 (N_1256,N_1123,N_1008);
xor U1257 (N_1257,N_1105,N_1113);
or U1258 (N_1258,N_1092,N_1115);
xnor U1259 (N_1259,N_1107,N_1110);
or U1260 (N_1260,N_1064,N_1022);
or U1261 (N_1261,N_1029,N_1171);
nand U1262 (N_1262,N_1109,N_1049);
or U1263 (N_1263,N_1014,N_1055);
xor U1264 (N_1264,N_1147,N_1103);
and U1265 (N_1265,N_1169,N_1181);
nor U1266 (N_1266,N_1170,N_1087);
nand U1267 (N_1267,N_1146,N_1104);
nand U1268 (N_1268,N_1141,N_1131);
or U1269 (N_1269,N_1183,N_1166);
nor U1270 (N_1270,N_1156,N_1125);
or U1271 (N_1271,N_1190,N_1136);
xor U1272 (N_1272,N_1102,N_1091);
nand U1273 (N_1273,N_1013,N_1174);
nor U1274 (N_1274,N_1157,N_1024);
nor U1275 (N_1275,N_1018,N_1002);
or U1276 (N_1276,N_1088,N_1120);
nand U1277 (N_1277,N_1186,N_1101);
nand U1278 (N_1278,N_1067,N_1086);
nor U1279 (N_1279,N_1161,N_1078);
or U1280 (N_1280,N_1011,N_1095);
and U1281 (N_1281,N_1192,N_1187);
nand U1282 (N_1282,N_1072,N_1145);
and U1283 (N_1283,N_1188,N_1070);
xnor U1284 (N_1284,N_1000,N_1074);
nand U1285 (N_1285,N_1165,N_1036);
nand U1286 (N_1286,N_1185,N_1004);
nor U1287 (N_1287,N_1158,N_1162);
and U1288 (N_1288,N_1118,N_1069);
xor U1289 (N_1289,N_1094,N_1176);
xor U1290 (N_1290,N_1106,N_1063);
xnor U1291 (N_1291,N_1160,N_1060);
or U1292 (N_1292,N_1054,N_1027);
nor U1293 (N_1293,N_1168,N_1178);
xnor U1294 (N_1294,N_1128,N_1196);
and U1295 (N_1295,N_1068,N_1112);
xnor U1296 (N_1296,N_1047,N_1052);
or U1297 (N_1297,N_1126,N_1177);
and U1298 (N_1298,N_1033,N_1197);
xnor U1299 (N_1299,N_1164,N_1003);
nand U1300 (N_1300,N_1176,N_1141);
or U1301 (N_1301,N_1159,N_1120);
nor U1302 (N_1302,N_1179,N_1015);
and U1303 (N_1303,N_1182,N_1034);
nor U1304 (N_1304,N_1017,N_1035);
nor U1305 (N_1305,N_1159,N_1093);
xor U1306 (N_1306,N_1091,N_1048);
xor U1307 (N_1307,N_1008,N_1051);
nand U1308 (N_1308,N_1075,N_1182);
or U1309 (N_1309,N_1025,N_1092);
and U1310 (N_1310,N_1047,N_1061);
nor U1311 (N_1311,N_1138,N_1132);
and U1312 (N_1312,N_1036,N_1060);
and U1313 (N_1313,N_1112,N_1153);
nor U1314 (N_1314,N_1049,N_1157);
and U1315 (N_1315,N_1109,N_1139);
or U1316 (N_1316,N_1009,N_1092);
xor U1317 (N_1317,N_1158,N_1108);
nor U1318 (N_1318,N_1150,N_1041);
nand U1319 (N_1319,N_1047,N_1119);
or U1320 (N_1320,N_1157,N_1048);
xor U1321 (N_1321,N_1003,N_1119);
or U1322 (N_1322,N_1065,N_1190);
nand U1323 (N_1323,N_1139,N_1169);
nor U1324 (N_1324,N_1087,N_1004);
nor U1325 (N_1325,N_1052,N_1132);
or U1326 (N_1326,N_1195,N_1027);
xnor U1327 (N_1327,N_1068,N_1022);
xnor U1328 (N_1328,N_1082,N_1064);
and U1329 (N_1329,N_1116,N_1059);
xor U1330 (N_1330,N_1113,N_1015);
nand U1331 (N_1331,N_1081,N_1052);
nor U1332 (N_1332,N_1032,N_1092);
nand U1333 (N_1333,N_1092,N_1019);
or U1334 (N_1334,N_1073,N_1056);
xor U1335 (N_1335,N_1174,N_1165);
and U1336 (N_1336,N_1109,N_1191);
xor U1337 (N_1337,N_1178,N_1103);
or U1338 (N_1338,N_1005,N_1146);
or U1339 (N_1339,N_1163,N_1111);
xnor U1340 (N_1340,N_1055,N_1022);
xor U1341 (N_1341,N_1187,N_1120);
xor U1342 (N_1342,N_1150,N_1171);
nand U1343 (N_1343,N_1156,N_1078);
xnor U1344 (N_1344,N_1044,N_1196);
nand U1345 (N_1345,N_1135,N_1033);
and U1346 (N_1346,N_1154,N_1086);
or U1347 (N_1347,N_1080,N_1065);
and U1348 (N_1348,N_1061,N_1073);
xor U1349 (N_1349,N_1144,N_1184);
xor U1350 (N_1350,N_1037,N_1078);
or U1351 (N_1351,N_1194,N_1153);
xnor U1352 (N_1352,N_1179,N_1051);
xnor U1353 (N_1353,N_1043,N_1178);
nand U1354 (N_1354,N_1109,N_1127);
nor U1355 (N_1355,N_1127,N_1105);
xor U1356 (N_1356,N_1124,N_1035);
nand U1357 (N_1357,N_1036,N_1083);
nand U1358 (N_1358,N_1051,N_1136);
or U1359 (N_1359,N_1008,N_1099);
nand U1360 (N_1360,N_1198,N_1187);
xor U1361 (N_1361,N_1174,N_1168);
or U1362 (N_1362,N_1159,N_1128);
or U1363 (N_1363,N_1005,N_1046);
and U1364 (N_1364,N_1179,N_1169);
nand U1365 (N_1365,N_1147,N_1159);
and U1366 (N_1366,N_1158,N_1090);
nor U1367 (N_1367,N_1076,N_1125);
and U1368 (N_1368,N_1063,N_1027);
nand U1369 (N_1369,N_1091,N_1021);
or U1370 (N_1370,N_1078,N_1041);
or U1371 (N_1371,N_1022,N_1101);
nand U1372 (N_1372,N_1155,N_1010);
xnor U1373 (N_1373,N_1142,N_1028);
and U1374 (N_1374,N_1199,N_1114);
nor U1375 (N_1375,N_1126,N_1123);
and U1376 (N_1376,N_1011,N_1158);
xnor U1377 (N_1377,N_1046,N_1108);
nor U1378 (N_1378,N_1009,N_1011);
xor U1379 (N_1379,N_1050,N_1067);
nor U1380 (N_1380,N_1194,N_1004);
or U1381 (N_1381,N_1003,N_1144);
or U1382 (N_1382,N_1104,N_1162);
and U1383 (N_1383,N_1020,N_1060);
or U1384 (N_1384,N_1158,N_1173);
nor U1385 (N_1385,N_1020,N_1061);
nor U1386 (N_1386,N_1039,N_1166);
xor U1387 (N_1387,N_1051,N_1127);
or U1388 (N_1388,N_1169,N_1077);
xnor U1389 (N_1389,N_1032,N_1161);
nor U1390 (N_1390,N_1150,N_1181);
and U1391 (N_1391,N_1085,N_1130);
nor U1392 (N_1392,N_1164,N_1032);
and U1393 (N_1393,N_1137,N_1069);
and U1394 (N_1394,N_1072,N_1069);
xor U1395 (N_1395,N_1174,N_1003);
xor U1396 (N_1396,N_1089,N_1106);
and U1397 (N_1397,N_1180,N_1167);
nand U1398 (N_1398,N_1115,N_1094);
xnor U1399 (N_1399,N_1013,N_1083);
and U1400 (N_1400,N_1317,N_1376);
nand U1401 (N_1401,N_1314,N_1291);
xnor U1402 (N_1402,N_1223,N_1265);
and U1403 (N_1403,N_1312,N_1390);
xnor U1404 (N_1404,N_1283,N_1246);
nor U1405 (N_1405,N_1386,N_1353);
xor U1406 (N_1406,N_1214,N_1228);
and U1407 (N_1407,N_1266,N_1289);
or U1408 (N_1408,N_1360,N_1329);
nor U1409 (N_1409,N_1320,N_1319);
xor U1410 (N_1410,N_1279,N_1315);
nand U1411 (N_1411,N_1292,N_1322);
or U1412 (N_1412,N_1389,N_1334);
and U1413 (N_1413,N_1299,N_1337);
nor U1414 (N_1414,N_1254,N_1395);
xor U1415 (N_1415,N_1318,N_1260);
and U1416 (N_1416,N_1234,N_1298);
xnor U1417 (N_1417,N_1288,N_1355);
xor U1418 (N_1418,N_1230,N_1392);
or U1419 (N_1419,N_1374,N_1364);
nor U1420 (N_1420,N_1216,N_1206);
xnor U1421 (N_1421,N_1211,N_1335);
xor U1422 (N_1422,N_1350,N_1370);
and U1423 (N_1423,N_1397,N_1294);
or U1424 (N_1424,N_1222,N_1250);
nor U1425 (N_1425,N_1371,N_1224);
nor U1426 (N_1426,N_1287,N_1356);
and U1427 (N_1427,N_1316,N_1278);
xor U1428 (N_1428,N_1351,N_1217);
or U1429 (N_1429,N_1380,N_1307);
or U1430 (N_1430,N_1375,N_1382);
and U1431 (N_1431,N_1241,N_1269);
nand U1432 (N_1432,N_1236,N_1237);
xnor U1433 (N_1433,N_1311,N_1306);
and U1434 (N_1434,N_1226,N_1367);
xnor U1435 (N_1435,N_1203,N_1282);
and U1436 (N_1436,N_1379,N_1385);
nand U1437 (N_1437,N_1251,N_1202);
nand U1438 (N_1438,N_1256,N_1340);
or U1439 (N_1439,N_1273,N_1247);
xnor U1440 (N_1440,N_1276,N_1277);
and U1441 (N_1441,N_1381,N_1387);
nor U1442 (N_1442,N_1394,N_1308);
and U1443 (N_1443,N_1272,N_1301);
nor U1444 (N_1444,N_1200,N_1391);
xor U1445 (N_1445,N_1366,N_1270);
or U1446 (N_1446,N_1255,N_1284);
and U1447 (N_1447,N_1285,N_1232);
nand U1448 (N_1448,N_1330,N_1238);
xor U1449 (N_1449,N_1264,N_1268);
and U1450 (N_1450,N_1348,N_1290);
nand U1451 (N_1451,N_1327,N_1243);
nand U1452 (N_1452,N_1369,N_1338);
nor U1453 (N_1453,N_1219,N_1281);
nand U1454 (N_1454,N_1296,N_1349);
and U1455 (N_1455,N_1305,N_1257);
nand U1456 (N_1456,N_1235,N_1336);
or U1457 (N_1457,N_1295,N_1297);
and U1458 (N_1458,N_1333,N_1332);
nor U1459 (N_1459,N_1212,N_1258);
nor U1460 (N_1460,N_1209,N_1262);
nor U1461 (N_1461,N_1384,N_1252);
nand U1462 (N_1462,N_1259,N_1229);
nor U1463 (N_1463,N_1242,N_1261);
and U1464 (N_1464,N_1221,N_1275);
nor U1465 (N_1465,N_1368,N_1293);
xnor U1466 (N_1466,N_1204,N_1205);
or U1467 (N_1467,N_1331,N_1398);
nand U1468 (N_1468,N_1267,N_1303);
or U1469 (N_1469,N_1325,N_1339);
or U1470 (N_1470,N_1358,N_1313);
nand U1471 (N_1471,N_1309,N_1324);
nand U1472 (N_1472,N_1342,N_1343);
nor U1473 (N_1473,N_1341,N_1207);
and U1474 (N_1474,N_1304,N_1245);
or U1475 (N_1475,N_1344,N_1365);
xnor U1476 (N_1476,N_1263,N_1399);
nand U1477 (N_1477,N_1328,N_1210);
nor U1478 (N_1478,N_1346,N_1218);
xor U1479 (N_1479,N_1326,N_1213);
and U1480 (N_1480,N_1363,N_1357);
xnor U1481 (N_1481,N_1244,N_1227);
nor U1482 (N_1482,N_1347,N_1373);
nor U1483 (N_1483,N_1396,N_1388);
or U1484 (N_1484,N_1359,N_1208);
nor U1485 (N_1485,N_1361,N_1215);
xor U1486 (N_1486,N_1372,N_1280);
xnor U1487 (N_1487,N_1393,N_1239);
or U1488 (N_1488,N_1248,N_1354);
and U1489 (N_1489,N_1286,N_1271);
nand U1490 (N_1490,N_1201,N_1231);
xor U1491 (N_1491,N_1225,N_1233);
nand U1492 (N_1492,N_1377,N_1378);
and U1493 (N_1493,N_1249,N_1383);
and U1494 (N_1494,N_1220,N_1321);
and U1495 (N_1495,N_1253,N_1302);
nand U1496 (N_1496,N_1362,N_1323);
nand U1497 (N_1497,N_1300,N_1345);
and U1498 (N_1498,N_1240,N_1352);
nand U1499 (N_1499,N_1274,N_1310);
and U1500 (N_1500,N_1377,N_1270);
nand U1501 (N_1501,N_1275,N_1395);
or U1502 (N_1502,N_1389,N_1204);
nand U1503 (N_1503,N_1260,N_1365);
nand U1504 (N_1504,N_1208,N_1368);
nor U1505 (N_1505,N_1368,N_1228);
and U1506 (N_1506,N_1294,N_1365);
xor U1507 (N_1507,N_1257,N_1256);
xor U1508 (N_1508,N_1326,N_1311);
nor U1509 (N_1509,N_1230,N_1235);
or U1510 (N_1510,N_1215,N_1228);
nor U1511 (N_1511,N_1385,N_1279);
and U1512 (N_1512,N_1296,N_1301);
nor U1513 (N_1513,N_1262,N_1330);
xor U1514 (N_1514,N_1347,N_1336);
nor U1515 (N_1515,N_1311,N_1249);
xor U1516 (N_1516,N_1265,N_1374);
or U1517 (N_1517,N_1316,N_1382);
nand U1518 (N_1518,N_1383,N_1216);
and U1519 (N_1519,N_1308,N_1330);
or U1520 (N_1520,N_1276,N_1379);
or U1521 (N_1521,N_1287,N_1216);
xnor U1522 (N_1522,N_1328,N_1313);
nor U1523 (N_1523,N_1321,N_1239);
and U1524 (N_1524,N_1285,N_1383);
nand U1525 (N_1525,N_1376,N_1218);
nor U1526 (N_1526,N_1386,N_1325);
nand U1527 (N_1527,N_1218,N_1384);
nand U1528 (N_1528,N_1256,N_1219);
and U1529 (N_1529,N_1277,N_1221);
or U1530 (N_1530,N_1248,N_1210);
and U1531 (N_1531,N_1268,N_1263);
xor U1532 (N_1532,N_1315,N_1398);
and U1533 (N_1533,N_1253,N_1380);
and U1534 (N_1534,N_1216,N_1397);
xnor U1535 (N_1535,N_1311,N_1263);
nor U1536 (N_1536,N_1349,N_1255);
xor U1537 (N_1537,N_1346,N_1377);
xor U1538 (N_1538,N_1242,N_1379);
nor U1539 (N_1539,N_1221,N_1351);
nand U1540 (N_1540,N_1297,N_1283);
xnor U1541 (N_1541,N_1241,N_1280);
xnor U1542 (N_1542,N_1293,N_1372);
and U1543 (N_1543,N_1357,N_1259);
nor U1544 (N_1544,N_1268,N_1230);
nand U1545 (N_1545,N_1229,N_1329);
xnor U1546 (N_1546,N_1364,N_1275);
or U1547 (N_1547,N_1207,N_1210);
or U1548 (N_1548,N_1346,N_1365);
xnor U1549 (N_1549,N_1208,N_1398);
nor U1550 (N_1550,N_1331,N_1277);
or U1551 (N_1551,N_1257,N_1347);
xor U1552 (N_1552,N_1202,N_1343);
or U1553 (N_1553,N_1362,N_1342);
and U1554 (N_1554,N_1229,N_1249);
and U1555 (N_1555,N_1383,N_1209);
or U1556 (N_1556,N_1253,N_1264);
nand U1557 (N_1557,N_1218,N_1265);
or U1558 (N_1558,N_1387,N_1226);
xnor U1559 (N_1559,N_1293,N_1274);
or U1560 (N_1560,N_1295,N_1311);
or U1561 (N_1561,N_1393,N_1263);
and U1562 (N_1562,N_1338,N_1269);
and U1563 (N_1563,N_1319,N_1333);
and U1564 (N_1564,N_1225,N_1215);
nand U1565 (N_1565,N_1398,N_1371);
nor U1566 (N_1566,N_1266,N_1310);
nor U1567 (N_1567,N_1224,N_1325);
nand U1568 (N_1568,N_1303,N_1399);
and U1569 (N_1569,N_1335,N_1218);
and U1570 (N_1570,N_1250,N_1344);
nor U1571 (N_1571,N_1304,N_1365);
xnor U1572 (N_1572,N_1303,N_1398);
or U1573 (N_1573,N_1365,N_1310);
nand U1574 (N_1574,N_1341,N_1236);
nand U1575 (N_1575,N_1215,N_1299);
nand U1576 (N_1576,N_1337,N_1242);
nand U1577 (N_1577,N_1251,N_1393);
xnor U1578 (N_1578,N_1358,N_1327);
nand U1579 (N_1579,N_1321,N_1356);
nor U1580 (N_1580,N_1390,N_1205);
nor U1581 (N_1581,N_1347,N_1296);
nor U1582 (N_1582,N_1268,N_1381);
xnor U1583 (N_1583,N_1381,N_1295);
xnor U1584 (N_1584,N_1365,N_1206);
nor U1585 (N_1585,N_1260,N_1381);
xor U1586 (N_1586,N_1272,N_1205);
or U1587 (N_1587,N_1230,N_1247);
nor U1588 (N_1588,N_1251,N_1292);
or U1589 (N_1589,N_1327,N_1217);
nand U1590 (N_1590,N_1229,N_1217);
or U1591 (N_1591,N_1267,N_1294);
nand U1592 (N_1592,N_1366,N_1364);
nand U1593 (N_1593,N_1227,N_1294);
nand U1594 (N_1594,N_1249,N_1395);
xor U1595 (N_1595,N_1365,N_1208);
xnor U1596 (N_1596,N_1242,N_1223);
nor U1597 (N_1597,N_1288,N_1325);
or U1598 (N_1598,N_1313,N_1316);
nand U1599 (N_1599,N_1253,N_1285);
or U1600 (N_1600,N_1558,N_1517);
nor U1601 (N_1601,N_1505,N_1570);
nor U1602 (N_1602,N_1457,N_1443);
nand U1603 (N_1603,N_1497,N_1516);
and U1604 (N_1604,N_1593,N_1592);
or U1605 (N_1605,N_1445,N_1458);
nor U1606 (N_1606,N_1486,N_1484);
and U1607 (N_1607,N_1571,N_1488);
nor U1608 (N_1608,N_1479,N_1544);
xor U1609 (N_1609,N_1524,N_1575);
and U1610 (N_1610,N_1401,N_1562);
xor U1611 (N_1611,N_1533,N_1491);
xor U1612 (N_1612,N_1446,N_1563);
and U1613 (N_1613,N_1549,N_1435);
and U1614 (N_1614,N_1480,N_1599);
nand U1615 (N_1615,N_1560,N_1509);
or U1616 (N_1616,N_1566,N_1522);
xor U1617 (N_1617,N_1536,N_1415);
and U1618 (N_1618,N_1559,N_1440);
xor U1619 (N_1619,N_1545,N_1568);
xor U1620 (N_1620,N_1438,N_1459);
nand U1621 (N_1621,N_1462,N_1402);
nor U1622 (N_1622,N_1431,N_1472);
and U1623 (N_1623,N_1535,N_1573);
xor U1624 (N_1624,N_1501,N_1555);
nand U1625 (N_1625,N_1531,N_1481);
xor U1626 (N_1626,N_1430,N_1450);
nand U1627 (N_1627,N_1574,N_1529);
or U1628 (N_1628,N_1520,N_1543);
nand U1629 (N_1629,N_1437,N_1478);
nor U1630 (N_1630,N_1589,N_1546);
xor U1631 (N_1631,N_1419,N_1407);
nor U1632 (N_1632,N_1406,N_1540);
nand U1633 (N_1633,N_1569,N_1539);
xnor U1634 (N_1634,N_1429,N_1493);
or U1635 (N_1635,N_1580,N_1565);
nand U1636 (N_1636,N_1495,N_1409);
nor U1637 (N_1637,N_1485,N_1477);
or U1638 (N_1638,N_1556,N_1586);
or U1639 (N_1639,N_1405,N_1578);
or U1640 (N_1640,N_1439,N_1494);
and U1641 (N_1641,N_1567,N_1417);
or U1642 (N_1642,N_1404,N_1500);
or U1643 (N_1643,N_1475,N_1428);
and U1644 (N_1644,N_1597,N_1548);
xnor U1645 (N_1645,N_1427,N_1499);
xnor U1646 (N_1646,N_1461,N_1526);
nand U1647 (N_1647,N_1518,N_1418);
and U1648 (N_1648,N_1442,N_1411);
nand U1649 (N_1649,N_1523,N_1420);
and U1650 (N_1650,N_1572,N_1421);
nand U1651 (N_1651,N_1508,N_1595);
nand U1652 (N_1652,N_1513,N_1576);
nand U1653 (N_1653,N_1554,N_1583);
nand U1654 (N_1654,N_1528,N_1542);
and U1655 (N_1655,N_1470,N_1504);
and U1656 (N_1656,N_1534,N_1482);
nor U1657 (N_1657,N_1553,N_1432);
nand U1658 (N_1658,N_1473,N_1521);
or U1659 (N_1659,N_1519,N_1577);
nand U1660 (N_1660,N_1424,N_1506);
nor U1661 (N_1661,N_1502,N_1403);
or U1662 (N_1662,N_1408,N_1483);
nand U1663 (N_1663,N_1468,N_1579);
or U1664 (N_1664,N_1551,N_1585);
nor U1665 (N_1665,N_1474,N_1465);
or U1666 (N_1666,N_1464,N_1448);
nand U1667 (N_1667,N_1423,N_1496);
nor U1668 (N_1668,N_1444,N_1591);
and U1669 (N_1669,N_1498,N_1489);
nand U1670 (N_1670,N_1453,N_1425);
and U1671 (N_1671,N_1532,N_1550);
xnor U1672 (N_1672,N_1564,N_1416);
and U1673 (N_1673,N_1503,N_1434);
or U1674 (N_1674,N_1525,N_1594);
xor U1675 (N_1675,N_1463,N_1512);
nand U1676 (N_1676,N_1584,N_1441);
or U1677 (N_1677,N_1460,N_1541);
or U1678 (N_1678,N_1452,N_1436);
xnor U1679 (N_1679,N_1487,N_1456);
and U1680 (N_1680,N_1414,N_1507);
or U1681 (N_1681,N_1582,N_1400);
nand U1682 (N_1682,N_1588,N_1537);
nand U1683 (N_1683,N_1467,N_1590);
nor U1684 (N_1684,N_1469,N_1596);
nand U1685 (N_1685,N_1547,N_1426);
and U1686 (N_1686,N_1492,N_1433);
and U1687 (N_1687,N_1581,N_1412);
and U1688 (N_1688,N_1413,N_1514);
nor U1689 (N_1689,N_1561,N_1476);
nand U1690 (N_1690,N_1587,N_1451);
or U1691 (N_1691,N_1538,N_1557);
xnor U1692 (N_1692,N_1422,N_1552);
xnor U1693 (N_1693,N_1510,N_1410);
nand U1694 (N_1694,N_1527,N_1454);
or U1695 (N_1695,N_1471,N_1515);
or U1696 (N_1696,N_1598,N_1449);
nor U1697 (N_1697,N_1530,N_1466);
xor U1698 (N_1698,N_1511,N_1490);
xor U1699 (N_1699,N_1447,N_1455);
nor U1700 (N_1700,N_1425,N_1516);
nand U1701 (N_1701,N_1439,N_1496);
nand U1702 (N_1702,N_1448,N_1405);
and U1703 (N_1703,N_1487,N_1435);
and U1704 (N_1704,N_1420,N_1490);
and U1705 (N_1705,N_1514,N_1478);
xor U1706 (N_1706,N_1468,N_1542);
and U1707 (N_1707,N_1468,N_1567);
nor U1708 (N_1708,N_1525,N_1515);
and U1709 (N_1709,N_1578,N_1580);
nor U1710 (N_1710,N_1411,N_1502);
nand U1711 (N_1711,N_1555,N_1486);
xor U1712 (N_1712,N_1569,N_1513);
xnor U1713 (N_1713,N_1427,N_1436);
nor U1714 (N_1714,N_1522,N_1598);
nor U1715 (N_1715,N_1462,N_1540);
or U1716 (N_1716,N_1456,N_1428);
xnor U1717 (N_1717,N_1518,N_1578);
xnor U1718 (N_1718,N_1551,N_1440);
or U1719 (N_1719,N_1594,N_1572);
nand U1720 (N_1720,N_1449,N_1423);
nand U1721 (N_1721,N_1400,N_1513);
nor U1722 (N_1722,N_1468,N_1524);
and U1723 (N_1723,N_1524,N_1567);
or U1724 (N_1724,N_1574,N_1487);
or U1725 (N_1725,N_1555,N_1432);
xor U1726 (N_1726,N_1424,N_1544);
and U1727 (N_1727,N_1438,N_1555);
nor U1728 (N_1728,N_1544,N_1541);
xor U1729 (N_1729,N_1537,N_1467);
and U1730 (N_1730,N_1592,N_1426);
or U1731 (N_1731,N_1489,N_1412);
xor U1732 (N_1732,N_1541,N_1492);
and U1733 (N_1733,N_1484,N_1489);
or U1734 (N_1734,N_1488,N_1449);
or U1735 (N_1735,N_1472,N_1461);
nor U1736 (N_1736,N_1535,N_1401);
nor U1737 (N_1737,N_1506,N_1590);
nor U1738 (N_1738,N_1439,N_1437);
and U1739 (N_1739,N_1482,N_1450);
or U1740 (N_1740,N_1513,N_1557);
xor U1741 (N_1741,N_1446,N_1498);
nand U1742 (N_1742,N_1495,N_1471);
or U1743 (N_1743,N_1474,N_1540);
xor U1744 (N_1744,N_1508,N_1485);
nand U1745 (N_1745,N_1402,N_1503);
and U1746 (N_1746,N_1571,N_1591);
and U1747 (N_1747,N_1540,N_1592);
nor U1748 (N_1748,N_1536,N_1599);
xor U1749 (N_1749,N_1510,N_1541);
nand U1750 (N_1750,N_1507,N_1494);
nand U1751 (N_1751,N_1525,N_1405);
or U1752 (N_1752,N_1520,N_1512);
nor U1753 (N_1753,N_1566,N_1504);
nand U1754 (N_1754,N_1436,N_1447);
nand U1755 (N_1755,N_1403,N_1450);
xor U1756 (N_1756,N_1565,N_1547);
or U1757 (N_1757,N_1563,N_1513);
nand U1758 (N_1758,N_1463,N_1452);
xor U1759 (N_1759,N_1403,N_1544);
and U1760 (N_1760,N_1544,N_1431);
nor U1761 (N_1761,N_1506,N_1584);
or U1762 (N_1762,N_1440,N_1535);
xnor U1763 (N_1763,N_1494,N_1470);
and U1764 (N_1764,N_1486,N_1574);
and U1765 (N_1765,N_1562,N_1579);
nand U1766 (N_1766,N_1409,N_1445);
and U1767 (N_1767,N_1534,N_1542);
nor U1768 (N_1768,N_1578,N_1441);
xor U1769 (N_1769,N_1411,N_1584);
nor U1770 (N_1770,N_1432,N_1440);
xor U1771 (N_1771,N_1465,N_1557);
nand U1772 (N_1772,N_1458,N_1473);
nand U1773 (N_1773,N_1546,N_1403);
nor U1774 (N_1774,N_1561,N_1527);
nand U1775 (N_1775,N_1491,N_1473);
and U1776 (N_1776,N_1523,N_1506);
nor U1777 (N_1777,N_1574,N_1458);
or U1778 (N_1778,N_1445,N_1419);
nand U1779 (N_1779,N_1483,N_1467);
or U1780 (N_1780,N_1477,N_1553);
xnor U1781 (N_1781,N_1559,N_1483);
xnor U1782 (N_1782,N_1447,N_1578);
or U1783 (N_1783,N_1573,N_1565);
xnor U1784 (N_1784,N_1453,N_1585);
nor U1785 (N_1785,N_1591,N_1442);
and U1786 (N_1786,N_1427,N_1584);
nand U1787 (N_1787,N_1484,N_1562);
nand U1788 (N_1788,N_1432,N_1488);
xnor U1789 (N_1789,N_1561,N_1405);
nand U1790 (N_1790,N_1558,N_1597);
nand U1791 (N_1791,N_1442,N_1514);
xor U1792 (N_1792,N_1485,N_1553);
or U1793 (N_1793,N_1485,N_1536);
or U1794 (N_1794,N_1414,N_1489);
and U1795 (N_1795,N_1513,N_1438);
or U1796 (N_1796,N_1535,N_1592);
nor U1797 (N_1797,N_1478,N_1598);
and U1798 (N_1798,N_1485,N_1479);
and U1799 (N_1799,N_1588,N_1527);
and U1800 (N_1800,N_1746,N_1619);
xor U1801 (N_1801,N_1623,N_1689);
or U1802 (N_1802,N_1693,N_1615);
or U1803 (N_1803,N_1650,N_1797);
xnor U1804 (N_1804,N_1699,N_1788);
or U1805 (N_1805,N_1755,N_1757);
or U1806 (N_1806,N_1708,N_1782);
xor U1807 (N_1807,N_1769,N_1696);
nor U1808 (N_1808,N_1784,N_1751);
nand U1809 (N_1809,N_1741,N_1601);
xnor U1810 (N_1810,N_1780,N_1799);
xor U1811 (N_1811,N_1733,N_1673);
and U1812 (N_1812,N_1743,N_1710);
and U1813 (N_1813,N_1632,N_1729);
nand U1814 (N_1814,N_1717,N_1759);
nand U1815 (N_1815,N_1770,N_1690);
nand U1816 (N_1816,N_1677,N_1613);
or U1817 (N_1817,N_1676,N_1672);
and U1818 (N_1818,N_1630,N_1791);
nand U1819 (N_1819,N_1728,N_1687);
nor U1820 (N_1820,N_1771,N_1698);
nor U1821 (N_1821,N_1686,N_1727);
and U1822 (N_1822,N_1656,N_1719);
xnor U1823 (N_1823,N_1684,N_1754);
or U1824 (N_1824,N_1787,N_1716);
or U1825 (N_1825,N_1685,N_1767);
or U1826 (N_1826,N_1622,N_1721);
xor U1827 (N_1827,N_1658,N_1645);
and U1828 (N_1828,N_1776,N_1709);
nor U1829 (N_1829,N_1660,N_1648);
nor U1830 (N_1830,N_1760,N_1665);
or U1831 (N_1831,N_1726,N_1705);
xnor U1832 (N_1832,N_1740,N_1643);
and U1833 (N_1833,N_1725,N_1775);
xor U1834 (N_1834,N_1627,N_1723);
and U1835 (N_1835,N_1704,N_1796);
nand U1836 (N_1836,N_1683,N_1611);
xnor U1837 (N_1837,N_1637,N_1793);
nor U1838 (N_1838,N_1764,N_1612);
xnor U1839 (N_1839,N_1748,N_1662);
nand U1840 (N_1840,N_1737,N_1608);
xnor U1841 (N_1841,N_1702,N_1634);
or U1842 (N_1842,N_1607,N_1681);
nand U1843 (N_1843,N_1640,N_1625);
xor U1844 (N_1844,N_1654,N_1605);
nand U1845 (N_1845,N_1786,N_1669);
and U1846 (N_1846,N_1688,N_1701);
or U1847 (N_1847,N_1626,N_1621);
and U1848 (N_1848,N_1715,N_1651);
nand U1849 (N_1849,N_1628,N_1659);
nor U1850 (N_1850,N_1722,N_1620);
or U1851 (N_1851,N_1629,N_1617);
nand U1852 (N_1852,N_1785,N_1778);
and U1853 (N_1853,N_1711,N_1609);
or U1854 (N_1854,N_1670,N_1649);
xor U1855 (N_1855,N_1739,N_1720);
xnor U1856 (N_1856,N_1795,N_1694);
or U1857 (N_1857,N_1638,N_1682);
or U1858 (N_1858,N_1730,N_1766);
and U1859 (N_1859,N_1697,N_1735);
and U1860 (N_1860,N_1783,N_1652);
nand U1861 (N_1861,N_1789,N_1745);
nand U1862 (N_1862,N_1762,N_1606);
xnor U1863 (N_1863,N_1792,N_1646);
nand U1864 (N_1864,N_1678,N_1765);
nand U1865 (N_1865,N_1674,N_1668);
or U1866 (N_1866,N_1761,N_1680);
xor U1867 (N_1867,N_1753,N_1604);
and U1868 (N_1868,N_1712,N_1758);
nor U1869 (N_1869,N_1706,N_1768);
nand U1870 (N_1870,N_1675,N_1616);
xor U1871 (N_1871,N_1664,N_1666);
nor U1872 (N_1872,N_1731,N_1714);
and U1873 (N_1873,N_1752,N_1653);
nand U1874 (N_1874,N_1631,N_1750);
or U1875 (N_1875,N_1772,N_1774);
nor U1876 (N_1876,N_1790,N_1661);
nand U1877 (N_1877,N_1713,N_1749);
nor U1878 (N_1878,N_1742,N_1647);
or U1879 (N_1879,N_1667,N_1779);
or U1880 (N_1880,N_1618,N_1614);
and U1881 (N_1881,N_1734,N_1600);
and U1882 (N_1882,N_1691,N_1657);
nand U1883 (N_1883,N_1692,N_1756);
nand U1884 (N_1884,N_1736,N_1707);
and U1885 (N_1885,N_1671,N_1624);
or U1886 (N_1886,N_1700,N_1738);
nand U1887 (N_1887,N_1703,N_1603);
nor U1888 (N_1888,N_1747,N_1777);
xor U1889 (N_1889,N_1794,N_1642);
xor U1890 (N_1890,N_1635,N_1724);
or U1891 (N_1891,N_1633,N_1655);
or U1892 (N_1892,N_1732,N_1602);
nor U1893 (N_1893,N_1798,N_1773);
nor U1894 (N_1894,N_1744,N_1636);
xor U1895 (N_1895,N_1695,N_1679);
nand U1896 (N_1896,N_1639,N_1781);
and U1897 (N_1897,N_1641,N_1610);
xor U1898 (N_1898,N_1644,N_1763);
xnor U1899 (N_1899,N_1663,N_1718);
nand U1900 (N_1900,N_1719,N_1798);
nor U1901 (N_1901,N_1658,N_1797);
nand U1902 (N_1902,N_1621,N_1784);
nand U1903 (N_1903,N_1675,N_1796);
nand U1904 (N_1904,N_1662,N_1797);
nor U1905 (N_1905,N_1602,N_1789);
nor U1906 (N_1906,N_1721,N_1725);
or U1907 (N_1907,N_1729,N_1615);
xnor U1908 (N_1908,N_1690,N_1627);
xnor U1909 (N_1909,N_1693,N_1612);
nand U1910 (N_1910,N_1623,N_1660);
nor U1911 (N_1911,N_1608,N_1702);
xnor U1912 (N_1912,N_1708,N_1679);
or U1913 (N_1913,N_1699,N_1679);
and U1914 (N_1914,N_1651,N_1702);
xnor U1915 (N_1915,N_1734,N_1616);
and U1916 (N_1916,N_1772,N_1669);
and U1917 (N_1917,N_1651,N_1602);
nor U1918 (N_1918,N_1778,N_1794);
nand U1919 (N_1919,N_1714,N_1779);
and U1920 (N_1920,N_1646,N_1720);
or U1921 (N_1921,N_1676,N_1716);
nand U1922 (N_1922,N_1619,N_1714);
and U1923 (N_1923,N_1722,N_1635);
nor U1924 (N_1924,N_1669,N_1613);
xnor U1925 (N_1925,N_1645,N_1716);
and U1926 (N_1926,N_1793,N_1727);
nor U1927 (N_1927,N_1794,N_1656);
nor U1928 (N_1928,N_1757,N_1751);
nand U1929 (N_1929,N_1669,N_1606);
and U1930 (N_1930,N_1750,N_1698);
and U1931 (N_1931,N_1707,N_1663);
or U1932 (N_1932,N_1677,N_1669);
nor U1933 (N_1933,N_1644,N_1758);
nor U1934 (N_1934,N_1649,N_1618);
nand U1935 (N_1935,N_1665,N_1613);
and U1936 (N_1936,N_1685,N_1795);
or U1937 (N_1937,N_1625,N_1649);
or U1938 (N_1938,N_1770,N_1651);
or U1939 (N_1939,N_1614,N_1607);
nor U1940 (N_1940,N_1695,N_1715);
and U1941 (N_1941,N_1738,N_1692);
and U1942 (N_1942,N_1768,N_1730);
nor U1943 (N_1943,N_1618,N_1796);
nand U1944 (N_1944,N_1776,N_1649);
nor U1945 (N_1945,N_1790,N_1748);
xnor U1946 (N_1946,N_1653,N_1618);
or U1947 (N_1947,N_1628,N_1790);
nor U1948 (N_1948,N_1660,N_1634);
and U1949 (N_1949,N_1637,N_1618);
nor U1950 (N_1950,N_1792,N_1681);
nand U1951 (N_1951,N_1668,N_1658);
xor U1952 (N_1952,N_1700,N_1616);
and U1953 (N_1953,N_1710,N_1654);
nor U1954 (N_1954,N_1753,N_1697);
or U1955 (N_1955,N_1793,N_1761);
nor U1956 (N_1956,N_1747,N_1785);
xor U1957 (N_1957,N_1689,N_1760);
and U1958 (N_1958,N_1617,N_1797);
xor U1959 (N_1959,N_1794,N_1741);
xor U1960 (N_1960,N_1720,N_1638);
nor U1961 (N_1961,N_1660,N_1732);
nand U1962 (N_1962,N_1623,N_1753);
or U1963 (N_1963,N_1661,N_1768);
nand U1964 (N_1964,N_1689,N_1766);
nand U1965 (N_1965,N_1700,N_1746);
nor U1966 (N_1966,N_1663,N_1626);
xnor U1967 (N_1967,N_1770,N_1782);
xor U1968 (N_1968,N_1791,N_1797);
xor U1969 (N_1969,N_1605,N_1647);
nand U1970 (N_1970,N_1669,N_1683);
nand U1971 (N_1971,N_1693,N_1710);
nand U1972 (N_1972,N_1651,N_1690);
nor U1973 (N_1973,N_1711,N_1668);
and U1974 (N_1974,N_1774,N_1712);
nor U1975 (N_1975,N_1768,N_1609);
and U1976 (N_1976,N_1657,N_1739);
nand U1977 (N_1977,N_1722,N_1703);
nor U1978 (N_1978,N_1607,N_1713);
nand U1979 (N_1979,N_1766,N_1618);
or U1980 (N_1980,N_1774,N_1626);
and U1981 (N_1981,N_1721,N_1675);
and U1982 (N_1982,N_1720,N_1747);
nand U1983 (N_1983,N_1690,N_1642);
nor U1984 (N_1984,N_1630,N_1739);
and U1985 (N_1985,N_1787,N_1694);
nor U1986 (N_1986,N_1693,N_1643);
nor U1987 (N_1987,N_1712,N_1785);
nand U1988 (N_1988,N_1757,N_1655);
nand U1989 (N_1989,N_1684,N_1621);
nor U1990 (N_1990,N_1721,N_1638);
or U1991 (N_1991,N_1748,N_1633);
nand U1992 (N_1992,N_1727,N_1628);
or U1993 (N_1993,N_1655,N_1763);
nor U1994 (N_1994,N_1757,N_1761);
nor U1995 (N_1995,N_1718,N_1602);
nand U1996 (N_1996,N_1634,N_1746);
nor U1997 (N_1997,N_1788,N_1620);
nor U1998 (N_1998,N_1677,N_1768);
and U1999 (N_1999,N_1652,N_1670);
nor U2000 (N_2000,N_1957,N_1913);
nand U2001 (N_2001,N_1988,N_1837);
nand U2002 (N_2002,N_1822,N_1918);
nand U2003 (N_2003,N_1896,N_1836);
nor U2004 (N_2004,N_1996,N_1926);
or U2005 (N_2005,N_1898,N_1857);
or U2006 (N_2006,N_1851,N_1911);
nor U2007 (N_2007,N_1844,N_1905);
or U2008 (N_2008,N_1801,N_1868);
xor U2009 (N_2009,N_1948,N_1906);
and U2010 (N_2010,N_1916,N_1874);
nor U2011 (N_2011,N_1934,N_1880);
xnor U2012 (N_2012,N_1807,N_1951);
nand U2013 (N_2013,N_1900,N_1902);
nand U2014 (N_2014,N_1929,N_1892);
xor U2015 (N_2015,N_1922,N_1802);
or U2016 (N_2016,N_1826,N_1921);
nand U2017 (N_2017,N_1998,N_1821);
and U2018 (N_2018,N_1897,N_1973);
and U2019 (N_2019,N_1971,N_1831);
nor U2020 (N_2020,N_1992,N_1842);
nor U2021 (N_2021,N_1838,N_1940);
and U2022 (N_2022,N_1977,N_1993);
xnor U2023 (N_2023,N_1869,N_1994);
nand U2024 (N_2024,N_1867,N_1811);
xor U2025 (N_2025,N_1887,N_1845);
nand U2026 (N_2026,N_1953,N_1979);
xor U2027 (N_2027,N_1866,N_1967);
nand U2028 (N_2028,N_1884,N_1894);
nor U2029 (N_2029,N_1817,N_1989);
or U2030 (N_2030,N_1871,N_1904);
nor U2031 (N_2031,N_1888,N_1968);
nand U2032 (N_2032,N_1827,N_1919);
nand U2033 (N_2033,N_1862,N_1819);
nor U2034 (N_2034,N_1877,N_1879);
or U2035 (N_2035,N_1864,N_1895);
xnor U2036 (N_2036,N_1834,N_1854);
and U2037 (N_2037,N_1901,N_1883);
xor U2038 (N_2038,N_1870,N_1936);
xnor U2039 (N_2039,N_1970,N_1985);
xor U2040 (N_2040,N_1991,N_1952);
xnor U2041 (N_2041,N_1853,N_1997);
nor U2042 (N_2042,N_1847,N_1825);
or U2043 (N_2043,N_1923,N_1806);
xnor U2044 (N_2044,N_1981,N_1984);
nor U2045 (N_2045,N_1975,N_1840);
nor U2046 (N_2046,N_1872,N_1959);
nor U2047 (N_2047,N_1875,N_1891);
nor U2048 (N_2048,N_1927,N_1805);
and U2049 (N_2049,N_1949,N_1890);
xor U2050 (N_2050,N_1976,N_1803);
xnor U2051 (N_2051,N_1958,N_1846);
nand U2052 (N_2052,N_1841,N_1933);
nor U2053 (N_2053,N_1815,N_1915);
nor U2054 (N_2054,N_1963,N_1947);
and U2055 (N_2055,N_1986,N_1859);
and U2056 (N_2056,N_1865,N_1983);
xor U2057 (N_2057,N_1928,N_1999);
nand U2058 (N_2058,N_1812,N_1804);
nand U2059 (N_2059,N_1850,N_1824);
nor U2060 (N_2060,N_1873,N_1830);
xnor U2061 (N_2061,N_1852,N_1954);
xnor U2062 (N_2062,N_1908,N_1848);
nand U2063 (N_2063,N_1964,N_1960);
nand U2064 (N_2064,N_1932,N_1858);
nor U2065 (N_2065,N_1849,N_1917);
nor U2066 (N_2066,N_1980,N_1843);
or U2067 (N_2067,N_1829,N_1925);
nand U2068 (N_2068,N_1818,N_1810);
nor U2069 (N_2069,N_1816,N_1878);
and U2070 (N_2070,N_1889,N_1939);
nor U2071 (N_2071,N_1863,N_1885);
nand U2072 (N_2072,N_1920,N_1876);
nor U2073 (N_2073,N_1974,N_1943);
or U2074 (N_2074,N_1814,N_1924);
nand U2075 (N_2075,N_1835,N_1950);
nor U2076 (N_2076,N_1942,N_1965);
xnor U2077 (N_2077,N_1944,N_1856);
or U2078 (N_2078,N_1938,N_1982);
or U2079 (N_2079,N_1935,N_1972);
and U2080 (N_2080,N_1808,N_1909);
and U2081 (N_2081,N_1886,N_1978);
xor U2082 (N_2082,N_1987,N_1966);
and U2083 (N_2083,N_1860,N_1893);
nor U2084 (N_2084,N_1910,N_1813);
nor U2085 (N_2085,N_1931,N_1820);
and U2086 (N_2086,N_1956,N_1961);
and U2087 (N_2087,N_1990,N_1882);
nor U2088 (N_2088,N_1937,N_1809);
nor U2089 (N_2089,N_1823,N_1941);
xnor U2090 (N_2090,N_1912,N_1946);
nand U2091 (N_2091,N_1907,N_1855);
and U2092 (N_2092,N_1969,N_1914);
nand U2093 (N_2093,N_1833,N_1832);
nor U2094 (N_2094,N_1800,N_1903);
and U2095 (N_2095,N_1945,N_1881);
and U2096 (N_2096,N_1962,N_1861);
xnor U2097 (N_2097,N_1995,N_1955);
xor U2098 (N_2098,N_1899,N_1930);
nor U2099 (N_2099,N_1839,N_1828);
xor U2100 (N_2100,N_1937,N_1824);
and U2101 (N_2101,N_1900,N_1963);
and U2102 (N_2102,N_1935,N_1989);
nor U2103 (N_2103,N_1830,N_1901);
or U2104 (N_2104,N_1888,N_1854);
and U2105 (N_2105,N_1814,N_1839);
or U2106 (N_2106,N_1855,N_1953);
and U2107 (N_2107,N_1924,N_1870);
nand U2108 (N_2108,N_1908,N_1811);
and U2109 (N_2109,N_1836,N_1994);
nand U2110 (N_2110,N_1862,N_1847);
or U2111 (N_2111,N_1995,N_1863);
nor U2112 (N_2112,N_1953,N_1985);
or U2113 (N_2113,N_1953,N_1834);
xor U2114 (N_2114,N_1865,N_1910);
nor U2115 (N_2115,N_1821,N_1903);
xnor U2116 (N_2116,N_1810,N_1992);
xor U2117 (N_2117,N_1914,N_1815);
nand U2118 (N_2118,N_1864,N_1803);
nand U2119 (N_2119,N_1966,N_1837);
xor U2120 (N_2120,N_1863,N_1981);
nand U2121 (N_2121,N_1877,N_1909);
and U2122 (N_2122,N_1889,N_1971);
xor U2123 (N_2123,N_1880,N_1928);
xor U2124 (N_2124,N_1995,N_1972);
and U2125 (N_2125,N_1873,N_1970);
nand U2126 (N_2126,N_1962,N_1869);
xnor U2127 (N_2127,N_1907,N_1970);
and U2128 (N_2128,N_1959,N_1887);
or U2129 (N_2129,N_1809,N_1863);
nor U2130 (N_2130,N_1815,N_1879);
or U2131 (N_2131,N_1853,N_1801);
and U2132 (N_2132,N_1914,N_1873);
nor U2133 (N_2133,N_1808,N_1961);
or U2134 (N_2134,N_1882,N_1941);
or U2135 (N_2135,N_1917,N_1850);
or U2136 (N_2136,N_1895,N_1961);
xnor U2137 (N_2137,N_1966,N_1835);
xnor U2138 (N_2138,N_1935,N_1889);
nor U2139 (N_2139,N_1933,N_1927);
nand U2140 (N_2140,N_1928,N_1890);
and U2141 (N_2141,N_1921,N_1914);
or U2142 (N_2142,N_1976,N_1828);
xor U2143 (N_2143,N_1803,N_1905);
xor U2144 (N_2144,N_1964,N_1913);
nor U2145 (N_2145,N_1948,N_1868);
nor U2146 (N_2146,N_1813,N_1992);
nor U2147 (N_2147,N_1928,N_1915);
xor U2148 (N_2148,N_1940,N_1956);
xor U2149 (N_2149,N_1809,N_1831);
nor U2150 (N_2150,N_1942,N_1922);
nor U2151 (N_2151,N_1967,N_1949);
nand U2152 (N_2152,N_1966,N_1827);
xor U2153 (N_2153,N_1953,N_1883);
or U2154 (N_2154,N_1829,N_1942);
nand U2155 (N_2155,N_1881,N_1910);
nor U2156 (N_2156,N_1995,N_1945);
nand U2157 (N_2157,N_1830,N_1948);
and U2158 (N_2158,N_1944,N_1901);
xnor U2159 (N_2159,N_1937,N_1865);
or U2160 (N_2160,N_1943,N_1961);
or U2161 (N_2161,N_1999,N_1975);
xnor U2162 (N_2162,N_1828,N_1956);
nand U2163 (N_2163,N_1819,N_1934);
xnor U2164 (N_2164,N_1971,N_1870);
and U2165 (N_2165,N_1892,N_1868);
nand U2166 (N_2166,N_1965,N_1978);
and U2167 (N_2167,N_1897,N_1883);
xnor U2168 (N_2168,N_1884,N_1976);
xor U2169 (N_2169,N_1884,N_1968);
or U2170 (N_2170,N_1924,N_1893);
nor U2171 (N_2171,N_1966,N_1982);
nor U2172 (N_2172,N_1960,N_1916);
nand U2173 (N_2173,N_1865,N_1820);
xor U2174 (N_2174,N_1983,N_1977);
and U2175 (N_2175,N_1983,N_1922);
xor U2176 (N_2176,N_1964,N_1848);
xor U2177 (N_2177,N_1923,N_1952);
or U2178 (N_2178,N_1850,N_1859);
nand U2179 (N_2179,N_1866,N_1887);
nand U2180 (N_2180,N_1883,N_1874);
or U2181 (N_2181,N_1951,N_1997);
nor U2182 (N_2182,N_1995,N_1827);
and U2183 (N_2183,N_1956,N_1845);
nand U2184 (N_2184,N_1995,N_1850);
and U2185 (N_2185,N_1893,N_1871);
or U2186 (N_2186,N_1991,N_1921);
xnor U2187 (N_2187,N_1916,N_1885);
nand U2188 (N_2188,N_1820,N_1980);
and U2189 (N_2189,N_1818,N_1978);
or U2190 (N_2190,N_1976,N_1811);
or U2191 (N_2191,N_1932,N_1966);
nor U2192 (N_2192,N_1900,N_1897);
xor U2193 (N_2193,N_1980,N_1914);
xnor U2194 (N_2194,N_1898,N_1834);
nand U2195 (N_2195,N_1945,N_1912);
or U2196 (N_2196,N_1957,N_1953);
or U2197 (N_2197,N_1876,N_1910);
xor U2198 (N_2198,N_1828,N_1808);
or U2199 (N_2199,N_1804,N_1832);
or U2200 (N_2200,N_2182,N_2080);
nor U2201 (N_2201,N_2118,N_2047);
nor U2202 (N_2202,N_2142,N_2100);
or U2203 (N_2203,N_2054,N_2145);
nor U2204 (N_2204,N_2191,N_2039);
xnor U2205 (N_2205,N_2075,N_2074);
or U2206 (N_2206,N_2156,N_2149);
and U2207 (N_2207,N_2048,N_2136);
nor U2208 (N_2208,N_2003,N_2058);
xnor U2209 (N_2209,N_2177,N_2186);
or U2210 (N_2210,N_2032,N_2181);
and U2211 (N_2211,N_2082,N_2139);
or U2212 (N_2212,N_2188,N_2031);
nor U2213 (N_2213,N_2183,N_2028);
xnor U2214 (N_2214,N_2130,N_2009);
or U2215 (N_2215,N_2107,N_2085);
and U2216 (N_2216,N_2042,N_2113);
or U2217 (N_2217,N_2012,N_2144);
or U2218 (N_2218,N_2024,N_2014);
nand U2219 (N_2219,N_2176,N_2120);
xnor U2220 (N_2220,N_2026,N_2180);
or U2221 (N_2221,N_2133,N_2061);
nand U2222 (N_2222,N_2089,N_2159);
nand U2223 (N_2223,N_2036,N_2006);
nor U2224 (N_2224,N_2148,N_2086);
or U2225 (N_2225,N_2005,N_2193);
and U2226 (N_2226,N_2132,N_2051);
nor U2227 (N_2227,N_2166,N_2063);
nor U2228 (N_2228,N_2093,N_2157);
xnor U2229 (N_2229,N_2110,N_2020);
and U2230 (N_2230,N_2083,N_2178);
nand U2231 (N_2231,N_2094,N_2000);
or U2232 (N_2232,N_2035,N_2084);
and U2233 (N_2233,N_2044,N_2053);
or U2234 (N_2234,N_2049,N_2114);
and U2235 (N_2235,N_2143,N_2165);
nand U2236 (N_2236,N_2038,N_2129);
and U2237 (N_2237,N_2041,N_2189);
nor U2238 (N_2238,N_2155,N_2174);
xnor U2239 (N_2239,N_2160,N_2116);
or U2240 (N_2240,N_2196,N_2168);
and U2241 (N_2241,N_2101,N_2119);
nand U2242 (N_2242,N_2018,N_2001);
nor U2243 (N_2243,N_2122,N_2173);
and U2244 (N_2244,N_2175,N_2138);
nor U2245 (N_2245,N_2109,N_2172);
or U2246 (N_2246,N_2135,N_2015);
nand U2247 (N_2247,N_2152,N_2077);
and U2248 (N_2248,N_2072,N_2103);
nand U2249 (N_2249,N_2106,N_2112);
xor U2250 (N_2250,N_2104,N_2069);
nand U2251 (N_2251,N_2187,N_2029);
and U2252 (N_2252,N_2016,N_2185);
nor U2253 (N_2253,N_2198,N_2030);
xnor U2254 (N_2254,N_2078,N_2154);
and U2255 (N_2255,N_2004,N_2199);
xor U2256 (N_2256,N_2197,N_2141);
nand U2257 (N_2257,N_2095,N_2096);
and U2258 (N_2258,N_2102,N_2153);
or U2259 (N_2259,N_2040,N_2127);
nand U2260 (N_2260,N_2194,N_2037);
nand U2261 (N_2261,N_2071,N_2195);
or U2262 (N_2262,N_2010,N_2081);
xor U2263 (N_2263,N_2060,N_2124);
and U2264 (N_2264,N_2052,N_2023);
nand U2265 (N_2265,N_2164,N_2192);
and U2266 (N_2266,N_2027,N_2163);
xor U2267 (N_2267,N_2073,N_2050);
and U2268 (N_2268,N_2151,N_2097);
xor U2269 (N_2269,N_2034,N_2140);
and U2270 (N_2270,N_2123,N_2179);
and U2271 (N_2271,N_2059,N_2017);
xnor U2272 (N_2272,N_2098,N_2167);
or U2273 (N_2273,N_2105,N_2126);
and U2274 (N_2274,N_2033,N_2066);
nand U2275 (N_2275,N_2079,N_2013);
and U2276 (N_2276,N_2171,N_2190);
and U2277 (N_2277,N_2091,N_2087);
and U2278 (N_2278,N_2070,N_2169);
and U2279 (N_2279,N_2043,N_2056);
nand U2280 (N_2280,N_2068,N_2076);
or U2281 (N_2281,N_2161,N_2021);
nand U2282 (N_2282,N_2011,N_2062);
or U2283 (N_2283,N_2146,N_2025);
or U2284 (N_2284,N_2088,N_2099);
nor U2285 (N_2285,N_2158,N_2150);
or U2286 (N_2286,N_2045,N_2131);
and U2287 (N_2287,N_2065,N_2067);
xor U2288 (N_2288,N_2002,N_2147);
or U2289 (N_2289,N_2057,N_2090);
and U2290 (N_2290,N_2111,N_2162);
or U2291 (N_2291,N_2022,N_2046);
or U2292 (N_2292,N_2117,N_2121);
or U2293 (N_2293,N_2137,N_2064);
and U2294 (N_2294,N_2125,N_2108);
xnor U2295 (N_2295,N_2170,N_2092);
xnor U2296 (N_2296,N_2115,N_2019);
and U2297 (N_2297,N_2128,N_2008);
and U2298 (N_2298,N_2184,N_2055);
xnor U2299 (N_2299,N_2134,N_2007);
and U2300 (N_2300,N_2030,N_2114);
xor U2301 (N_2301,N_2104,N_2180);
and U2302 (N_2302,N_2097,N_2138);
or U2303 (N_2303,N_2098,N_2186);
nand U2304 (N_2304,N_2007,N_2151);
and U2305 (N_2305,N_2049,N_2102);
and U2306 (N_2306,N_2189,N_2024);
xor U2307 (N_2307,N_2121,N_2101);
or U2308 (N_2308,N_2054,N_2059);
xnor U2309 (N_2309,N_2179,N_2063);
or U2310 (N_2310,N_2172,N_2176);
xor U2311 (N_2311,N_2126,N_2179);
or U2312 (N_2312,N_2178,N_2097);
or U2313 (N_2313,N_2180,N_2107);
or U2314 (N_2314,N_2127,N_2101);
nand U2315 (N_2315,N_2138,N_2046);
or U2316 (N_2316,N_2084,N_2046);
nor U2317 (N_2317,N_2188,N_2100);
xor U2318 (N_2318,N_2166,N_2097);
and U2319 (N_2319,N_2091,N_2116);
and U2320 (N_2320,N_2118,N_2155);
and U2321 (N_2321,N_2098,N_2091);
nor U2322 (N_2322,N_2075,N_2186);
nor U2323 (N_2323,N_2070,N_2101);
nand U2324 (N_2324,N_2176,N_2056);
xnor U2325 (N_2325,N_2106,N_2147);
and U2326 (N_2326,N_2190,N_2033);
nor U2327 (N_2327,N_2007,N_2089);
nand U2328 (N_2328,N_2051,N_2015);
nor U2329 (N_2329,N_2074,N_2144);
nor U2330 (N_2330,N_2144,N_2043);
and U2331 (N_2331,N_2106,N_2145);
xnor U2332 (N_2332,N_2081,N_2181);
nor U2333 (N_2333,N_2127,N_2188);
or U2334 (N_2334,N_2197,N_2191);
nand U2335 (N_2335,N_2083,N_2127);
and U2336 (N_2336,N_2102,N_2026);
nand U2337 (N_2337,N_2180,N_2033);
or U2338 (N_2338,N_2028,N_2188);
nand U2339 (N_2339,N_2002,N_2084);
and U2340 (N_2340,N_2008,N_2077);
nor U2341 (N_2341,N_2155,N_2011);
xnor U2342 (N_2342,N_2001,N_2110);
nand U2343 (N_2343,N_2114,N_2084);
or U2344 (N_2344,N_2158,N_2131);
xnor U2345 (N_2345,N_2051,N_2178);
or U2346 (N_2346,N_2082,N_2054);
xor U2347 (N_2347,N_2056,N_2039);
nor U2348 (N_2348,N_2137,N_2027);
nand U2349 (N_2349,N_2124,N_2104);
or U2350 (N_2350,N_2047,N_2058);
or U2351 (N_2351,N_2113,N_2163);
xnor U2352 (N_2352,N_2098,N_2119);
nand U2353 (N_2353,N_2144,N_2009);
nand U2354 (N_2354,N_2050,N_2055);
and U2355 (N_2355,N_2068,N_2175);
or U2356 (N_2356,N_2009,N_2122);
or U2357 (N_2357,N_2146,N_2051);
nand U2358 (N_2358,N_2179,N_2094);
xor U2359 (N_2359,N_2059,N_2009);
or U2360 (N_2360,N_2179,N_2092);
nor U2361 (N_2361,N_2011,N_2158);
nand U2362 (N_2362,N_2181,N_2003);
xor U2363 (N_2363,N_2160,N_2189);
nand U2364 (N_2364,N_2123,N_2054);
nor U2365 (N_2365,N_2130,N_2174);
nand U2366 (N_2366,N_2138,N_2079);
xor U2367 (N_2367,N_2004,N_2114);
nand U2368 (N_2368,N_2034,N_2195);
or U2369 (N_2369,N_2030,N_2063);
xor U2370 (N_2370,N_2100,N_2034);
xor U2371 (N_2371,N_2035,N_2079);
or U2372 (N_2372,N_2083,N_2102);
xnor U2373 (N_2373,N_2051,N_2166);
or U2374 (N_2374,N_2172,N_2047);
and U2375 (N_2375,N_2154,N_2132);
nand U2376 (N_2376,N_2150,N_2112);
and U2377 (N_2377,N_2102,N_2136);
nor U2378 (N_2378,N_2100,N_2070);
xor U2379 (N_2379,N_2103,N_2178);
xnor U2380 (N_2380,N_2147,N_2009);
xnor U2381 (N_2381,N_2040,N_2181);
nand U2382 (N_2382,N_2087,N_2163);
or U2383 (N_2383,N_2035,N_2193);
nor U2384 (N_2384,N_2025,N_2090);
nand U2385 (N_2385,N_2171,N_2180);
or U2386 (N_2386,N_2109,N_2140);
xnor U2387 (N_2387,N_2078,N_2039);
and U2388 (N_2388,N_2013,N_2139);
nand U2389 (N_2389,N_2074,N_2096);
nand U2390 (N_2390,N_2175,N_2033);
or U2391 (N_2391,N_2110,N_2152);
or U2392 (N_2392,N_2122,N_2099);
nor U2393 (N_2393,N_2071,N_2022);
and U2394 (N_2394,N_2127,N_2107);
and U2395 (N_2395,N_2184,N_2000);
and U2396 (N_2396,N_2051,N_2113);
and U2397 (N_2397,N_2051,N_2165);
and U2398 (N_2398,N_2029,N_2099);
nor U2399 (N_2399,N_2179,N_2030);
nand U2400 (N_2400,N_2363,N_2320);
xnor U2401 (N_2401,N_2375,N_2233);
or U2402 (N_2402,N_2225,N_2369);
and U2403 (N_2403,N_2350,N_2308);
and U2404 (N_2404,N_2314,N_2278);
or U2405 (N_2405,N_2344,N_2274);
or U2406 (N_2406,N_2330,N_2231);
or U2407 (N_2407,N_2389,N_2374);
or U2408 (N_2408,N_2244,N_2255);
and U2409 (N_2409,N_2354,N_2391);
xor U2410 (N_2410,N_2318,N_2239);
xor U2411 (N_2411,N_2220,N_2340);
nand U2412 (N_2412,N_2297,N_2379);
or U2413 (N_2413,N_2356,N_2224);
and U2414 (N_2414,N_2305,N_2201);
nand U2415 (N_2415,N_2212,N_2282);
nand U2416 (N_2416,N_2321,N_2202);
nand U2417 (N_2417,N_2392,N_2217);
xnor U2418 (N_2418,N_2246,N_2262);
xor U2419 (N_2419,N_2264,N_2381);
nand U2420 (N_2420,N_2345,N_2315);
and U2421 (N_2421,N_2336,N_2347);
nand U2422 (N_2422,N_2250,N_2309);
nor U2423 (N_2423,N_2329,N_2307);
nor U2424 (N_2424,N_2215,N_2322);
or U2425 (N_2425,N_2259,N_2251);
xnor U2426 (N_2426,N_2298,N_2371);
xnor U2427 (N_2427,N_2341,N_2205);
and U2428 (N_2428,N_2261,N_2326);
and U2429 (N_2429,N_2333,N_2204);
nor U2430 (N_2430,N_2208,N_2284);
or U2431 (N_2431,N_2324,N_2325);
and U2432 (N_2432,N_2200,N_2388);
and U2433 (N_2433,N_2241,N_2351);
nand U2434 (N_2434,N_2252,N_2238);
nand U2435 (N_2435,N_2221,N_2273);
or U2436 (N_2436,N_2258,N_2260);
xnor U2437 (N_2437,N_2218,N_2370);
and U2438 (N_2438,N_2206,N_2397);
and U2439 (N_2439,N_2236,N_2245);
or U2440 (N_2440,N_2243,N_2288);
nand U2441 (N_2441,N_2293,N_2384);
xnor U2442 (N_2442,N_2294,N_2285);
nand U2443 (N_2443,N_2365,N_2272);
or U2444 (N_2444,N_2378,N_2346);
nor U2445 (N_2445,N_2292,N_2368);
or U2446 (N_2446,N_2210,N_2376);
nor U2447 (N_2447,N_2248,N_2317);
xnor U2448 (N_2448,N_2242,N_2234);
or U2449 (N_2449,N_2240,N_2228);
nand U2450 (N_2450,N_2316,N_2364);
nand U2451 (N_2451,N_2271,N_2373);
xor U2452 (N_2452,N_2339,N_2253);
and U2453 (N_2453,N_2319,N_2280);
nor U2454 (N_2454,N_2267,N_2349);
nand U2455 (N_2455,N_2394,N_2366);
or U2456 (N_2456,N_2396,N_2304);
nand U2457 (N_2457,N_2377,N_2289);
xor U2458 (N_2458,N_2380,N_2355);
and U2459 (N_2459,N_2306,N_2343);
nor U2460 (N_2460,N_2303,N_2279);
or U2461 (N_2461,N_2287,N_2361);
or U2462 (N_2462,N_2219,N_2227);
nand U2463 (N_2463,N_2290,N_2256);
nand U2464 (N_2464,N_2372,N_2277);
nor U2465 (N_2465,N_2313,N_2265);
nor U2466 (N_2466,N_2257,N_2276);
xor U2467 (N_2467,N_2353,N_2203);
xnor U2468 (N_2468,N_2295,N_2254);
nor U2469 (N_2469,N_2399,N_2332);
nand U2470 (N_2470,N_2263,N_2390);
and U2471 (N_2471,N_2395,N_2266);
nand U2472 (N_2472,N_2232,N_2362);
nor U2473 (N_2473,N_2357,N_2327);
nor U2474 (N_2474,N_2331,N_2235);
or U2475 (N_2475,N_2360,N_2383);
or U2476 (N_2476,N_2342,N_2398);
and U2477 (N_2477,N_2300,N_2301);
nor U2478 (N_2478,N_2310,N_2275);
nor U2479 (N_2479,N_2348,N_2367);
and U2480 (N_2480,N_2323,N_2249);
or U2481 (N_2481,N_2299,N_2358);
xnor U2482 (N_2482,N_2207,N_2296);
or U2483 (N_2483,N_2283,N_2214);
or U2484 (N_2484,N_2338,N_2222);
nand U2485 (N_2485,N_2335,N_2230);
nor U2486 (N_2486,N_2302,N_2382);
and U2487 (N_2487,N_2213,N_2393);
xnor U2488 (N_2488,N_2209,N_2216);
nor U2489 (N_2489,N_2268,N_2281);
and U2490 (N_2490,N_2352,N_2291);
and U2491 (N_2491,N_2223,N_2385);
or U2492 (N_2492,N_2387,N_2226);
or U2493 (N_2493,N_2312,N_2269);
nor U2494 (N_2494,N_2270,N_2337);
nor U2495 (N_2495,N_2237,N_2286);
xnor U2496 (N_2496,N_2311,N_2386);
and U2497 (N_2497,N_2247,N_2328);
and U2498 (N_2498,N_2211,N_2229);
nor U2499 (N_2499,N_2359,N_2334);
nor U2500 (N_2500,N_2214,N_2348);
xor U2501 (N_2501,N_2329,N_2247);
nor U2502 (N_2502,N_2207,N_2357);
nor U2503 (N_2503,N_2336,N_2397);
and U2504 (N_2504,N_2371,N_2279);
and U2505 (N_2505,N_2261,N_2216);
and U2506 (N_2506,N_2379,N_2342);
nand U2507 (N_2507,N_2292,N_2288);
nand U2508 (N_2508,N_2219,N_2272);
or U2509 (N_2509,N_2333,N_2313);
xor U2510 (N_2510,N_2394,N_2235);
nor U2511 (N_2511,N_2259,N_2303);
and U2512 (N_2512,N_2362,N_2261);
nand U2513 (N_2513,N_2383,N_2249);
and U2514 (N_2514,N_2236,N_2293);
and U2515 (N_2515,N_2225,N_2254);
or U2516 (N_2516,N_2244,N_2394);
nand U2517 (N_2517,N_2227,N_2366);
nand U2518 (N_2518,N_2318,N_2291);
nor U2519 (N_2519,N_2229,N_2346);
nand U2520 (N_2520,N_2273,N_2378);
xor U2521 (N_2521,N_2267,N_2317);
and U2522 (N_2522,N_2254,N_2330);
and U2523 (N_2523,N_2338,N_2349);
or U2524 (N_2524,N_2322,N_2332);
or U2525 (N_2525,N_2392,N_2352);
nor U2526 (N_2526,N_2373,N_2317);
and U2527 (N_2527,N_2244,N_2264);
xor U2528 (N_2528,N_2229,N_2381);
and U2529 (N_2529,N_2379,N_2374);
and U2530 (N_2530,N_2381,N_2311);
xor U2531 (N_2531,N_2395,N_2267);
nor U2532 (N_2532,N_2301,N_2252);
and U2533 (N_2533,N_2250,N_2272);
xnor U2534 (N_2534,N_2379,N_2271);
and U2535 (N_2535,N_2385,N_2326);
and U2536 (N_2536,N_2380,N_2366);
and U2537 (N_2537,N_2311,N_2245);
xor U2538 (N_2538,N_2208,N_2383);
and U2539 (N_2539,N_2202,N_2342);
nor U2540 (N_2540,N_2297,N_2205);
xor U2541 (N_2541,N_2398,N_2288);
and U2542 (N_2542,N_2271,N_2218);
or U2543 (N_2543,N_2317,N_2315);
or U2544 (N_2544,N_2320,N_2348);
xnor U2545 (N_2545,N_2313,N_2269);
nor U2546 (N_2546,N_2369,N_2232);
or U2547 (N_2547,N_2316,N_2254);
and U2548 (N_2548,N_2296,N_2286);
or U2549 (N_2549,N_2301,N_2312);
nor U2550 (N_2550,N_2346,N_2348);
or U2551 (N_2551,N_2258,N_2339);
nor U2552 (N_2552,N_2340,N_2352);
or U2553 (N_2553,N_2265,N_2301);
or U2554 (N_2554,N_2257,N_2356);
xnor U2555 (N_2555,N_2298,N_2340);
xnor U2556 (N_2556,N_2313,N_2277);
nand U2557 (N_2557,N_2393,N_2367);
nor U2558 (N_2558,N_2294,N_2257);
nand U2559 (N_2559,N_2374,N_2356);
and U2560 (N_2560,N_2372,N_2290);
and U2561 (N_2561,N_2363,N_2270);
nor U2562 (N_2562,N_2264,N_2303);
nand U2563 (N_2563,N_2279,N_2314);
nand U2564 (N_2564,N_2211,N_2210);
or U2565 (N_2565,N_2365,N_2216);
xor U2566 (N_2566,N_2282,N_2296);
nand U2567 (N_2567,N_2279,N_2220);
and U2568 (N_2568,N_2263,N_2392);
and U2569 (N_2569,N_2344,N_2265);
and U2570 (N_2570,N_2340,N_2282);
and U2571 (N_2571,N_2270,N_2318);
and U2572 (N_2572,N_2306,N_2353);
or U2573 (N_2573,N_2384,N_2339);
or U2574 (N_2574,N_2262,N_2238);
and U2575 (N_2575,N_2261,N_2375);
xnor U2576 (N_2576,N_2205,N_2335);
nand U2577 (N_2577,N_2388,N_2363);
and U2578 (N_2578,N_2320,N_2311);
xnor U2579 (N_2579,N_2311,N_2339);
and U2580 (N_2580,N_2214,N_2279);
nor U2581 (N_2581,N_2206,N_2314);
xor U2582 (N_2582,N_2304,N_2266);
or U2583 (N_2583,N_2203,N_2275);
and U2584 (N_2584,N_2305,N_2274);
and U2585 (N_2585,N_2306,N_2223);
nor U2586 (N_2586,N_2303,N_2217);
or U2587 (N_2587,N_2355,N_2391);
nand U2588 (N_2588,N_2393,N_2387);
nand U2589 (N_2589,N_2338,N_2303);
xnor U2590 (N_2590,N_2281,N_2272);
or U2591 (N_2591,N_2269,N_2242);
or U2592 (N_2592,N_2320,N_2248);
nand U2593 (N_2593,N_2372,N_2227);
nand U2594 (N_2594,N_2231,N_2337);
or U2595 (N_2595,N_2393,N_2304);
nand U2596 (N_2596,N_2337,N_2309);
and U2597 (N_2597,N_2213,N_2259);
nand U2598 (N_2598,N_2235,N_2304);
and U2599 (N_2599,N_2210,N_2312);
nor U2600 (N_2600,N_2470,N_2451);
and U2601 (N_2601,N_2507,N_2407);
xnor U2602 (N_2602,N_2596,N_2461);
and U2603 (N_2603,N_2439,N_2421);
nand U2604 (N_2604,N_2588,N_2503);
xnor U2605 (N_2605,N_2545,N_2559);
nor U2606 (N_2606,N_2478,N_2531);
nand U2607 (N_2607,N_2415,N_2414);
xor U2608 (N_2608,N_2513,N_2575);
nand U2609 (N_2609,N_2447,N_2413);
nand U2610 (N_2610,N_2568,N_2405);
or U2611 (N_2611,N_2573,N_2410);
nand U2612 (N_2612,N_2592,N_2479);
or U2613 (N_2613,N_2565,N_2549);
nand U2614 (N_2614,N_2408,N_2480);
or U2615 (N_2615,N_2482,N_2540);
or U2616 (N_2616,N_2420,N_2584);
and U2617 (N_2617,N_2489,N_2435);
nor U2618 (N_2618,N_2591,N_2467);
nor U2619 (N_2619,N_2550,N_2578);
nand U2620 (N_2620,N_2494,N_2430);
or U2621 (N_2621,N_2424,N_2416);
and U2622 (N_2622,N_2535,N_2576);
and U2623 (N_2623,N_2598,N_2562);
xor U2624 (N_2624,N_2590,N_2506);
xor U2625 (N_2625,N_2541,N_2446);
and U2626 (N_2626,N_2476,N_2577);
nor U2627 (N_2627,N_2533,N_2516);
nand U2628 (N_2628,N_2417,N_2496);
xnor U2629 (N_2629,N_2589,N_2501);
nand U2630 (N_2630,N_2574,N_2555);
and U2631 (N_2631,N_2436,N_2442);
nand U2632 (N_2632,N_2460,N_2581);
or U2633 (N_2633,N_2428,N_2566);
and U2634 (N_2634,N_2542,N_2412);
nand U2635 (N_2635,N_2561,N_2409);
and U2636 (N_2636,N_2492,N_2418);
or U2637 (N_2637,N_2486,N_2457);
or U2638 (N_2638,N_2406,N_2563);
or U2639 (N_2639,N_2403,N_2499);
and U2640 (N_2640,N_2534,N_2468);
and U2641 (N_2641,N_2572,N_2569);
xnor U2642 (N_2642,N_2471,N_2517);
nand U2643 (N_2643,N_2510,N_2431);
nand U2644 (N_2644,N_2469,N_2437);
nand U2645 (N_2645,N_2466,N_2521);
nand U2646 (N_2646,N_2434,N_2583);
or U2647 (N_2647,N_2595,N_2465);
and U2648 (N_2648,N_2487,N_2498);
xnor U2649 (N_2649,N_2536,N_2538);
or U2650 (N_2650,N_2473,N_2526);
nor U2651 (N_2651,N_2481,N_2548);
nand U2652 (N_2652,N_2475,N_2557);
nand U2653 (N_2653,N_2554,N_2462);
nand U2654 (N_2654,N_2522,N_2530);
or U2655 (N_2655,N_2452,N_2432);
xnor U2656 (N_2656,N_2593,N_2456);
or U2657 (N_2657,N_2525,N_2441);
and U2658 (N_2658,N_2580,N_2449);
nand U2659 (N_2659,N_2422,N_2458);
nor U2660 (N_2660,N_2532,N_2527);
nand U2661 (N_2661,N_2438,N_2445);
or U2662 (N_2662,N_2401,N_2474);
xor U2663 (N_2663,N_2539,N_2579);
and U2664 (N_2664,N_2485,N_2443);
or U2665 (N_2665,N_2484,N_2423);
nor U2666 (N_2666,N_2508,N_2491);
nor U2667 (N_2667,N_2433,N_2426);
and U2668 (N_2668,N_2518,N_2523);
nor U2669 (N_2669,N_2520,N_2552);
and U2670 (N_2670,N_2400,N_2515);
and U2671 (N_2671,N_2488,N_2490);
or U2672 (N_2672,N_2495,N_2505);
or U2673 (N_2673,N_2528,N_2463);
nand U2674 (N_2674,N_2504,N_2453);
and U2675 (N_2675,N_2543,N_2511);
nor U2676 (N_2676,N_2570,N_2448);
xor U2677 (N_2677,N_2444,N_2402);
nor U2678 (N_2678,N_2546,N_2477);
nand U2679 (N_2679,N_2537,N_2586);
nand U2680 (N_2680,N_2594,N_2571);
nand U2681 (N_2681,N_2459,N_2454);
nor U2682 (N_2682,N_2599,N_2547);
and U2683 (N_2683,N_2560,N_2553);
or U2684 (N_2684,N_2558,N_2425);
and U2685 (N_2685,N_2524,N_2497);
and U2686 (N_2686,N_2404,N_2450);
xor U2687 (N_2687,N_2411,N_2483);
xor U2688 (N_2688,N_2519,N_2514);
or U2689 (N_2689,N_2587,N_2493);
or U2690 (N_2690,N_2585,N_2500);
xor U2691 (N_2691,N_2502,N_2472);
nor U2692 (N_2692,N_2427,N_2512);
nand U2693 (N_2693,N_2556,N_2582);
or U2694 (N_2694,N_2567,N_2429);
nor U2695 (N_2695,N_2509,N_2464);
nand U2696 (N_2696,N_2564,N_2529);
and U2697 (N_2697,N_2551,N_2597);
nor U2698 (N_2698,N_2544,N_2455);
xor U2699 (N_2699,N_2440,N_2419);
and U2700 (N_2700,N_2551,N_2520);
xnor U2701 (N_2701,N_2436,N_2475);
nor U2702 (N_2702,N_2486,N_2518);
xor U2703 (N_2703,N_2463,N_2466);
nor U2704 (N_2704,N_2558,N_2490);
xor U2705 (N_2705,N_2580,N_2469);
or U2706 (N_2706,N_2425,N_2490);
nand U2707 (N_2707,N_2451,N_2529);
and U2708 (N_2708,N_2433,N_2465);
nand U2709 (N_2709,N_2599,N_2528);
xor U2710 (N_2710,N_2433,N_2417);
nor U2711 (N_2711,N_2567,N_2557);
nor U2712 (N_2712,N_2429,N_2472);
nand U2713 (N_2713,N_2431,N_2513);
nand U2714 (N_2714,N_2405,N_2424);
or U2715 (N_2715,N_2505,N_2534);
nand U2716 (N_2716,N_2492,N_2533);
nor U2717 (N_2717,N_2407,N_2404);
and U2718 (N_2718,N_2507,N_2535);
nor U2719 (N_2719,N_2453,N_2409);
xnor U2720 (N_2720,N_2540,N_2497);
xor U2721 (N_2721,N_2474,N_2468);
xnor U2722 (N_2722,N_2500,N_2597);
and U2723 (N_2723,N_2474,N_2574);
xnor U2724 (N_2724,N_2529,N_2504);
or U2725 (N_2725,N_2486,N_2426);
or U2726 (N_2726,N_2463,N_2594);
nor U2727 (N_2727,N_2508,N_2423);
xnor U2728 (N_2728,N_2563,N_2540);
or U2729 (N_2729,N_2525,N_2451);
and U2730 (N_2730,N_2402,N_2507);
and U2731 (N_2731,N_2409,N_2571);
nand U2732 (N_2732,N_2578,N_2495);
and U2733 (N_2733,N_2581,N_2535);
nor U2734 (N_2734,N_2548,N_2462);
or U2735 (N_2735,N_2588,N_2447);
or U2736 (N_2736,N_2454,N_2444);
or U2737 (N_2737,N_2586,N_2514);
and U2738 (N_2738,N_2437,N_2598);
nand U2739 (N_2739,N_2471,N_2414);
or U2740 (N_2740,N_2567,N_2556);
xnor U2741 (N_2741,N_2559,N_2577);
nand U2742 (N_2742,N_2442,N_2555);
xor U2743 (N_2743,N_2517,N_2467);
and U2744 (N_2744,N_2554,N_2477);
or U2745 (N_2745,N_2419,N_2476);
or U2746 (N_2746,N_2455,N_2459);
or U2747 (N_2747,N_2509,N_2489);
nand U2748 (N_2748,N_2519,N_2525);
nand U2749 (N_2749,N_2457,N_2459);
nor U2750 (N_2750,N_2484,N_2561);
and U2751 (N_2751,N_2578,N_2476);
or U2752 (N_2752,N_2477,N_2466);
xnor U2753 (N_2753,N_2419,N_2591);
nand U2754 (N_2754,N_2541,N_2426);
nor U2755 (N_2755,N_2558,N_2556);
nand U2756 (N_2756,N_2443,N_2406);
nand U2757 (N_2757,N_2589,N_2490);
xor U2758 (N_2758,N_2501,N_2424);
nand U2759 (N_2759,N_2425,N_2536);
nor U2760 (N_2760,N_2477,N_2562);
nand U2761 (N_2761,N_2522,N_2479);
or U2762 (N_2762,N_2526,N_2462);
nor U2763 (N_2763,N_2500,N_2584);
or U2764 (N_2764,N_2496,N_2499);
xor U2765 (N_2765,N_2500,N_2400);
nand U2766 (N_2766,N_2553,N_2566);
nor U2767 (N_2767,N_2546,N_2547);
xor U2768 (N_2768,N_2524,N_2442);
xor U2769 (N_2769,N_2504,N_2471);
or U2770 (N_2770,N_2504,N_2423);
nand U2771 (N_2771,N_2569,N_2456);
or U2772 (N_2772,N_2563,N_2482);
or U2773 (N_2773,N_2402,N_2411);
or U2774 (N_2774,N_2587,N_2548);
or U2775 (N_2775,N_2446,N_2484);
and U2776 (N_2776,N_2537,N_2569);
xor U2777 (N_2777,N_2511,N_2498);
xnor U2778 (N_2778,N_2581,N_2410);
nor U2779 (N_2779,N_2535,N_2532);
nand U2780 (N_2780,N_2424,N_2530);
nand U2781 (N_2781,N_2406,N_2525);
nor U2782 (N_2782,N_2451,N_2559);
xor U2783 (N_2783,N_2422,N_2530);
nand U2784 (N_2784,N_2404,N_2492);
xnor U2785 (N_2785,N_2567,N_2423);
xor U2786 (N_2786,N_2408,N_2582);
nand U2787 (N_2787,N_2561,N_2535);
or U2788 (N_2788,N_2580,N_2425);
or U2789 (N_2789,N_2595,N_2570);
or U2790 (N_2790,N_2487,N_2583);
nor U2791 (N_2791,N_2546,N_2536);
nand U2792 (N_2792,N_2419,N_2477);
nand U2793 (N_2793,N_2591,N_2547);
or U2794 (N_2794,N_2467,N_2404);
and U2795 (N_2795,N_2456,N_2509);
or U2796 (N_2796,N_2593,N_2488);
xnor U2797 (N_2797,N_2583,N_2548);
and U2798 (N_2798,N_2529,N_2456);
xnor U2799 (N_2799,N_2485,N_2594);
nand U2800 (N_2800,N_2757,N_2681);
or U2801 (N_2801,N_2671,N_2632);
nor U2802 (N_2802,N_2621,N_2688);
and U2803 (N_2803,N_2696,N_2690);
nor U2804 (N_2804,N_2680,N_2736);
and U2805 (N_2805,N_2722,N_2756);
nand U2806 (N_2806,N_2619,N_2734);
nor U2807 (N_2807,N_2789,N_2629);
nor U2808 (N_2808,N_2635,N_2617);
xnor U2809 (N_2809,N_2695,N_2731);
nor U2810 (N_2810,N_2684,N_2606);
and U2811 (N_2811,N_2618,N_2720);
nand U2812 (N_2812,N_2780,N_2763);
nand U2813 (N_2813,N_2770,N_2624);
and U2814 (N_2814,N_2602,N_2796);
nand U2815 (N_2815,N_2742,N_2768);
and U2816 (N_2816,N_2764,N_2612);
or U2817 (N_2817,N_2758,N_2639);
or U2818 (N_2818,N_2740,N_2773);
and U2819 (N_2819,N_2750,N_2663);
nor U2820 (N_2820,N_2775,N_2609);
nor U2821 (N_2821,N_2652,N_2751);
xnor U2822 (N_2822,N_2672,N_2753);
or U2823 (N_2823,N_2797,N_2600);
xor U2824 (N_2824,N_2719,N_2739);
xor U2825 (N_2825,N_2712,N_2691);
and U2826 (N_2826,N_2779,N_2748);
nand U2827 (N_2827,N_2657,N_2747);
xnor U2828 (N_2828,N_2707,N_2642);
or U2829 (N_2829,N_2646,N_2608);
nand U2830 (N_2830,N_2708,N_2648);
nor U2831 (N_2831,N_2737,N_2728);
and U2832 (N_2832,N_2792,N_2638);
and U2833 (N_2833,N_2794,N_2721);
and U2834 (N_2834,N_2603,N_2611);
and U2835 (N_2835,N_2741,N_2631);
or U2836 (N_2836,N_2760,N_2769);
and U2837 (N_2837,N_2662,N_2774);
nand U2838 (N_2838,N_2656,N_2613);
and U2839 (N_2839,N_2706,N_2653);
xor U2840 (N_2840,N_2647,N_2676);
or U2841 (N_2841,N_2749,N_2715);
nor U2842 (N_2842,N_2645,N_2733);
or U2843 (N_2843,N_2700,N_2738);
or U2844 (N_2844,N_2687,N_2704);
nor U2845 (N_2845,N_2667,N_2767);
and U2846 (N_2846,N_2746,N_2776);
nor U2847 (N_2847,N_2795,N_2660);
and U2848 (N_2848,N_2670,N_2701);
or U2849 (N_2849,N_2730,N_2655);
nand U2850 (N_2850,N_2729,N_2685);
and U2851 (N_2851,N_2714,N_2743);
nor U2852 (N_2852,N_2786,N_2709);
and U2853 (N_2853,N_2703,N_2636);
and U2854 (N_2854,N_2772,N_2759);
nand U2855 (N_2855,N_2744,N_2785);
xnor U2856 (N_2856,N_2614,N_2735);
nand U2857 (N_2857,N_2790,N_2761);
or U2858 (N_2858,N_2783,N_2683);
nor U2859 (N_2859,N_2713,N_2661);
xor U2860 (N_2860,N_2766,N_2745);
nand U2861 (N_2861,N_2651,N_2674);
nor U2862 (N_2862,N_2610,N_2615);
or U2863 (N_2863,N_2771,N_2787);
xor U2864 (N_2864,N_2673,N_2732);
nand U2865 (N_2865,N_2702,N_2798);
or U2866 (N_2866,N_2623,N_2716);
or U2867 (N_2867,N_2699,N_2625);
and U2868 (N_2868,N_2601,N_2778);
nand U2869 (N_2869,N_2765,N_2755);
xor U2870 (N_2870,N_2643,N_2634);
xor U2871 (N_2871,N_2799,N_2658);
or U2872 (N_2872,N_2644,N_2633);
xnor U2873 (N_2873,N_2607,N_2641);
xnor U2874 (N_2874,N_2689,N_2664);
and U2875 (N_2875,N_2637,N_2675);
nand U2876 (N_2876,N_2630,N_2781);
and U2877 (N_2877,N_2725,N_2668);
xnor U2878 (N_2878,N_2666,N_2604);
nand U2879 (N_2879,N_2727,N_2654);
nor U2880 (N_2880,N_2724,N_2710);
nor U2881 (N_2881,N_2622,N_2782);
nor U2882 (N_2882,N_2686,N_2605);
and U2883 (N_2883,N_2705,N_2788);
nand U2884 (N_2884,N_2777,N_2698);
or U2885 (N_2885,N_2649,N_2723);
nor U2886 (N_2886,N_2665,N_2678);
nor U2887 (N_2887,N_2694,N_2793);
or U2888 (N_2888,N_2752,N_2718);
nand U2889 (N_2889,N_2754,N_2711);
xnor U2890 (N_2890,N_2669,N_2626);
and U2891 (N_2891,N_2784,N_2697);
nor U2892 (N_2892,N_2693,N_2677);
or U2893 (N_2893,N_2717,N_2640);
or U2894 (N_2894,N_2682,N_2627);
nor U2895 (N_2895,N_2791,N_2692);
nand U2896 (N_2896,N_2762,N_2620);
and U2897 (N_2897,N_2679,N_2726);
and U2898 (N_2898,N_2659,N_2650);
or U2899 (N_2899,N_2628,N_2616);
and U2900 (N_2900,N_2744,N_2687);
nor U2901 (N_2901,N_2727,N_2680);
nand U2902 (N_2902,N_2699,N_2785);
and U2903 (N_2903,N_2712,N_2658);
nand U2904 (N_2904,N_2791,N_2777);
and U2905 (N_2905,N_2673,N_2744);
nor U2906 (N_2906,N_2738,N_2649);
nor U2907 (N_2907,N_2785,N_2735);
nor U2908 (N_2908,N_2740,N_2686);
xor U2909 (N_2909,N_2669,N_2790);
or U2910 (N_2910,N_2702,N_2780);
nand U2911 (N_2911,N_2623,N_2624);
xnor U2912 (N_2912,N_2648,N_2771);
nand U2913 (N_2913,N_2734,N_2771);
xnor U2914 (N_2914,N_2604,N_2611);
nor U2915 (N_2915,N_2740,N_2682);
and U2916 (N_2916,N_2774,N_2767);
xnor U2917 (N_2917,N_2717,N_2615);
or U2918 (N_2918,N_2614,N_2765);
nor U2919 (N_2919,N_2734,N_2673);
and U2920 (N_2920,N_2778,N_2773);
and U2921 (N_2921,N_2731,N_2751);
and U2922 (N_2922,N_2604,N_2709);
nand U2923 (N_2923,N_2659,N_2694);
or U2924 (N_2924,N_2724,N_2634);
and U2925 (N_2925,N_2736,N_2612);
and U2926 (N_2926,N_2655,N_2614);
nor U2927 (N_2927,N_2700,N_2623);
or U2928 (N_2928,N_2712,N_2772);
and U2929 (N_2929,N_2730,N_2666);
or U2930 (N_2930,N_2727,N_2789);
or U2931 (N_2931,N_2713,N_2745);
or U2932 (N_2932,N_2774,N_2742);
nor U2933 (N_2933,N_2686,N_2756);
nand U2934 (N_2934,N_2798,N_2602);
xor U2935 (N_2935,N_2626,N_2630);
xor U2936 (N_2936,N_2790,N_2741);
nor U2937 (N_2937,N_2795,N_2753);
and U2938 (N_2938,N_2685,N_2677);
xor U2939 (N_2939,N_2618,N_2705);
nand U2940 (N_2940,N_2745,N_2763);
nor U2941 (N_2941,N_2753,N_2681);
or U2942 (N_2942,N_2743,N_2672);
and U2943 (N_2943,N_2771,N_2694);
nand U2944 (N_2944,N_2618,N_2646);
nor U2945 (N_2945,N_2732,N_2644);
xnor U2946 (N_2946,N_2684,N_2679);
and U2947 (N_2947,N_2606,N_2643);
or U2948 (N_2948,N_2700,N_2691);
or U2949 (N_2949,N_2648,N_2717);
or U2950 (N_2950,N_2679,N_2756);
nand U2951 (N_2951,N_2741,N_2794);
xnor U2952 (N_2952,N_2777,N_2732);
nand U2953 (N_2953,N_2755,N_2641);
or U2954 (N_2954,N_2623,N_2693);
and U2955 (N_2955,N_2727,N_2705);
and U2956 (N_2956,N_2757,N_2693);
nand U2957 (N_2957,N_2673,N_2759);
xnor U2958 (N_2958,N_2631,N_2740);
nor U2959 (N_2959,N_2634,N_2731);
nand U2960 (N_2960,N_2718,N_2670);
and U2961 (N_2961,N_2733,N_2608);
xor U2962 (N_2962,N_2699,N_2696);
and U2963 (N_2963,N_2708,N_2730);
or U2964 (N_2964,N_2741,N_2766);
or U2965 (N_2965,N_2703,N_2791);
nand U2966 (N_2966,N_2716,N_2784);
and U2967 (N_2967,N_2658,N_2686);
xor U2968 (N_2968,N_2745,N_2668);
or U2969 (N_2969,N_2753,N_2609);
nor U2970 (N_2970,N_2677,N_2682);
nand U2971 (N_2971,N_2625,N_2785);
and U2972 (N_2972,N_2689,N_2757);
xnor U2973 (N_2973,N_2735,N_2739);
and U2974 (N_2974,N_2682,N_2600);
xnor U2975 (N_2975,N_2712,N_2755);
and U2976 (N_2976,N_2770,N_2632);
and U2977 (N_2977,N_2635,N_2778);
and U2978 (N_2978,N_2602,N_2647);
nand U2979 (N_2979,N_2754,N_2696);
and U2980 (N_2980,N_2712,N_2745);
nor U2981 (N_2981,N_2775,N_2625);
or U2982 (N_2982,N_2799,N_2767);
and U2983 (N_2983,N_2716,N_2612);
nor U2984 (N_2984,N_2667,N_2650);
and U2985 (N_2985,N_2747,N_2712);
nor U2986 (N_2986,N_2665,N_2613);
xor U2987 (N_2987,N_2785,N_2615);
or U2988 (N_2988,N_2645,N_2789);
nor U2989 (N_2989,N_2710,N_2741);
or U2990 (N_2990,N_2676,N_2788);
nand U2991 (N_2991,N_2794,N_2777);
or U2992 (N_2992,N_2671,N_2641);
and U2993 (N_2993,N_2766,N_2738);
xor U2994 (N_2994,N_2790,N_2630);
or U2995 (N_2995,N_2692,N_2721);
or U2996 (N_2996,N_2644,N_2694);
nor U2997 (N_2997,N_2675,N_2784);
and U2998 (N_2998,N_2707,N_2677);
nor U2999 (N_2999,N_2662,N_2710);
xor UO_0 (O_0,N_2825,N_2851);
xor UO_1 (O_1,N_2921,N_2878);
nand UO_2 (O_2,N_2885,N_2804);
xor UO_3 (O_3,N_2953,N_2920);
and UO_4 (O_4,N_2992,N_2984);
or UO_5 (O_5,N_2810,N_2861);
nor UO_6 (O_6,N_2905,N_2989);
nand UO_7 (O_7,N_2858,N_2894);
and UO_8 (O_8,N_2855,N_2958);
nand UO_9 (O_9,N_2819,N_2866);
nand UO_10 (O_10,N_2967,N_2979);
nand UO_11 (O_11,N_2927,N_2814);
or UO_12 (O_12,N_2933,N_2808);
or UO_13 (O_13,N_2838,N_2978);
and UO_14 (O_14,N_2892,N_2987);
xnor UO_15 (O_15,N_2834,N_2983);
xor UO_16 (O_16,N_2897,N_2818);
and UO_17 (O_17,N_2908,N_2898);
or UO_18 (O_18,N_2880,N_2988);
nor UO_19 (O_19,N_2928,N_2854);
and UO_20 (O_20,N_2845,N_2950);
nand UO_21 (O_21,N_2900,N_2852);
nor UO_22 (O_22,N_2969,N_2930);
nor UO_23 (O_23,N_2912,N_2977);
xor UO_24 (O_24,N_2824,N_2888);
xnor UO_25 (O_25,N_2879,N_2887);
or UO_26 (O_26,N_2823,N_2999);
nor UO_27 (O_27,N_2996,N_2981);
nor UO_28 (O_28,N_2847,N_2993);
and UO_29 (O_29,N_2980,N_2839);
and UO_30 (O_30,N_2807,N_2954);
nand UO_31 (O_31,N_2849,N_2947);
xor UO_32 (O_32,N_2955,N_2917);
nor UO_33 (O_33,N_2929,N_2995);
nor UO_34 (O_34,N_2835,N_2886);
and UO_35 (O_35,N_2938,N_2925);
nor UO_36 (O_36,N_2826,N_2811);
or UO_37 (O_37,N_2973,N_2964);
nand UO_38 (O_38,N_2812,N_2890);
xnor UO_39 (O_39,N_2840,N_2815);
or UO_40 (O_40,N_2831,N_2919);
nor UO_41 (O_41,N_2837,N_2971);
xnor UO_42 (O_42,N_2903,N_2957);
or UO_43 (O_43,N_2830,N_2809);
or UO_44 (O_44,N_2956,N_2800);
xnor UO_45 (O_45,N_2922,N_2939);
nand UO_46 (O_46,N_2934,N_2867);
nor UO_47 (O_47,N_2870,N_2871);
nand UO_48 (O_48,N_2961,N_2937);
and UO_49 (O_49,N_2959,N_2943);
and UO_50 (O_50,N_2990,N_2962);
xor UO_51 (O_51,N_2926,N_2899);
nand UO_52 (O_52,N_2881,N_2806);
and UO_53 (O_53,N_2915,N_2844);
xnor UO_54 (O_54,N_2802,N_2828);
or UO_55 (O_55,N_2803,N_2902);
nor UO_56 (O_56,N_2972,N_2949);
nor UO_57 (O_57,N_2931,N_2813);
nand UO_58 (O_58,N_2982,N_2856);
and UO_59 (O_59,N_2891,N_2850);
nand UO_60 (O_60,N_2960,N_2864);
xor UO_61 (O_61,N_2948,N_2986);
nand UO_62 (O_62,N_2843,N_2994);
or UO_63 (O_63,N_2918,N_2966);
nor UO_64 (O_64,N_2822,N_2841);
xnor UO_65 (O_65,N_2907,N_2863);
nand UO_66 (O_66,N_2889,N_2942);
nand UO_67 (O_67,N_2991,N_2935);
xor UO_68 (O_68,N_2936,N_2869);
xnor UO_69 (O_69,N_2883,N_2976);
xnor UO_70 (O_70,N_2944,N_2884);
nand UO_71 (O_71,N_2945,N_2997);
and UO_72 (O_72,N_2901,N_2868);
or UO_73 (O_73,N_2801,N_2848);
nor UO_74 (O_74,N_2853,N_2941);
nand UO_75 (O_75,N_2909,N_2985);
xor UO_76 (O_76,N_2827,N_2963);
nor UO_77 (O_77,N_2873,N_2893);
nand UO_78 (O_78,N_2875,N_2951);
nor UO_79 (O_79,N_2968,N_2874);
nand UO_80 (O_80,N_2859,N_2829);
xor UO_81 (O_81,N_2846,N_2895);
or UO_82 (O_82,N_2916,N_2975);
nor UO_83 (O_83,N_2816,N_2842);
xor UO_84 (O_84,N_2860,N_2946);
or UO_85 (O_85,N_2940,N_2877);
nor UO_86 (O_86,N_2833,N_2817);
nor UO_87 (O_87,N_2911,N_2836);
xnor UO_88 (O_88,N_2906,N_2872);
and UO_89 (O_89,N_2965,N_2970);
xor UO_90 (O_90,N_2924,N_2904);
or UO_91 (O_91,N_2910,N_2952);
nor UO_92 (O_92,N_2805,N_2862);
or UO_93 (O_93,N_2820,N_2865);
nor UO_94 (O_94,N_2998,N_2832);
nor UO_95 (O_95,N_2932,N_2857);
xor UO_96 (O_96,N_2974,N_2913);
nor UO_97 (O_97,N_2923,N_2876);
and UO_98 (O_98,N_2896,N_2914);
or UO_99 (O_99,N_2882,N_2821);
or UO_100 (O_100,N_2849,N_2843);
xor UO_101 (O_101,N_2890,N_2853);
xnor UO_102 (O_102,N_2941,N_2982);
nor UO_103 (O_103,N_2870,N_2851);
or UO_104 (O_104,N_2838,N_2982);
and UO_105 (O_105,N_2948,N_2873);
and UO_106 (O_106,N_2868,N_2922);
and UO_107 (O_107,N_2800,N_2869);
nand UO_108 (O_108,N_2898,N_2887);
xor UO_109 (O_109,N_2927,N_2819);
nand UO_110 (O_110,N_2908,N_2980);
xnor UO_111 (O_111,N_2806,N_2866);
nor UO_112 (O_112,N_2990,N_2816);
nor UO_113 (O_113,N_2964,N_2934);
and UO_114 (O_114,N_2994,N_2888);
nor UO_115 (O_115,N_2877,N_2858);
xnor UO_116 (O_116,N_2973,N_2831);
nand UO_117 (O_117,N_2984,N_2919);
or UO_118 (O_118,N_2969,N_2880);
or UO_119 (O_119,N_2954,N_2893);
and UO_120 (O_120,N_2806,N_2973);
or UO_121 (O_121,N_2849,N_2889);
nand UO_122 (O_122,N_2817,N_2860);
nor UO_123 (O_123,N_2808,N_2866);
nand UO_124 (O_124,N_2887,N_2871);
and UO_125 (O_125,N_2985,N_2894);
xor UO_126 (O_126,N_2880,N_2816);
nor UO_127 (O_127,N_2963,N_2891);
nand UO_128 (O_128,N_2878,N_2913);
and UO_129 (O_129,N_2938,N_2988);
nand UO_130 (O_130,N_2923,N_2884);
nor UO_131 (O_131,N_2809,N_2954);
or UO_132 (O_132,N_2960,N_2999);
xor UO_133 (O_133,N_2813,N_2934);
nor UO_134 (O_134,N_2822,N_2816);
nand UO_135 (O_135,N_2918,N_2823);
nor UO_136 (O_136,N_2962,N_2853);
nor UO_137 (O_137,N_2818,N_2899);
or UO_138 (O_138,N_2930,N_2885);
xnor UO_139 (O_139,N_2947,N_2926);
or UO_140 (O_140,N_2907,N_2964);
and UO_141 (O_141,N_2976,N_2932);
and UO_142 (O_142,N_2819,N_2834);
and UO_143 (O_143,N_2896,N_2968);
and UO_144 (O_144,N_2937,N_2967);
nor UO_145 (O_145,N_2915,N_2924);
and UO_146 (O_146,N_2910,N_2931);
or UO_147 (O_147,N_2992,N_2811);
and UO_148 (O_148,N_2964,N_2886);
xnor UO_149 (O_149,N_2885,N_2843);
nand UO_150 (O_150,N_2856,N_2901);
or UO_151 (O_151,N_2962,N_2991);
or UO_152 (O_152,N_2959,N_2962);
or UO_153 (O_153,N_2863,N_2834);
and UO_154 (O_154,N_2837,N_2948);
or UO_155 (O_155,N_2818,N_2831);
or UO_156 (O_156,N_2960,N_2975);
nor UO_157 (O_157,N_2961,N_2960);
xnor UO_158 (O_158,N_2857,N_2868);
or UO_159 (O_159,N_2833,N_2960);
or UO_160 (O_160,N_2843,N_2857);
and UO_161 (O_161,N_2923,N_2831);
nand UO_162 (O_162,N_2821,N_2992);
nor UO_163 (O_163,N_2809,N_2821);
or UO_164 (O_164,N_2954,N_2957);
xor UO_165 (O_165,N_2941,N_2932);
xnor UO_166 (O_166,N_2875,N_2923);
and UO_167 (O_167,N_2860,N_2883);
and UO_168 (O_168,N_2970,N_2979);
nand UO_169 (O_169,N_2967,N_2864);
nor UO_170 (O_170,N_2832,N_2892);
or UO_171 (O_171,N_2842,N_2985);
xnor UO_172 (O_172,N_2829,N_2879);
nor UO_173 (O_173,N_2833,N_2970);
nand UO_174 (O_174,N_2895,N_2861);
and UO_175 (O_175,N_2992,N_2993);
nand UO_176 (O_176,N_2833,N_2820);
or UO_177 (O_177,N_2925,N_2872);
nor UO_178 (O_178,N_2842,N_2829);
nor UO_179 (O_179,N_2973,N_2914);
and UO_180 (O_180,N_2834,N_2966);
nand UO_181 (O_181,N_2803,N_2924);
or UO_182 (O_182,N_2868,N_2939);
nand UO_183 (O_183,N_2838,N_2812);
nand UO_184 (O_184,N_2950,N_2825);
and UO_185 (O_185,N_2995,N_2956);
nand UO_186 (O_186,N_2992,N_2869);
nor UO_187 (O_187,N_2811,N_2988);
xnor UO_188 (O_188,N_2826,N_2901);
or UO_189 (O_189,N_2844,N_2801);
and UO_190 (O_190,N_2852,N_2899);
nor UO_191 (O_191,N_2852,N_2842);
and UO_192 (O_192,N_2859,N_2961);
nor UO_193 (O_193,N_2863,N_2989);
nor UO_194 (O_194,N_2856,N_2965);
nand UO_195 (O_195,N_2932,N_2995);
xor UO_196 (O_196,N_2837,N_2953);
or UO_197 (O_197,N_2956,N_2894);
nor UO_198 (O_198,N_2866,N_2985);
nand UO_199 (O_199,N_2826,N_2963);
nand UO_200 (O_200,N_2875,N_2933);
nand UO_201 (O_201,N_2898,N_2858);
nand UO_202 (O_202,N_2982,N_2918);
nand UO_203 (O_203,N_2957,N_2882);
xor UO_204 (O_204,N_2974,N_2946);
nand UO_205 (O_205,N_2934,N_2937);
or UO_206 (O_206,N_2965,N_2868);
nand UO_207 (O_207,N_2893,N_2840);
xor UO_208 (O_208,N_2807,N_2879);
or UO_209 (O_209,N_2923,N_2930);
or UO_210 (O_210,N_2901,N_2976);
nor UO_211 (O_211,N_2933,N_2810);
nand UO_212 (O_212,N_2973,N_2853);
nand UO_213 (O_213,N_2944,N_2894);
nor UO_214 (O_214,N_2828,N_2849);
and UO_215 (O_215,N_2846,N_2861);
or UO_216 (O_216,N_2902,N_2868);
nor UO_217 (O_217,N_2950,N_2907);
or UO_218 (O_218,N_2937,N_2884);
and UO_219 (O_219,N_2880,N_2933);
or UO_220 (O_220,N_2917,N_2879);
or UO_221 (O_221,N_2833,N_2992);
xor UO_222 (O_222,N_2875,N_2872);
and UO_223 (O_223,N_2977,N_2844);
xor UO_224 (O_224,N_2834,N_2876);
and UO_225 (O_225,N_2964,N_2855);
nand UO_226 (O_226,N_2858,N_2967);
xnor UO_227 (O_227,N_2969,N_2809);
nand UO_228 (O_228,N_2971,N_2804);
and UO_229 (O_229,N_2889,N_2918);
nor UO_230 (O_230,N_2838,N_2956);
and UO_231 (O_231,N_2979,N_2835);
xnor UO_232 (O_232,N_2832,N_2982);
nand UO_233 (O_233,N_2893,N_2980);
and UO_234 (O_234,N_2988,N_2911);
nand UO_235 (O_235,N_2814,N_2851);
xnor UO_236 (O_236,N_2914,N_2933);
or UO_237 (O_237,N_2935,N_2920);
and UO_238 (O_238,N_2969,N_2954);
or UO_239 (O_239,N_2879,N_2897);
and UO_240 (O_240,N_2976,N_2859);
nand UO_241 (O_241,N_2929,N_2947);
nand UO_242 (O_242,N_2839,N_2993);
nor UO_243 (O_243,N_2966,N_2911);
or UO_244 (O_244,N_2942,N_2825);
or UO_245 (O_245,N_2821,N_2945);
or UO_246 (O_246,N_2839,N_2889);
and UO_247 (O_247,N_2984,N_2985);
or UO_248 (O_248,N_2862,N_2855);
nand UO_249 (O_249,N_2991,N_2821);
nand UO_250 (O_250,N_2837,N_2984);
nand UO_251 (O_251,N_2948,N_2834);
or UO_252 (O_252,N_2809,N_2831);
nor UO_253 (O_253,N_2814,N_2967);
nor UO_254 (O_254,N_2916,N_2929);
xnor UO_255 (O_255,N_2987,N_2907);
xnor UO_256 (O_256,N_2840,N_2813);
xnor UO_257 (O_257,N_2941,N_2987);
xor UO_258 (O_258,N_2918,N_2957);
nand UO_259 (O_259,N_2969,N_2942);
or UO_260 (O_260,N_2827,N_2926);
nand UO_261 (O_261,N_2844,N_2962);
and UO_262 (O_262,N_2826,N_2966);
or UO_263 (O_263,N_2892,N_2818);
and UO_264 (O_264,N_2914,N_2820);
and UO_265 (O_265,N_2913,N_2955);
and UO_266 (O_266,N_2854,N_2841);
xnor UO_267 (O_267,N_2831,N_2943);
and UO_268 (O_268,N_2928,N_2931);
nor UO_269 (O_269,N_2857,N_2909);
xor UO_270 (O_270,N_2969,N_2876);
and UO_271 (O_271,N_2858,N_2862);
and UO_272 (O_272,N_2828,N_2811);
nand UO_273 (O_273,N_2928,N_2847);
and UO_274 (O_274,N_2808,N_2953);
nor UO_275 (O_275,N_2992,N_2972);
nand UO_276 (O_276,N_2860,N_2911);
nand UO_277 (O_277,N_2973,N_2946);
and UO_278 (O_278,N_2952,N_2977);
nand UO_279 (O_279,N_2952,N_2837);
xnor UO_280 (O_280,N_2931,N_2929);
nor UO_281 (O_281,N_2980,N_2810);
nor UO_282 (O_282,N_2944,N_2914);
and UO_283 (O_283,N_2972,N_2806);
and UO_284 (O_284,N_2994,N_2814);
nand UO_285 (O_285,N_2985,N_2992);
nand UO_286 (O_286,N_2864,N_2917);
or UO_287 (O_287,N_2903,N_2849);
nand UO_288 (O_288,N_2839,N_2973);
xnor UO_289 (O_289,N_2860,N_2801);
and UO_290 (O_290,N_2840,N_2819);
nor UO_291 (O_291,N_2816,N_2942);
nand UO_292 (O_292,N_2811,N_2860);
nor UO_293 (O_293,N_2942,N_2813);
and UO_294 (O_294,N_2970,N_2940);
xnor UO_295 (O_295,N_2911,N_2995);
and UO_296 (O_296,N_2913,N_2977);
and UO_297 (O_297,N_2851,N_2961);
xor UO_298 (O_298,N_2986,N_2979);
or UO_299 (O_299,N_2827,N_2901);
or UO_300 (O_300,N_2954,N_2914);
xor UO_301 (O_301,N_2806,N_2849);
xnor UO_302 (O_302,N_2810,N_2990);
xnor UO_303 (O_303,N_2841,N_2806);
nand UO_304 (O_304,N_2872,N_2968);
and UO_305 (O_305,N_2907,N_2917);
and UO_306 (O_306,N_2947,N_2903);
nor UO_307 (O_307,N_2965,N_2914);
and UO_308 (O_308,N_2884,N_2973);
nor UO_309 (O_309,N_2808,N_2878);
xor UO_310 (O_310,N_2975,N_2854);
and UO_311 (O_311,N_2818,N_2808);
and UO_312 (O_312,N_2992,N_2800);
or UO_313 (O_313,N_2882,N_2901);
or UO_314 (O_314,N_2835,N_2958);
xnor UO_315 (O_315,N_2817,N_2839);
nor UO_316 (O_316,N_2842,N_2954);
or UO_317 (O_317,N_2989,N_2957);
xnor UO_318 (O_318,N_2839,N_2807);
xor UO_319 (O_319,N_2929,N_2982);
nand UO_320 (O_320,N_2979,N_2841);
nand UO_321 (O_321,N_2984,N_2910);
nand UO_322 (O_322,N_2847,N_2889);
nand UO_323 (O_323,N_2891,N_2867);
and UO_324 (O_324,N_2844,N_2997);
nand UO_325 (O_325,N_2996,N_2891);
or UO_326 (O_326,N_2825,N_2992);
and UO_327 (O_327,N_2938,N_2992);
xnor UO_328 (O_328,N_2936,N_2939);
or UO_329 (O_329,N_2878,N_2938);
xnor UO_330 (O_330,N_2964,N_2819);
xor UO_331 (O_331,N_2800,N_2947);
nor UO_332 (O_332,N_2879,N_2811);
or UO_333 (O_333,N_2912,N_2860);
and UO_334 (O_334,N_2889,N_2955);
nor UO_335 (O_335,N_2828,N_2814);
or UO_336 (O_336,N_2866,N_2829);
xor UO_337 (O_337,N_2969,N_2956);
and UO_338 (O_338,N_2905,N_2863);
xnor UO_339 (O_339,N_2976,N_2996);
nor UO_340 (O_340,N_2843,N_2841);
or UO_341 (O_341,N_2968,N_2928);
or UO_342 (O_342,N_2823,N_2871);
or UO_343 (O_343,N_2960,N_2900);
nand UO_344 (O_344,N_2871,N_2845);
nor UO_345 (O_345,N_2883,N_2931);
xnor UO_346 (O_346,N_2867,N_2948);
nor UO_347 (O_347,N_2849,N_2863);
and UO_348 (O_348,N_2818,N_2804);
or UO_349 (O_349,N_2879,N_2849);
xnor UO_350 (O_350,N_2894,N_2990);
and UO_351 (O_351,N_2861,N_2881);
and UO_352 (O_352,N_2839,N_2835);
or UO_353 (O_353,N_2865,N_2830);
nand UO_354 (O_354,N_2963,N_2925);
or UO_355 (O_355,N_2978,N_2845);
nor UO_356 (O_356,N_2917,N_2856);
nor UO_357 (O_357,N_2808,N_2951);
nand UO_358 (O_358,N_2829,N_2823);
nor UO_359 (O_359,N_2965,N_2964);
and UO_360 (O_360,N_2996,N_2861);
nor UO_361 (O_361,N_2858,N_2951);
nor UO_362 (O_362,N_2823,N_2882);
nor UO_363 (O_363,N_2827,N_2842);
and UO_364 (O_364,N_2979,N_2897);
nor UO_365 (O_365,N_2827,N_2840);
xor UO_366 (O_366,N_2843,N_2984);
nand UO_367 (O_367,N_2983,N_2989);
and UO_368 (O_368,N_2975,N_2936);
and UO_369 (O_369,N_2819,N_2828);
nor UO_370 (O_370,N_2860,N_2835);
and UO_371 (O_371,N_2895,N_2823);
and UO_372 (O_372,N_2823,N_2988);
nor UO_373 (O_373,N_2994,N_2981);
xor UO_374 (O_374,N_2971,N_2894);
nand UO_375 (O_375,N_2840,N_2973);
nor UO_376 (O_376,N_2903,N_2864);
nand UO_377 (O_377,N_2877,N_2936);
nand UO_378 (O_378,N_2894,N_2981);
or UO_379 (O_379,N_2859,N_2875);
nor UO_380 (O_380,N_2842,N_2917);
xnor UO_381 (O_381,N_2845,N_2861);
xnor UO_382 (O_382,N_2903,N_2939);
nor UO_383 (O_383,N_2922,N_2869);
nor UO_384 (O_384,N_2869,N_2948);
xor UO_385 (O_385,N_2819,N_2886);
nor UO_386 (O_386,N_2836,N_2976);
nor UO_387 (O_387,N_2905,N_2960);
nand UO_388 (O_388,N_2964,N_2861);
or UO_389 (O_389,N_2932,N_2895);
nor UO_390 (O_390,N_2878,N_2940);
nor UO_391 (O_391,N_2934,N_2870);
xnor UO_392 (O_392,N_2966,N_2849);
nor UO_393 (O_393,N_2840,N_2990);
xor UO_394 (O_394,N_2857,N_2871);
or UO_395 (O_395,N_2886,N_2979);
and UO_396 (O_396,N_2849,N_2943);
nand UO_397 (O_397,N_2973,N_2860);
or UO_398 (O_398,N_2858,N_2834);
xor UO_399 (O_399,N_2936,N_2871);
nand UO_400 (O_400,N_2955,N_2981);
or UO_401 (O_401,N_2822,N_2981);
nand UO_402 (O_402,N_2851,N_2897);
or UO_403 (O_403,N_2887,N_2953);
and UO_404 (O_404,N_2829,N_2996);
and UO_405 (O_405,N_2899,N_2820);
nor UO_406 (O_406,N_2875,N_2844);
xor UO_407 (O_407,N_2809,N_2909);
and UO_408 (O_408,N_2885,N_2919);
and UO_409 (O_409,N_2948,N_2811);
or UO_410 (O_410,N_2964,N_2900);
or UO_411 (O_411,N_2957,N_2922);
or UO_412 (O_412,N_2876,N_2808);
nand UO_413 (O_413,N_2845,N_2942);
or UO_414 (O_414,N_2907,N_2826);
or UO_415 (O_415,N_2864,N_2878);
nand UO_416 (O_416,N_2837,N_2934);
or UO_417 (O_417,N_2808,N_2861);
or UO_418 (O_418,N_2901,N_2832);
nor UO_419 (O_419,N_2829,N_2991);
nor UO_420 (O_420,N_2925,N_2882);
nand UO_421 (O_421,N_2918,N_2869);
nor UO_422 (O_422,N_2872,N_2949);
nor UO_423 (O_423,N_2959,N_2945);
nor UO_424 (O_424,N_2810,N_2973);
xor UO_425 (O_425,N_2821,N_2895);
or UO_426 (O_426,N_2960,N_2964);
xnor UO_427 (O_427,N_2985,N_2818);
or UO_428 (O_428,N_2848,N_2962);
xor UO_429 (O_429,N_2822,N_2927);
and UO_430 (O_430,N_2916,N_2876);
and UO_431 (O_431,N_2842,N_2825);
xnor UO_432 (O_432,N_2851,N_2869);
and UO_433 (O_433,N_2851,N_2936);
and UO_434 (O_434,N_2876,N_2981);
xnor UO_435 (O_435,N_2974,N_2816);
and UO_436 (O_436,N_2827,N_2934);
nand UO_437 (O_437,N_2957,N_2907);
and UO_438 (O_438,N_2891,N_2815);
nor UO_439 (O_439,N_2876,N_2831);
nor UO_440 (O_440,N_2936,N_2914);
or UO_441 (O_441,N_2991,N_2948);
and UO_442 (O_442,N_2900,N_2908);
xor UO_443 (O_443,N_2894,N_2856);
xor UO_444 (O_444,N_2958,N_2952);
or UO_445 (O_445,N_2947,N_2931);
or UO_446 (O_446,N_2878,N_2891);
nor UO_447 (O_447,N_2967,N_2923);
nand UO_448 (O_448,N_2860,N_2830);
nand UO_449 (O_449,N_2969,N_2840);
nor UO_450 (O_450,N_2942,N_2904);
nand UO_451 (O_451,N_2954,N_2864);
nand UO_452 (O_452,N_2998,N_2966);
nor UO_453 (O_453,N_2971,N_2865);
nand UO_454 (O_454,N_2931,N_2839);
and UO_455 (O_455,N_2818,N_2916);
nand UO_456 (O_456,N_2809,N_2825);
nor UO_457 (O_457,N_2838,N_2874);
xor UO_458 (O_458,N_2970,N_2911);
nand UO_459 (O_459,N_2962,N_2887);
nor UO_460 (O_460,N_2958,N_2977);
nand UO_461 (O_461,N_2890,N_2964);
xnor UO_462 (O_462,N_2935,N_2802);
and UO_463 (O_463,N_2972,N_2836);
xnor UO_464 (O_464,N_2919,N_2815);
nand UO_465 (O_465,N_2998,N_2840);
and UO_466 (O_466,N_2834,N_2972);
xnor UO_467 (O_467,N_2865,N_2837);
nor UO_468 (O_468,N_2989,N_2932);
xnor UO_469 (O_469,N_2826,N_2931);
xor UO_470 (O_470,N_2822,N_2835);
nor UO_471 (O_471,N_2993,N_2982);
or UO_472 (O_472,N_2857,N_2812);
nor UO_473 (O_473,N_2832,N_2860);
xor UO_474 (O_474,N_2992,N_2810);
and UO_475 (O_475,N_2819,N_2813);
nand UO_476 (O_476,N_2973,N_2978);
xor UO_477 (O_477,N_2880,N_2999);
and UO_478 (O_478,N_2900,N_2808);
nor UO_479 (O_479,N_2864,N_2854);
or UO_480 (O_480,N_2930,N_2811);
or UO_481 (O_481,N_2834,N_2900);
xor UO_482 (O_482,N_2892,N_2808);
and UO_483 (O_483,N_2919,N_2929);
xnor UO_484 (O_484,N_2957,N_2935);
and UO_485 (O_485,N_2988,N_2869);
nor UO_486 (O_486,N_2998,N_2899);
and UO_487 (O_487,N_2972,N_2865);
or UO_488 (O_488,N_2811,N_2966);
and UO_489 (O_489,N_2958,N_2863);
nand UO_490 (O_490,N_2961,N_2953);
nor UO_491 (O_491,N_2844,N_2874);
nand UO_492 (O_492,N_2868,N_2960);
nand UO_493 (O_493,N_2994,N_2940);
nand UO_494 (O_494,N_2868,N_2813);
and UO_495 (O_495,N_2990,N_2890);
nand UO_496 (O_496,N_2893,N_2836);
and UO_497 (O_497,N_2962,N_2918);
nor UO_498 (O_498,N_2887,N_2836);
nor UO_499 (O_499,N_2866,N_2939);
endmodule