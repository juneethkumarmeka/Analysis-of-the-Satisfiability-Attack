module basic_500_3000_500_4_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_78,In_208);
nor U1 (N_1,In_414,In_117);
and U2 (N_2,In_236,In_231);
and U3 (N_3,In_308,In_366);
and U4 (N_4,In_454,In_88);
or U5 (N_5,In_399,In_199);
nand U6 (N_6,In_242,In_22);
nor U7 (N_7,In_371,In_135);
nand U8 (N_8,In_447,In_28);
or U9 (N_9,In_138,In_426);
nand U10 (N_10,In_52,In_184);
nand U11 (N_11,In_380,In_268);
nor U12 (N_12,In_172,In_329);
nand U13 (N_13,In_266,In_243);
nand U14 (N_14,In_37,In_79);
nor U15 (N_15,In_216,In_108);
nand U16 (N_16,In_171,In_48);
xnor U17 (N_17,In_407,In_474);
and U18 (N_18,In_444,In_360);
nand U19 (N_19,In_433,In_265);
or U20 (N_20,In_470,In_343);
nor U21 (N_21,In_60,In_2);
or U22 (N_22,In_259,In_30);
or U23 (N_23,In_167,In_304);
or U24 (N_24,In_123,In_29);
nor U25 (N_25,In_333,In_347);
and U26 (N_26,In_73,In_84);
or U27 (N_27,In_315,In_13);
or U28 (N_28,In_132,In_173);
xnor U29 (N_29,In_211,In_6);
nand U30 (N_30,In_194,In_203);
xnor U31 (N_31,In_481,In_449);
or U32 (N_32,In_480,In_381);
nand U33 (N_33,In_128,In_295);
or U34 (N_34,In_363,In_321);
or U35 (N_35,In_392,In_465);
and U36 (N_36,In_400,In_302);
or U37 (N_37,In_74,In_107);
nor U38 (N_38,In_182,In_374);
nand U39 (N_39,In_262,In_458);
nand U40 (N_40,In_386,In_334);
nor U41 (N_41,In_376,In_101);
nand U42 (N_42,In_403,In_353);
nand U43 (N_43,In_402,In_387);
or U44 (N_44,In_174,In_16);
xor U45 (N_45,In_46,In_65);
or U46 (N_46,In_1,In_87);
nor U47 (N_47,In_18,In_396);
nor U48 (N_48,In_346,In_168);
nand U49 (N_49,In_111,In_326);
nand U50 (N_50,In_336,In_264);
and U51 (N_51,In_148,In_330);
and U52 (N_52,In_252,In_340);
nor U53 (N_53,In_254,In_328);
and U54 (N_54,In_141,In_115);
and U55 (N_55,In_8,In_357);
or U56 (N_56,In_42,In_450);
nor U57 (N_57,In_446,In_122);
nand U58 (N_58,In_9,In_318);
nor U59 (N_59,In_187,In_200);
and U60 (N_60,In_472,In_440);
nand U61 (N_61,In_384,In_225);
nand U62 (N_62,In_142,In_105);
nor U63 (N_63,In_218,In_70);
xor U64 (N_64,In_11,In_473);
nor U65 (N_65,In_395,In_139);
xnor U66 (N_66,In_124,In_322);
xnor U67 (N_67,In_398,In_202);
and U68 (N_68,In_244,In_405);
or U69 (N_69,In_298,In_147);
and U70 (N_70,In_417,In_99);
or U71 (N_71,In_114,In_325);
and U72 (N_72,In_209,In_475);
nor U73 (N_73,In_483,In_119);
nand U74 (N_74,In_319,In_485);
or U75 (N_75,In_198,In_61);
or U76 (N_76,In_255,In_62);
and U77 (N_77,In_14,In_4);
nor U78 (N_78,In_97,In_226);
nor U79 (N_79,In_300,In_44);
nand U80 (N_80,In_248,In_435);
nor U81 (N_81,In_453,In_206);
xnor U82 (N_82,In_489,In_156);
nand U83 (N_83,In_331,In_320);
nand U84 (N_84,In_288,In_462);
nand U85 (N_85,In_256,In_219);
or U86 (N_86,In_3,In_423);
nand U87 (N_87,In_327,In_19);
nand U88 (N_88,In_136,In_188);
or U89 (N_89,In_192,In_281);
nand U90 (N_90,In_36,In_146);
nand U91 (N_91,In_478,In_234);
nor U92 (N_92,In_116,In_134);
xor U93 (N_93,In_212,In_246);
nand U94 (N_94,In_272,In_348);
or U95 (N_95,In_409,In_176);
and U96 (N_96,In_373,In_283);
or U97 (N_97,In_185,In_238);
xor U98 (N_98,In_408,In_130);
xnor U99 (N_99,In_422,In_229);
or U100 (N_100,In_496,In_7);
nand U101 (N_101,In_245,In_190);
nand U102 (N_102,In_120,In_152);
xnor U103 (N_103,In_487,In_72);
or U104 (N_104,In_493,In_227);
xor U105 (N_105,In_210,In_32);
nor U106 (N_106,In_498,In_388);
xor U107 (N_107,In_488,In_314);
or U108 (N_108,In_436,In_367);
xnor U109 (N_109,In_249,In_232);
and U110 (N_110,In_239,In_193);
or U111 (N_111,In_466,In_75);
nand U112 (N_112,In_230,In_150);
nor U113 (N_113,In_307,In_279);
or U114 (N_114,In_362,In_67);
nand U115 (N_115,In_175,In_179);
xor U116 (N_116,In_448,In_165);
or U117 (N_117,In_10,In_497);
nor U118 (N_118,In_154,In_424);
or U119 (N_119,In_47,In_297);
xnor U120 (N_120,In_170,In_253);
xnor U121 (N_121,In_349,In_499);
nor U122 (N_122,In_34,In_484);
and U123 (N_123,In_278,In_76);
nand U124 (N_124,In_80,In_186);
or U125 (N_125,In_23,In_197);
and U126 (N_126,In_109,In_207);
or U127 (N_127,In_35,In_391);
nand U128 (N_128,In_385,In_15);
and U129 (N_129,In_393,In_121);
xor U130 (N_130,In_394,In_181);
xnor U131 (N_131,In_151,In_439);
or U132 (N_132,In_241,In_91);
and U133 (N_133,In_103,In_416);
or U134 (N_134,In_258,In_351);
xnor U135 (N_135,In_270,In_89);
xor U136 (N_136,In_93,In_276);
nor U137 (N_137,In_277,In_341);
nor U138 (N_138,In_289,In_419);
nor U139 (N_139,In_406,In_285);
xnor U140 (N_140,In_335,In_378);
nor U141 (N_141,In_204,In_57);
nor U142 (N_142,In_482,In_303);
nand U143 (N_143,In_126,In_25);
nand U144 (N_144,In_369,In_0);
and U145 (N_145,In_260,In_411);
xnor U146 (N_146,In_309,In_251);
nor U147 (N_147,In_45,In_443);
nand U148 (N_148,In_191,In_460);
or U149 (N_149,In_477,In_316);
or U150 (N_150,In_180,In_90);
and U151 (N_151,In_274,In_292);
nand U152 (N_152,In_293,In_494);
or U153 (N_153,In_112,In_31);
or U154 (N_154,In_461,In_77);
xor U155 (N_155,In_178,In_306);
nand U156 (N_156,In_442,In_476);
xnor U157 (N_157,In_43,In_40);
nor U158 (N_158,In_222,In_468);
xnor U159 (N_159,In_213,In_413);
nand U160 (N_160,In_305,In_269);
xor U161 (N_161,In_20,In_323);
nor U162 (N_162,In_158,In_492);
xor U163 (N_163,In_183,In_273);
nand U164 (N_164,In_317,In_166);
nor U165 (N_165,In_479,In_12);
or U166 (N_166,In_250,In_368);
and U167 (N_167,In_286,In_127);
or U168 (N_168,In_54,In_137);
nand U169 (N_169,In_104,In_92);
or U170 (N_170,In_415,In_235);
xor U171 (N_171,In_163,In_100);
and U172 (N_172,In_71,In_355);
and U173 (N_173,In_358,In_189);
and U174 (N_174,In_467,In_177);
nand U175 (N_175,In_196,In_275);
and U176 (N_176,In_421,In_294);
nand U177 (N_177,In_296,In_490);
xor U178 (N_178,In_162,In_427);
xor U179 (N_179,In_233,In_214);
xnor U180 (N_180,In_313,In_431);
nor U181 (N_181,In_459,In_401);
xor U182 (N_182,In_350,In_159);
nand U183 (N_183,In_464,In_83);
and U184 (N_184,In_469,In_471);
nor U185 (N_185,In_430,In_56);
and U186 (N_186,In_157,In_261);
nor U187 (N_187,In_94,In_133);
xnor U188 (N_188,In_66,In_257);
xnor U189 (N_189,In_145,In_339);
and U190 (N_190,In_342,In_98);
or U191 (N_191,In_379,In_50);
nor U192 (N_192,In_457,In_224);
and U193 (N_193,In_33,In_110);
or U194 (N_194,In_68,In_228);
nor U195 (N_195,In_425,In_53);
nand U196 (N_196,In_332,In_397);
nand U197 (N_197,In_280,In_438);
nand U198 (N_198,In_24,In_445);
xnor U199 (N_199,In_284,In_85);
or U200 (N_200,In_95,In_389);
and U201 (N_201,In_164,In_5);
xor U202 (N_202,In_361,In_82);
nand U203 (N_203,In_59,In_131);
nand U204 (N_204,In_161,In_51);
or U205 (N_205,In_352,In_21);
nor U206 (N_206,In_129,In_382);
nand U207 (N_207,In_486,In_372);
or U208 (N_208,In_437,In_432);
nand U209 (N_209,In_324,In_377);
or U210 (N_210,In_160,In_220);
or U211 (N_211,In_410,In_38);
and U212 (N_212,In_299,In_365);
and U213 (N_213,In_429,In_282);
nand U214 (N_214,In_420,In_215);
or U215 (N_215,In_149,In_310);
or U216 (N_216,In_412,In_271);
nand U217 (N_217,In_375,In_301);
or U218 (N_218,In_143,In_456);
nor U219 (N_219,In_370,In_337);
nand U220 (N_220,In_41,In_153);
or U221 (N_221,In_217,In_63);
and U222 (N_222,In_247,In_81);
or U223 (N_223,In_64,In_263);
or U224 (N_224,In_201,In_495);
or U225 (N_225,In_345,In_451);
or U226 (N_226,In_155,In_390);
xor U227 (N_227,In_195,In_39);
nand U228 (N_228,In_27,In_96);
and U229 (N_229,In_452,In_26);
nor U230 (N_230,In_338,In_354);
nor U231 (N_231,In_383,In_205);
nand U232 (N_232,In_58,In_434);
xnor U233 (N_233,In_364,In_237);
nor U234 (N_234,In_356,In_491);
nand U235 (N_235,In_311,In_441);
or U236 (N_236,In_118,In_240);
xor U237 (N_237,In_140,In_404);
xor U238 (N_238,In_291,In_17);
nor U239 (N_239,In_455,In_463);
nand U240 (N_240,In_267,In_287);
xor U241 (N_241,In_169,In_49);
nand U242 (N_242,In_125,In_55);
nor U243 (N_243,In_428,In_223);
or U244 (N_244,In_359,In_113);
and U245 (N_245,In_106,In_221);
xnor U246 (N_246,In_344,In_290);
nand U247 (N_247,In_102,In_144);
or U248 (N_248,In_418,In_312);
or U249 (N_249,In_69,In_86);
nand U250 (N_250,In_309,In_422);
and U251 (N_251,In_96,In_408);
xor U252 (N_252,In_277,In_27);
or U253 (N_253,In_277,In_25);
and U254 (N_254,In_293,In_278);
or U255 (N_255,In_380,In_342);
nand U256 (N_256,In_487,In_453);
xor U257 (N_257,In_9,In_161);
xnor U258 (N_258,In_26,In_149);
xnor U259 (N_259,In_191,In_208);
nand U260 (N_260,In_4,In_491);
xor U261 (N_261,In_435,In_2);
xnor U262 (N_262,In_30,In_334);
and U263 (N_263,In_65,In_430);
or U264 (N_264,In_419,In_331);
xor U265 (N_265,In_166,In_55);
xnor U266 (N_266,In_182,In_275);
nor U267 (N_267,In_10,In_481);
nor U268 (N_268,In_431,In_399);
and U269 (N_269,In_8,In_288);
xor U270 (N_270,In_132,In_8);
and U271 (N_271,In_477,In_253);
xnor U272 (N_272,In_389,In_73);
and U273 (N_273,In_76,In_274);
xor U274 (N_274,In_489,In_235);
nand U275 (N_275,In_199,In_362);
nand U276 (N_276,In_432,In_269);
nand U277 (N_277,In_377,In_221);
nand U278 (N_278,In_479,In_297);
nand U279 (N_279,In_291,In_479);
nor U280 (N_280,In_39,In_0);
or U281 (N_281,In_224,In_349);
xor U282 (N_282,In_180,In_93);
nor U283 (N_283,In_77,In_332);
or U284 (N_284,In_127,In_468);
and U285 (N_285,In_12,In_50);
or U286 (N_286,In_285,In_116);
xor U287 (N_287,In_487,In_450);
or U288 (N_288,In_274,In_32);
or U289 (N_289,In_396,In_175);
nor U290 (N_290,In_287,In_412);
nor U291 (N_291,In_22,In_406);
and U292 (N_292,In_164,In_206);
and U293 (N_293,In_209,In_5);
nor U294 (N_294,In_94,In_227);
xnor U295 (N_295,In_328,In_402);
and U296 (N_296,In_473,In_9);
xor U297 (N_297,In_326,In_208);
xnor U298 (N_298,In_189,In_237);
nand U299 (N_299,In_451,In_302);
or U300 (N_300,In_247,In_217);
nor U301 (N_301,In_321,In_449);
and U302 (N_302,In_273,In_100);
nand U303 (N_303,In_45,In_89);
xor U304 (N_304,In_161,In_55);
nand U305 (N_305,In_119,In_66);
and U306 (N_306,In_3,In_272);
nor U307 (N_307,In_72,In_365);
or U308 (N_308,In_472,In_239);
or U309 (N_309,In_449,In_282);
or U310 (N_310,In_225,In_377);
xor U311 (N_311,In_432,In_259);
or U312 (N_312,In_38,In_323);
nand U313 (N_313,In_378,In_483);
nand U314 (N_314,In_483,In_130);
nand U315 (N_315,In_185,In_313);
and U316 (N_316,In_373,In_54);
nor U317 (N_317,In_267,In_183);
nand U318 (N_318,In_28,In_319);
xor U319 (N_319,In_482,In_128);
nand U320 (N_320,In_463,In_493);
nand U321 (N_321,In_308,In_166);
nor U322 (N_322,In_42,In_294);
nor U323 (N_323,In_496,In_437);
nand U324 (N_324,In_376,In_279);
nand U325 (N_325,In_161,In_94);
and U326 (N_326,In_274,In_141);
xor U327 (N_327,In_193,In_59);
nand U328 (N_328,In_134,In_443);
nand U329 (N_329,In_207,In_203);
xor U330 (N_330,In_487,In_161);
or U331 (N_331,In_266,In_389);
xor U332 (N_332,In_388,In_87);
nor U333 (N_333,In_217,In_268);
xnor U334 (N_334,In_427,In_206);
nand U335 (N_335,In_86,In_374);
nand U336 (N_336,In_374,In_486);
nand U337 (N_337,In_460,In_42);
and U338 (N_338,In_1,In_408);
nand U339 (N_339,In_483,In_452);
xor U340 (N_340,In_248,In_270);
nand U341 (N_341,In_93,In_136);
nor U342 (N_342,In_369,In_167);
and U343 (N_343,In_39,In_132);
nand U344 (N_344,In_432,In_478);
xnor U345 (N_345,In_10,In_361);
and U346 (N_346,In_339,In_64);
or U347 (N_347,In_397,In_440);
nor U348 (N_348,In_351,In_138);
xor U349 (N_349,In_398,In_316);
nand U350 (N_350,In_43,In_23);
xnor U351 (N_351,In_393,In_221);
xnor U352 (N_352,In_13,In_398);
xnor U353 (N_353,In_449,In_370);
or U354 (N_354,In_24,In_319);
nand U355 (N_355,In_143,In_103);
nand U356 (N_356,In_243,In_41);
nor U357 (N_357,In_485,In_418);
or U358 (N_358,In_22,In_44);
and U359 (N_359,In_141,In_496);
nand U360 (N_360,In_359,In_443);
and U361 (N_361,In_468,In_25);
or U362 (N_362,In_300,In_149);
and U363 (N_363,In_441,In_65);
nor U364 (N_364,In_287,In_76);
and U365 (N_365,In_339,In_482);
nor U366 (N_366,In_37,In_373);
nand U367 (N_367,In_391,In_137);
nand U368 (N_368,In_206,In_358);
nor U369 (N_369,In_450,In_11);
and U370 (N_370,In_348,In_76);
nor U371 (N_371,In_368,In_271);
and U372 (N_372,In_415,In_123);
xor U373 (N_373,In_321,In_113);
or U374 (N_374,In_384,In_130);
xor U375 (N_375,In_240,In_78);
nand U376 (N_376,In_68,In_499);
or U377 (N_377,In_296,In_373);
or U378 (N_378,In_111,In_363);
and U379 (N_379,In_286,In_260);
nand U380 (N_380,In_240,In_197);
and U381 (N_381,In_199,In_167);
nand U382 (N_382,In_263,In_130);
xor U383 (N_383,In_227,In_29);
nand U384 (N_384,In_33,In_57);
or U385 (N_385,In_371,In_310);
nor U386 (N_386,In_226,In_345);
nand U387 (N_387,In_64,In_18);
or U388 (N_388,In_271,In_66);
nor U389 (N_389,In_231,In_295);
nand U390 (N_390,In_36,In_168);
nand U391 (N_391,In_55,In_315);
xnor U392 (N_392,In_116,In_135);
nor U393 (N_393,In_236,In_482);
or U394 (N_394,In_409,In_356);
nor U395 (N_395,In_443,In_468);
xor U396 (N_396,In_167,In_97);
and U397 (N_397,In_471,In_281);
or U398 (N_398,In_424,In_492);
or U399 (N_399,In_88,In_414);
or U400 (N_400,In_391,In_413);
or U401 (N_401,In_324,In_253);
xnor U402 (N_402,In_102,In_485);
or U403 (N_403,In_112,In_303);
xor U404 (N_404,In_470,In_120);
nand U405 (N_405,In_3,In_91);
xor U406 (N_406,In_118,In_23);
nor U407 (N_407,In_225,In_97);
or U408 (N_408,In_87,In_113);
nand U409 (N_409,In_46,In_350);
xor U410 (N_410,In_491,In_273);
and U411 (N_411,In_166,In_291);
or U412 (N_412,In_447,In_44);
and U413 (N_413,In_441,In_436);
nand U414 (N_414,In_495,In_465);
or U415 (N_415,In_345,In_190);
and U416 (N_416,In_213,In_184);
nor U417 (N_417,In_31,In_276);
nand U418 (N_418,In_383,In_117);
xnor U419 (N_419,In_34,In_278);
or U420 (N_420,In_494,In_213);
xnor U421 (N_421,In_314,In_274);
or U422 (N_422,In_283,In_493);
nand U423 (N_423,In_211,In_226);
and U424 (N_424,In_489,In_105);
nor U425 (N_425,In_178,In_14);
nor U426 (N_426,In_129,In_225);
nor U427 (N_427,In_238,In_466);
xor U428 (N_428,In_307,In_323);
nor U429 (N_429,In_225,In_93);
nor U430 (N_430,In_57,In_366);
nand U431 (N_431,In_30,In_213);
or U432 (N_432,In_67,In_315);
or U433 (N_433,In_26,In_461);
nor U434 (N_434,In_162,In_130);
or U435 (N_435,In_438,In_254);
nor U436 (N_436,In_358,In_46);
or U437 (N_437,In_404,In_92);
and U438 (N_438,In_434,In_30);
nor U439 (N_439,In_203,In_344);
or U440 (N_440,In_72,In_431);
or U441 (N_441,In_345,In_57);
nand U442 (N_442,In_351,In_423);
xor U443 (N_443,In_0,In_69);
or U444 (N_444,In_276,In_288);
xnor U445 (N_445,In_231,In_368);
nand U446 (N_446,In_279,In_138);
nor U447 (N_447,In_37,In_321);
or U448 (N_448,In_26,In_170);
or U449 (N_449,In_376,In_86);
nor U450 (N_450,In_44,In_223);
nor U451 (N_451,In_155,In_151);
xor U452 (N_452,In_1,In_437);
or U453 (N_453,In_81,In_77);
xor U454 (N_454,In_243,In_180);
or U455 (N_455,In_244,In_365);
nor U456 (N_456,In_110,In_11);
nor U457 (N_457,In_65,In_206);
and U458 (N_458,In_381,In_41);
nor U459 (N_459,In_161,In_380);
and U460 (N_460,In_141,In_197);
xor U461 (N_461,In_418,In_478);
or U462 (N_462,In_233,In_313);
and U463 (N_463,In_93,In_363);
nand U464 (N_464,In_416,In_9);
nand U465 (N_465,In_228,In_160);
or U466 (N_466,In_201,In_254);
xnor U467 (N_467,In_336,In_464);
and U468 (N_468,In_30,In_0);
xor U469 (N_469,In_69,In_379);
nor U470 (N_470,In_490,In_432);
and U471 (N_471,In_40,In_479);
nor U472 (N_472,In_231,In_351);
and U473 (N_473,In_462,In_23);
xor U474 (N_474,In_184,In_16);
xnor U475 (N_475,In_223,In_63);
nand U476 (N_476,In_141,In_25);
xnor U477 (N_477,In_235,In_112);
or U478 (N_478,In_132,In_363);
nand U479 (N_479,In_159,In_188);
nor U480 (N_480,In_213,In_317);
and U481 (N_481,In_154,In_499);
nand U482 (N_482,In_56,In_123);
xor U483 (N_483,In_275,In_227);
nand U484 (N_484,In_196,In_266);
or U485 (N_485,In_158,In_354);
xor U486 (N_486,In_389,In_361);
and U487 (N_487,In_117,In_191);
and U488 (N_488,In_439,In_240);
nor U489 (N_489,In_493,In_226);
xnor U490 (N_490,In_449,In_142);
nor U491 (N_491,In_65,In_389);
xor U492 (N_492,In_164,In_354);
nor U493 (N_493,In_102,In_478);
or U494 (N_494,In_478,In_392);
nand U495 (N_495,In_157,In_162);
nor U496 (N_496,In_158,In_476);
xor U497 (N_497,In_343,In_468);
and U498 (N_498,In_355,In_66);
nand U499 (N_499,In_485,In_215);
nor U500 (N_500,In_34,In_142);
and U501 (N_501,In_321,In_333);
or U502 (N_502,In_347,In_173);
and U503 (N_503,In_15,In_336);
nor U504 (N_504,In_163,In_139);
and U505 (N_505,In_43,In_312);
and U506 (N_506,In_123,In_389);
or U507 (N_507,In_25,In_339);
nor U508 (N_508,In_369,In_382);
and U509 (N_509,In_108,In_125);
and U510 (N_510,In_133,In_47);
and U511 (N_511,In_467,In_250);
xor U512 (N_512,In_302,In_171);
nand U513 (N_513,In_330,In_453);
or U514 (N_514,In_57,In_352);
or U515 (N_515,In_412,In_207);
nor U516 (N_516,In_303,In_435);
nand U517 (N_517,In_75,In_435);
xnor U518 (N_518,In_135,In_417);
xor U519 (N_519,In_336,In_102);
nand U520 (N_520,In_406,In_348);
nor U521 (N_521,In_189,In_216);
xnor U522 (N_522,In_247,In_21);
nand U523 (N_523,In_71,In_270);
xnor U524 (N_524,In_440,In_452);
and U525 (N_525,In_402,In_252);
xnor U526 (N_526,In_168,In_213);
xor U527 (N_527,In_46,In_237);
or U528 (N_528,In_371,In_46);
nor U529 (N_529,In_0,In_89);
xnor U530 (N_530,In_319,In_191);
and U531 (N_531,In_111,In_239);
xor U532 (N_532,In_292,In_27);
nor U533 (N_533,In_89,In_401);
nand U534 (N_534,In_324,In_66);
or U535 (N_535,In_258,In_127);
xnor U536 (N_536,In_334,In_105);
or U537 (N_537,In_161,In_258);
xor U538 (N_538,In_125,In_22);
or U539 (N_539,In_1,In_265);
or U540 (N_540,In_236,In_237);
nor U541 (N_541,In_138,In_404);
xor U542 (N_542,In_175,In_4);
nor U543 (N_543,In_342,In_268);
nor U544 (N_544,In_163,In_230);
or U545 (N_545,In_218,In_280);
xor U546 (N_546,In_334,In_165);
nand U547 (N_547,In_16,In_398);
nor U548 (N_548,In_301,In_292);
xnor U549 (N_549,In_180,In_496);
nand U550 (N_550,In_47,In_27);
or U551 (N_551,In_4,In_311);
xnor U552 (N_552,In_270,In_378);
or U553 (N_553,In_195,In_177);
nor U554 (N_554,In_88,In_485);
or U555 (N_555,In_79,In_126);
nor U556 (N_556,In_153,In_364);
nand U557 (N_557,In_473,In_331);
xor U558 (N_558,In_26,In_489);
or U559 (N_559,In_45,In_410);
and U560 (N_560,In_22,In_312);
nand U561 (N_561,In_444,In_157);
nand U562 (N_562,In_180,In_425);
nand U563 (N_563,In_0,In_331);
nor U564 (N_564,In_423,In_425);
and U565 (N_565,In_385,In_405);
nor U566 (N_566,In_403,In_138);
nor U567 (N_567,In_150,In_12);
or U568 (N_568,In_392,In_311);
and U569 (N_569,In_419,In_310);
and U570 (N_570,In_44,In_205);
xnor U571 (N_571,In_312,In_289);
nor U572 (N_572,In_70,In_319);
nor U573 (N_573,In_214,In_455);
nor U574 (N_574,In_297,In_293);
and U575 (N_575,In_110,In_0);
xor U576 (N_576,In_104,In_368);
nor U577 (N_577,In_108,In_66);
and U578 (N_578,In_379,In_22);
nor U579 (N_579,In_287,In_13);
nor U580 (N_580,In_397,In_367);
nand U581 (N_581,In_397,In_102);
nand U582 (N_582,In_315,In_136);
and U583 (N_583,In_97,In_151);
or U584 (N_584,In_496,In_194);
nand U585 (N_585,In_305,In_217);
xnor U586 (N_586,In_444,In_372);
nand U587 (N_587,In_311,In_239);
and U588 (N_588,In_294,In_270);
and U589 (N_589,In_121,In_190);
nor U590 (N_590,In_242,In_64);
and U591 (N_591,In_148,In_189);
xnor U592 (N_592,In_430,In_187);
or U593 (N_593,In_224,In_482);
nor U594 (N_594,In_210,In_439);
and U595 (N_595,In_242,In_54);
or U596 (N_596,In_149,In_232);
nand U597 (N_597,In_350,In_143);
nor U598 (N_598,In_273,In_71);
nor U599 (N_599,In_490,In_357);
nand U600 (N_600,In_420,In_493);
nor U601 (N_601,In_188,In_371);
nor U602 (N_602,In_330,In_479);
xnor U603 (N_603,In_68,In_149);
or U604 (N_604,In_234,In_260);
or U605 (N_605,In_452,In_216);
nand U606 (N_606,In_428,In_365);
or U607 (N_607,In_353,In_357);
xnor U608 (N_608,In_14,In_43);
or U609 (N_609,In_163,In_31);
nor U610 (N_610,In_153,In_76);
and U611 (N_611,In_160,In_73);
and U612 (N_612,In_498,In_402);
nand U613 (N_613,In_219,In_285);
nor U614 (N_614,In_200,In_397);
nand U615 (N_615,In_63,In_154);
nand U616 (N_616,In_419,In_293);
nor U617 (N_617,In_14,In_433);
nor U618 (N_618,In_437,In_393);
nand U619 (N_619,In_419,In_479);
and U620 (N_620,In_493,In_280);
nor U621 (N_621,In_59,In_453);
nand U622 (N_622,In_129,In_22);
nor U623 (N_623,In_450,In_434);
nor U624 (N_624,In_106,In_128);
and U625 (N_625,In_345,In_444);
xnor U626 (N_626,In_477,In_304);
and U627 (N_627,In_269,In_0);
nand U628 (N_628,In_486,In_60);
xor U629 (N_629,In_467,In_457);
nor U630 (N_630,In_132,In_251);
nand U631 (N_631,In_65,In_302);
nand U632 (N_632,In_405,In_72);
nor U633 (N_633,In_373,In_357);
or U634 (N_634,In_124,In_137);
and U635 (N_635,In_224,In_33);
nor U636 (N_636,In_309,In_495);
and U637 (N_637,In_309,In_275);
or U638 (N_638,In_200,In_311);
xnor U639 (N_639,In_247,In_452);
nand U640 (N_640,In_20,In_47);
xor U641 (N_641,In_467,In_180);
xor U642 (N_642,In_78,In_133);
nand U643 (N_643,In_191,In_206);
or U644 (N_644,In_495,In_244);
nand U645 (N_645,In_462,In_353);
and U646 (N_646,In_49,In_325);
xnor U647 (N_647,In_265,In_438);
nor U648 (N_648,In_50,In_174);
or U649 (N_649,In_395,In_142);
nor U650 (N_650,In_344,In_12);
nand U651 (N_651,In_85,In_410);
xor U652 (N_652,In_115,In_474);
or U653 (N_653,In_322,In_283);
or U654 (N_654,In_414,In_246);
nand U655 (N_655,In_392,In_448);
and U656 (N_656,In_191,In_184);
nand U657 (N_657,In_225,In_1);
and U658 (N_658,In_273,In_325);
and U659 (N_659,In_429,In_203);
xor U660 (N_660,In_331,In_338);
nand U661 (N_661,In_407,In_176);
nor U662 (N_662,In_277,In_352);
and U663 (N_663,In_49,In_435);
or U664 (N_664,In_119,In_355);
nor U665 (N_665,In_118,In_282);
xor U666 (N_666,In_363,In_169);
or U667 (N_667,In_101,In_220);
nand U668 (N_668,In_306,In_81);
nor U669 (N_669,In_452,In_124);
xor U670 (N_670,In_436,In_299);
xor U671 (N_671,In_454,In_451);
and U672 (N_672,In_133,In_375);
nand U673 (N_673,In_61,In_178);
nor U674 (N_674,In_358,In_362);
nand U675 (N_675,In_133,In_142);
xor U676 (N_676,In_317,In_203);
nor U677 (N_677,In_83,In_318);
and U678 (N_678,In_141,In_300);
and U679 (N_679,In_108,In_60);
nand U680 (N_680,In_471,In_171);
or U681 (N_681,In_84,In_417);
xnor U682 (N_682,In_343,In_281);
xnor U683 (N_683,In_84,In_460);
xor U684 (N_684,In_107,In_285);
nor U685 (N_685,In_411,In_113);
nand U686 (N_686,In_124,In_403);
and U687 (N_687,In_299,In_494);
nor U688 (N_688,In_338,In_116);
nand U689 (N_689,In_211,In_145);
nand U690 (N_690,In_399,In_434);
or U691 (N_691,In_142,In_452);
nor U692 (N_692,In_351,In_94);
nor U693 (N_693,In_402,In_323);
xor U694 (N_694,In_271,In_203);
nor U695 (N_695,In_191,In_17);
xor U696 (N_696,In_275,In_413);
nand U697 (N_697,In_294,In_106);
nand U698 (N_698,In_95,In_78);
nand U699 (N_699,In_419,In_376);
or U700 (N_700,In_412,In_9);
nand U701 (N_701,In_476,In_235);
nor U702 (N_702,In_368,In_321);
nor U703 (N_703,In_63,In_404);
and U704 (N_704,In_316,In_208);
or U705 (N_705,In_122,In_471);
nor U706 (N_706,In_480,In_227);
nand U707 (N_707,In_77,In_315);
nand U708 (N_708,In_304,In_373);
xor U709 (N_709,In_452,In_332);
or U710 (N_710,In_470,In_388);
nand U711 (N_711,In_348,In_282);
or U712 (N_712,In_449,In_49);
or U713 (N_713,In_355,In_360);
and U714 (N_714,In_420,In_408);
and U715 (N_715,In_187,In_434);
or U716 (N_716,In_416,In_168);
nand U717 (N_717,In_15,In_61);
nand U718 (N_718,In_368,In_46);
nand U719 (N_719,In_137,In_324);
xor U720 (N_720,In_404,In_136);
nor U721 (N_721,In_253,In_4);
and U722 (N_722,In_157,In_374);
nand U723 (N_723,In_221,In_305);
nor U724 (N_724,In_457,In_335);
xor U725 (N_725,In_361,In_115);
and U726 (N_726,In_102,In_455);
nand U727 (N_727,In_101,In_234);
or U728 (N_728,In_377,In_271);
and U729 (N_729,In_255,In_254);
nand U730 (N_730,In_313,In_103);
nand U731 (N_731,In_222,In_115);
nor U732 (N_732,In_481,In_480);
nand U733 (N_733,In_84,In_214);
nor U734 (N_734,In_242,In_23);
nor U735 (N_735,In_271,In_392);
nand U736 (N_736,In_367,In_231);
or U737 (N_737,In_46,In_112);
and U738 (N_738,In_277,In_85);
nor U739 (N_739,In_280,In_137);
nor U740 (N_740,In_89,In_321);
and U741 (N_741,In_172,In_114);
or U742 (N_742,In_417,In_393);
and U743 (N_743,In_446,In_336);
nand U744 (N_744,In_223,In_144);
nor U745 (N_745,In_275,In_3);
and U746 (N_746,In_355,In_396);
nor U747 (N_747,In_345,In_303);
xnor U748 (N_748,In_295,In_499);
and U749 (N_749,In_438,In_80);
xnor U750 (N_750,N_10,N_394);
or U751 (N_751,N_336,N_132);
or U752 (N_752,N_662,N_640);
xor U753 (N_753,N_602,N_643);
nor U754 (N_754,N_749,N_223);
and U755 (N_755,N_212,N_139);
nor U756 (N_756,N_387,N_495);
nand U757 (N_757,N_689,N_275);
and U758 (N_758,N_197,N_573);
nor U759 (N_759,N_681,N_24);
xnor U760 (N_760,N_235,N_352);
or U761 (N_761,N_242,N_55);
xnor U762 (N_762,N_106,N_99);
and U763 (N_763,N_327,N_489);
nor U764 (N_764,N_150,N_627);
xnor U765 (N_765,N_628,N_422);
or U766 (N_766,N_375,N_193);
and U767 (N_767,N_202,N_335);
nand U768 (N_768,N_700,N_737);
nor U769 (N_769,N_326,N_463);
or U770 (N_770,N_511,N_88);
and U771 (N_771,N_187,N_119);
and U772 (N_772,N_151,N_38);
nor U773 (N_773,N_87,N_78);
or U774 (N_774,N_588,N_559);
or U775 (N_775,N_736,N_62);
nand U776 (N_776,N_431,N_654);
nand U777 (N_777,N_490,N_22);
xor U778 (N_778,N_478,N_144);
nand U779 (N_779,N_597,N_137);
and U780 (N_780,N_60,N_469);
nor U781 (N_781,N_158,N_286);
and U782 (N_782,N_484,N_444);
nor U783 (N_783,N_111,N_102);
nand U784 (N_784,N_488,N_441);
nand U785 (N_785,N_25,N_466);
xnor U786 (N_786,N_405,N_86);
or U787 (N_787,N_708,N_694);
nor U788 (N_788,N_474,N_679);
and U789 (N_789,N_477,N_259);
xor U790 (N_790,N_255,N_531);
nand U791 (N_791,N_362,N_126);
nor U792 (N_792,N_575,N_346);
nor U793 (N_793,N_682,N_297);
xnor U794 (N_794,N_677,N_644);
nand U795 (N_795,N_639,N_157);
and U796 (N_796,N_353,N_181);
xnor U797 (N_797,N_131,N_35);
nand U798 (N_798,N_623,N_434);
nor U799 (N_799,N_527,N_211);
and U800 (N_800,N_101,N_250);
xor U801 (N_801,N_166,N_717);
and U802 (N_802,N_670,N_520);
nand U803 (N_803,N_134,N_214);
nor U804 (N_804,N_746,N_601);
or U805 (N_805,N_70,N_403);
nor U806 (N_806,N_625,N_200);
nand U807 (N_807,N_709,N_620);
or U808 (N_808,N_500,N_284);
or U809 (N_809,N_687,N_50);
nor U810 (N_810,N_153,N_7);
or U811 (N_811,N_8,N_536);
and U812 (N_812,N_622,N_430);
nor U813 (N_813,N_381,N_46);
nor U814 (N_814,N_376,N_438);
xnor U815 (N_815,N_747,N_369);
and U816 (N_816,N_159,N_428);
and U817 (N_817,N_548,N_5);
nand U818 (N_818,N_311,N_169);
or U819 (N_819,N_452,N_554);
xnor U820 (N_820,N_518,N_162);
or U821 (N_821,N_94,N_537);
and U822 (N_822,N_322,N_39);
nor U823 (N_823,N_269,N_615);
nor U824 (N_824,N_388,N_419);
nor U825 (N_825,N_341,N_613);
xnor U826 (N_826,N_26,N_517);
and U827 (N_827,N_324,N_423);
nor U828 (N_828,N_278,N_456);
nor U829 (N_829,N_174,N_237);
or U830 (N_830,N_658,N_95);
nor U831 (N_831,N_268,N_260);
or U832 (N_832,N_112,N_15);
or U833 (N_833,N_674,N_528);
xor U834 (N_834,N_450,N_233);
nand U835 (N_835,N_649,N_692);
and U836 (N_836,N_199,N_265);
and U837 (N_837,N_49,N_522);
nor U838 (N_838,N_105,N_343);
and U839 (N_839,N_263,N_164);
or U840 (N_840,N_98,N_12);
xor U841 (N_841,N_551,N_421);
nor U842 (N_842,N_535,N_704);
or U843 (N_843,N_392,N_114);
nand U844 (N_844,N_360,N_509);
nor U845 (N_845,N_671,N_180);
or U846 (N_846,N_184,N_266);
nand U847 (N_847,N_308,N_406);
or U848 (N_848,N_440,N_523);
xor U849 (N_849,N_110,N_72);
and U850 (N_850,N_225,N_271);
or U851 (N_851,N_247,N_465);
and U852 (N_852,N_67,N_203);
nor U853 (N_853,N_118,N_274);
or U854 (N_854,N_635,N_107);
xor U855 (N_855,N_296,N_366);
and U856 (N_856,N_619,N_479);
or U857 (N_857,N_222,N_560);
or U858 (N_858,N_226,N_426);
nor U859 (N_859,N_331,N_29);
nor U860 (N_860,N_312,N_541);
nor U861 (N_861,N_128,N_384);
xor U862 (N_862,N_443,N_345);
or U863 (N_863,N_748,N_614);
nor U864 (N_864,N_1,N_143);
nor U865 (N_865,N_349,N_84);
nand U866 (N_866,N_486,N_14);
or U867 (N_867,N_257,N_719);
nand U868 (N_868,N_267,N_437);
or U869 (N_869,N_244,N_665);
and U870 (N_870,N_585,N_612);
and U871 (N_871,N_580,N_40);
nor U872 (N_872,N_172,N_314);
or U873 (N_873,N_165,N_329);
or U874 (N_874,N_395,N_75);
nor U875 (N_875,N_241,N_688);
nand U876 (N_876,N_294,N_348);
and U877 (N_877,N_552,N_653);
or U878 (N_878,N_122,N_82);
xor U879 (N_879,N_476,N_501);
and U880 (N_880,N_496,N_538);
or U881 (N_881,N_213,N_705);
nand U882 (N_882,N_90,N_487);
nor U883 (N_883,N_81,N_215);
nand U884 (N_884,N_481,N_564);
nor U885 (N_885,N_634,N_393);
nor U886 (N_886,N_351,N_636);
xnor U887 (N_887,N_328,N_66);
and U888 (N_888,N_707,N_549);
nor U889 (N_889,N_617,N_177);
nor U890 (N_890,N_660,N_371);
or U891 (N_891,N_383,N_224);
or U892 (N_892,N_546,N_230);
nor U893 (N_893,N_347,N_148);
or U894 (N_894,N_273,N_338);
and U895 (N_895,N_20,N_333);
nand U896 (N_896,N_120,N_11);
xor U897 (N_897,N_485,N_295);
or U898 (N_898,N_725,N_0);
and U899 (N_899,N_567,N_36);
nor U900 (N_900,N_377,N_616);
or U901 (N_901,N_133,N_594);
and U902 (N_902,N_716,N_251);
nor U903 (N_903,N_695,N_140);
nor U904 (N_904,N_404,N_53);
nor U905 (N_905,N_599,N_115);
and U906 (N_906,N_711,N_100);
nor U907 (N_907,N_397,N_684);
or U908 (N_908,N_93,N_80);
xor U909 (N_909,N_73,N_589);
and U910 (N_910,N_23,N_651);
and U911 (N_911,N_261,N_483);
and U912 (N_912,N_370,N_3);
or U913 (N_913,N_491,N_79);
or U914 (N_914,N_661,N_621);
nand U915 (N_915,N_647,N_252);
or U916 (N_916,N_410,N_4);
or U917 (N_917,N_583,N_603);
or U918 (N_918,N_323,N_21);
nor U919 (N_919,N_141,N_109);
nor U920 (N_920,N_590,N_432);
nand U921 (N_921,N_570,N_386);
nand U922 (N_922,N_642,N_697);
nor U923 (N_923,N_188,N_71);
nor U924 (N_924,N_154,N_355);
or U925 (N_925,N_445,N_731);
xor U926 (N_926,N_412,N_638);
nand U927 (N_927,N_339,N_506);
xnor U928 (N_928,N_192,N_680);
and U929 (N_929,N_89,N_396);
and U930 (N_930,N_675,N_156);
or U931 (N_931,N_291,N_280);
and U932 (N_932,N_641,N_703);
or U933 (N_933,N_659,N_701);
xor U934 (N_934,N_206,N_16);
xor U935 (N_935,N_142,N_666);
or U936 (N_936,N_33,N_47);
xor U937 (N_937,N_686,N_702);
nand U938 (N_938,N_401,N_306);
and U939 (N_939,N_685,N_530);
or U940 (N_940,N_494,N_63);
nor U941 (N_941,N_553,N_354);
or U942 (N_942,N_626,N_318);
and U943 (N_943,N_399,N_744);
or U944 (N_944,N_372,N_582);
nor U945 (N_945,N_359,N_710);
and U946 (N_946,N_418,N_356);
nand U947 (N_947,N_28,N_210);
or U948 (N_948,N_713,N_698);
nor U949 (N_949,N_637,N_497);
and U950 (N_950,N_103,N_358);
and U951 (N_951,N_390,N_44);
or U952 (N_952,N_52,N_631);
nand U953 (N_953,N_69,N_43);
xnor U954 (N_954,N_454,N_59);
and U955 (N_955,N_729,N_6);
and U956 (N_956,N_379,N_198);
xnor U957 (N_957,N_715,N_357);
or U958 (N_958,N_467,N_340);
nor U959 (N_959,N_730,N_473);
nand U960 (N_960,N_555,N_216);
or U961 (N_961,N_720,N_108);
and U962 (N_962,N_342,N_436);
and U963 (N_963,N_524,N_556);
or U964 (N_964,N_85,N_526);
or U965 (N_965,N_185,N_457);
nor U966 (N_966,N_163,N_217);
and U967 (N_967,N_58,N_27);
nor U968 (N_968,N_17,N_232);
and U969 (N_969,N_293,N_482);
nand U970 (N_970,N_600,N_676);
nand U971 (N_971,N_533,N_305);
or U972 (N_972,N_236,N_303);
nor U973 (N_973,N_309,N_170);
and U974 (N_974,N_595,N_258);
nor U975 (N_975,N_249,N_461);
and U976 (N_976,N_195,N_718);
or U977 (N_977,N_632,N_34);
and U978 (N_978,N_565,N_168);
xor U979 (N_979,N_529,N_194);
nor U980 (N_980,N_167,N_310);
xor U981 (N_981,N_499,N_571);
and U982 (N_982,N_502,N_30);
and U983 (N_983,N_240,N_732);
or U984 (N_984,N_179,N_657);
xor U985 (N_985,N_544,N_596);
and U986 (N_986,N_664,N_146);
and U987 (N_987,N_219,N_65);
and U988 (N_988,N_130,N_283);
nor U989 (N_989,N_51,N_734);
and U990 (N_990,N_584,N_429);
nor U991 (N_991,N_451,N_407);
or U992 (N_992,N_319,N_385);
nand U993 (N_993,N_735,N_498);
nand U994 (N_994,N_175,N_545);
nor U995 (N_995,N_389,N_712);
xor U996 (N_996,N_667,N_147);
and U997 (N_997,N_514,N_97);
nand U998 (N_998,N_54,N_42);
and U999 (N_999,N_447,N_609);
nor U1000 (N_1000,N_2,N_453);
nand U1001 (N_1001,N_209,N_152);
xnor U1002 (N_1002,N_516,N_364);
nand U1003 (N_1003,N_227,N_299);
nand U1004 (N_1004,N_254,N_424);
nand U1005 (N_1005,N_380,N_563);
xor U1006 (N_1006,N_276,N_205);
and U1007 (N_1007,N_513,N_591);
and U1008 (N_1008,N_646,N_663);
nand U1009 (N_1009,N_733,N_231);
nand U1010 (N_1010,N_672,N_307);
xnor U1011 (N_1011,N_74,N_367);
xor U1012 (N_1012,N_547,N_178);
and U1013 (N_1013,N_18,N_234);
and U1014 (N_1014,N_160,N_690);
nand U1015 (N_1015,N_543,N_539);
nand U1016 (N_1016,N_460,N_577);
or U1017 (N_1017,N_41,N_427);
and U1018 (N_1018,N_204,N_525);
and U1019 (N_1019,N_442,N_745);
nand U1020 (N_1020,N_155,N_208);
xor U1021 (N_1021,N_723,N_532);
nor U1022 (N_1022,N_714,N_721);
or U1023 (N_1023,N_726,N_724);
xor U1024 (N_1024,N_183,N_699);
nor U1025 (N_1025,N_459,N_604);
xor U1026 (N_1026,N_201,N_587);
nand U1027 (N_1027,N_648,N_398);
nand U1028 (N_1028,N_425,N_610);
and U1029 (N_1029,N_470,N_13);
xnor U1030 (N_1030,N_400,N_361);
or U1031 (N_1031,N_321,N_61);
nor U1032 (N_1032,N_693,N_507);
nand U1033 (N_1033,N_416,N_334);
and U1034 (N_1034,N_607,N_569);
nor U1035 (N_1035,N_540,N_253);
xor U1036 (N_1036,N_92,N_542);
nor U1037 (N_1037,N_298,N_382);
and U1038 (N_1038,N_138,N_218);
and U1039 (N_1039,N_37,N_618);
nor U1040 (N_1040,N_277,N_455);
or U1041 (N_1041,N_678,N_673);
or U1042 (N_1042,N_316,N_557);
nand U1043 (N_1043,N_696,N_550);
nor U1044 (N_1044,N_449,N_468);
nor U1045 (N_1045,N_691,N_239);
or U1046 (N_1046,N_471,N_503);
nand U1047 (N_1047,N_365,N_189);
or U1048 (N_1048,N_207,N_534);
and U1049 (N_1049,N_127,N_743);
xnor U1050 (N_1050,N_413,N_301);
and U1051 (N_1051,N_581,N_578);
xnor U1052 (N_1052,N_45,N_281);
or U1053 (N_1053,N_124,N_629);
nand U1054 (N_1054,N_608,N_264);
nor U1055 (N_1055,N_519,N_568);
or U1056 (N_1056,N_579,N_56);
nand U1057 (N_1057,N_722,N_191);
or U1058 (N_1058,N_290,N_439);
and U1059 (N_1059,N_408,N_173);
nor U1060 (N_1060,N_475,N_562);
xor U1061 (N_1061,N_561,N_669);
nand U1062 (N_1062,N_123,N_121);
xor U1063 (N_1063,N_350,N_287);
xor U1064 (N_1064,N_593,N_113);
and U1065 (N_1065,N_317,N_136);
nor U1066 (N_1066,N_320,N_727);
or U1067 (N_1067,N_282,N_262);
nand U1068 (N_1068,N_330,N_464);
nor U1069 (N_1069,N_129,N_19);
xor U1070 (N_1070,N_728,N_145);
nor U1071 (N_1071,N_521,N_221);
xor U1072 (N_1072,N_472,N_652);
or U1073 (N_1073,N_337,N_741);
nor U1074 (N_1074,N_433,N_611);
and U1075 (N_1075,N_586,N_480);
xnor U1076 (N_1076,N_446,N_592);
xnor U1077 (N_1077,N_272,N_373);
nor U1078 (N_1078,N_76,N_64);
and U1079 (N_1079,N_116,N_31);
nor U1080 (N_1080,N_125,N_83);
nor U1081 (N_1081,N_368,N_409);
nand U1082 (N_1082,N_302,N_344);
nor U1083 (N_1083,N_558,N_515);
xor U1084 (N_1084,N_505,N_650);
and U1085 (N_1085,N_462,N_414);
or U1086 (N_1086,N_572,N_238);
nor U1087 (N_1087,N_96,N_633);
and U1088 (N_1088,N_279,N_668);
nor U1089 (N_1089,N_315,N_292);
or U1090 (N_1090,N_492,N_228);
or U1091 (N_1091,N_32,N_304);
nand U1092 (N_1092,N_566,N_220);
nor U1093 (N_1093,N_458,N_186);
xor U1094 (N_1094,N_493,N_598);
and U1095 (N_1095,N_448,N_182);
or U1096 (N_1096,N_417,N_740);
and U1097 (N_1097,N_288,N_508);
xnor U1098 (N_1098,N_229,N_739);
nor U1099 (N_1099,N_510,N_683);
nor U1100 (N_1100,N_742,N_504);
nand U1101 (N_1101,N_68,N_332);
or U1102 (N_1102,N_91,N_325);
nor U1103 (N_1103,N_246,N_270);
and U1104 (N_1104,N_378,N_104);
nor U1105 (N_1105,N_77,N_176);
xnor U1106 (N_1106,N_402,N_300);
xor U1107 (N_1107,N_243,N_435);
nand U1108 (N_1108,N_57,N_630);
xnor U1109 (N_1109,N_576,N_645);
and U1110 (N_1110,N_624,N_289);
nor U1111 (N_1111,N_196,N_656);
nor U1112 (N_1112,N_391,N_285);
or U1113 (N_1113,N_245,N_48);
or U1114 (N_1114,N_655,N_149);
xor U1115 (N_1115,N_411,N_374);
nor U1116 (N_1116,N_313,N_135);
xor U1117 (N_1117,N_256,N_363);
and U1118 (N_1118,N_9,N_415);
xnor U1119 (N_1119,N_738,N_512);
xor U1120 (N_1120,N_605,N_161);
nand U1121 (N_1121,N_574,N_190);
or U1122 (N_1122,N_420,N_706);
xor U1123 (N_1123,N_606,N_248);
xor U1124 (N_1124,N_117,N_171);
or U1125 (N_1125,N_303,N_293);
nand U1126 (N_1126,N_259,N_452);
xor U1127 (N_1127,N_153,N_346);
and U1128 (N_1128,N_172,N_709);
xor U1129 (N_1129,N_679,N_345);
nand U1130 (N_1130,N_586,N_427);
and U1131 (N_1131,N_33,N_669);
or U1132 (N_1132,N_610,N_401);
nand U1133 (N_1133,N_585,N_695);
and U1134 (N_1134,N_624,N_489);
xnor U1135 (N_1135,N_345,N_242);
xnor U1136 (N_1136,N_241,N_323);
or U1137 (N_1137,N_514,N_3);
and U1138 (N_1138,N_110,N_414);
nand U1139 (N_1139,N_219,N_439);
and U1140 (N_1140,N_692,N_705);
nor U1141 (N_1141,N_256,N_342);
or U1142 (N_1142,N_164,N_22);
nor U1143 (N_1143,N_396,N_569);
and U1144 (N_1144,N_222,N_239);
nor U1145 (N_1145,N_544,N_395);
and U1146 (N_1146,N_190,N_657);
nand U1147 (N_1147,N_86,N_177);
or U1148 (N_1148,N_173,N_699);
or U1149 (N_1149,N_251,N_698);
or U1150 (N_1150,N_315,N_694);
nand U1151 (N_1151,N_141,N_312);
nor U1152 (N_1152,N_316,N_4);
nor U1153 (N_1153,N_704,N_94);
or U1154 (N_1154,N_13,N_571);
or U1155 (N_1155,N_670,N_139);
nand U1156 (N_1156,N_126,N_289);
and U1157 (N_1157,N_525,N_602);
nand U1158 (N_1158,N_588,N_205);
xnor U1159 (N_1159,N_373,N_424);
and U1160 (N_1160,N_506,N_64);
nor U1161 (N_1161,N_741,N_745);
xnor U1162 (N_1162,N_510,N_671);
xnor U1163 (N_1163,N_36,N_464);
nor U1164 (N_1164,N_539,N_28);
nor U1165 (N_1165,N_674,N_108);
xor U1166 (N_1166,N_162,N_251);
nand U1167 (N_1167,N_711,N_358);
or U1168 (N_1168,N_659,N_702);
nand U1169 (N_1169,N_548,N_338);
xnor U1170 (N_1170,N_34,N_455);
and U1171 (N_1171,N_311,N_346);
or U1172 (N_1172,N_339,N_266);
and U1173 (N_1173,N_675,N_539);
or U1174 (N_1174,N_651,N_364);
xor U1175 (N_1175,N_393,N_554);
nand U1176 (N_1176,N_306,N_423);
and U1177 (N_1177,N_142,N_420);
nand U1178 (N_1178,N_664,N_509);
nand U1179 (N_1179,N_349,N_288);
xnor U1180 (N_1180,N_732,N_618);
or U1181 (N_1181,N_443,N_439);
or U1182 (N_1182,N_308,N_437);
and U1183 (N_1183,N_533,N_291);
xnor U1184 (N_1184,N_410,N_403);
xor U1185 (N_1185,N_636,N_287);
nor U1186 (N_1186,N_431,N_730);
xnor U1187 (N_1187,N_390,N_635);
nand U1188 (N_1188,N_363,N_160);
or U1189 (N_1189,N_49,N_683);
and U1190 (N_1190,N_412,N_27);
and U1191 (N_1191,N_108,N_68);
or U1192 (N_1192,N_309,N_25);
or U1193 (N_1193,N_418,N_245);
xnor U1194 (N_1194,N_507,N_106);
nand U1195 (N_1195,N_355,N_87);
nand U1196 (N_1196,N_652,N_657);
nand U1197 (N_1197,N_743,N_565);
nor U1198 (N_1198,N_406,N_289);
nor U1199 (N_1199,N_117,N_235);
or U1200 (N_1200,N_536,N_269);
and U1201 (N_1201,N_219,N_131);
nor U1202 (N_1202,N_15,N_714);
xnor U1203 (N_1203,N_341,N_99);
nor U1204 (N_1204,N_340,N_264);
nand U1205 (N_1205,N_470,N_165);
nand U1206 (N_1206,N_100,N_386);
nor U1207 (N_1207,N_197,N_114);
xor U1208 (N_1208,N_121,N_338);
and U1209 (N_1209,N_381,N_9);
or U1210 (N_1210,N_371,N_517);
xor U1211 (N_1211,N_597,N_269);
or U1212 (N_1212,N_653,N_64);
nand U1213 (N_1213,N_113,N_595);
or U1214 (N_1214,N_530,N_632);
or U1215 (N_1215,N_596,N_220);
nand U1216 (N_1216,N_667,N_488);
or U1217 (N_1217,N_84,N_482);
nor U1218 (N_1218,N_730,N_198);
nor U1219 (N_1219,N_360,N_122);
and U1220 (N_1220,N_201,N_220);
and U1221 (N_1221,N_614,N_8);
xnor U1222 (N_1222,N_652,N_520);
nor U1223 (N_1223,N_160,N_397);
nor U1224 (N_1224,N_617,N_550);
and U1225 (N_1225,N_727,N_636);
nand U1226 (N_1226,N_672,N_172);
and U1227 (N_1227,N_682,N_656);
and U1228 (N_1228,N_636,N_327);
and U1229 (N_1229,N_580,N_132);
and U1230 (N_1230,N_308,N_148);
or U1231 (N_1231,N_703,N_55);
xnor U1232 (N_1232,N_35,N_415);
and U1233 (N_1233,N_409,N_355);
nand U1234 (N_1234,N_616,N_503);
or U1235 (N_1235,N_415,N_115);
xor U1236 (N_1236,N_586,N_723);
or U1237 (N_1237,N_565,N_483);
and U1238 (N_1238,N_636,N_739);
or U1239 (N_1239,N_176,N_342);
nand U1240 (N_1240,N_142,N_91);
nand U1241 (N_1241,N_351,N_583);
xor U1242 (N_1242,N_607,N_37);
nor U1243 (N_1243,N_211,N_20);
and U1244 (N_1244,N_203,N_389);
or U1245 (N_1245,N_265,N_240);
nor U1246 (N_1246,N_125,N_583);
nor U1247 (N_1247,N_60,N_345);
nand U1248 (N_1248,N_260,N_553);
nand U1249 (N_1249,N_77,N_748);
nor U1250 (N_1250,N_715,N_645);
xor U1251 (N_1251,N_560,N_743);
nand U1252 (N_1252,N_5,N_591);
nand U1253 (N_1253,N_138,N_412);
nand U1254 (N_1254,N_550,N_148);
nand U1255 (N_1255,N_460,N_477);
nand U1256 (N_1256,N_282,N_288);
and U1257 (N_1257,N_344,N_269);
and U1258 (N_1258,N_734,N_239);
and U1259 (N_1259,N_517,N_416);
xor U1260 (N_1260,N_421,N_125);
xnor U1261 (N_1261,N_532,N_747);
xor U1262 (N_1262,N_726,N_244);
xor U1263 (N_1263,N_284,N_517);
and U1264 (N_1264,N_77,N_417);
and U1265 (N_1265,N_19,N_165);
xnor U1266 (N_1266,N_478,N_673);
or U1267 (N_1267,N_522,N_303);
and U1268 (N_1268,N_747,N_188);
nand U1269 (N_1269,N_407,N_488);
or U1270 (N_1270,N_426,N_721);
nand U1271 (N_1271,N_580,N_739);
nor U1272 (N_1272,N_166,N_317);
nor U1273 (N_1273,N_197,N_29);
and U1274 (N_1274,N_28,N_679);
or U1275 (N_1275,N_286,N_574);
nor U1276 (N_1276,N_94,N_664);
and U1277 (N_1277,N_606,N_141);
and U1278 (N_1278,N_216,N_390);
or U1279 (N_1279,N_559,N_331);
or U1280 (N_1280,N_191,N_473);
nand U1281 (N_1281,N_723,N_362);
nor U1282 (N_1282,N_732,N_189);
or U1283 (N_1283,N_181,N_314);
nor U1284 (N_1284,N_463,N_664);
nor U1285 (N_1285,N_11,N_56);
xnor U1286 (N_1286,N_277,N_614);
xnor U1287 (N_1287,N_264,N_358);
nor U1288 (N_1288,N_572,N_95);
nand U1289 (N_1289,N_83,N_533);
nor U1290 (N_1290,N_618,N_132);
xnor U1291 (N_1291,N_131,N_85);
and U1292 (N_1292,N_422,N_473);
xnor U1293 (N_1293,N_353,N_510);
xnor U1294 (N_1294,N_413,N_61);
nand U1295 (N_1295,N_497,N_376);
nand U1296 (N_1296,N_44,N_690);
and U1297 (N_1297,N_0,N_83);
or U1298 (N_1298,N_494,N_479);
nand U1299 (N_1299,N_476,N_722);
xor U1300 (N_1300,N_128,N_355);
or U1301 (N_1301,N_132,N_86);
nor U1302 (N_1302,N_421,N_2);
nand U1303 (N_1303,N_366,N_233);
and U1304 (N_1304,N_89,N_659);
nand U1305 (N_1305,N_341,N_410);
nor U1306 (N_1306,N_652,N_39);
or U1307 (N_1307,N_407,N_559);
xnor U1308 (N_1308,N_304,N_244);
nand U1309 (N_1309,N_130,N_654);
xor U1310 (N_1310,N_540,N_115);
nand U1311 (N_1311,N_148,N_461);
nand U1312 (N_1312,N_544,N_444);
or U1313 (N_1313,N_183,N_86);
and U1314 (N_1314,N_483,N_669);
or U1315 (N_1315,N_496,N_470);
nand U1316 (N_1316,N_700,N_283);
and U1317 (N_1317,N_53,N_70);
and U1318 (N_1318,N_125,N_730);
and U1319 (N_1319,N_122,N_729);
and U1320 (N_1320,N_660,N_62);
nor U1321 (N_1321,N_707,N_487);
or U1322 (N_1322,N_181,N_705);
or U1323 (N_1323,N_537,N_109);
xor U1324 (N_1324,N_506,N_108);
nand U1325 (N_1325,N_563,N_97);
nand U1326 (N_1326,N_253,N_418);
nor U1327 (N_1327,N_537,N_383);
nand U1328 (N_1328,N_704,N_736);
and U1329 (N_1329,N_261,N_85);
xnor U1330 (N_1330,N_271,N_82);
or U1331 (N_1331,N_554,N_298);
or U1332 (N_1332,N_675,N_708);
xnor U1333 (N_1333,N_527,N_298);
or U1334 (N_1334,N_584,N_728);
nor U1335 (N_1335,N_197,N_566);
nor U1336 (N_1336,N_180,N_518);
xnor U1337 (N_1337,N_733,N_490);
xor U1338 (N_1338,N_214,N_346);
xnor U1339 (N_1339,N_74,N_687);
or U1340 (N_1340,N_5,N_449);
xor U1341 (N_1341,N_18,N_500);
nand U1342 (N_1342,N_148,N_358);
nand U1343 (N_1343,N_512,N_559);
nand U1344 (N_1344,N_733,N_58);
and U1345 (N_1345,N_294,N_686);
xor U1346 (N_1346,N_211,N_421);
and U1347 (N_1347,N_530,N_382);
or U1348 (N_1348,N_5,N_613);
and U1349 (N_1349,N_394,N_386);
nor U1350 (N_1350,N_630,N_398);
and U1351 (N_1351,N_39,N_521);
and U1352 (N_1352,N_575,N_72);
xnor U1353 (N_1353,N_739,N_677);
or U1354 (N_1354,N_230,N_160);
or U1355 (N_1355,N_503,N_696);
nor U1356 (N_1356,N_341,N_73);
nor U1357 (N_1357,N_14,N_669);
nand U1358 (N_1358,N_426,N_251);
xnor U1359 (N_1359,N_192,N_311);
nor U1360 (N_1360,N_274,N_136);
nor U1361 (N_1361,N_143,N_48);
or U1362 (N_1362,N_664,N_377);
and U1363 (N_1363,N_237,N_385);
or U1364 (N_1364,N_202,N_171);
xor U1365 (N_1365,N_210,N_213);
xor U1366 (N_1366,N_172,N_262);
nor U1367 (N_1367,N_498,N_250);
or U1368 (N_1368,N_551,N_408);
xnor U1369 (N_1369,N_718,N_437);
xor U1370 (N_1370,N_723,N_346);
or U1371 (N_1371,N_475,N_30);
nand U1372 (N_1372,N_348,N_244);
and U1373 (N_1373,N_508,N_111);
nor U1374 (N_1374,N_119,N_478);
and U1375 (N_1375,N_207,N_613);
or U1376 (N_1376,N_112,N_88);
nand U1377 (N_1377,N_593,N_451);
xnor U1378 (N_1378,N_245,N_615);
nand U1379 (N_1379,N_35,N_382);
xor U1380 (N_1380,N_259,N_497);
or U1381 (N_1381,N_355,N_576);
or U1382 (N_1382,N_475,N_50);
nor U1383 (N_1383,N_738,N_53);
xnor U1384 (N_1384,N_560,N_507);
or U1385 (N_1385,N_645,N_65);
or U1386 (N_1386,N_135,N_579);
xor U1387 (N_1387,N_276,N_165);
nor U1388 (N_1388,N_565,N_396);
nand U1389 (N_1389,N_188,N_102);
nand U1390 (N_1390,N_29,N_745);
nand U1391 (N_1391,N_605,N_505);
xor U1392 (N_1392,N_232,N_527);
nand U1393 (N_1393,N_578,N_112);
nand U1394 (N_1394,N_696,N_402);
or U1395 (N_1395,N_582,N_458);
or U1396 (N_1396,N_112,N_535);
and U1397 (N_1397,N_389,N_628);
or U1398 (N_1398,N_648,N_394);
nand U1399 (N_1399,N_5,N_31);
xnor U1400 (N_1400,N_228,N_61);
xnor U1401 (N_1401,N_65,N_179);
nand U1402 (N_1402,N_130,N_417);
nand U1403 (N_1403,N_414,N_239);
and U1404 (N_1404,N_356,N_483);
and U1405 (N_1405,N_571,N_466);
nand U1406 (N_1406,N_409,N_380);
xnor U1407 (N_1407,N_166,N_457);
xnor U1408 (N_1408,N_562,N_185);
nand U1409 (N_1409,N_224,N_691);
nand U1410 (N_1410,N_311,N_172);
and U1411 (N_1411,N_651,N_54);
and U1412 (N_1412,N_75,N_46);
and U1413 (N_1413,N_77,N_326);
and U1414 (N_1414,N_213,N_159);
or U1415 (N_1415,N_646,N_5);
nor U1416 (N_1416,N_20,N_150);
nor U1417 (N_1417,N_408,N_341);
and U1418 (N_1418,N_702,N_225);
or U1419 (N_1419,N_641,N_418);
and U1420 (N_1420,N_272,N_412);
and U1421 (N_1421,N_681,N_101);
nor U1422 (N_1422,N_441,N_83);
nor U1423 (N_1423,N_496,N_100);
xor U1424 (N_1424,N_418,N_313);
and U1425 (N_1425,N_685,N_499);
and U1426 (N_1426,N_695,N_592);
or U1427 (N_1427,N_226,N_650);
nor U1428 (N_1428,N_366,N_560);
nand U1429 (N_1429,N_67,N_142);
and U1430 (N_1430,N_728,N_0);
xnor U1431 (N_1431,N_317,N_385);
nor U1432 (N_1432,N_531,N_558);
or U1433 (N_1433,N_537,N_137);
xor U1434 (N_1434,N_682,N_603);
nand U1435 (N_1435,N_395,N_506);
xor U1436 (N_1436,N_258,N_69);
xor U1437 (N_1437,N_311,N_240);
xor U1438 (N_1438,N_403,N_171);
nor U1439 (N_1439,N_347,N_288);
or U1440 (N_1440,N_203,N_623);
and U1441 (N_1441,N_409,N_713);
xnor U1442 (N_1442,N_158,N_240);
and U1443 (N_1443,N_712,N_409);
xor U1444 (N_1444,N_243,N_488);
nand U1445 (N_1445,N_267,N_582);
nor U1446 (N_1446,N_112,N_675);
and U1447 (N_1447,N_56,N_257);
nor U1448 (N_1448,N_450,N_51);
xnor U1449 (N_1449,N_412,N_231);
and U1450 (N_1450,N_481,N_9);
nor U1451 (N_1451,N_280,N_645);
xnor U1452 (N_1452,N_252,N_480);
nor U1453 (N_1453,N_453,N_573);
xor U1454 (N_1454,N_371,N_130);
and U1455 (N_1455,N_30,N_75);
and U1456 (N_1456,N_649,N_319);
or U1457 (N_1457,N_259,N_543);
and U1458 (N_1458,N_701,N_232);
or U1459 (N_1459,N_404,N_519);
xor U1460 (N_1460,N_717,N_313);
nand U1461 (N_1461,N_406,N_301);
and U1462 (N_1462,N_527,N_320);
or U1463 (N_1463,N_510,N_220);
nand U1464 (N_1464,N_491,N_370);
xor U1465 (N_1465,N_63,N_390);
nor U1466 (N_1466,N_742,N_364);
or U1467 (N_1467,N_531,N_8);
xnor U1468 (N_1468,N_546,N_42);
nand U1469 (N_1469,N_412,N_42);
and U1470 (N_1470,N_508,N_728);
and U1471 (N_1471,N_176,N_556);
nand U1472 (N_1472,N_288,N_556);
nand U1473 (N_1473,N_658,N_198);
nand U1474 (N_1474,N_32,N_8);
and U1475 (N_1475,N_363,N_359);
nor U1476 (N_1476,N_545,N_223);
or U1477 (N_1477,N_654,N_30);
or U1478 (N_1478,N_93,N_45);
nand U1479 (N_1479,N_521,N_365);
nor U1480 (N_1480,N_639,N_159);
nand U1481 (N_1481,N_385,N_152);
and U1482 (N_1482,N_260,N_4);
xnor U1483 (N_1483,N_6,N_107);
nand U1484 (N_1484,N_418,N_581);
nand U1485 (N_1485,N_651,N_424);
and U1486 (N_1486,N_518,N_71);
or U1487 (N_1487,N_454,N_660);
nor U1488 (N_1488,N_470,N_716);
nand U1489 (N_1489,N_218,N_582);
or U1490 (N_1490,N_562,N_615);
xnor U1491 (N_1491,N_471,N_638);
and U1492 (N_1492,N_355,N_578);
and U1493 (N_1493,N_403,N_268);
nor U1494 (N_1494,N_519,N_452);
and U1495 (N_1495,N_248,N_444);
or U1496 (N_1496,N_29,N_252);
or U1497 (N_1497,N_737,N_319);
nand U1498 (N_1498,N_698,N_196);
xnor U1499 (N_1499,N_250,N_115);
or U1500 (N_1500,N_1432,N_1428);
nand U1501 (N_1501,N_1497,N_1458);
nand U1502 (N_1502,N_940,N_1258);
nand U1503 (N_1503,N_1046,N_1347);
xor U1504 (N_1504,N_984,N_1254);
and U1505 (N_1505,N_1020,N_1293);
nor U1506 (N_1506,N_1282,N_771);
nor U1507 (N_1507,N_1337,N_1405);
nand U1508 (N_1508,N_843,N_1033);
xnor U1509 (N_1509,N_822,N_900);
xnor U1510 (N_1510,N_1461,N_1292);
xnor U1511 (N_1511,N_787,N_1081);
or U1512 (N_1512,N_1335,N_1499);
xnor U1513 (N_1513,N_1099,N_1010);
nand U1514 (N_1514,N_1225,N_1174);
nand U1515 (N_1515,N_1267,N_1249);
or U1516 (N_1516,N_781,N_1275);
xor U1517 (N_1517,N_1440,N_1086);
xor U1518 (N_1518,N_1131,N_1412);
nand U1519 (N_1519,N_1236,N_850);
nor U1520 (N_1520,N_773,N_1318);
nand U1521 (N_1521,N_1492,N_1379);
xor U1522 (N_1522,N_1392,N_1423);
nor U1523 (N_1523,N_963,N_1052);
xnor U1524 (N_1524,N_1083,N_1127);
nand U1525 (N_1525,N_942,N_1111);
nand U1526 (N_1526,N_955,N_1448);
xnor U1527 (N_1527,N_1303,N_837);
nand U1528 (N_1528,N_1186,N_1212);
nand U1529 (N_1529,N_758,N_859);
and U1530 (N_1530,N_829,N_1168);
and U1531 (N_1531,N_1334,N_1073);
nand U1532 (N_1532,N_795,N_925);
nor U1533 (N_1533,N_1313,N_941);
xnor U1534 (N_1534,N_928,N_1351);
xnor U1535 (N_1535,N_782,N_968);
or U1536 (N_1536,N_1365,N_1358);
and U1537 (N_1537,N_1354,N_1382);
nand U1538 (N_1538,N_1326,N_969);
xnor U1539 (N_1539,N_977,N_1253);
xor U1540 (N_1540,N_1203,N_993);
and U1541 (N_1541,N_1281,N_1116);
or U1542 (N_1542,N_1134,N_1418);
and U1543 (N_1543,N_912,N_1399);
or U1544 (N_1544,N_1336,N_1150);
nand U1545 (N_1545,N_1393,N_1265);
xor U1546 (N_1546,N_1179,N_750);
nand U1547 (N_1547,N_897,N_1145);
nand U1548 (N_1548,N_798,N_1343);
or U1549 (N_1549,N_1471,N_1012);
or U1550 (N_1550,N_1095,N_1284);
or U1551 (N_1551,N_1328,N_1390);
and U1552 (N_1552,N_863,N_1270);
xnor U1553 (N_1553,N_943,N_1064);
and U1554 (N_1554,N_1210,N_1307);
nor U1555 (N_1555,N_842,N_1325);
or U1556 (N_1556,N_1066,N_1297);
nand U1557 (N_1557,N_905,N_820);
and U1558 (N_1558,N_1115,N_865);
nand U1559 (N_1559,N_869,N_1030);
nand U1560 (N_1560,N_1202,N_1463);
and U1561 (N_1561,N_929,N_1079);
nor U1562 (N_1562,N_1386,N_828);
nand U1563 (N_1563,N_777,N_1108);
or U1564 (N_1564,N_1072,N_906);
or U1565 (N_1565,N_1170,N_1209);
or U1566 (N_1566,N_1451,N_1213);
nand U1567 (N_1567,N_1027,N_1067);
nor U1568 (N_1568,N_967,N_1457);
or U1569 (N_1569,N_1375,N_1415);
xnor U1570 (N_1570,N_1479,N_1402);
nand U1571 (N_1571,N_910,N_803);
nor U1572 (N_1572,N_792,N_805);
nor U1573 (N_1573,N_919,N_1446);
xnor U1574 (N_1574,N_1107,N_1201);
or U1575 (N_1575,N_1369,N_1009);
and U1576 (N_1576,N_1319,N_1105);
xnor U1577 (N_1577,N_1345,N_1187);
nor U1578 (N_1578,N_946,N_1207);
and U1579 (N_1579,N_997,N_961);
or U1580 (N_1580,N_1262,N_1023);
nand U1581 (N_1581,N_834,N_809);
or U1582 (N_1582,N_1443,N_1288);
or U1583 (N_1583,N_1407,N_938);
nor U1584 (N_1584,N_838,N_1389);
nand U1585 (N_1585,N_1192,N_1077);
and U1586 (N_1586,N_1000,N_1024);
and U1587 (N_1587,N_1229,N_880);
xor U1588 (N_1588,N_1406,N_867);
xnor U1589 (N_1589,N_1005,N_1339);
and U1590 (N_1590,N_1039,N_960);
or U1591 (N_1591,N_995,N_1093);
or U1592 (N_1592,N_1460,N_1472);
nand U1593 (N_1593,N_1333,N_1287);
nand U1594 (N_1594,N_918,N_1200);
or U1595 (N_1595,N_1036,N_1342);
nand U1596 (N_1596,N_879,N_1137);
nand U1597 (N_1597,N_807,N_1427);
nand U1598 (N_1598,N_1422,N_1260);
or U1599 (N_1599,N_1188,N_1006);
or U1600 (N_1600,N_1181,N_889);
and U1601 (N_1601,N_1147,N_904);
or U1602 (N_1602,N_1104,N_931);
and U1603 (N_1603,N_1372,N_896);
and U1604 (N_1604,N_770,N_1491);
nor U1605 (N_1605,N_1165,N_1082);
xor U1606 (N_1606,N_1241,N_1435);
xor U1607 (N_1607,N_887,N_1196);
nand U1608 (N_1608,N_1475,N_1214);
nor U1609 (N_1609,N_1255,N_1444);
nand U1610 (N_1610,N_1374,N_1465);
nand U1611 (N_1611,N_785,N_1110);
nand U1612 (N_1612,N_1172,N_1280);
or U1613 (N_1613,N_893,N_1143);
or U1614 (N_1614,N_1273,N_1154);
nor U1615 (N_1615,N_1349,N_1166);
xor U1616 (N_1616,N_1447,N_1118);
and U1617 (N_1617,N_1388,N_835);
nor U1618 (N_1618,N_1032,N_878);
nor U1619 (N_1619,N_1062,N_965);
and U1620 (N_1620,N_1332,N_1261);
nor U1621 (N_1621,N_826,N_877);
or U1622 (N_1622,N_1121,N_907);
and U1623 (N_1623,N_1409,N_934);
or U1624 (N_1624,N_1431,N_1051);
and U1625 (N_1625,N_1139,N_1157);
nor U1626 (N_1626,N_1160,N_884);
or U1627 (N_1627,N_1259,N_866);
nor U1628 (N_1628,N_913,N_1123);
or U1629 (N_1629,N_1194,N_1411);
nor U1630 (N_1630,N_830,N_1169);
xor U1631 (N_1631,N_839,N_1494);
and U1632 (N_1632,N_1290,N_1218);
nor U1633 (N_1633,N_761,N_1119);
nand U1634 (N_1634,N_936,N_1237);
nor U1635 (N_1635,N_851,N_808);
nor U1636 (N_1636,N_767,N_1245);
or U1637 (N_1637,N_1314,N_1294);
and U1638 (N_1638,N_1059,N_1408);
nor U1639 (N_1639,N_1084,N_1252);
nor U1640 (N_1640,N_1430,N_1204);
and U1641 (N_1641,N_799,N_1383);
nor U1642 (N_1642,N_760,N_1025);
nand U1643 (N_1643,N_1173,N_1381);
or U1644 (N_1644,N_1056,N_1128);
xor U1645 (N_1645,N_1223,N_1308);
nor U1646 (N_1646,N_1346,N_1161);
and U1647 (N_1647,N_1243,N_1031);
nand U1648 (N_1648,N_915,N_1164);
nand U1649 (N_1649,N_999,N_1352);
and U1650 (N_1650,N_847,N_778);
nand U1651 (N_1651,N_939,N_1331);
nor U1652 (N_1652,N_1060,N_914);
nand U1653 (N_1653,N_1038,N_1410);
or U1654 (N_1654,N_1050,N_890);
xor U1655 (N_1655,N_844,N_860);
or U1656 (N_1656,N_1055,N_1271);
and U1657 (N_1657,N_1250,N_895);
and U1658 (N_1658,N_1348,N_1124);
xor U1659 (N_1659,N_1324,N_875);
xnor U1660 (N_1660,N_1268,N_1026);
nor U1661 (N_1661,N_762,N_1011);
nor U1662 (N_1662,N_956,N_1106);
or U1663 (N_1663,N_1125,N_814);
and U1664 (N_1664,N_1103,N_901);
xor U1665 (N_1665,N_1069,N_924);
or U1666 (N_1666,N_1433,N_797);
xnor U1667 (N_1667,N_786,N_796);
nor U1668 (N_1668,N_979,N_1498);
nor U1669 (N_1669,N_1016,N_1013);
and U1670 (N_1670,N_983,N_1053);
xor U1671 (N_1671,N_1248,N_1340);
xnor U1672 (N_1672,N_1305,N_1378);
or U1673 (N_1673,N_1240,N_1112);
or U1674 (N_1674,N_1075,N_1063);
nand U1675 (N_1675,N_923,N_1100);
nand U1676 (N_1676,N_794,N_861);
nand U1677 (N_1677,N_1442,N_1473);
xor U1678 (N_1678,N_886,N_1163);
xnor U1679 (N_1679,N_802,N_998);
xor U1680 (N_1680,N_751,N_1138);
nor U1681 (N_1681,N_1384,N_789);
xor U1682 (N_1682,N_1436,N_1074);
or U1683 (N_1683,N_1306,N_1417);
nand U1684 (N_1684,N_1329,N_1048);
nand U1685 (N_1685,N_1373,N_1330);
and U1686 (N_1686,N_817,N_1396);
and U1687 (N_1687,N_1395,N_823);
nand U1688 (N_1688,N_1028,N_1061);
nor U1689 (N_1689,N_1485,N_1449);
nand U1690 (N_1690,N_1316,N_1088);
xnor U1691 (N_1691,N_1301,N_1017);
nor U1692 (N_1692,N_892,N_1155);
nand U1693 (N_1693,N_1018,N_1320);
xnor U1694 (N_1694,N_874,N_945);
xor U1695 (N_1695,N_1247,N_1054);
xnor U1696 (N_1696,N_972,N_981);
nor U1697 (N_1697,N_811,N_1311);
nand U1698 (N_1698,N_1178,N_1175);
xnor U1699 (N_1699,N_1357,N_1456);
nor U1700 (N_1700,N_1484,N_849);
xnor U1701 (N_1701,N_1226,N_1129);
or U1702 (N_1702,N_1044,N_898);
and U1703 (N_1703,N_780,N_1003);
and U1704 (N_1704,N_793,N_1257);
and U1705 (N_1705,N_1263,N_756);
xor U1706 (N_1706,N_1092,N_916);
nor U1707 (N_1707,N_1397,N_1487);
and U1708 (N_1708,N_1199,N_985);
xnor U1709 (N_1709,N_894,N_1219);
and U1710 (N_1710,N_1228,N_1158);
and U1711 (N_1711,N_1042,N_1264);
and U1712 (N_1712,N_774,N_1398);
and U1713 (N_1713,N_1424,N_824);
nand U1714 (N_1714,N_818,N_1058);
xor U1715 (N_1715,N_1438,N_1477);
nor U1716 (N_1716,N_1437,N_1285);
xnor U1717 (N_1717,N_1327,N_1295);
xor U1718 (N_1718,N_765,N_954);
nand U1719 (N_1719,N_806,N_1117);
nand U1720 (N_1720,N_1312,N_1216);
or U1721 (N_1721,N_1470,N_1286);
or U1722 (N_1722,N_821,N_1230);
nand U1723 (N_1723,N_1356,N_1221);
nand U1724 (N_1724,N_1101,N_813);
xnor U1725 (N_1725,N_926,N_1183);
or U1726 (N_1726,N_958,N_982);
or U1727 (N_1727,N_1469,N_949);
nand U1728 (N_1728,N_1246,N_1141);
or U1729 (N_1729,N_1146,N_920);
nand U1730 (N_1730,N_1120,N_973);
nand U1731 (N_1731,N_1135,N_902);
and U1732 (N_1732,N_976,N_1231);
nor U1733 (N_1733,N_1495,N_975);
xor U1734 (N_1734,N_1377,N_1490);
nor U1735 (N_1735,N_1130,N_930);
nand U1736 (N_1736,N_853,N_921);
nor U1737 (N_1737,N_856,N_1300);
and U1738 (N_1738,N_1162,N_812);
nand U1739 (N_1739,N_1021,N_841);
and U1740 (N_1740,N_1047,N_991);
xor U1741 (N_1741,N_1208,N_1310);
nand U1742 (N_1742,N_827,N_1233);
and U1743 (N_1743,N_1489,N_1114);
xor U1744 (N_1744,N_1113,N_980);
nand U1745 (N_1745,N_953,N_840);
nand U1746 (N_1746,N_1291,N_1482);
xor U1747 (N_1747,N_1467,N_864);
nor U1748 (N_1748,N_1171,N_1279);
or U1749 (N_1749,N_957,N_784);
and U1750 (N_1750,N_833,N_1454);
nor U1751 (N_1751,N_882,N_810);
and U1752 (N_1752,N_1420,N_1078);
or U1753 (N_1753,N_1429,N_801);
xor U1754 (N_1754,N_752,N_1401);
and U1755 (N_1755,N_1122,N_1140);
and U1756 (N_1756,N_816,N_1272);
nand U1757 (N_1757,N_1015,N_1296);
nor U1758 (N_1758,N_1387,N_854);
and U1759 (N_1759,N_962,N_764);
xnor U1760 (N_1760,N_1089,N_1197);
nand U1761 (N_1761,N_911,N_1496);
nor U1762 (N_1762,N_1205,N_988);
xor U1763 (N_1763,N_870,N_1190);
xor U1764 (N_1764,N_1298,N_1156);
nor U1765 (N_1765,N_964,N_927);
nor U1766 (N_1766,N_768,N_1421);
nor U1767 (N_1767,N_1302,N_1283);
xnor U1768 (N_1768,N_1317,N_757);
and U1769 (N_1769,N_951,N_868);
nand U1770 (N_1770,N_1152,N_1222);
or U1771 (N_1771,N_1094,N_1315);
or U1772 (N_1772,N_1189,N_947);
xnor U1773 (N_1773,N_1468,N_881);
nor U1774 (N_1774,N_1353,N_1483);
nor U1775 (N_1775,N_1344,N_832);
and U1776 (N_1776,N_1478,N_1211);
and U1777 (N_1777,N_800,N_852);
nor U1778 (N_1778,N_1364,N_1041);
nand U1779 (N_1779,N_948,N_1142);
and U1780 (N_1780,N_888,N_1238);
nand U1781 (N_1781,N_1109,N_1087);
nor U1782 (N_1782,N_873,N_1256);
nor U1783 (N_1783,N_1195,N_876);
nor U1784 (N_1784,N_1459,N_990);
xor U1785 (N_1785,N_1132,N_944);
or U1786 (N_1786,N_1151,N_974);
and U1787 (N_1787,N_1480,N_1363);
and U1788 (N_1788,N_1425,N_755);
nor U1789 (N_1789,N_1450,N_1413);
and U1790 (N_1790,N_1133,N_1476);
nor U1791 (N_1791,N_825,N_1419);
and U1792 (N_1792,N_1414,N_1445);
xor U1793 (N_1793,N_1278,N_1182);
nor U1794 (N_1794,N_1368,N_763);
nand U1795 (N_1795,N_1338,N_1350);
xnor U1796 (N_1796,N_788,N_1167);
xnor U1797 (N_1797,N_804,N_1251);
xnor U1798 (N_1798,N_1136,N_885);
xor U1799 (N_1799,N_971,N_1085);
nor U1800 (N_1800,N_1266,N_848);
nor U1801 (N_1801,N_1191,N_1304);
and U1802 (N_1802,N_1022,N_1014);
nand U1803 (N_1803,N_1455,N_1098);
nand U1804 (N_1804,N_1299,N_1486);
and U1805 (N_1805,N_1068,N_1391);
nand U1806 (N_1806,N_1323,N_1227);
xor U1807 (N_1807,N_855,N_1462);
nand U1808 (N_1808,N_922,N_1040);
and U1809 (N_1809,N_754,N_1466);
or U1810 (N_1810,N_909,N_1370);
and U1811 (N_1811,N_753,N_1359);
or U1812 (N_1812,N_1217,N_1057);
or U1813 (N_1813,N_1361,N_1269);
xor U1814 (N_1814,N_772,N_1090);
xor U1815 (N_1815,N_1309,N_1070);
or U1816 (N_1816,N_1439,N_917);
xor U1817 (N_1817,N_1185,N_1234);
or U1818 (N_1818,N_1376,N_1274);
or U1819 (N_1819,N_836,N_858);
xnor U1820 (N_1820,N_1224,N_1242);
or U1821 (N_1821,N_862,N_1341);
nor U1822 (N_1822,N_1276,N_1091);
or U1823 (N_1823,N_1029,N_1159);
nand U1824 (N_1824,N_1096,N_1180);
xnor U1825 (N_1825,N_1474,N_1049);
xor U1826 (N_1826,N_908,N_883);
and U1827 (N_1827,N_1277,N_1148);
and U1828 (N_1828,N_1235,N_1004);
xnor U1829 (N_1829,N_1034,N_1404);
or U1830 (N_1830,N_989,N_1453);
nand U1831 (N_1831,N_769,N_1035);
and U1832 (N_1832,N_1400,N_1321);
or U1833 (N_1833,N_1367,N_1403);
xnor U1834 (N_1834,N_791,N_1149);
nand U1835 (N_1835,N_1193,N_1394);
and U1836 (N_1836,N_966,N_1097);
and U1837 (N_1837,N_857,N_831);
nand U1838 (N_1838,N_1488,N_790);
xnor U1839 (N_1839,N_950,N_1289);
and U1840 (N_1840,N_1215,N_846);
and U1841 (N_1841,N_986,N_1080);
nand U1842 (N_1842,N_1076,N_1206);
or U1843 (N_1843,N_1362,N_933);
or U1844 (N_1844,N_1037,N_766);
or U1845 (N_1845,N_1198,N_935);
and U1846 (N_1846,N_1385,N_819);
and U1847 (N_1847,N_1019,N_1001);
or U1848 (N_1848,N_970,N_1452);
and U1849 (N_1849,N_959,N_937);
xnor U1850 (N_1850,N_903,N_1232);
and U1851 (N_1851,N_1481,N_815);
or U1852 (N_1852,N_994,N_1002);
xnor U1853 (N_1853,N_776,N_872);
nand U1854 (N_1854,N_779,N_1007);
or U1855 (N_1855,N_1008,N_1102);
xnor U1856 (N_1856,N_1360,N_1220);
and U1857 (N_1857,N_1153,N_932);
nand U1858 (N_1858,N_759,N_1366);
or U1859 (N_1859,N_775,N_1464);
xor U1860 (N_1860,N_1176,N_899);
or U1861 (N_1861,N_1355,N_1045);
nor U1862 (N_1862,N_1144,N_1184);
or U1863 (N_1863,N_1177,N_978);
nand U1864 (N_1864,N_783,N_871);
or U1865 (N_1865,N_987,N_1244);
nand U1866 (N_1866,N_1426,N_1239);
or U1867 (N_1867,N_845,N_1071);
nand U1868 (N_1868,N_1043,N_1434);
nand U1869 (N_1869,N_1065,N_1126);
nand U1870 (N_1870,N_1416,N_992);
nand U1871 (N_1871,N_1371,N_1380);
and U1872 (N_1872,N_1441,N_996);
and U1873 (N_1873,N_1493,N_952);
xor U1874 (N_1874,N_891,N_1322);
and U1875 (N_1875,N_1027,N_1066);
nor U1876 (N_1876,N_926,N_1162);
nor U1877 (N_1877,N_1321,N_841);
xnor U1878 (N_1878,N_1390,N_1150);
and U1879 (N_1879,N_1328,N_1114);
nor U1880 (N_1880,N_872,N_1160);
xnor U1881 (N_1881,N_932,N_1100);
xnor U1882 (N_1882,N_1284,N_882);
and U1883 (N_1883,N_1221,N_1425);
nor U1884 (N_1884,N_1066,N_805);
nor U1885 (N_1885,N_1178,N_1307);
and U1886 (N_1886,N_1273,N_1291);
xnor U1887 (N_1887,N_870,N_1110);
nand U1888 (N_1888,N_1450,N_964);
nor U1889 (N_1889,N_1406,N_1126);
xnor U1890 (N_1890,N_1416,N_1273);
xnor U1891 (N_1891,N_831,N_1163);
xnor U1892 (N_1892,N_1330,N_1188);
or U1893 (N_1893,N_1302,N_1441);
xor U1894 (N_1894,N_1452,N_1292);
nor U1895 (N_1895,N_1270,N_1074);
nand U1896 (N_1896,N_758,N_1308);
nand U1897 (N_1897,N_925,N_1064);
nor U1898 (N_1898,N_884,N_1233);
and U1899 (N_1899,N_843,N_801);
or U1900 (N_1900,N_1173,N_967);
xor U1901 (N_1901,N_946,N_1176);
and U1902 (N_1902,N_923,N_1038);
xor U1903 (N_1903,N_1408,N_1355);
nand U1904 (N_1904,N_917,N_998);
xnor U1905 (N_1905,N_1094,N_820);
or U1906 (N_1906,N_1323,N_1124);
and U1907 (N_1907,N_893,N_1272);
xnor U1908 (N_1908,N_1191,N_1447);
xnor U1909 (N_1909,N_826,N_1066);
nor U1910 (N_1910,N_1206,N_1042);
xnor U1911 (N_1911,N_1200,N_1279);
xnor U1912 (N_1912,N_1033,N_1165);
nor U1913 (N_1913,N_1344,N_1161);
nor U1914 (N_1914,N_892,N_1229);
or U1915 (N_1915,N_1092,N_1372);
and U1916 (N_1916,N_750,N_1235);
nand U1917 (N_1917,N_1085,N_1143);
xnor U1918 (N_1918,N_776,N_815);
nand U1919 (N_1919,N_1156,N_1401);
or U1920 (N_1920,N_1212,N_1410);
xor U1921 (N_1921,N_1294,N_1496);
nand U1922 (N_1922,N_1211,N_1173);
xor U1923 (N_1923,N_873,N_1347);
nor U1924 (N_1924,N_1484,N_787);
and U1925 (N_1925,N_958,N_802);
nor U1926 (N_1926,N_1451,N_1340);
xnor U1927 (N_1927,N_915,N_867);
xor U1928 (N_1928,N_929,N_1025);
xor U1929 (N_1929,N_1181,N_911);
nand U1930 (N_1930,N_1072,N_1411);
nand U1931 (N_1931,N_1119,N_1160);
xnor U1932 (N_1932,N_1224,N_877);
or U1933 (N_1933,N_1408,N_1260);
or U1934 (N_1934,N_1192,N_1333);
nor U1935 (N_1935,N_1300,N_860);
xnor U1936 (N_1936,N_1039,N_1280);
xor U1937 (N_1937,N_1142,N_1144);
nand U1938 (N_1938,N_1332,N_969);
xor U1939 (N_1939,N_943,N_827);
nand U1940 (N_1940,N_1007,N_1157);
or U1941 (N_1941,N_1250,N_1230);
and U1942 (N_1942,N_1212,N_1382);
nand U1943 (N_1943,N_1376,N_1062);
nor U1944 (N_1944,N_878,N_862);
nand U1945 (N_1945,N_991,N_1098);
and U1946 (N_1946,N_1068,N_986);
nor U1947 (N_1947,N_965,N_1390);
and U1948 (N_1948,N_1121,N_1377);
or U1949 (N_1949,N_1339,N_1146);
xnor U1950 (N_1950,N_1369,N_1137);
or U1951 (N_1951,N_1313,N_1355);
nand U1952 (N_1952,N_952,N_997);
nor U1953 (N_1953,N_1353,N_1294);
or U1954 (N_1954,N_1343,N_784);
nand U1955 (N_1955,N_1170,N_1302);
and U1956 (N_1956,N_1242,N_1356);
nor U1957 (N_1957,N_1151,N_1382);
nand U1958 (N_1958,N_947,N_1458);
and U1959 (N_1959,N_1373,N_1139);
nand U1960 (N_1960,N_785,N_918);
and U1961 (N_1961,N_860,N_1374);
or U1962 (N_1962,N_916,N_857);
or U1963 (N_1963,N_889,N_990);
and U1964 (N_1964,N_1087,N_1431);
nand U1965 (N_1965,N_821,N_971);
nor U1966 (N_1966,N_1031,N_914);
or U1967 (N_1967,N_889,N_1375);
nand U1968 (N_1968,N_882,N_1441);
nand U1969 (N_1969,N_965,N_1350);
and U1970 (N_1970,N_986,N_973);
xor U1971 (N_1971,N_1374,N_1229);
nor U1972 (N_1972,N_806,N_1009);
and U1973 (N_1973,N_1325,N_759);
nand U1974 (N_1974,N_1476,N_1251);
xor U1975 (N_1975,N_867,N_896);
or U1976 (N_1976,N_769,N_984);
or U1977 (N_1977,N_1458,N_977);
nand U1978 (N_1978,N_830,N_1165);
nand U1979 (N_1979,N_796,N_1176);
or U1980 (N_1980,N_1136,N_1249);
xor U1981 (N_1981,N_852,N_799);
or U1982 (N_1982,N_861,N_1483);
nor U1983 (N_1983,N_1077,N_780);
xor U1984 (N_1984,N_983,N_794);
nor U1985 (N_1985,N_1304,N_873);
xor U1986 (N_1986,N_1152,N_1209);
or U1987 (N_1987,N_1099,N_1309);
or U1988 (N_1988,N_887,N_1064);
or U1989 (N_1989,N_992,N_1394);
nand U1990 (N_1990,N_1088,N_951);
nand U1991 (N_1991,N_1013,N_1252);
or U1992 (N_1992,N_1226,N_791);
nor U1993 (N_1993,N_1116,N_1143);
and U1994 (N_1994,N_780,N_1052);
nor U1995 (N_1995,N_1122,N_1383);
xor U1996 (N_1996,N_757,N_1426);
xor U1997 (N_1997,N_1100,N_1493);
and U1998 (N_1998,N_1336,N_1306);
nor U1999 (N_1999,N_922,N_960);
nor U2000 (N_2000,N_1120,N_906);
or U2001 (N_2001,N_897,N_759);
or U2002 (N_2002,N_827,N_1017);
or U2003 (N_2003,N_1395,N_839);
nand U2004 (N_2004,N_1137,N_1259);
nor U2005 (N_2005,N_1243,N_764);
or U2006 (N_2006,N_1060,N_1351);
and U2007 (N_2007,N_1315,N_1323);
or U2008 (N_2008,N_997,N_931);
nor U2009 (N_2009,N_1264,N_1162);
or U2010 (N_2010,N_782,N_783);
xnor U2011 (N_2011,N_1294,N_1407);
nor U2012 (N_2012,N_1405,N_1463);
or U2013 (N_2013,N_1288,N_1209);
nand U2014 (N_2014,N_861,N_759);
and U2015 (N_2015,N_875,N_1004);
and U2016 (N_2016,N_1315,N_1101);
or U2017 (N_2017,N_1324,N_815);
and U2018 (N_2018,N_1204,N_1069);
nand U2019 (N_2019,N_757,N_1356);
xnor U2020 (N_2020,N_1288,N_824);
and U2021 (N_2021,N_1154,N_1186);
nor U2022 (N_2022,N_1430,N_1180);
xnor U2023 (N_2023,N_1206,N_1463);
xor U2024 (N_2024,N_1097,N_1098);
nor U2025 (N_2025,N_1152,N_1242);
nand U2026 (N_2026,N_1149,N_1325);
and U2027 (N_2027,N_914,N_1198);
xnor U2028 (N_2028,N_1376,N_1407);
xor U2029 (N_2029,N_1052,N_1201);
nand U2030 (N_2030,N_1475,N_1498);
nor U2031 (N_2031,N_929,N_1423);
nand U2032 (N_2032,N_797,N_1480);
nand U2033 (N_2033,N_790,N_761);
nand U2034 (N_2034,N_1219,N_1280);
nand U2035 (N_2035,N_1222,N_984);
nor U2036 (N_2036,N_824,N_804);
nand U2037 (N_2037,N_1377,N_1334);
nor U2038 (N_2038,N_1476,N_857);
and U2039 (N_2039,N_1088,N_1300);
and U2040 (N_2040,N_1496,N_872);
nor U2041 (N_2041,N_1305,N_1106);
and U2042 (N_2042,N_1033,N_856);
nand U2043 (N_2043,N_1244,N_1211);
and U2044 (N_2044,N_1417,N_972);
and U2045 (N_2045,N_1092,N_1393);
and U2046 (N_2046,N_753,N_863);
nand U2047 (N_2047,N_1483,N_859);
xor U2048 (N_2048,N_1050,N_1393);
and U2049 (N_2049,N_1179,N_1083);
xnor U2050 (N_2050,N_1151,N_1327);
nand U2051 (N_2051,N_952,N_1322);
or U2052 (N_2052,N_1320,N_937);
nor U2053 (N_2053,N_1090,N_1220);
or U2054 (N_2054,N_900,N_1414);
nor U2055 (N_2055,N_1356,N_1220);
xor U2056 (N_2056,N_1122,N_779);
or U2057 (N_2057,N_1160,N_1431);
and U2058 (N_2058,N_1372,N_1179);
or U2059 (N_2059,N_1241,N_1278);
or U2060 (N_2060,N_1489,N_1194);
or U2061 (N_2061,N_1446,N_910);
xor U2062 (N_2062,N_1240,N_959);
and U2063 (N_2063,N_1455,N_942);
nand U2064 (N_2064,N_1367,N_1156);
or U2065 (N_2065,N_1134,N_1445);
nand U2066 (N_2066,N_1028,N_1270);
nor U2067 (N_2067,N_1218,N_1338);
nor U2068 (N_2068,N_859,N_1176);
and U2069 (N_2069,N_1140,N_1467);
nor U2070 (N_2070,N_820,N_1225);
xnor U2071 (N_2071,N_987,N_1102);
and U2072 (N_2072,N_850,N_780);
nor U2073 (N_2073,N_1022,N_1271);
xor U2074 (N_2074,N_1186,N_1036);
xnor U2075 (N_2075,N_853,N_753);
xnor U2076 (N_2076,N_1243,N_1251);
xnor U2077 (N_2077,N_1442,N_1385);
nand U2078 (N_2078,N_926,N_1137);
nor U2079 (N_2079,N_1473,N_892);
nand U2080 (N_2080,N_1367,N_1494);
xor U2081 (N_2081,N_873,N_974);
nor U2082 (N_2082,N_756,N_1325);
xor U2083 (N_2083,N_1341,N_1303);
nand U2084 (N_2084,N_1434,N_979);
nor U2085 (N_2085,N_1196,N_951);
and U2086 (N_2086,N_934,N_1128);
nand U2087 (N_2087,N_765,N_1445);
nor U2088 (N_2088,N_1473,N_999);
nor U2089 (N_2089,N_858,N_1385);
and U2090 (N_2090,N_783,N_1231);
nand U2091 (N_2091,N_1196,N_1224);
and U2092 (N_2092,N_974,N_1406);
nor U2093 (N_2093,N_1265,N_1467);
or U2094 (N_2094,N_1396,N_1311);
or U2095 (N_2095,N_1320,N_1170);
and U2096 (N_2096,N_788,N_1010);
and U2097 (N_2097,N_1092,N_990);
and U2098 (N_2098,N_761,N_1374);
nor U2099 (N_2099,N_910,N_1229);
and U2100 (N_2100,N_993,N_1048);
or U2101 (N_2101,N_1423,N_916);
nor U2102 (N_2102,N_779,N_1038);
nor U2103 (N_2103,N_1078,N_826);
and U2104 (N_2104,N_1225,N_1446);
xnor U2105 (N_2105,N_1412,N_1313);
or U2106 (N_2106,N_814,N_1176);
xnor U2107 (N_2107,N_1410,N_1389);
nand U2108 (N_2108,N_1196,N_878);
or U2109 (N_2109,N_1211,N_1280);
and U2110 (N_2110,N_794,N_1340);
or U2111 (N_2111,N_1251,N_1265);
and U2112 (N_2112,N_1195,N_1158);
xnor U2113 (N_2113,N_1318,N_907);
and U2114 (N_2114,N_1409,N_1007);
or U2115 (N_2115,N_751,N_832);
and U2116 (N_2116,N_1179,N_1440);
nor U2117 (N_2117,N_1097,N_1245);
xor U2118 (N_2118,N_916,N_1468);
xnor U2119 (N_2119,N_1408,N_1428);
or U2120 (N_2120,N_1295,N_1415);
and U2121 (N_2121,N_1396,N_1044);
xnor U2122 (N_2122,N_1438,N_1295);
nor U2123 (N_2123,N_1049,N_1489);
nor U2124 (N_2124,N_1194,N_967);
xnor U2125 (N_2125,N_1293,N_841);
nor U2126 (N_2126,N_1062,N_853);
xnor U2127 (N_2127,N_1045,N_798);
xnor U2128 (N_2128,N_1417,N_957);
and U2129 (N_2129,N_983,N_810);
nor U2130 (N_2130,N_983,N_835);
and U2131 (N_2131,N_808,N_770);
or U2132 (N_2132,N_822,N_1336);
nand U2133 (N_2133,N_1175,N_1418);
nor U2134 (N_2134,N_1367,N_1082);
or U2135 (N_2135,N_1098,N_1182);
and U2136 (N_2136,N_1345,N_1248);
and U2137 (N_2137,N_762,N_1469);
or U2138 (N_2138,N_1251,N_1220);
or U2139 (N_2139,N_963,N_948);
nor U2140 (N_2140,N_1363,N_1165);
nand U2141 (N_2141,N_1082,N_796);
nor U2142 (N_2142,N_879,N_917);
xor U2143 (N_2143,N_836,N_1468);
nand U2144 (N_2144,N_1434,N_1199);
or U2145 (N_2145,N_1301,N_1069);
nor U2146 (N_2146,N_1241,N_1058);
xor U2147 (N_2147,N_1090,N_803);
nor U2148 (N_2148,N_831,N_829);
nor U2149 (N_2149,N_1139,N_792);
or U2150 (N_2150,N_818,N_1138);
and U2151 (N_2151,N_1074,N_1135);
nand U2152 (N_2152,N_1273,N_1290);
nor U2153 (N_2153,N_1427,N_892);
and U2154 (N_2154,N_1012,N_1193);
and U2155 (N_2155,N_1097,N_1290);
nor U2156 (N_2156,N_1299,N_951);
xnor U2157 (N_2157,N_947,N_1005);
nand U2158 (N_2158,N_1403,N_1192);
xor U2159 (N_2159,N_884,N_1282);
xor U2160 (N_2160,N_1311,N_1439);
nor U2161 (N_2161,N_1482,N_1090);
xnor U2162 (N_2162,N_1262,N_751);
nand U2163 (N_2163,N_1004,N_1311);
nand U2164 (N_2164,N_906,N_884);
nor U2165 (N_2165,N_985,N_1377);
nand U2166 (N_2166,N_1124,N_1095);
xnor U2167 (N_2167,N_951,N_1202);
xnor U2168 (N_2168,N_873,N_1040);
nor U2169 (N_2169,N_1014,N_1486);
nor U2170 (N_2170,N_1009,N_1285);
or U2171 (N_2171,N_940,N_1470);
and U2172 (N_2172,N_1320,N_1190);
xor U2173 (N_2173,N_752,N_1292);
nor U2174 (N_2174,N_762,N_1308);
and U2175 (N_2175,N_935,N_773);
nand U2176 (N_2176,N_1054,N_1151);
nand U2177 (N_2177,N_780,N_1438);
or U2178 (N_2178,N_1126,N_1327);
nand U2179 (N_2179,N_1045,N_822);
nor U2180 (N_2180,N_1217,N_1330);
xnor U2181 (N_2181,N_1269,N_1321);
xnor U2182 (N_2182,N_911,N_763);
xnor U2183 (N_2183,N_1278,N_927);
nand U2184 (N_2184,N_1131,N_773);
nand U2185 (N_2185,N_885,N_983);
xor U2186 (N_2186,N_1253,N_1224);
or U2187 (N_2187,N_1205,N_1321);
or U2188 (N_2188,N_933,N_981);
nand U2189 (N_2189,N_776,N_1067);
nand U2190 (N_2190,N_1099,N_1424);
or U2191 (N_2191,N_1411,N_966);
and U2192 (N_2192,N_1231,N_1447);
xor U2193 (N_2193,N_887,N_797);
xnor U2194 (N_2194,N_1317,N_956);
xnor U2195 (N_2195,N_872,N_1378);
xnor U2196 (N_2196,N_1029,N_1415);
or U2197 (N_2197,N_1008,N_1351);
or U2198 (N_2198,N_1200,N_1063);
and U2199 (N_2199,N_1287,N_830);
xnor U2200 (N_2200,N_926,N_1481);
or U2201 (N_2201,N_1190,N_1084);
nand U2202 (N_2202,N_1000,N_1448);
and U2203 (N_2203,N_1409,N_1142);
nor U2204 (N_2204,N_816,N_929);
nand U2205 (N_2205,N_1136,N_794);
nor U2206 (N_2206,N_817,N_1149);
nand U2207 (N_2207,N_1205,N_1326);
nor U2208 (N_2208,N_1348,N_1051);
xor U2209 (N_2209,N_1202,N_771);
nor U2210 (N_2210,N_1028,N_1292);
and U2211 (N_2211,N_1221,N_1152);
and U2212 (N_2212,N_1151,N_1101);
or U2213 (N_2213,N_814,N_922);
nand U2214 (N_2214,N_996,N_1427);
xor U2215 (N_2215,N_1396,N_1336);
xor U2216 (N_2216,N_1031,N_1440);
and U2217 (N_2217,N_1064,N_840);
and U2218 (N_2218,N_1300,N_1217);
and U2219 (N_2219,N_1005,N_803);
nand U2220 (N_2220,N_1343,N_958);
nand U2221 (N_2221,N_1245,N_1459);
nor U2222 (N_2222,N_1162,N_1422);
nand U2223 (N_2223,N_1323,N_875);
nand U2224 (N_2224,N_1349,N_1237);
and U2225 (N_2225,N_994,N_1214);
and U2226 (N_2226,N_1118,N_820);
nand U2227 (N_2227,N_1232,N_998);
and U2228 (N_2228,N_751,N_1140);
xor U2229 (N_2229,N_1441,N_1398);
and U2230 (N_2230,N_1461,N_884);
or U2231 (N_2231,N_913,N_1433);
or U2232 (N_2232,N_1299,N_1079);
and U2233 (N_2233,N_1201,N_1335);
nor U2234 (N_2234,N_1304,N_1157);
nor U2235 (N_2235,N_1352,N_763);
nand U2236 (N_2236,N_1393,N_1483);
or U2237 (N_2237,N_1485,N_1226);
nor U2238 (N_2238,N_1349,N_1180);
and U2239 (N_2239,N_1404,N_1255);
nor U2240 (N_2240,N_1192,N_1035);
and U2241 (N_2241,N_1156,N_759);
and U2242 (N_2242,N_1320,N_1303);
nor U2243 (N_2243,N_1324,N_1289);
nand U2244 (N_2244,N_873,N_935);
nor U2245 (N_2245,N_1324,N_1016);
xnor U2246 (N_2246,N_1407,N_1161);
or U2247 (N_2247,N_1232,N_1411);
nor U2248 (N_2248,N_906,N_946);
nand U2249 (N_2249,N_1488,N_908);
or U2250 (N_2250,N_2069,N_2240);
nand U2251 (N_2251,N_1954,N_2208);
xor U2252 (N_2252,N_1836,N_2138);
xor U2253 (N_2253,N_1701,N_2155);
and U2254 (N_2254,N_1830,N_1748);
nor U2255 (N_2255,N_2246,N_1851);
xor U2256 (N_2256,N_1734,N_1964);
and U2257 (N_2257,N_1772,N_1525);
nand U2258 (N_2258,N_1846,N_1580);
and U2259 (N_2259,N_1704,N_1604);
xor U2260 (N_2260,N_1583,N_1940);
xnor U2261 (N_2261,N_2065,N_1688);
xor U2262 (N_2262,N_1803,N_1901);
nor U2263 (N_2263,N_1922,N_1596);
nor U2264 (N_2264,N_2095,N_2093);
xor U2265 (N_2265,N_1721,N_1700);
xnor U2266 (N_2266,N_1632,N_2144);
and U2267 (N_2267,N_2014,N_2153);
nor U2268 (N_2268,N_1880,N_1729);
or U2269 (N_2269,N_1902,N_1832);
nor U2270 (N_2270,N_2146,N_1656);
nor U2271 (N_2271,N_1741,N_1963);
or U2272 (N_2272,N_1614,N_1816);
nand U2273 (N_2273,N_2171,N_1641);
and U2274 (N_2274,N_1731,N_2131);
nor U2275 (N_2275,N_1548,N_2159);
or U2276 (N_2276,N_1989,N_2060);
nor U2277 (N_2277,N_1648,N_1707);
nor U2278 (N_2278,N_2202,N_1978);
xor U2279 (N_2279,N_1988,N_1626);
and U2280 (N_2280,N_1782,N_1802);
nor U2281 (N_2281,N_2126,N_1679);
or U2282 (N_2282,N_2086,N_2218);
and U2283 (N_2283,N_1603,N_2206);
nor U2284 (N_2284,N_1853,N_1594);
xor U2285 (N_2285,N_1588,N_1864);
xnor U2286 (N_2286,N_2191,N_2213);
nor U2287 (N_2287,N_1541,N_1736);
or U2288 (N_2288,N_1900,N_2006);
xor U2289 (N_2289,N_2104,N_2166);
or U2290 (N_2290,N_1983,N_2228);
or U2291 (N_2291,N_2168,N_2132);
nor U2292 (N_2292,N_1818,N_1638);
and U2293 (N_2293,N_2128,N_1757);
and U2294 (N_2294,N_1821,N_2230);
and U2295 (N_2295,N_1814,N_1623);
or U2296 (N_2296,N_1998,N_1810);
or U2297 (N_2297,N_2081,N_1589);
xor U2298 (N_2298,N_1709,N_1886);
or U2299 (N_2299,N_1778,N_1920);
and U2300 (N_2300,N_1654,N_1724);
and U2301 (N_2301,N_1783,N_2140);
xor U2302 (N_2302,N_1697,N_1575);
nor U2303 (N_2303,N_2116,N_2048);
nand U2304 (N_2304,N_2204,N_1765);
or U2305 (N_2305,N_1667,N_1610);
nor U2306 (N_2306,N_1970,N_1934);
nand U2307 (N_2307,N_2067,N_1912);
nand U2308 (N_2308,N_1758,N_1696);
and U2309 (N_2309,N_2198,N_1711);
xor U2310 (N_2310,N_1767,N_1618);
and U2311 (N_2311,N_1677,N_1749);
nor U2312 (N_2312,N_1935,N_1595);
xor U2313 (N_2313,N_1825,N_1811);
xor U2314 (N_2314,N_1761,N_1671);
or U2315 (N_2315,N_2013,N_1508);
xor U2316 (N_2316,N_1943,N_2039);
xor U2317 (N_2317,N_1552,N_2125);
and U2318 (N_2318,N_2192,N_1511);
or U2319 (N_2319,N_1518,N_1655);
nor U2320 (N_2320,N_1725,N_1553);
xor U2321 (N_2321,N_1564,N_2111);
nand U2322 (N_2322,N_2018,N_1567);
nor U2323 (N_2323,N_1965,N_1652);
or U2324 (N_2324,N_2053,N_1666);
and U2325 (N_2325,N_1766,N_1789);
and U2326 (N_2326,N_2118,N_2187);
nand U2327 (N_2327,N_1530,N_2100);
xnor U2328 (N_2328,N_2249,N_2112);
or U2329 (N_2329,N_1670,N_1608);
or U2330 (N_2330,N_1539,N_1826);
xnor U2331 (N_2331,N_1545,N_2079);
nand U2332 (N_2332,N_2143,N_1873);
nor U2333 (N_2333,N_1947,N_1999);
or U2334 (N_2334,N_2108,N_2003);
nand U2335 (N_2335,N_1703,N_2227);
xor U2336 (N_2336,N_1537,N_1764);
and U2337 (N_2337,N_2139,N_1733);
or U2338 (N_2338,N_1584,N_1566);
and U2339 (N_2339,N_1885,N_1571);
or U2340 (N_2340,N_1513,N_1891);
or U2341 (N_2341,N_1787,N_1946);
nor U2342 (N_2342,N_2148,N_2169);
nor U2343 (N_2343,N_1865,N_2123);
xor U2344 (N_2344,N_1684,N_2222);
and U2345 (N_2345,N_1611,N_1939);
nor U2346 (N_2346,N_2034,N_1848);
and U2347 (N_2347,N_1805,N_1624);
or U2348 (N_2348,N_2154,N_1505);
and U2349 (N_2349,N_1630,N_1898);
nor U2350 (N_2350,N_1834,N_1637);
nor U2351 (N_2351,N_1607,N_2219);
or U2352 (N_2352,N_2133,N_2084);
nand U2353 (N_2353,N_2130,N_1977);
xor U2354 (N_2354,N_1658,N_1650);
or U2355 (N_2355,N_1907,N_1953);
xor U2356 (N_2356,N_1689,N_1519);
and U2357 (N_2357,N_1890,N_1936);
xnor U2358 (N_2358,N_1823,N_1516);
or U2359 (N_2359,N_1585,N_1639);
and U2360 (N_2360,N_1502,N_1923);
and U2361 (N_2361,N_1872,N_1510);
nand U2362 (N_2362,N_2186,N_2041);
nand U2363 (N_2363,N_2064,N_1629);
or U2364 (N_2364,N_1841,N_1822);
nor U2365 (N_2365,N_1877,N_1889);
nand U2366 (N_2366,N_2244,N_1905);
nor U2367 (N_2367,N_1888,N_1617);
and U2368 (N_2368,N_2174,N_1961);
xnor U2369 (N_2369,N_1957,N_1723);
nor U2370 (N_2370,N_1599,N_1887);
or U2371 (N_2371,N_2181,N_1913);
or U2372 (N_2372,N_1556,N_2045);
or U2373 (N_2373,N_2021,N_1842);
nand U2374 (N_2374,N_1839,N_2040);
nor U2375 (N_2375,N_2110,N_1625);
nand U2376 (N_2376,N_1949,N_1928);
and U2377 (N_2377,N_1561,N_1906);
nand U2378 (N_2378,N_2050,N_2190);
xnor U2379 (N_2379,N_1966,N_1806);
and U2380 (N_2380,N_1560,N_2054);
or U2381 (N_2381,N_1793,N_2152);
nor U2382 (N_2382,N_2070,N_1535);
or U2383 (N_2383,N_1770,N_1859);
nand U2384 (N_2384,N_2059,N_2151);
nand U2385 (N_2385,N_2092,N_2073);
xor U2386 (N_2386,N_1874,N_2077);
nor U2387 (N_2387,N_1693,N_1742);
nor U2388 (N_2388,N_1959,N_1929);
nand U2389 (N_2389,N_1911,N_2197);
xnor U2390 (N_2390,N_1531,N_1676);
and U2391 (N_2391,N_2231,N_2033);
and U2392 (N_2392,N_1815,N_1615);
nor U2393 (N_2393,N_2245,N_2184);
or U2394 (N_2394,N_2141,N_1634);
nand U2395 (N_2395,N_1692,N_1753);
or U2396 (N_2396,N_1549,N_1601);
and U2397 (N_2397,N_1645,N_1820);
xnor U2398 (N_2398,N_1523,N_1570);
nand U2399 (N_2399,N_1771,N_1643);
xor U2400 (N_2400,N_2164,N_2150);
nor U2401 (N_2401,N_1948,N_1909);
nand U2402 (N_2402,N_2234,N_1892);
nand U2403 (N_2403,N_1587,N_1665);
or U2404 (N_2404,N_1554,N_2149);
nand U2405 (N_2405,N_1745,N_1675);
xor U2406 (N_2406,N_1555,N_1717);
and U2407 (N_2407,N_2000,N_2221);
or U2408 (N_2408,N_1956,N_1857);
nand U2409 (N_2409,N_1660,N_1792);
nor U2410 (N_2410,N_1609,N_1651);
xor U2411 (N_2411,N_2176,N_1706);
nor U2412 (N_2412,N_1718,N_1780);
nor U2413 (N_2413,N_2012,N_1582);
xnor U2414 (N_2414,N_1878,N_1881);
and U2415 (N_2415,N_1534,N_2109);
and U2416 (N_2416,N_1992,N_2010);
nand U2417 (N_2417,N_1845,N_1715);
and U2418 (N_2418,N_1691,N_2119);
and U2419 (N_2419,N_1997,N_1526);
nor U2420 (N_2420,N_1524,N_1850);
nor U2421 (N_2421,N_1600,N_1543);
nand U2422 (N_2422,N_1790,N_1503);
nor U2423 (N_2423,N_1875,N_2072);
nand U2424 (N_2424,N_2124,N_1659);
and U2425 (N_2425,N_1747,N_2101);
nor U2426 (N_2426,N_1819,N_1685);
xor U2427 (N_2427,N_1572,N_1722);
or U2428 (N_2428,N_1663,N_2165);
nand U2429 (N_2429,N_1507,N_2099);
xor U2430 (N_2430,N_1960,N_1969);
or U2431 (N_2431,N_1788,N_2002);
nor U2432 (N_2432,N_1708,N_2063);
nand U2433 (N_2433,N_1581,N_2005);
or U2434 (N_2434,N_1628,N_1786);
and U2435 (N_2435,N_1972,N_2019);
nor U2436 (N_2436,N_2178,N_1574);
and U2437 (N_2437,N_1833,N_1680);
nor U2438 (N_2438,N_2177,N_1759);
and U2439 (N_2439,N_2106,N_2029);
xor U2440 (N_2440,N_2170,N_1515);
xnor U2441 (N_2441,N_1514,N_1699);
xnor U2442 (N_2442,N_1807,N_1904);
nor U2443 (N_2443,N_2032,N_2097);
xor U2444 (N_2444,N_1565,N_2031);
and U2445 (N_2445,N_1784,N_2238);
and U2446 (N_2446,N_1678,N_1591);
and U2447 (N_2447,N_1797,N_1991);
and U2448 (N_2448,N_1592,N_1569);
xor U2449 (N_2449,N_1835,N_1698);
nand U2450 (N_2450,N_1727,N_1536);
and U2451 (N_2451,N_1871,N_2121);
nand U2452 (N_2452,N_2022,N_1687);
and U2453 (N_2453,N_1795,N_1751);
nand U2454 (N_2454,N_1995,N_1924);
nand U2455 (N_2455,N_2188,N_2136);
nand U2456 (N_2456,N_1750,N_2102);
xor U2457 (N_2457,N_1631,N_2237);
and U2458 (N_2458,N_2026,N_1719);
xnor U2459 (N_2459,N_2137,N_1903);
or U2460 (N_2460,N_2062,N_1915);
xor U2461 (N_2461,N_2017,N_1527);
xor U2462 (N_2462,N_2113,N_2057);
xnor U2463 (N_2463,N_2117,N_2223);
xor U2464 (N_2464,N_1635,N_2247);
and U2465 (N_2465,N_2134,N_2142);
nor U2466 (N_2466,N_2157,N_1577);
or U2467 (N_2467,N_1776,N_2196);
xor U2468 (N_2468,N_2229,N_1775);
or U2469 (N_2469,N_2158,N_1768);
or U2470 (N_2470,N_2078,N_2211);
nand U2471 (N_2471,N_2199,N_1602);
xor U2472 (N_2472,N_1763,N_1504);
nor U2473 (N_2473,N_2147,N_1895);
or U2474 (N_2474,N_1796,N_2056);
nor U2475 (N_2475,N_2127,N_1683);
nor U2476 (N_2476,N_2129,N_1984);
or U2477 (N_2477,N_1674,N_1740);
xnor U2478 (N_2478,N_1612,N_1506);
and U2479 (N_2479,N_1967,N_1798);
nor U2480 (N_2480,N_1551,N_1883);
or U2481 (N_2481,N_1528,N_2200);
or U2482 (N_2482,N_1546,N_2207);
nand U2483 (N_2483,N_1686,N_1661);
and U2484 (N_2484,N_1840,N_1868);
xor U2485 (N_2485,N_1668,N_1996);
xor U2486 (N_2486,N_1973,N_1917);
nor U2487 (N_2487,N_2089,N_1653);
xor U2488 (N_2488,N_1829,N_2183);
xnor U2489 (N_2489,N_1843,N_1705);
or U2490 (N_2490,N_1993,N_1662);
or U2491 (N_2491,N_1925,N_1938);
xor U2492 (N_2492,N_1897,N_2226);
or U2493 (N_2493,N_1914,N_1756);
or U2494 (N_2494,N_1918,N_2043);
and U2495 (N_2495,N_1644,N_2074);
nand U2496 (N_2496,N_1713,N_1896);
xnor U2497 (N_2497,N_1509,N_2058);
xor U2498 (N_2498,N_1616,N_1562);
and U2499 (N_2499,N_1739,N_1694);
nand U2500 (N_2500,N_1547,N_1952);
nand U2501 (N_2501,N_2044,N_2114);
and U2502 (N_2502,N_1971,N_1559);
xor U2503 (N_2503,N_1737,N_1590);
and U2504 (N_2504,N_1844,N_1870);
and U2505 (N_2505,N_1861,N_2224);
xor U2506 (N_2506,N_2135,N_2236);
or U2507 (N_2507,N_1542,N_2161);
nor U2508 (N_2508,N_2076,N_1712);
and U2509 (N_2509,N_2009,N_1933);
and U2510 (N_2510,N_2087,N_1578);
nor U2511 (N_2511,N_1919,N_1894);
nand U2512 (N_2512,N_2212,N_1828);
nand U2513 (N_2513,N_1837,N_1944);
and U2514 (N_2514,N_1801,N_2215);
nand U2515 (N_2515,N_1974,N_2047);
nor U2516 (N_2516,N_2001,N_1831);
xor U2517 (N_2517,N_1808,N_2046);
and U2518 (N_2518,N_2209,N_2172);
and U2519 (N_2519,N_1867,N_1517);
and U2520 (N_2520,N_1852,N_1576);
and U2521 (N_2521,N_1520,N_2080);
nand U2522 (N_2522,N_1994,N_2233);
xor U2523 (N_2523,N_1533,N_1827);
or U2524 (N_2524,N_1744,N_1926);
nor U2525 (N_2525,N_1856,N_1858);
or U2526 (N_2526,N_2105,N_1538);
or U2527 (N_2527,N_2232,N_2241);
and U2528 (N_2528,N_1695,N_2094);
xor U2529 (N_2529,N_1951,N_2028);
nor U2530 (N_2530,N_1664,N_2225);
or U2531 (N_2531,N_1968,N_1647);
nand U2532 (N_2532,N_1855,N_1521);
or U2533 (N_2533,N_2201,N_2055);
nand U2534 (N_2534,N_2107,N_1550);
nand U2535 (N_2535,N_1910,N_2007);
xor U2536 (N_2536,N_1681,N_1669);
xnor U2537 (N_2537,N_1942,N_1762);
nand U2538 (N_2538,N_2160,N_2096);
nor U2539 (N_2539,N_1975,N_1893);
nor U2540 (N_2540,N_1899,N_2122);
nand U2541 (N_2541,N_1673,N_1755);
nor U2542 (N_2542,N_1779,N_1573);
and U2543 (N_2543,N_1710,N_1781);
and U2544 (N_2544,N_1813,N_2035);
nor U2545 (N_2545,N_2194,N_1791);
or U2546 (N_2546,N_1649,N_2205);
or U2547 (N_2547,N_1838,N_1500);
nand U2548 (N_2548,N_1950,N_1847);
xnor U2549 (N_2549,N_1882,N_1908);
nand U2550 (N_2550,N_2023,N_1743);
nand U2551 (N_2551,N_2243,N_1849);
or U2552 (N_2552,N_2030,N_1812);
nand U2553 (N_2553,N_1622,N_1777);
and U2554 (N_2554,N_2248,N_1785);
xnor U2555 (N_2555,N_1854,N_1800);
xnor U2556 (N_2556,N_1937,N_1876);
nand U2557 (N_2557,N_2085,N_2068);
nor U2558 (N_2558,N_2195,N_1540);
xnor U2559 (N_2559,N_1532,N_1985);
nor U2560 (N_2560,N_1732,N_1979);
nand U2561 (N_2561,N_2027,N_2162);
xor U2562 (N_2562,N_1804,N_1672);
nor U2563 (N_2563,N_1636,N_1916);
nor U2564 (N_2564,N_1930,N_1501);
and U2565 (N_2565,N_2015,N_1774);
nand U2566 (N_2566,N_1931,N_2011);
xor U2567 (N_2567,N_2091,N_1606);
nand U2568 (N_2568,N_1529,N_2051);
and U2569 (N_2569,N_1642,N_2180);
nor U2570 (N_2570,N_1613,N_2179);
nand U2571 (N_2571,N_1932,N_1769);
xnor U2572 (N_2572,N_1728,N_1976);
nor U2573 (N_2573,N_1633,N_2061);
xnor U2574 (N_2574,N_2115,N_1927);
nand U2575 (N_2575,N_1760,N_1619);
xor U2576 (N_2576,N_1863,N_2193);
nor U2577 (N_2577,N_2004,N_2016);
nand U2578 (N_2578,N_1726,N_1557);
nand U2579 (N_2579,N_1640,N_1958);
and U2580 (N_2580,N_2025,N_1605);
and U2581 (N_2581,N_1884,N_2052);
or U2582 (N_2582,N_1980,N_1646);
nand U2583 (N_2583,N_1579,N_1752);
or U2584 (N_2584,N_1702,N_1568);
or U2585 (N_2585,N_1512,N_1738);
or U2586 (N_2586,N_2075,N_1522);
nor U2587 (N_2587,N_1773,N_1598);
xor U2588 (N_2588,N_1730,N_2173);
xnor U2589 (N_2589,N_2156,N_1714);
and U2590 (N_2590,N_2083,N_1955);
nor U2591 (N_2591,N_2239,N_1860);
xor U2592 (N_2592,N_1817,N_2082);
or U2593 (N_2593,N_1593,N_2098);
nand U2594 (N_2594,N_2042,N_2037);
or U2595 (N_2595,N_2210,N_1990);
nand U2596 (N_2596,N_2182,N_2024);
nand U2597 (N_2597,N_1558,N_2020);
and U2598 (N_2598,N_2145,N_1690);
or U2599 (N_2599,N_2036,N_1986);
or U2600 (N_2600,N_1981,N_1735);
nand U2601 (N_2601,N_2203,N_2167);
and U2602 (N_2602,N_1862,N_2088);
xor U2603 (N_2603,N_1824,N_2090);
nor U2604 (N_2604,N_2216,N_1746);
or U2605 (N_2605,N_1544,N_2189);
xnor U2606 (N_2606,N_1866,N_1962);
nand U2607 (N_2607,N_2214,N_2217);
and U2608 (N_2608,N_1799,N_2220);
or U2609 (N_2609,N_1945,N_2242);
xor U2610 (N_2610,N_2103,N_2175);
xor U2611 (N_2611,N_1720,N_2185);
xor U2612 (N_2612,N_1921,N_2071);
xor U2613 (N_2613,N_2008,N_1879);
and U2614 (N_2614,N_1597,N_1563);
xnor U2615 (N_2615,N_1620,N_2163);
and U2616 (N_2616,N_1586,N_1657);
or U2617 (N_2617,N_2235,N_1941);
xnor U2618 (N_2618,N_2049,N_2038);
nor U2619 (N_2619,N_2120,N_1809);
or U2620 (N_2620,N_1987,N_1869);
nand U2621 (N_2621,N_1627,N_1754);
nor U2622 (N_2622,N_1716,N_1682);
nor U2623 (N_2623,N_1621,N_2066);
and U2624 (N_2624,N_1794,N_1982);
or U2625 (N_2625,N_2229,N_1506);
nor U2626 (N_2626,N_1716,N_2246);
and U2627 (N_2627,N_2140,N_1522);
nor U2628 (N_2628,N_2191,N_1712);
xnor U2629 (N_2629,N_1804,N_1951);
nor U2630 (N_2630,N_1803,N_2041);
and U2631 (N_2631,N_1506,N_1865);
nor U2632 (N_2632,N_1728,N_1511);
xor U2633 (N_2633,N_1788,N_2035);
nor U2634 (N_2634,N_1945,N_1794);
or U2635 (N_2635,N_1536,N_1820);
nand U2636 (N_2636,N_1689,N_1930);
nor U2637 (N_2637,N_2232,N_2041);
and U2638 (N_2638,N_2022,N_1912);
xor U2639 (N_2639,N_1511,N_2005);
xnor U2640 (N_2640,N_2200,N_1885);
nand U2641 (N_2641,N_1889,N_2080);
or U2642 (N_2642,N_2149,N_1950);
nor U2643 (N_2643,N_2038,N_1703);
or U2644 (N_2644,N_1908,N_1807);
nand U2645 (N_2645,N_1972,N_2010);
and U2646 (N_2646,N_2205,N_1582);
nor U2647 (N_2647,N_1801,N_2050);
xnor U2648 (N_2648,N_2206,N_1773);
nor U2649 (N_2649,N_1730,N_1929);
nand U2650 (N_2650,N_1761,N_2214);
nor U2651 (N_2651,N_1680,N_1593);
and U2652 (N_2652,N_1831,N_1670);
xor U2653 (N_2653,N_2222,N_1998);
xnor U2654 (N_2654,N_1535,N_1720);
nor U2655 (N_2655,N_1510,N_2240);
xor U2656 (N_2656,N_1755,N_2205);
xnor U2657 (N_2657,N_1764,N_1952);
nor U2658 (N_2658,N_2212,N_1951);
or U2659 (N_2659,N_1545,N_1595);
xnor U2660 (N_2660,N_1778,N_1521);
nand U2661 (N_2661,N_2175,N_2207);
and U2662 (N_2662,N_1638,N_2156);
nand U2663 (N_2663,N_2020,N_1616);
nor U2664 (N_2664,N_1878,N_1512);
or U2665 (N_2665,N_1825,N_1822);
nor U2666 (N_2666,N_1947,N_1771);
nor U2667 (N_2667,N_1767,N_1681);
xor U2668 (N_2668,N_2166,N_1929);
and U2669 (N_2669,N_1566,N_1916);
nand U2670 (N_2670,N_1538,N_1926);
nand U2671 (N_2671,N_1642,N_2005);
or U2672 (N_2672,N_1752,N_1744);
nand U2673 (N_2673,N_1795,N_2060);
nor U2674 (N_2674,N_1889,N_1653);
nand U2675 (N_2675,N_1775,N_2128);
and U2676 (N_2676,N_2219,N_1727);
and U2677 (N_2677,N_1761,N_1795);
xor U2678 (N_2678,N_1639,N_1511);
xnor U2679 (N_2679,N_2055,N_1840);
nand U2680 (N_2680,N_2149,N_2124);
and U2681 (N_2681,N_2212,N_1532);
nand U2682 (N_2682,N_1794,N_2089);
or U2683 (N_2683,N_1649,N_2144);
xnor U2684 (N_2684,N_1792,N_2095);
or U2685 (N_2685,N_1939,N_1896);
or U2686 (N_2686,N_1898,N_1891);
or U2687 (N_2687,N_1984,N_1500);
xor U2688 (N_2688,N_1530,N_1792);
xnor U2689 (N_2689,N_1530,N_1688);
and U2690 (N_2690,N_1946,N_1961);
and U2691 (N_2691,N_1742,N_1812);
and U2692 (N_2692,N_2164,N_1629);
or U2693 (N_2693,N_1662,N_2195);
nor U2694 (N_2694,N_1892,N_2130);
or U2695 (N_2695,N_1850,N_1805);
or U2696 (N_2696,N_1625,N_1746);
nor U2697 (N_2697,N_1783,N_2063);
and U2698 (N_2698,N_1509,N_2176);
and U2699 (N_2699,N_2056,N_1684);
nand U2700 (N_2700,N_2140,N_1689);
nand U2701 (N_2701,N_1991,N_1681);
nand U2702 (N_2702,N_1593,N_1721);
nor U2703 (N_2703,N_1646,N_1729);
or U2704 (N_2704,N_1631,N_1619);
xnor U2705 (N_2705,N_1992,N_1817);
and U2706 (N_2706,N_2169,N_1973);
and U2707 (N_2707,N_1599,N_1957);
xnor U2708 (N_2708,N_1995,N_1722);
or U2709 (N_2709,N_1789,N_2134);
xor U2710 (N_2710,N_2060,N_1995);
nor U2711 (N_2711,N_2041,N_1527);
nand U2712 (N_2712,N_1617,N_1731);
and U2713 (N_2713,N_1601,N_2051);
nand U2714 (N_2714,N_1905,N_1828);
or U2715 (N_2715,N_1522,N_1783);
nand U2716 (N_2716,N_1943,N_1984);
and U2717 (N_2717,N_2204,N_2234);
xor U2718 (N_2718,N_1616,N_1952);
and U2719 (N_2719,N_1996,N_1717);
and U2720 (N_2720,N_1763,N_2132);
xnor U2721 (N_2721,N_1704,N_1550);
nor U2722 (N_2722,N_1649,N_1752);
nand U2723 (N_2723,N_1947,N_1662);
xor U2724 (N_2724,N_2175,N_2123);
or U2725 (N_2725,N_1965,N_1785);
nor U2726 (N_2726,N_1758,N_2030);
and U2727 (N_2727,N_1584,N_2236);
nand U2728 (N_2728,N_2112,N_2190);
nand U2729 (N_2729,N_1674,N_1924);
xor U2730 (N_2730,N_1525,N_1533);
or U2731 (N_2731,N_1903,N_2191);
and U2732 (N_2732,N_1527,N_1995);
nand U2733 (N_2733,N_1643,N_2113);
xor U2734 (N_2734,N_1519,N_1923);
or U2735 (N_2735,N_1955,N_1854);
xnor U2736 (N_2736,N_2025,N_1584);
xnor U2737 (N_2737,N_1893,N_2072);
nor U2738 (N_2738,N_1901,N_1681);
nor U2739 (N_2739,N_2111,N_1995);
xnor U2740 (N_2740,N_1957,N_1564);
nand U2741 (N_2741,N_1932,N_1779);
and U2742 (N_2742,N_1853,N_2220);
nand U2743 (N_2743,N_1704,N_2160);
nor U2744 (N_2744,N_1882,N_1615);
nand U2745 (N_2745,N_1685,N_1671);
nor U2746 (N_2746,N_1955,N_1613);
or U2747 (N_2747,N_1889,N_1825);
xnor U2748 (N_2748,N_2077,N_2027);
xor U2749 (N_2749,N_2133,N_1708);
or U2750 (N_2750,N_1683,N_2197);
nor U2751 (N_2751,N_2102,N_1800);
or U2752 (N_2752,N_1556,N_1968);
nor U2753 (N_2753,N_2091,N_1845);
or U2754 (N_2754,N_2158,N_2137);
or U2755 (N_2755,N_1978,N_1725);
xor U2756 (N_2756,N_1728,N_1905);
nor U2757 (N_2757,N_2126,N_1683);
or U2758 (N_2758,N_1772,N_2239);
or U2759 (N_2759,N_2191,N_1737);
nor U2760 (N_2760,N_1879,N_1534);
nor U2761 (N_2761,N_1719,N_1728);
nor U2762 (N_2762,N_2167,N_1906);
nor U2763 (N_2763,N_1646,N_1990);
xnor U2764 (N_2764,N_1683,N_1718);
nor U2765 (N_2765,N_1541,N_2174);
xor U2766 (N_2766,N_2109,N_1538);
nor U2767 (N_2767,N_1766,N_1709);
nand U2768 (N_2768,N_2181,N_1629);
and U2769 (N_2769,N_1796,N_1967);
xnor U2770 (N_2770,N_1668,N_1746);
or U2771 (N_2771,N_1774,N_1825);
xor U2772 (N_2772,N_2184,N_1553);
nand U2773 (N_2773,N_2159,N_1828);
or U2774 (N_2774,N_1699,N_1911);
and U2775 (N_2775,N_1724,N_2092);
or U2776 (N_2776,N_2097,N_2100);
xnor U2777 (N_2777,N_1966,N_2235);
or U2778 (N_2778,N_2241,N_1953);
xor U2779 (N_2779,N_2224,N_1956);
nor U2780 (N_2780,N_1516,N_1872);
nor U2781 (N_2781,N_1757,N_1894);
and U2782 (N_2782,N_1537,N_1668);
or U2783 (N_2783,N_2007,N_1664);
xor U2784 (N_2784,N_1630,N_1800);
xnor U2785 (N_2785,N_1791,N_2040);
and U2786 (N_2786,N_2106,N_1581);
nor U2787 (N_2787,N_1726,N_2184);
and U2788 (N_2788,N_1643,N_1917);
nor U2789 (N_2789,N_1507,N_2232);
or U2790 (N_2790,N_2185,N_1672);
nor U2791 (N_2791,N_1661,N_1764);
nand U2792 (N_2792,N_1958,N_1540);
nor U2793 (N_2793,N_1553,N_1694);
nor U2794 (N_2794,N_1942,N_2206);
or U2795 (N_2795,N_2006,N_1611);
nor U2796 (N_2796,N_1907,N_1933);
xnor U2797 (N_2797,N_2027,N_1659);
xor U2798 (N_2798,N_1895,N_1668);
nand U2799 (N_2799,N_2247,N_2015);
xnor U2800 (N_2800,N_1580,N_2078);
nand U2801 (N_2801,N_2137,N_1600);
or U2802 (N_2802,N_2091,N_1578);
and U2803 (N_2803,N_2062,N_1992);
nand U2804 (N_2804,N_1624,N_1695);
or U2805 (N_2805,N_1644,N_1771);
and U2806 (N_2806,N_1590,N_1559);
and U2807 (N_2807,N_1766,N_1934);
nand U2808 (N_2808,N_1586,N_1543);
xnor U2809 (N_2809,N_2042,N_1657);
and U2810 (N_2810,N_2096,N_1825);
xnor U2811 (N_2811,N_2144,N_1682);
xnor U2812 (N_2812,N_2159,N_2197);
nand U2813 (N_2813,N_1829,N_2036);
nand U2814 (N_2814,N_1962,N_1930);
or U2815 (N_2815,N_1852,N_1835);
nor U2816 (N_2816,N_1921,N_1650);
nor U2817 (N_2817,N_1819,N_1673);
nand U2818 (N_2818,N_1663,N_1542);
nor U2819 (N_2819,N_2249,N_2164);
and U2820 (N_2820,N_1779,N_2078);
xor U2821 (N_2821,N_1799,N_2226);
xor U2822 (N_2822,N_1534,N_1703);
nor U2823 (N_2823,N_2155,N_2084);
and U2824 (N_2824,N_1917,N_2057);
nand U2825 (N_2825,N_1988,N_1732);
and U2826 (N_2826,N_2171,N_1669);
and U2827 (N_2827,N_2080,N_2165);
or U2828 (N_2828,N_2117,N_1615);
nor U2829 (N_2829,N_1572,N_1640);
xor U2830 (N_2830,N_2064,N_2091);
nor U2831 (N_2831,N_2169,N_2173);
or U2832 (N_2832,N_1721,N_1930);
nand U2833 (N_2833,N_1515,N_2106);
or U2834 (N_2834,N_2215,N_1905);
and U2835 (N_2835,N_2160,N_1504);
nor U2836 (N_2836,N_2083,N_1784);
or U2837 (N_2837,N_2095,N_1992);
nor U2838 (N_2838,N_2169,N_1946);
and U2839 (N_2839,N_1547,N_1818);
xnor U2840 (N_2840,N_1566,N_1513);
nand U2841 (N_2841,N_1930,N_1590);
nand U2842 (N_2842,N_1564,N_1540);
xor U2843 (N_2843,N_1840,N_2088);
nand U2844 (N_2844,N_1959,N_1594);
and U2845 (N_2845,N_2076,N_1543);
and U2846 (N_2846,N_1631,N_1783);
or U2847 (N_2847,N_2045,N_1956);
or U2848 (N_2848,N_1764,N_2003);
nand U2849 (N_2849,N_2003,N_1584);
xnor U2850 (N_2850,N_1869,N_2011);
xor U2851 (N_2851,N_1860,N_2140);
xnor U2852 (N_2852,N_1962,N_2031);
nor U2853 (N_2853,N_1533,N_2028);
nand U2854 (N_2854,N_2043,N_1793);
nand U2855 (N_2855,N_1923,N_2214);
and U2856 (N_2856,N_2192,N_1685);
and U2857 (N_2857,N_1804,N_1705);
nand U2858 (N_2858,N_1820,N_1947);
and U2859 (N_2859,N_2229,N_1961);
and U2860 (N_2860,N_2123,N_1996);
xnor U2861 (N_2861,N_1542,N_2000);
and U2862 (N_2862,N_1522,N_1887);
and U2863 (N_2863,N_2153,N_2103);
or U2864 (N_2864,N_2040,N_1716);
and U2865 (N_2865,N_1897,N_1772);
nor U2866 (N_2866,N_2064,N_1834);
nor U2867 (N_2867,N_1553,N_1722);
or U2868 (N_2868,N_1501,N_1568);
xor U2869 (N_2869,N_1933,N_2003);
and U2870 (N_2870,N_1695,N_1719);
or U2871 (N_2871,N_2037,N_2229);
and U2872 (N_2872,N_1693,N_1673);
nand U2873 (N_2873,N_1522,N_2174);
xnor U2874 (N_2874,N_1810,N_1624);
xor U2875 (N_2875,N_1712,N_1614);
xor U2876 (N_2876,N_1963,N_1605);
xnor U2877 (N_2877,N_1707,N_1706);
and U2878 (N_2878,N_1788,N_1676);
and U2879 (N_2879,N_1939,N_1622);
or U2880 (N_2880,N_2002,N_1905);
xnor U2881 (N_2881,N_1687,N_1986);
or U2882 (N_2882,N_1732,N_1733);
nor U2883 (N_2883,N_1975,N_1609);
xnor U2884 (N_2884,N_1898,N_1776);
or U2885 (N_2885,N_2240,N_2114);
xor U2886 (N_2886,N_2198,N_1878);
or U2887 (N_2887,N_2082,N_1812);
nand U2888 (N_2888,N_1962,N_1987);
nand U2889 (N_2889,N_1589,N_1542);
xor U2890 (N_2890,N_1743,N_1893);
nand U2891 (N_2891,N_1914,N_1832);
nor U2892 (N_2892,N_2125,N_2029);
xnor U2893 (N_2893,N_1775,N_1957);
nand U2894 (N_2894,N_1713,N_1502);
xor U2895 (N_2895,N_2247,N_1627);
nand U2896 (N_2896,N_1920,N_1566);
xor U2897 (N_2897,N_1997,N_1707);
nand U2898 (N_2898,N_1519,N_2151);
xnor U2899 (N_2899,N_1562,N_1566);
nor U2900 (N_2900,N_1578,N_1978);
nand U2901 (N_2901,N_1836,N_2049);
nand U2902 (N_2902,N_1788,N_1987);
xor U2903 (N_2903,N_1781,N_2002);
and U2904 (N_2904,N_1890,N_1718);
nand U2905 (N_2905,N_1933,N_1677);
xnor U2906 (N_2906,N_1828,N_2142);
nand U2907 (N_2907,N_2061,N_1700);
xnor U2908 (N_2908,N_1907,N_1789);
nor U2909 (N_2909,N_1527,N_1777);
or U2910 (N_2910,N_1681,N_1758);
nand U2911 (N_2911,N_1617,N_1993);
xor U2912 (N_2912,N_1875,N_1938);
nor U2913 (N_2913,N_1675,N_2225);
xor U2914 (N_2914,N_1533,N_1561);
nor U2915 (N_2915,N_1839,N_1673);
and U2916 (N_2916,N_2088,N_1517);
nor U2917 (N_2917,N_2105,N_1982);
and U2918 (N_2918,N_1825,N_2155);
or U2919 (N_2919,N_2133,N_1961);
xnor U2920 (N_2920,N_2226,N_1757);
nand U2921 (N_2921,N_2081,N_1620);
nor U2922 (N_2922,N_2115,N_1793);
xor U2923 (N_2923,N_1758,N_2221);
xor U2924 (N_2924,N_2006,N_1599);
or U2925 (N_2925,N_1915,N_1577);
xor U2926 (N_2926,N_1629,N_2126);
nor U2927 (N_2927,N_1642,N_1807);
nand U2928 (N_2928,N_1876,N_1867);
or U2929 (N_2929,N_1913,N_1702);
xnor U2930 (N_2930,N_1933,N_1777);
nand U2931 (N_2931,N_1876,N_1945);
nand U2932 (N_2932,N_1782,N_1599);
xnor U2933 (N_2933,N_2136,N_1850);
and U2934 (N_2934,N_2059,N_1899);
nor U2935 (N_2935,N_2136,N_2213);
nor U2936 (N_2936,N_1688,N_1559);
nor U2937 (N_2937,N_2173,N_1854);
nor U2938 (N_2938,N_1539,N_2100);
and U2939 (N_2939,N_2204,N_1649);
xor U2940 (N_2940,N_1586,N_1948);
nor U2941 (N_2941,N_2159,N_1559);
xor U2942 (N_2942,N_1828,N_1825);
nand U2943 (N_2943,N_1620,N_1873);
nor U2944 (N_2944,N_1776,N_1789);
and U2945 (N_2945,N_1505,N_1524);
and U2946 (N_2946,N_2187,N_2113);
xnor U2947 (N_2947,N_2150,N_1913);
xor U2948 (N_2948,N_1620,N_1669);
xnor U2949 (N_2949,N_2186,N_1565);
and U2950 (N_2950,N_2068,N_1655);
xor U2951 (N_2951,N_1920,N_2039);
xnor U2952 (N_2952,N_1699,N_1897);
xnor U2953 (N_2953,N_1564,N_1989);
nor U2954 (N_2954,N_1668,N_1634);
nand U2955 (N_2955,N_1650,N_1580);
and U2956 (N_2956,N_2145,N_2124);
xor U2957 (N_2957,N_2170,N_1830);
nor U2958 (N_2958,N_1940,N_2091);
or U2959 (N_2959,N_1524,N_1838);
nor U2960 (N_2960,N_1933,N_1809);
xnor U2961 (N_2961,N_1604,N_2174);
or U2962 (N_2962,N_2054,N_1573);
xnor U2963 (N_2963,N_1605,N_1562);
and U2964 (N_2964,N_1606,N_1852);
nand U2965 (N_2965,N_1860,N_2210);
and U2966 (N_2966,N_2192,N_1740);
nor U2967 (N_2967,N_1751,N_2238);
nand U2968 (N_2968,N_1877,N_1726);
or U2969 (N_2969,N_1930,N_1967);
and U2970 (N_2970,N_2133,N_1548);
nor U2971 (N_2971,N_2038,N_1854);
nand U2972 (N_2972,N_2049,N_1760);
xnor U2973 (N_2973,N_1861,N_1726);
nor U2974 (N_2974,N_1630,N_1759);
nand U2975 (N_2975,N_2173,N_2148);
and U2976 (N_2976,N_1699,N_1641);
nand U2977 (N_2977,N_1801,N_2224);
and U2978 (N_2978,N_2196,N_1843);
nor U2979 (N_2979,N_1843,N_1850);
nand U2980 (N_2980,N_2158,N_2076);
xor U2981 (N_2981,N_2238,N_2244);
or U2982 (N_2982,N_1668,N_2034);
xnor U2983 (N_2983,N_2098,N_1518);
or U2984 (N_2984,N_1970,N_1623);
nand U2985 (N_2985,N_1921,N_2182);
xnor U2986 (N_2986,N_2046,N_2135);
nor U2987 (N_2987,N_1877,N_2147);
or U2988 (N_2988,N_1555,N_2132);
nor U2989 (N_2989,N_1774,N_1648);
xor U2990 (N_2990,N_2206,N_1914);
or U2991 (N_2991,N_2215,N_1744);
xnor U2992 (N_2992,N_1596,N_2180);
nand U2993 (N_2993,N_1576,N_1699);
nand U2994 (N_2994,N_2007,N_1775);
nor U2995 (N_2995,N_1742,N_1559);
nand U2996 (N_2996,N_2038,N_1732);
nand U2997 (N_2997,N_2030,N_1788);
nand U2998 (N_2998,N_1847,N_2205);
or U2999 (N_2999,N_1586,N_2075);
nor UO_0 (O_0,N_2876,N_2888);
nor UO_1 (O_1,N_2405,N_2644);
nor UO_2 (O_2,N_2348,N_2687);
and UO_3 (O_3,N_2514,N_2276);
nand UO_4 (O_4,N_2866,N_2670);
nand UO_5 (O_5,N_2333,N_2338);
xnor UO_6 (O_6,N_2287,N_2800);
nand UO_7 (O_7,N_2836,N_2335);
nand UO_8 (O_8,N_2921,N_2395);
nor UO_9 (O_9,N_2994,N_2343);
nor UO_10 (O_10,N_2812,N_2359);
and UO_11 (O_11,N_2816,N_2599);
xor UO_12 (O_12,N_2721,N_2488);
and UO_13 (O_13,N_2879,N_2317);
and UO_14 (O_14,N_2542,N_2367);
xnor UO_15 (O_15,N_2320,N_2718);
xnor UO_16 (O_16,N_2482,N_2511);
or UO_17 (O_17,N_2944,N_2328);
xnor UO_18 (O_18,N_2749,N_2590);
or UO_19 (O_19,N_2856,N_2517);
nor UO_20 (O_20,N_2289,N_2272);
or UO_21 (O_21,N_2956,N_2733);
xor UO_22 (O_22,N_2336,N_2327);
nor UO_23 (O_23,N_2660,N_2356);
nand UO_24 (O_24,N_2665,N_2398);
and UO_25 (O_25,N_2776,N_2652);
nor UO_26 (O_26,N_2429,N_2406);
or UO_27 (O_27,N_2403,N_2522);
xnor UO_28 (O_28,N_2720,N_2539);
xor UO_29 (O_29,N_2266,N_2691);
and UO_30 (O_30,N_2420,N_2910);
or UO_31 (O_31,N_2834,N_2515);
nand UO_32 (O_32,N_2679,N_2702);
or UO_33 (O_33,N_2917,N_2578);
and UO_34 (O_34,N_2468,N_2388);
nor UO_35 (O_35,N_2843,N_2851);
or UO_36 (O_36,N_2635,N_2678);
xnor UO_37 (O_37,N_2307,N_2825);
nor UO_38 (O_38,N_2999,N_2439);
and UO_39 (O_39,N_2778,N_2970);
and UO_40 (O_40,N_2774,N_2273);
and UO_41 (O_41,N_2625,N_2919);
xnor UO_42 (O_42,N_2380,N_2638);
xnor UO_43 (O_43,N_2714,N_2346);
and UO_44 (O_44,N_2407,N_2996);
or UO_45 (O_45,N_2770,N_2832);
nand UO_46 (O_46,N_2941,N_2586);
and UO_47 (O_47,N_2736,N_2848);
nand UO_48 (O_48,N_2989,N_2427);
nand UO_49 (O_49,N_2805,N_2837);
xor UO_50 (O_50,N_2576,N_2732);
nor UO_51 (O_51,N_2467,N_2309);
xor UO_52 (O_52,N_2797,N_2601);
xnor UO_53 (O_53,N_2557,N_2294);
nor UO_54 (O_54,N_2788,N_2345);
and UO_55 (O_55,N_2389,N_2842);
nand UO_56 (O_56,N_2632,N_2622);
and UO_57 (O_57,N_2486,N_2293);
nand UO_58 (O_58,N_2755,N_2377);
and UO_59 (O_59,N_2803,N_2719);
and UO_60 (O_60,N_2779,N_2822);
or UO_61 (O_61,N_2763,N_2870);
and UO_62 (O_62,N_2920,N_2386);
nand UO_63 (O_63,N_2823,N_2869);
nor UO_64 (O_64,N_2591,N_2344);
nand UO_65 (O_65,N_2551,N_2936);
xor UO_66 (O_66,N_2971,N_2484);
or UO_67 (O_67,N_2260,N_2833);
nand UO_68 (O_68,N_2904,N_2623);
nor UO_69 (O_69,N_2878,N_2559);
nor UO_70 (O_70,N_2606,N_2533);
nand UO_71 (O_71,N_2705,N_2311);
or UO_72 (O_72,N_2525,N_2499);
or UO_73 (O_73,N_2791,N_2914);
nor UO_74 (O_74,N_2594,N_2751);
or UO_75 (O_75,N_2686,N_2497);
and UO_76 (O_76,N_2713,N_2577);
and UO_77 (O_77,N_2628,N_2383);
xnor UO_78 (O_78,N_2663,N_2912);
and UO_79 (O_79,N_2545,N_2364);
nor UO_80 (O_80,N_2980,N_2384);
or UO_81 (O_81,N_2711,N_2505);
nor UO_82 (O_82,N_2761,N_2846);
xnor UO_83 (O_83,N_2664,N_2408);
nor UO_84 (O_84,N_2444,N_2618);
xor UO_85 (O_85,N_2865,N_2790);
nor UO_86 (O_86,N_2454,N_2772);
nand UO_87 (O_87,N_2759,N_2813);
and UO_88 (O_88,N_2633,N_2789);
nor UO_89 (O_89,N_2830,N_2990);
and UO_90 (O_90,N_2821,N_2321);
xor UO_91 (O_91,N_2935,N_2933);
nor UO_92 (O_92,N_2458,N_2529);
xor UO_93 (O_93,N_2826,N_2681);
nor UO_94 (O_94,N_2643,N_2948);
xor UO_95 (O_95,N_2654,N_2569);
nand UO_96 (O_96,N_2758,N_2510);
xor UO_97 (O_97,N_2326,N_2741);
nor UO_98 (O_98,N_2438,N_2563);
nor UO_99 (O_99,N_2891,N_2685);
and UO_100 (O_100,N_2672,N_2564);
xor UO_101 (O_101,N_2674,N_2903);
nor UO_102 (O_102,N_2414,N_2491);
xor UO_103 (O_103,N_2587,N_2949);
xor UO_104 (O_104,N_2259,N_2602);
xnor UO_105 (O_105,N_2548,N_2739);
xor UO_106 (O_106,N_2417,N_2655);
nand UO_107 (O_107,N_2595,N_2441);
nand UO_108 (O_108,N_2967,N_2984);
nor UO_109 (O_109,N_2730,N_2598);
nor UO_110 (O_110,N_2583,N_2490);
xnor UO_111 (O_111,N_2561,N_2331);
nand UO_112 (O_112,N_2735,N_2503);
and UO_113 (O_113,N_2396,N_2554);
nor UO_114 (O_114,N_2820,N_2908);
nand UO_115 (O_115,N_2611,N_2526);
nor UO_116 (O_116,N_2337,N_2962);
or UO_117 (O_117,N_2649,N_2316);
nand UO_118 (O_118,N_2659,N_2430);
nor UO_119 (O_119,N_2859,N_2983);
nand UO_120 (O_120,N_2571,N_2905);
xnor UO_121 (O_121,N_2267,N_2811);
xor UO_122 (O_122,N_2762,N_2462);
nor UO_123 (O_123,N_2552,N_2470);
nor UO_124 (O_124,N_2447,N_2916);
nor UO_125 (O_125,N_2558,N_2712);
and UO_126 (O_126,N_2880,N_2324);
or UO_127 (O_127,N_2974,N_2613);
and UO_128 (O_128,N_2780,N_2899);
nand UO_129 (O_129,N_2262,N_2708);
nand UO_130 (O_130,N_2620,N_2945);
and UO_131 (O_131,N_2371,N_2565);
nor UO_132 (O_132,N_2781,N_2902);
and UO_133 (O_133,N_2802,N_2640);
and UO_134 (O_134,N_2881,N_2656);
and UO_135 (O_135,N_2255,N_2303);
nand UO_136 (O_136,N_2284,N_2305);
or UO_137 (O_137,N_2524,N_2951);
xnor UO_138 (O_138,N_2516,N_2302);
and UO_139 (O_139,N_2955,N_2254);
nand UO_140 (O_140,N_2471,N_2634);
and UO_141 (O_141,N_2639,N_2617);
or UO_142 (O_142,N_2434,N_2319);
xnor UO_143 (O_143,N_2332,N_2753);
or UO_144 (O_144,N_2412,N_2932);
nor UO_145 (O_145,N_2960,N_2306);
or UO_146 (O_146,N_2894,N_2715);
nor UO_147 (O_147,N_2693,N_2804);
xnor UO_148 (O_148,N_2357,N_2862);
or UO_149 (O_149,N_2278,N_2415);
nor UO_150 (O_150,N_2279,N_2815);
and UO_151 (O_151,N_2323,N_2523);
xnor UO_152 (O_152,N_2858,N_2473);
xor UO_153 (O_153,N_2745,N_2647);
and UO_154 (O_154,N_2299,N_2729);
or UO_155 (O_155,N_2442,N_2330);
and UO_156 (O_156,N_2992,N_2263);
xor UO_157 (O_157,N_2728,N_2322);
nand UO_158 (O_158,N_2425,N_2924);
nand UO_159 (O_159,N_2703,N_2373);
xor UO_160 (O_160,N_2394,N_2677);
or UO_161 (O_161,N_2304,N_2694);
xor UO_162 (O_162,N_2937,N_2286);
nor UO_163 (O_163,N_2431,N_2630);
and UO_164 (O_164,N_2401,N_2968);
nand UO_165 (O_165,N_2883,N_2291);
nand UO_166 (O_166,N_2814,N_2661);
xnor UO_167 (O_167,N_2997,N_2926);
nand UO_168 (O_168,N_2740,N_2609);
or UO_169 (O_169,N_2852,N_2795);
or UO_170 (O_170,N_2385,N_2727);
and UO_171 (O_171,N_2621,N_2452);
xnor UO_172 (O_172,N_2958,N_2969);
and UO_173 (O_173,N_2965,N_2280);
and UO_174 (O_174,N_2939,N_2701);
nor UO_175 (O_175,N_2864,N_2954);
nor UO_176 (O_176,N_2459,N_2349);
nand UO_177 (O_177,N_2413,N_2987);
nand UO_178 (O_178,N_2483,N_2596);
xnor UO_179 (O_179,N_2556,N_2301);
nand UO_180 (O_180,N_2637,N_2895);
xor UO_181 (O_181,N_2509,N_2886);
nor UO_182 (O_182,N_2746,N_2614);
nand UO_183 (O_183,N_2250,N_2750);
and UO_184 (O_184,N_2867,N_2629);
nand UO_185 (O_185,N_2979,N_2648);
xnor UO_186 (O_186,N_2872,N_2900);
nor UO_187 (O_187,N_2544,N_2698);
nor UO_188 (O_188,N_2379,N_2453);
or UO_189 (O_189,N_2950,N_2363);
or UO_190 (O_190,N_2756,N_2940);
nor UO_191 (O_191,N_2798,N_2451);
or UO_192 (O_192,N_2873,N_2566);
or UO_193 (O_193,N_2794,N_2251);
and UO_194 (O_194,N_2946,N_2972);
nor UO_195 (O_195,N_2487,N_2771);
and UO_196 (O_196,N_2570,N_2847);
nor UO_197 (O_197,N_2773,N_2799);
and UO_198 (O_198,N_2699,N_2671);
or UO_199 (O_199,N_2722,N_2754);
xor UO_200 (O_200,N_2313,N_2877);
nand UO_201 (O_201,N_2710,N_2424);
nor UO_202 (O_202,N_2976,N_2393);
xor UO_203 (O_203,N_2423,N_2502);
and UO_204 (O_204,N_2476,N_2546);
and UO_205 (O_205,N_2769,N_2519);
xor UO_206 (O_206,N_2675,N_2726);
xor UO_207 (O_207,N_2624,N_2572);
xor UO_208 (O_208,N_2818,N_2456);
nand UO_209 (O_209,N_2582,N_2469);
and UO_210 (O_210,N_2448,N_2314);
and UO_211 (O_211,N_2959,N_2861);
or UO_212 (O_212,N_2562,N_2391);
nor UO_213 (O_213,N_2261,N_2928);
xor UO_214 (O_214,N_2929,N_2603);
nor UO_215 (O_215,N_2450,N_2466);
and UO_216 (O_216,N_2695,N_2810);
nor UO_217 (O_217,N_2964,N_2354);
nor UO_218 (O_218,N_2353,N_2270);
nand UO_219 (O_219,N_2528,N_2288);
and UO_220 (O_220,N_2376,N_2874);
nand UO_221 (O_221,N_2436,N_2352);
or UO_222 (O_222,N_2475,N_2807);
xnor UO_223 (O_223,N_2839,N_2474);
or UO_224 (O_224,N_2890,N_2700);
nand UO_225 (O_225,N_2374,N_2446);
xor UO_226 (O_226,N_2966,N_2930);
or UO_227 (O_227,N_2860,N_2579);
nand UO_228 (O_228,N_2938,N_2692);
or UO_229 (O_229,N_2824,N_2642);
xor UO_230 (O_230,N_2518,N_2428);
and UO_231 (O_231,N_2706,N_2738);
xor UO_232 (O_232,N_2896,N_2600);
and UO_233 (O_233,N_2682,N_2366);
nor UO_234 (O_234,N_2985,N_2308);
xor UO_235 (O_235,N_2724,N_2585);
or UO_236 (O_236,N_2943,N_2485);
nand UO_237 (O_237,N_2257,N_2889);
xnor UO_238 (O_238,N_2381,N_2378);
or UO_239 (O_239,N_2828,N_2597);
xnor UO_240 (O_240,N_2443,N_2775);
nor UO_241 (O_241,N_2295,N_2574);
xnor UO_242 (O_242,N_2478,N_2455);
or UO_243 (O_243,N_2689,N_2553);
or UO_244 (O_244,N_2651,N_2657);
nand UO_245 (O_245,N_2827,N_2748);
nor UO_246 (O_246,N_2666,N_2426);
and UO_247 (O_247,N_2673,N_2290);
and UO_248 (O_248,N_2285,N_2809);
xnor UO_249 (O_249,N_2543,N_2717);
nor UO_250 (O_250,N_2942,N_2785);
nand UO_251 (O_251,N_2680,N_2765);
nor UO_252 (O_252,N_2907,N_2977);
or UO_253 (O_253,N_2885,N_2683);
nor UO_254 (O_254,N_2555,N_2645);
nand UO_255 (O_255,N_2787,N_2350);
xnor UO_256 (O_256,N_2537,N_2991);
nor UO_257 (O_257,N_2339,N_2786);
nor UO_258 (O_258,N_2422,N_2658);
nor UO_259 (O_259,N_2747,N_2777);
and UO_260 (O_260,N_2281,N_2995);
and UO_261 (O_261,N_2981,N_2646);
nor UO_262 (O_262,N_2461,N_2538);
or UO_263 (O_263,N_2315,N_2341);
or UO_264 (O_264,N_2690,N_2766);
and UO_265 (O_265,N_2922,N_2342);
xnor UO_266 (O_266,N_2871,N_2909);
nand UO_267 (O_267,N_2863,N_2684);
xor UO_268 (O_268,N_2831,N_2957);
xnor UO_269 (O_269,N_2952,N_2560);
nor UO_270 (O_270,N_2806,N_2540);
or UO_271 (O_271,N_2530,N_2392);
nor UO_272 (O_272,N_2709,N_2667);
xor UO_273 (O_273,N_2688,N_2887);
nor UO_274 (O_274,N_2998,N_2399);
nor UO_275 (O_275,N_2849,N_2744);
xor UO_276 (O_276,N_2498,N_2449);
nand UO_277 (O_277,N_2404,N_2662);
nand UO_278 (O_278,N_2963,N_2913);
or UO_279 (O_279,N_2927,N_2841);
nor UO_280 (O_280,N_2782,N_2676);
nor UO_281 (O_281,N_2588,N_2256);
xnor UO_282 (O_282,N_2854,N_2764);
xnor UO_283 (O_283,N_2608,N_2931);
nand UO_284 (O_284,N_2589,N_2882);
xor UO_285 (O_285,N_2535,N_2734);
nor UO_286 (O_286,N_2725,N_2743);
nor UO_287 (O_287,N_2868,N_2362);
nand UO_288 (O_288,N_2875,N_2521);
nor UO_289 (O_289,N_2500,N_2568);
nor UO_290 (O_290,N_2495,N_2653);
and UO_291 (O_291,N_2402,N_2419);
nand UO_292 (O_292,N_2612,N_2416);
nand UO_293 (O_293,N_2465,N_2440);
and UO_294 (O_294,N_2477,N_2650);
and UO_295 (O_295,N_2372,N_2271);
and UO_296 (O_296,N_2619,N_2507);
or UO_297 (O_297,N_2737,N_2707);
xor UO_298 (O_298,N_2752,N_2541);
or UO_299 (O_299,N_2855,N_2840);
nand UO_300 (O_300,N_2796,N_2369);
or UO_301 (O_301,N_2370,N_2573);
xor UO_302 (O_302,N_2897,N_2906);
or UO_303 (O_303,N_2433,N_2463);
and UO_304 (O_304,N_2636,N_2567);
xnor UO_305 (O_305,N_2527,N_2547);
nor UO_306 (O_306,N_2742,N_2584);
nand UO_307 (O_307,N_2923,N_2480);
nand UO_308 (O_308,N_2973,N_2550);
or UO_309 (O_309,N_2975,N_2580);
and UO_310 (O_310,N_2704,N_2808);
and UO_311 (O_311,N_2911,N_2829);
xnor UO_312 (O_312,N_2925,N_2953);
xor UO_313 (O_313,N_2387,N_2592);
nor UO_314 (O_314,N_2610,N_2496);
nand UO_315 (O_315,N_2631,N_2892);
nand UO_316 (O_316,N_2898,N_2801);
xor UO_317 (O_317,N_2275,N_2947);
or UO_318 (O_318,N_2616,N_2605);
xor UO_319 (O_319,N_2397,N_2768);
and UO_320 (O_320,N_2575,N_2626);
or UO_321 (O_321,N_2844,N_2534);
or UO_322 (O_322,N_2993,N_2986);
xor UO_323 (O_323,N_2934,N_2784);
nand UO_324 (O_324,N_2838,N_2258);
nor UO_325 (O_325,N_2421,N_2792);
and UO_326 (O_326,N_2549,N_2767);
xnor UO_327 (O_327,N_2382,N_2593);
and UO_328 (O_328,N_2504,N_2501);
nand UO_329 (O_329,N_2731,N_2669);
nand UO_330 (O_330,N_2437,N_2520);
or UO_331 (O_331,N_2268,N_2358);
nand UO_332 (O_332,N_2893,N_2978);
nand UO_333 (O_333,N_2982,N_2696);
xor UO_334 (O_334,N_2296,N_2400);
nor UO_335 (O_335,N_2489,N_2508);
and UO_336 (O_336,N_2292,N_2988);
nand UO_337 (O_337,N_2347,N_2265);
nand UO_338 (O_338,N_2783,N_2264);
nand UO_339 (O_339,N_2411,N_2340);
nor UO_340 (O_340,N_2512,N_2581);
and UO_341 (O_341,N_2457,N_2531);
or UO_342 (O_342,N_2850,N_2697);
xor UO_343 (O_343,N_2435,N_2375);
and UO_344 (O_344,N_2368,N_2760);
or UO_345 (O_345,N_2918,N_2493);
and UO_346 (O_346,N_2334,N_2460);
nand UO_347 (O_347,N_2835,N_2318);
nor UO_348 (O_348,N_2464,N_2274);
or UO_349 (O_349,N_2604,N_2819);
or UO_350 (O_350,N_2409,N_2723);
and UO_351 (O_351,N_2300,N_2627);
nor UO_352 (O_352,N_2481,N_2961);
nor UO_353 (O_353,N_2492,N_2418);
xnor UO_354 (O_354,N_2360,N_2310);
nand UO_355 (O_355,N_2325,N_2901);
xor UO_356 (O_356,N_2277,N_2506);
or UO_357 (O_357,N_2390,N_2361);
nor UO_358 (O_358,N_2252,N_2536);
nor UO_359 (O_359,N_2432,N_2853);
nor UO_360 (O_360,N_2351,N_2857);
nand UO_361 (O_361,N_2793,N_2845);
nand UO_362 (O_362,N_2298,N_2329);
and UO_363 (O_363,N_2716,N_2269);
xnor UO_364 (O_364,N_2513,N_2282);
and UO_365 (O_365,N_2472,N_2312);
and UO_366 (O_366,N_2607,N_2757);
xor UO_367 (O_367,N_2410,N_2365);
nor UO_368 (O_368,N_2297,N_2283);
xor UO_369 (O_369,N_2668,N_2445);
and UO_370 (O_370,N_2479,N_2532);
nand UO_371 (O_371,N_2641,N_2615);
or UO_372 (O_372,N_2817,N_2253);
xor UO_373 (O_373,N_2884,N_2355);
and UO_374 (O_374,N_2915,N_2494);
nand UO_375 (O_375,N_2695,N_2816);
or UO_376 (O_376,N_2821,N_2500);
nor UO_377 (O_377,N_2539,N_2447);
xor UO_378 (O_378,N_2826,N_2287);
nor UO_379 (O_379,N_2591,N_2523);
or UO_380 (O_380,N_2496,N_2792);
nand UO_381 (O_381,N_2659,N_2271);
nor UO_382 (O_382,N_2740,N_2706);
xor UO_383 (O_383,N_2757,N_2317);
nand UO_384 (O_384,N_2756,N_2394);
xnor UO_385 (O_385,N_2929,N_2684);
xnor UO_386 (O_386,N_2927,N_2703);
xor UO_387 (O_387,N_2729,N_2885);
and UO_388 (O_388,N_2328,N_2809);
nor UO_389 (O_389,N_2421,N_2509);
xor UO_390 (O_390,N_2963,N_2571);
or UO_391 (O_391,N_2587,N_2713);
or UO_392 (O_392,N_2689,N_2507);
or UO_393 (O_393,N_2403,N_2880);
or UO_394 (O_394,N_2848,N_2583);
and UO_395 (O_395,N_2893,N_2955);
and UO_396 (O_396,N_2562,N_2379);
or UO_397 (O_397,N_2460,N_2905);
xor UO_398 (O_398,N_2439,N_2361);
nand UO_399 (O_399,N_2576,N_2433);
nand UO_400 (O_400,N_2905,N_2670);
xor UO_401 (O_401,N_2881,N_2312);
and UO_402 (O_402,N_2414,N_2407);
and UO_403 (O_403,N_2651,N_2285);
and UO_404 (O_404,N_2982,N_2334);
xnor UO_405 (O_405,N_2478,N_2517);
and UO_406 (O_406,N_2717,N_2556);
nand UO_407 (O_407,N_2560,N_2562);
xor UO_408 (O_408,N_2352,N_2774);
nor UO_409 (O_409,N_2937,N_2293);
nand UO_410 (O_410,N_2491,N_2353);
xnor UO_411 (O_411,N_2795,N_2473);
and UO_412 (O_412,N_2627,N_2635);
and UO_413 (O_413,N_2411,N_2613);
and UO_414 (O_414,N_2937,N_2739);
xor UO_415 (O_415,N_2764,N_2369);
or UO_416 (O_416,N_2715,N_2818);
nand UO_417 (O_417,N_2864,N_2420);
or UO_418 (O_418,N_2278,N_2385);
xnor UO_419 (O_419,N_2769,N_2862);
or UO_420 (O_420,N_2364,N_2609);
nand UO_421 (O_421,N_2877,N_2592);
nor UO_422 (O_422,N_2625,N_2808);
or UO_423 (O_423,N_2646,N_2886);
and UO_424 (O_424,N_2858,N_2359);
or UO_425 (O_425,N_2782,N_2898);
and UO_426 (O_426,N_2314,N_2521);
nand UO_427 (O_427,N_2279,N_2434);
nor UO_428 (O_428,N_2619,N_2628);
and UO_429 (O_429,N_2717,N_2690);
and UO_430 (O_430,N_2889,N_2262);
nor UO_431 (O_431,N_2972,N_2904);
or UO_432 (O_432,N_2712,N_2474);
xor UO_433 (O_433,N_2449,N_2712);
or UO_434 (O_434,N_2420,N_2389);
nand UO_435 (O_435,N_2754,N_2795);
or UO_436 (O_436,N_2288,N_2861);
and UO_437 (O_437,N_2807,N_2907);
or UO_438 (O_438,N_2316,N_2320);
nor UO_439 (O_439,N_2710,N_2645);
nor UO_440 (O_440,N_2434,N_2370);
nor UO_441 (O_441,N_2813,N_2614);
nand UO_442 (O_442,N_2937,N_2800);
or UO_443 (O_443,N_2537,N_2598);
xnor UO_444 (O_444,N_2328,N_2600);
nor UO_445 (O_445,N_2808,N_2775);
nor UO_446 (O_446,N_2795,N_2474);
or UO_447 (O_447,N_2742,N_2355);
and UO_448 (O_448,N_2592,N_2495);
and UO_449 (O_449,N_2276,N_2729);
and UO_450 (O_450,N_2267,N_2740);
and UO_451 (O_451,N_2428,N_2809);
nand UO_452 (O_452,N_2380,N_2991);
and UO_453 (O_453,N_2403,N_2656);
or UO_454 (O_454,N_2605,N_2644);
or UO_455 (O_455,N_2800,N_2608);
nor UO_456 (O_456,N_2450,N_2571);
or UO_457 (O_457,N_2343,N_2325);
xnor UO_458 (O_458,N_2756,N_2771);
or UO_459 (O_459,N_2323,N_2470);
and UO_460 (O_460,N_2460,N_2434);
nor UO_461 (O_461,N_2513,N_2507);
or UO_462 (O_462,N_2389,N_2830);
nor UO_463 (O_463,N_2576,N_2746);
xnor UO_464 (O_464,N_2311,N_2486);
or UO_465 (O_465,N_2946,N_2958);
nor UO_466 (O_466,N_2997,N_2896);
nand UO_467 (O_467,N_2481,N_2308);
nor UO_468 (O_468,N_2731,N_2816);
or UO_469 (O_469,N_2656,N_2978);
or UO_470 (O_470,N_2435,N_2393);
nand UO_471 (O_471,N_2253,N_2992);
nor UO_472 (O_472,N_2405,N_2916);
xor UO_473 (O_473,N_2478,N_2730);
nand UO_474 (O_474,N_2908,N_2663);
nor UO_475 (O_475,N_2465,N_2705);
nand UO_476 (O_476,N_2318,N_2387);
nor UO_477 (O_477,N_2426,N_2681);
and UO_478 (O_478,N_2689,N_2279);
or UO_479 (O_479,N_2721,N_2795);
xor UO_480 (O_480,N_2481,N_2325);
nand UO_481 (O_481,N_2931,N_2433);
or UO_482 (O_482,N_2380,N_2932);
and UO_483 (O_483,N_2431,N_2829);
xnor UO_484 (O_484,N_2581,N_2451);
nand UO_485 (O_485,N_2531,N_2576);
xnor UO_486 (O_486,N_2970,N_2378);
and UO_487 (O_487,N_2862,N_2675);
nand UO_488 (O_488,N_2454,N_2697);
xor UO_489 (O_489,N_2701,N_2256);
nand UO_490 (O_490,N_2400,N_2554);
xor UO_491 (O_491,N_2896,N_2334);
xor UO_492 (O_492,N_2619,N_2823);
nand UO_493 (O_493,N_2835,N_2359);
or UO_494 (O_494,N_2563,N_2859);
xnor UO_495 (O_495,N_2494,N_2646);
and UO_496 (O_496,N_2629,N_2563);
nand UO_497 (O_497,N_2354,N_2811);
and UO_498 (O_498,N_2278,N_2772);
and UO_499 (O_499,N_2798,N_2865);
endmodule