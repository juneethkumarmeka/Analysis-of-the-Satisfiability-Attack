module basic_500_3000_500_3_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_211,In_239);
xnor U1 (N_1,In_416,In_489);
nand U2 (N_2,In_354,In_132);
xor U3 (N_3,In_279,In_126);
nand U4 (N_4,In_454,In_66);
xor U5 (N_5,In_178,In_165);
xor U6 (N_6,In_161,In_310);
nor U7 (N_7,In_380,In_272);
and U8 (N_8,In_363,In_192);
xor U9 (N_9,In_460,In_295);
or U10 (N_10,In_313,In_494);
xor U11 (N_11,In_248,In_333);
nand U12 (N_12,In_458,In_6);
xnor U13 (N_13,In_235,In_409);
xnor U14 (N_14,In_260,In_332);
or U15 (N_15,In_434,In_375);
and U16 (N_16,In_207,In_309);
and U17 (N_17,In_120,In_254);
and U18 (N_18,In_155,In_73);
xnor U19 (N_19,In_92,In_237);
and U20 (N_20,In_480,In_497);
nor U21 (N_21,In_232,In_338);
xor U22 (N_22,In_361,In_17);
nor U23 (N_23,In_439,In_445);
xor U24 (N_24,In_205,In_326);
nor U25 (N_25,In_209,In_60);
xnor U26 (N_26,In_9,In_459);
nor U27 (N_27,In_321,In_101);
or U28 (N_28,In_187,In_369);
xor U29 (N_29,In_122,In_371);
or U30 (N_30,In_173,In_314);
nor U31 (N_31,In_399,In_418);
xnor U32 (N_32,In_202,In_44);
nand U33 (N_33,In_72,In_374);
nor U34 (N_34,In_137,In_322);
and U35 (N_35,In_293,In_53);
xor U36 (N_36,In_340,In_87);
and U37 (N_37,In_141,In_258);
xnor U38 (N_38,In_482,In_164);
and U39 (N_39,In_347,In_378);
or U40 (N_40,In_426,In_135);
and U41 (N_41,In_413,In_140);
nor U42 (N_42,In_414,In_197);
xnor U43 (N_43,In_407,In_10);
or U44 (N_44,In_220,In_107);
nand U45 (N_45,In_334,In_465);
nor U46 (N_46,In_269,In_475);
or U47 (N_47,In_70,In_134);
xnor U48 (N_48,In_429,In_243);
nor U49 (N_49,In_64,In_149);
or U50 (N_50,In_303,In_224);
nand U51 (N_51,In_447,In_163);
and U52 (N_52,In_34,In_183);
and U53 (N_53,In_46,In_138);
or U54 (N_54,In_204,In_170);
xor U55 (N_55,In_136,In_95);
nand U56 (N_56,In_198,In_287);
or U57 (N_57,In_49,In_75);
xnor U58 (N_58,In_125,In_423);
nor U59 (N_59,In_194,In_278);
or U60 (N_60,In_487,In_167);
xnor U61 (N_61,In_115,In_233);
nand U62 (N_62,In_308,In_388);
nor U63 (N_63,In_244,In_365);
or U64 (N_64,In_415,In_306);
or U65 (N_65,In_346,In_215);
nor U66 (N_66,In_495,In_417);
and U67 (N_67,In_223,In_474);
xnor U68 (N_68,In_39,In_370);
and U69 (N_69,In_214,In_102);
and U70 (N_70,In_411,In_216);
xnor U71 (N_71,In_16,In_21);
nand U72 (N_72,In_477,In_284);
nor U73 (N_73,In_291,In_432);
nor U74 (N_74,In_241,In_180);
nor U75 (N_75,In_320,In_276);
and U76 (N_76,In_142,In_103);
xor U77 (N_77,In_43,In_403);
or U78 (N_78,In_355,In_47);
xor U79 (N_79,In_182,In_315);
nor U80 (N_80,In_491,In_41);
xor U81 (N_81,In_82,In_33);
xnor U82 (N_82,In_419,In_457);
nor U83 (N_83,In_30,In_225);
nor U84 (N_84,In_357,In_240);
and U85 (N_85,In_430,In_36);
xor U86 (N_86,In_290,In_106);
nand U87 (N_87,In_468,In_257);
nor U88 (N_88,In_174,In_345);
or U89 (N_89,In_473,In_159);
xnor U90 (N_90,In_461,In_234);
xor U91 (N_91,In_379,In_110);
nand U92 (N_92,In_440,In_448);
and U93 (N_93,In_443,In_302);
and U94 (N_94,In_230,In_61);
or U95 (N_95,In_130,In_266);
xor U96 (N_96,In_329,In_63);
nor U97 (N_97,In_1,In_492);
nor U98 (N_98,In_65,In_146);
xnor U99 (N_99,In_152,In_50);
and U100 (N_100,In_376,In_394);
nand U101 (N_101,In_40,In_263);
and U102 (N_102,In_479,In_2);
or U103 (N_103,In_78,In_79);
xnor U104 (N_104,In_26,In_97);
or U105 (N_105,In_188,In_435);
and U106 (N_106,In_160,In_20);
or U107 (N_107,In_285,In_493);
or U108 (N_108,In_350,In_496);
nor U109 (N_109,In_166,In_108);
or U110 (N_110,In_386,In_499);
nand U111 (N_111,In_292,In_286);
and U112 (N_112,In_307,In_94);
nor U113 (N_113,In_297,In_13);
or U114 (N_114,In_123,In_294);
nor U115 (N_115,In_451,In_362);
xnor U116 (N_116,In_245,In_219);
or U117 (N_117,In_452,In_169);
nor U118 (N_118,In_498,In_264);
xnor U119 (N_119,In_100,In_90);
xor U120 (N_120,In_19,In_481);
xor U121 (N_121,In_31,In_368);
xor U122 (N_122,In_151,In_144);
xnor U123 (N_123,In_217,In_88);
nor U124 (N_124,In_444,In_406);
and U125 (N_125,In_80,In_55);
xnor U126 (N_126,In_181,In_441);
or U127 (N_127,In_324,In_208);
nand U128 (N_128,In_238,In_171);
xnor U129 (N_129,In_450,In_62);
xnor U130 (N_130,In_466,In_341);
xnor U131 (N_131,In_54,In_401);
or U132 (N_132,In_277,In_455);
nand U133 (N_133,In_304,In_8);
nor U134 (N_134,In_328,In_358);
or U135 (N_135,In_133,In_176);
nor U136 (N_136,In_390,In_471);
nand U137 (N_137,In_112,In_428);
or U138 (N_138,In_89,In_131);
nor U139 (N_139,In_23,In_317);
and U140 (N_140,In_425,In_145);
xor U141 (N_141,In_15,In_400);
and U142 (N_142,In_117,In_300);
nand U143 (N_143,In_18,In_256);
or U144 (N_144,In_372,In_190);
or U145 (N_145,In_484,In_253);
or U146 (N_146,In_154,In_476);
nor U147 (N_147,In_381,In_335);
xor U148 (N_148,In_349,In_485);
nor U149 (N_149,In_218,In_37);
nand U150 (N_150,In_360,In_305);
or U151 (N_151,In_195,In_25);
or U152 (N_152,In_121,In_29);
and U153 (N_153,In_456,In_299);
or U154 (N_154,In_177,In_339);
xnor U155 (N_155,In_453,In_81);
xor U156 (N_156,In_38,In_283);
nor U157 (N_157,In_472,In_311);
xor U158 (N_158,In_77,In_255);
xnor U159 (N_159,In_270,In_199);
nor U160 (N_160,In_228,In_249);
and U161 (N_161,In_402,In_221);
nand U162 (N_162,In_464,In_196);
nor U163 (N_163,In_420,In_282);
nand U164 (N_164,In_325,In_5);
nor U165 (N_165,In_252,In_84);
or U166 (N_166,In_113,In_442);
or U167 (N_167,In_93,In_373);
xnor U168 (N_168,In_393,In_236);
and U169 (N_169,In_344,In_86);
and U170 (N_170,In_446,In_56);
nor U171 (N_171,In_438,In_377);
and U172 (N_172,In_470,In_143);
or U173 (N_173,In_449,In_312);
or U174 (N_174,In_437,In_210);
nor U175 (N_175,In_391,In_27);
nor U176 (N_176,In_229,In_383);
and U177 (N_177,In_222,In_227);
xor U178 (N_178,In_319,In_127);
and U179 (N_179,In_323,In_3);
or U180 (N_180,In_273,In_488);
or U181 (N_181,In_71,In_268);
nand U182 (N_182,In_280,In_42);
nor U183 (N_183,In_261,In_316);
xnor U184 (N_184,In_35,In_109);
nor U185 (N_185,In_367,In_68);
nand U186 (N_186,In_99,In_343);
nor U187 (N_187,In_118,In_69);
and U188 (N_188,In_247,In_433);
nor U189 (N_189,In_184,In_342);
or U190 (N_190,In_150,In_246);
or U191 (N_191,In_168,In_7);
and U192 (N_192,In_111,In_147);
xnor U193 (N_193,In_327,In_22);
and U194 (N_194,In_0,In_395);
or U195 (N_195,In_116,In_410);
xor U196 (N_196,In_201,In_348);
and U197 (N_197,In_124,In_296);
and U198 (N_198,In_431,In_436);
nor U199 (N_199,In_271,In_486);
or U200 (N_200,In_11,In_179);
nand U201 (N_201,In_148,In_74);
and U202 (N_202,In_212,In_250);
nor U203 (N_203,In_59,In_45);
xnor U204 (N_204,In_4,In_231);
xnor U205 (N_205,In_265,In_189);
or U206 (N_206,In_424,In_397);
xor U207 (N_207,In_356,In_289);
nand U208 (N_208,In_337,In_104);
and U209 (N_209,In_387,In_83);
or U210 (N_210,In_96,In_427);
or U211 (N_211,In_193,In_382);
xor U212 (N_212,In_421,In_364);
xor U213 (N_213,In_408,In_359);
xnor U214 (N_214,In_12,In_274);
xnor U215 (N_215,In_259,In_412);
nand U216 (N_216,In_331,In_404);
xnor U217 (N_217,In_288,In_52);
nor U218 (N_218,In_389,In_275);
or U219 (N_219,In_251,In_162);
and U220 (N_220,In_85,In_483);
xor U221 (N_221,In_200,In_58);
and U222 (N_222,In_298,In_114);
nor U223 (N_223,In_24,In_191);
xor U224 (N_224,In_213,In_185);
xnor U225 (N_225,In_186,In_281);
and U226 (N_226,In_462,In_128);
nand U227 (N_227,In_14,In_139);
nand U228 (N_228,In_330,In_384);
xor U229 (N_229,In_156,In_385);
nor U230 (N_230,In_352,In_105);
or U231 (N_231,In_76,In_175);
nand U232 (N_232,In_467,In_203);
and U233 (N_233,In_336,In_153);
nor U234 (N_234,In_48,In_463);
or U235 (N_235,In_98,In_32);
nand U236 (N_236,In_398,In_469);
and U237 (N_237,In_67,In_158);
or U238 (N_238,In_119,In_262);
nand U239 (N_239,In_366,In_51);
nand U240 (N_240,In_422,In_392);
nand U241 (N_241,In_157,In_490);
nand U242 (N_242,In_478,In_405);
nor U243 (N_243,In_91,In_318);
nor U244 (N_244,In_267,In_301);
nor U245 (N_245,In_226,In_28);
or U246 (N_246,In_129,In_206);
nor U247 (N_247,In_396,In_242);
nor U248 (N_248,In_353,In_351);
xnor U249 (N_249,In_57,In_172);
and U250 (N_250,In_202,In_329);
and U251 (N_251,In_175,In_399);
xor U252 (N_252,In_92,In_355);
xor U253 (N_253,In_136,In_259);
nor U254 (N_254,In_378,In_448);
nor U255 (N_255,In_447,In_134);
nand U256 (N_256,In_240,In_232);
or U257 (N_257,In_175,In_80);
or U258 (N_258,In_329,In_444);
and U259 (N_259,In_261,In_302);
nor U260 (N_260,In_123,In_188);
nor U261 (N_261,In_129,In_172);
or U262 (N_262,In_121,In_144);
xor U263 (N_263,In_493,In_31);
and U264 (N_264,In_43,In_100);
nor U265 (N_265,In_212,In_39);
or U266 (N_266,In_37,In_349);
and U267 (N_267,In_320,In_364);
or U268 (N_268,In_382,In_12);
or U269 (N_269,In_404,In_296);
and U270 (N_270,In_181,In_220);
nor U271 (N_271,In_217,In_28);
xnor U272 (N_272,In_344,In_92);
nand U273 (N_273,In_472,In_405);
xor U274 (N_274,In_1,In_284);
nand U275 (N_275,In_363,In_479);
nand U276 (N_276,In_195,In_143);
xor U277 (N_277,In_422,In_205);
nor U278 (N_278,In_498,In_1);
xor U279 (N_279,In_451,In_438);
and U280 (N_280,In_225,In_224);
xnor U281 (N_281,In_385,In_458);
or U282 (N_282,In_350,In_155);
nand U283 (N_283,In_32,In_279);
xnor U284 (N_284,In_96,In_322);
nand U285 (N_285,In_479,In_38);
nand U286 (N_286,In_79,In_145);
nor U287 (N_287,In_90,In_480);
or U288 (N_288,In_299,In_441);
and U289 (N_289,In_42,In_485);
xnor U290 (N_290,In_430,In_416);
nor U291 (N_291,In_314,In_2);
or U292 (N_292,In_388,In_279);
or U293 (N_293,In_7,In_164);
nand U294 (N_294,In_68,In_290);
nor U295 (N_295,In_161,In_172);
and U296 (N_296,In_157,In_161);
and U297 (N_297,In_89,In_413);
xnor U298 (N_298,In_343,In_427);
and U299 (N_299,In_179,In_104);
and U300 (N_300,In_171,In_409);
xnor U301 (N_301,In_312,In_74);
or U302 (N_302,In_229,In_160);
or U303 (N_303,In_436,In_119);
xnor U304 (N_304,In_61,In_177);
nor U305 (N_305,In_293,In_189);
nor U306 (N_306,In_25,In_40);
and U307 (N_307,In_214,In_2);
or U308 (N_308,In_285,In_151);
nand U309 (N_309,In_492,In_378);
and U310 (N_310,In_200,In_347);
or U311 (N_311,In_473,In_166);
nor U312 (N_312,In_228,In_20);
nand U313 (N_313,In_369,In_443);
and U314 (N_314,In_492,In_288);
and U315 (N_315,In_135,In_365);
xor U316 (N_316,In_285,In_149);
nand U317 (N_317,In_97,In_25);
xor U318 (N_318,In_476,In_41);
nor U319 (N_319,In_97,In_232);
xor U320 (N_320,In_350,In_67);
nor U321 (N_321,In_156,In_483);
and U322 (N_322,In_51,In_389);
xnor U323 (N_323,In_388,In_115);
nand U324 (N_324,In_75,In_323);
nand U325 (N_325,In_431,In_494);
xor U326 (N_326,In_449,In_253);
and U327 (N_327,In_410,In_419);
xnor U328 (N_328,In_275,In_258);
or U329 (N_329,In_398,In_145);
xor U330 (N_330,In_95,In_217);
xor U331 (N_331,In_493,In_62);
nor U332 (N_332,In_497,In_221);
xnor U333 (N_333,In_456,In_118);
or U334 (N_334,In_307,In_478);
and U335 (N_335,In_137,In_328);
nor U336 (N_336,In_466,In_286);
and U337 (N_337,In_214,In_133);
and U338 (N_338,In_121,In_186);
or U339 (N_339,In_257,In_52);
or U340 (N_340,In_115,In_415);
nand U341 (N_341,In_38,In_455);
and U342 (N_342,In_368,In_3);
or U343 (N_343,In_252,In_186);
and U344 (N_344,In_196,In_269);
and U345 (N_345,In_190,In_84);
nand U346 (N_346,In_35,In_264);
and U347 (N_347,In_148,In_9);
or U348 (N_348,In_211,In_322);
and U349 (N_349,In_344,In_48);
or U350 (N_350,In_260,In_274);
nor U351 (N_351,In_25,In_349);
xor U352 (N_352,In_450,In_221);
nand U353 (N_353,In_159,In_91);
or U354 (N_354,In_171,In_493);
nor U355 (N_355,In_342,In_378);
nor U356 (N_356,In_363,In_471);
nor U357 (N_357,In_97,In_118);
and U358 (N_358,In_12,In_3);
and U359 (N_359,In_341,In_241);
nand U360 (N_360,In_190,In_155);
and U361 (N_361,In_106,In_307);
and U362 (N_362,In_449,In_302);
nand U363 (N_363,In_446,In_70);
or U364 (N_364,In_67,In_490);
and U365 (N_365,In_133,In_404);
or U366 (N_366,In_35,In_195);
and U367 (N_367,In_240,In_109);
and U368 (N_368,In_167,In_405);
nor U369 (N_369,In_353,In_152);
nor U370 (N_370,In_123,In_485);
xor U371 (N_371,In_154,In_171);
nand U372 (N_372,In_439,In_21);
or U373 (N_373,In_78,In_402);
or U374 (N_374,In_138,In_384);
nor U375 (N_375,In_64,In_37);
nor U376 (N_376,In_440,In_23);
nand U377 (N_377,In_262,In_292);
nor U378 (N_378,In_302,In_162);
nor U379 (N_379,In_464,In_41);
nor U380 (N_380,In_21,In_163);
xnor U381 (N_381,In_227,In_78);
nand U382 (N_382,In_360,In_292);
nand U383 (N_383,In_90,In_175);
nand U384 (N_384,In_67,In_56);
xnor U385 (N_385,In_363,In_433);
nor U386 (N_386,In_26,In_299);
nor U387 (N_387,In_102,In_205);
nor U388 (N_388,In_341,In_203);
nor U389 (N_389,In_473,In_368);
and U390 (N_390,In_261,In_156);
or U391 (N_391,In_276,In_347);
nand U392 (N_392,In_371,In_133);
and U393 (N_393,In_306,In_98);
xnor U394 (N_394,In_444,In_421);
nand U395 (N_395,In_196,In_366);
nor U396 (N_396,In_369,In_132);
nor U397 (N_397,In_129,In_188);
xnor U398 (N_398,In_154,In_312);
nor U399 (N_399,In_106,In_367);
xor U400 (N_400,In_486,In_277);
or U401 (N_401,In_376,In_322);
and U402 (N_402,In_347,In_210);
or U403 (N_403,In_229,In_245);
and U404 (N_404,In_446,In_352);
nand U405 (N_405,In_495,In_244);
xnor U406 (N_406,In_258,In_154);
and U407 (N_407,In_254,In_229);
nand U408 (N_408,In_386,In_238);
xor U409 (N_409,In_232,In_332);
and U410 (N_410,In_21,In_405);
xnor U411 (N_411,In_287,In_85);
nand U412 (N_412,In_149,In_138);
nand U413 (N_413,In_388,In_233);
and U414 (N_414,In_271,In_249);
or U415 (N_415,In_63,In_125);
nand U416 (N_416,In_343,In_180);
and U417 (N_417,In_158,In_486);
or U418 (N_418,In_427,In_208);
nand U419 (N_419,In_229,In_205);
or U420 (N_420,In_65,In_104);
or U421 (N_421,In_193,In_346);
and U422 (N_422,In_227,In_323);
nand U423 (N_423,In_401,In_274);
or U424 (N_424,In_459,In_100);
or U425 (N_425,In_165,In_410);
nand U426 (N_426,In_498,In_153);
and U427 (N_427,In_481,In_89);
or U428 (N_428,In_359,In_254);
and U429 (N_429,In_184,In_313);
xnor U430 (N_430,In_240,In_468);
nand U431 (N_431,In_263,In_463);
nand U432 (N_432,In_245,In_232);
xnor U433 (N_433,In_408,In_499);
nand U434 (N_434,In_385,In_403);
nand U435 (N_435,In_208,In_458);
xnor U436 (N_436,In_83,In_99);
nand U437 (N_437,In_260,In_402);
or U438 (N_438,In_166,In_319);
and U439 (N_439,In_440,In_306);
xor U440 (N_440,In_331,In_496);
xnor U441 (N_441,In_298,In_368);
xnor U442 (N_442,In_126,In_407);
nor U443 (N_443,In_119,In_449);
or U444 (N_444,In_417,In_118);
and U445 (N_445,In_400,In_422);
or U446 (N_446,In_449,In_431);
or U447 (N_447,In_447,In_129);
and U448 (N_448,In_70,In_445);
nor U449 (N_449,In_167,In_484);
nor U450 (N_450,In_412,In_15);
xor U451 (N_451,In_236,In_60);
and U452 (N_452,In_468,In_229);
nor U453 (N_453,In_451,In_421);
xor U454 (N_454,In_344,In_24);
or U455 (N_455,In_231,In_498);
or U456 (N_456,In_274,In_453);
and U457 (N_457,In_50,In_127);
and U458 (N_458,In_409,In_323);
nor U459 (N_459,In_328,In_7);
nand U460 (N_460,In_268,In_347);
nor U461 (N_461,In_212,In_73);
nor U462 (N_462,In_352,In_231);
nor U463 (N_463,In_399,In_410);
and U464 (N_464,In_445,In_199);
xor U465 (N_465,In_342,In_447);
nand U466 (N_466,In_311,In_179);
nand U467 (N_467,In_89,In_164);
nand U468 (N_468,In_414,In_90);
xor U469 (N_469,In_154,In_67);
or U470 (N_470,In_31,In_83);
or U471 (N_471,In_97,In_298);
or U472 (N_472,In_169,In_58);
and U473 (N_473,In_274,In_498);
or U474 (N_474,In_107,In_265);
nor U475 (N_475,In_253,In_336);
and U476 (N_476,In_389,In_396);
or U477 (N_477,In_239,In_452);
or U478 (N_478,In_226,In_50);
nor U479 (N_479,In_98,In_217);
nand U480 (N_480,In_236,In_368);
and U481 (N_481,In_35,In_219);
or U482 (N_482,In_473,In_493);
nand U483 (N_483,In_212,In_36);
and U484 (N_484,In_277,In_249);
nand U485 (N_485,In_296,In_175);
and U486 (N_486,In_214,In_410);
nand U487 (N_487,In_393,In_6);
and U488 (N_488,In_453,In_260);
nor U489 (N_489,In_382,In_402);
xnor U490 (N_490,In_5,In_464);
and U491 (N_491,In_344,In_306);
nand U492 (N_492,In_462,In_190);
nand U493 (N_493,In_48,In_474);
nor U494 (N_494,In_366,In_53);
nor U495 (N_495,In_246,In_369);
or U496 (N_496,In_41,In_481);
or U497 (N_497,In_132,In_151);
xnor U498 (N_498,In_288,In_468);
xor U499 (N_499,In_119,In_317);
xnor U500 (N_500,In_40,In_360);
nor U501 (N_501,In_94,In_433);
xnor U502 (N_502,In_46,In_277);
nor U503 (N_503,In_262,In_163);
and U504 (N_504,In_5,In_179);
xnor U505 (N_505,In_151,In_112);
or U506 (N_506,In_62,In_142);
and U507 (N_507,In_49,In_203);
nor U508 (N_508,In_22,In_324);
and U509 (N_509,In_464,In_368);
and U510 (N_510,In_325,In_131);
or U511 (N_511,In_19,In_60);
nand U512 (N_512,In_490,In_28);
xnor U513 (N_513,In_234,In_394);
nor U514 (N_514,In_267,In_156);
nand U515 (N_515,In_389,In_305);
or U516 (N_516,In_331,In_3);
xnor U517 (N_517,In_462,In_19);
xnor U518 (N_518,In_160,In_486);
nor U519 (N_519,In_63,In_96);
and U520 (N_520,In_126,In_35);
nand U521 (N_521,In_408,In_151);
nand U522 (N_522,In_227,In_239);
xnor U523 (N_523,In_218,In_331);
or U524 (N_524,In_246,In_235);
xor U525 (N_525,In_483,In_212);
and U526 (N_526,In_363,In_494);
or U527 (N_527,In_80,In_47);
nor U528 (N_528,In_465,In_321);
nor U529 (N_529,In_369,In_330);
xor U530 (N_530,In_321,In_368);
nor U531 (N_531,In_268,In_439);
xor U532 (N_532,In_318,In_376);
nand U533 (N_533,In_189,In_498);
and U534 (N_534,In_364,In_344);
nand U535 (N_535,In_74,In_78);
or U536 (N_536,In_120,In_218);
or U537 (N_537,In_165,In_281);
xnor U538 (N_538,In_149,In_333);
xor U539 (N_539,In_95,In_67);
and U540 (N_540,In_159,In_33);
or U541 (N_541,In_395,In_228);
and U542 (N_542,In_290,In_233);
nand U543 (N_543,In_25,In_228);
nor U544 (N_544,In_270,In_182);
nand U545 (N_545,In_4,In_178);
or U546 (N_546,In_438,In_93);
nand U547 (N_547,In_496,In_451);
nand U548 (N_548,In_302,In_255);
and U549 (N_549,In_400,In_372);
or U550 (N_550,In_124,In_415);
xor U551 (N_551,In_54,In_199);
or U552 (N_552,In_371,In_375);
nand U553 (N_553,In_225,In_221);
xor U554 (N_554,In_231,In_234);
and U555 (N_555,In_422,In_488);
and U556 (N_556,In_480,In_163);
or U557 (N_557,In_149,In_402);
nand U558 (N_558,In_80,In_62);
nor U559 (N_559,In_397,In_224);
and U560 (N_560,In_207,In_341);
nor U561 (N_561,In_128,In_56);
and U562 (N_562,In_44,In_382);
or U563 (N_563,In_149,In_190);
nand U564 (N_564,In_122,In_217);
nand U565 (N_565,In_395,In_57);
nor U566 (N_566,In_221,In_301);
and U567 (N_567,In_90,In_72);
nand U568 (N_568,In_318,In_467);
nand U569 (N_569,In_285,In_29);
and U570 (N_570,In_360,In_285);
nor U571 (N_571,In_268,In_372);
xor U572 (N_572,In_79,In_412);
nor U573 (N_573,In_38,In_30);
and U574 (N_574,In_90,In_473);
or U575 (N_575,In_397,In_208);
nand U576 (N_576,In_206,In_71);
nor U577 (N_577,In_164,In_311);
or U578 (N_578,In_237,In_116);
or U579 (N_579,In_485,In_457);
nor U580 (N_580,In_428,In_247);
or U581 (N_581,In_144,In_185);
nor U582 (N_582,In_162,In_46);
and U583 (N_583,In_218,In_232);
nand U584 (N_584,In_432,In_277);
and U585 (N_585,In_333,In_222);
nor U586 (N_586,In_4,In_416);
nand U587 (N_587,In_254,In_496);
nand U588 (N_588,In_318,In_377);
and U589 (N_589,In_425,In_279);
xnor U590 (N_590,In_386,In_132);
and U591 (N_591,In_36,In_112);
and U592 (N_592,In_228,In_125);
or U593 (N_593,In_47,In_186);
and U594 (N_594,In_362,In_32);
nor U595 (N_595,In_399,In_243);
nor U596 (N_596,In_215,In_452);
xor U597 (N_597,In_260,In_223);
nor U598 (N_598,In_79,In_77);
or U599 (N_599,In_144,In_111);
or U600 (N_600,In_265,In_455);
nand U601 (N_601,In_245,In_293);
xnor U602 (N_602,In_311,In_361);
or U603 (N_603,In_97,In_267);
and U604 (N_604,In_291,In_427);
xnor U605 (N_605,In_118,In_221);
and U606 (N_606,In_141,In_31);
xor U607 (N_607,In_273,In_444);
or U608 (N_608,In_365,In_387);
nand U609 (N_609,In_391,In_190);
and U610 (N_610,In_406,In_17);
and U611 (N_611,In_421,In_231);
or U612 (N_612,In_139,In_4);
xor U613 (N_613,In_384,In_80);
and U614 (N_614,In_343,In_267);
or U615 (N_615,In_465,In_487);
nand U616 (N_616,In_344,In_141);
or U617 (N_617,In_182,In_220);
xnor U618 (N_618,In_100,In_279);
and U619 (N_619,In_477,In_388);
nand U620 (N_620,In_369,In_225);
nor U621 (N_621,In_332,In_138);
and U622 (N_622,In_243,In_442);
and U623 (N_623,In_207,In_318);
or U624 (N_624,In_22,In_194);
or U625 (N_625,In_486,In_208);
nand U626 (N_626,In_389,In_211);
and U627 (N_627,In_223,In_370);
nor U628 (N_628,In_497,In_133);
nand U629 (N_629,In_436,In_59);
xor U630 (N_630,In_45,In_131);
and U631 (N_631,In_106,In_348);
nand U632 (N_632,In_471,In_244);
xor U633 (N_633,In_366,In_223);
nor U634 (N_634,In_147,In_107);
xnor U635 (N_635,In_180,In_2);
or U636 (N_636,In_427,In_148);
or U637 (N_637,In_273,In_80);
or U638 (N_638,In_335,In_492);
nor U639 (N_639,In_16,In_215);
xnor U640 (N_640,In_337,In_290);
nor U641 (N_641,In_126,In_97);
and U642 (N_642,In_421,In_17);
nor U643 (N_643,In_474,In_360);
xnor U644 (N_644,In_343,In_330);
nand U645 (N_645,In_270,In_458);
xor U646 (N_646,In_489,In_303);
and U647 (N_647,In_169,In_264);
xor U648 (N_648,In_349,In_470);
xnor U649 (N_649,In_157,In_472);
and U650 (N_650,In_25,In_114);
nor U651 (N_651,In_203,In_8);
nor U652 (N_652,In_174,In_44);
and U653 (N_653,In_12,In_324);
and U654 (N_654,In_262,In_96);
or U655 (N_655,In_77,In_125);
xor U656 (N_656,In_392,In_245);
and U657 (N_657,In_281,In_31);
nor U658 (N_658,In_195,In_52);
nand U659 (N_659,In_78,In_331);
nor U660 (N_660,In_460,In_81);
or U661 (N_661,In_90,In_417);
or U662 (N_662,In_371,In_252);
nand U663 (N_663,In_73,In_486);
nor U664 (N_664,In_436,In_230);
nand U665 (N_665,In_482,In_343);
xnor U666 (N_666,In_185,In_442);
nand U667 (N_667,In_425,In_199);
xnor U668 (N_668,In_455,In_127);
xnor U669 (N_669,In_430,In_4);
or U670 (N_670,In_197,In_469);
xnor U671 (N_671,In_265,In_462);
xnor U672 (N_672,In_115,In_3);
nand U673 (N_673,In_132,In_75);
nand U674 (N_674,In_420,In_37);
xnor U675 (N_675,In_448,In_134);
nor U676 (N_676,In_373,In_135);
nor U677 (N_677,In_87,In_421);
or U678 (N_678,In_274,In_56);
and U679 (N_679,In_472,In_179);
or U680 (N_680,In_49,In_139);
or U681 (N_681,In_4,In_475);
or U682 (N_682,In_240,In_410);
and U683 (N_683,In_424,In_414);
or U684 (N_684,In_268,In_499);
nor U685 (N_685,In_320,In_442);
nor U686 (N_686,In_286,In_329);
or U687 (N_687,In_19,In_207);
nand U688 (N_688,In_272,In_314);
xor U689 (N_689,In_381,In_200);
nor U690 (N_690,In_227,In_71);
and U691 (N_691,In_202,In_42);
nand U692 (N_692,In_315,In_325);
or U693 (N_693,In_66,In_428);
nand U694 (N_694,In_154,In_163);
or U695 (N_695,In_430,In_187);
xor U696 (N_696,In_172,In_462);
nand U697 (N_697,In_218,In_341);
nand U698 (N_698,In_34,In_353);
or U699 (N_699,In_178,In_18);
xor U700 (N_700,In_388,In_218);
nor U701 (N_701,In_377,In_470);
xnor U702 (N_702,In_181,In_457);
nand U703 (N_703,In_146,In_466);
or U704 (N_704,In_244,In_212);
or U705 (N_705,In_357,In_59);
nand U706 (N_706,In_115,In_426);
or U707 (N_707,In_262,In_177);
or U708 (N_708,In_383,In_442);
and U709 (N_709,In_369,In_361);
xor U710 (N_710,In_77,In_141);
or U711 (N_711,In_280,In_293);
or U712 (N_712,In_4,In_376);
nor U713 (N_713,In_188,In_361);
or U714 (N_714,In_334,In_98);
and U715 (N_715,In_388,In_204);
nor U716 (N_716,In_425,In_18);
nor U717 (N_717,In_408,In_158);
and U718 (N_718,In_172,In_215);
or U719 (N_719,In_90,In_82);
xor U720 (N_720,In_135,In_460);
xor U721 (N_721,In_284,In_385);
and U722 (N_722,In_445,In_420);
nand U723 (N_723,In_388,In_341);
or U724 (N_724,In_349,In_399);
xnor U725 (N_725,In_186,In_114);
nand U726 (N_726,In_431,In_295);
and U727 (N_727,In_340,In_81);
nand U728 (N_728,In_140,In_157);
nand U729 (N_729,In_393,In_375);
and U730 (N_730,In_96,In_401);
nand U731 (N_731,In_405,In_227);
and U732 (N_732,In_46,In_383);
nand U733 (N_733,In_480,In_28);
nand U734 (N_734,In_114,In_202);
or U735 (N_735,In_253,In_10);
nand U736 (N_736,In_214,In_60);
or U737 (N_737,In_305,In_41);
and U738 (N_738,In_487,In_485);
or U739 (N_739,In_342,In_203);
or U740 (N_740,In_439,In_35);
xnor U741 (N_741,In_107,In_304);
and U742 (N_742,In_54,In_368);
nand U743 (N_743,In_43,In_159);
nand U744 (N_744,In_127,In_184);
nand U745 (N_745,In_258,In_384);
xnor U746 (N_746,In_288,In_477);
xor U747 (N_747,In_278,In_17);
nor U748 (N_748,In_399,In_165);
nor U749 (N_749,In_406,In_302);
nand U750 (N_750,In_43,In_157);
or U751 (N_751,In_30,In_430);
or U752 (N_752,In_243,In_16);
and U753 (N_753,In_459,In_15);
or U754 (N_754,In_148,In_155);
nor U755 (N_755,In_62,In_234);
nor U756 (N_756,In_11,In_39);
and U757 (N_757,In_304,In_111);
or U758 (N_758,In_297,In_368);
nor U759 (N_759,In_52,In_494);
nor U760 (N_760,In_415,In_390);
xnor U761 (N_761,In_464,In_143);
xor U762 (N_762,In_183,In_229);
nor U763 (N_763,In_355,In_127);
or U764 (N_764,In_457,In_204);
nor U765 (N_765,In_421,In_456);
or U766 (N_766,In_154,In_49);
nand U767 (N_767,In_111,In_432);
nor U768 (N_768,In_48,In_496);
nor U769 (N_769,In_306,In_387);
xor U770 (N_770,In_434,In_420);
nor U771 (N_771,In_285,In_177);
nand U772 (N_772,In_490,In_72);
nand U773 (N_773,In_221,In_36);
xnor U774 (N_774,In_122,In_79);
xnor U775 (N_775,In_309,In_219);
or U776 (N_776,In_495,In_106);
and U777 (N_777,In_234,In_418);
nand U778 (N_778,In_229,In_460);
xor U779 (N_779,In_160,In_464);
xor U780 (N_780,In_434,In_102);
and U781 (N_781,In_422,In_64);
xnor U782 (N_782,In_69,In_21);
or U783 (N_783,In_91,In_52);
xnor U784 (N_784,In_134,In_35);
and U785 (N_785,In_81,In_6);
nor U786 (N_786,In_192,In_179);
and U787 (N_787,In_139,In_326);
nand U788 (N_788,In_74,In_1);
nor U789 (N_789,In_101,In_350);
or U790 (N_790,In_481,In_177);
or U791 (N_791,In_104,In_266);
nand U792 (N_792,In_389,In_170);
xor U793 (N_793,In_372,In_275);
and U794 (N_794,In_56,In_26);
xor U795 (N_795,In_430,In_361);
or U796 (N_796,In_104,In_453);
nor U797 (N_797,In_183,In_94);
and U798 (N_798,In_121,In_101);
nor U799 (N_799,In_145,In_407);
and U800 (N_800,In_479,In_204);
nand U801 (N_801,In_273,In_348);
and U802 (N_802,In_185,In_239);
and U803 (N_803,In_497,In_99);
xor U804 (N_804,In_340,In_198);
nor U805 (N_805,In_344,In_166);
and U806 (N_806,In_232,In_164);
or U807 (N_807,In_17,In_182);
nand U808 (N_808,In_9,In_247);
nand U809 (N_809,In_33,In_202);
or U810 (N_810,In_329,In_431);
xor U811 (N_811,In_89,In_300);
and U812 (N_812,In_422,In_44);
nor U813 (N_813,In_296,In_236);
or U814 (N_814,In_115,In_460);
nor U815 (N_815,In_154,In_7);
nor U816 (N_816,In_452,In_165);
nand U817 (N_817,In_215,In_445);
and U818 (N_818,In_16,In_269);
nand U819 (N_819,In_145,In_69);
nand U820 (N_820,In_193,In_192);
and U821 (N_821,In_185,In_447);
and U822 (N_822,In_256,In_421);
or U823 (N_823,In_147,In_182);
nand U824 (N_824,In_276,In_265);
xnor U825 (N_825,In_252,In_99);
nand U826 (N_826,In_369,In_58);
nand U827 (N_827,In_298,In_184);
or U828 (N_828,In_362,In_324);
and U829 (N_829,In_325,In_364);
nor U830 (N_830,In_414,In_215);
and U831 (N_831,In_69,In_317);
xnor U832 (N_832,In_70,In_465);
or U833 (N_833,In_297,In_67);
and U834 (N_834,In_132,In_430);
nand U835 (N_835,In_290,In_267);
nor U836 (N_836,In_156,In_65);
nand U837 (N_837,In_425,In_79);
nor U838 (N_838,In_220,In_342);
and U839 (N_839,In_482,In_303);
xor U840 (N_840,In_172,In_233);
nand U841 (N_841,In_209,In_49);
and U842 (N_842,In_214,In_207);
and U843 (N_843,In_316,In_491);
xor U844 (N_844,In_141,In_361);
xnor U845 (N_845,In_89,In_231);
and U846 (N_846,In_429,In_32);
xnor U847 (N_847,In_91,In_155);
and U848 (N_848,In_28,In_289);
nand U849 (N_849,In_75,In_254);
and U850 (N_850,In_214,In_5);
nor U851 (N_851,In_195,In_71);
and U852 (N_852,In_325,In_188);
or U853 (N_853,In_193,In_433);
and U854 (N_854,In_22,In_70);
or U855 (N_855,In_39,In_311);
xnor U856 (N_856,In_19,In_27);
or U857 (N_857,In_332,In_102);
or U858 (N_858,In_384,In_213);
or U859 (N_859,In_137,In_141);
nor U860 (N_860,In_461,In_83);
nand U861 (N_861,In_341,In_421);
xnor U862 (N_862,In_20,In_190);
nor U863 (N_863,In_11,In_136);
xnor U864 (N_864,In_45,In_71);
xnor U865 (N_865,In_224,In_104);
or U866 (N_866,In_452,In_284);
xor U867 (N_867,In_51,In_301);
or U868 (N_868,In_250,In_73);
nor U869 (N_869,In_7,In_160);
xnor U870 (N_870,In_95,In_375);
nand U871 (N_871,In_210,In_291);
or U872 (N_872,In_492,In_441);
or U873 (N_873,In_65,In_475);
and U874 (N_874,In_60,In_198);
nand U875 (N_875,In_21,In_352);
and U876 (N_876,In_152,In_100);
xor U877 (N_877,In_298,In_252);
nand U878 (N_878,In_29,In_67);
nand U879 (N_879,In_222,In_239);
and U880 (N_880,In_81,In_386);
and U881 (N_881,In_318,In_192);
or U882 (N_882,In_20,In_58);
nor U883 (N_883,In_42,In_310);
nand U884 (N_884,In_233,In_469);
xnor U885 (N_885,In_39,In_391);
xnor U886 (N_886,In_196,In_163);
and U887 (N_887,In_291,In_349);
and U888 (N_888,In_208,In_151);
and U889 (N_889,In_200,In_257);
or U890 (N_890,In_139,In_89);
or U891 (N_891,In_305,In_403);
nor U892 (N_892,In_2,In_163);
nand U893 (N_893,In_319,In_208);
xor U894 (N_894,In_476,In_119);
or U895 (N_895,In_61,In_44);
or U896 (N_896,In_156,In_448);
nand U897 (N_897,In_319,In_362);
nand U898 (N_898,In_260,In_127);
xnor U899 (N_899,In_481,In_465);
nor U900 (N_900,In_452,In_273);
and U901 (N_901,In_375,In_286);
nor U902 (N_902,In_61,In_88);
nor U903 (N_903,In_339,In_199);
nand U904 (N_904,In_117,In_155);
nand U905 (N_905,In_244,In_121);
nor U906 (N_906,In_450,In_172);
and U907 (N_907,In_270,In_422);
xnor U908 (N_908,In_179,In_20);
xnor U909 (N_909,In_8,In_393);
nand U910 (N_910,In_476,In_424);
nand U911 (N_911,In_111,In_393);
or U912 (N_912,In_70,In_65);
nor U913 (N_913,In_25,In_464);
or U914 (N_914,In_408,In_253);
nor U915 (N_915,In_387,In_106);
nand U916 (N_916,In_56,In_73);
nand U917 (N_917,In_330,In_56);
and U918 (N_918,In_492,In_63);
and U919 (N_919,In_376,In_189);
xor U920 (N_920,In_228,In_384);
nor U921 (N_921,In_205,In_75);
xor U922 (N_922,In_1,In_349);
nor U923 (N_923,In_204,In_341);
or U924 (N_924,In_29,In_66);
nand U925 (N_925,In_55,In_84);
and U926 (N_926,In_74,In_221);
xnor U927 (N_927,In_127,In_129);
xor U928 (N_928,In_296,In_66);
nand U929 (N_929,In_372,In_289);
xor U930 (N_930,In_39,In_195);
nor U931 (N_931,In_185,In_246);
and U932 (N_932,In_112,In_317);
or U933 (N_933,In_88,In_181);
or U934 (N_934,In_393,In_280);
nand U935 (N_935,In_291,In_252);
and U936 (N_936,In_219,In_345);
or U937 (N_937,In_235,In_9);
nor U938 (N_938,In_117,In_390);
nor U939 (N_939,In_42,In_473);
and U940 (N_940,In_240,In_498);
xnor U941 (N_941,In_231,In_230);
nand U942 (N_942,In_60,In_298);
xnor U943 (N_943,In_226,In_330);
nand U944 (N_944,In_321,In_166);
and U945 (N_945,In_150,In_144);
nand U946 (N_946,In_29,In_398);
or U947 (N_947,In_43,In_448);
nor U948 (N_948,In_407,In_284);
xnor U949 (N_949,In_68,In_374);
nand U950 (N_950,In_283,In_455);
nor U951 (N_951,In_118,In_146);
nand U952 (N_952,In_176,In_153);
nand U953 (N_953,In_230,In_98);
nor U954 (N_954,In_302,In_207);
or U955 (N_955,In_169,In_4);
nand U956 (N_956,In_4,In_44);
nor U957 (N_957,In_217,In_158);
and U958 (N_958,In_73,In_243);
xor U959 (N_959,In_65,In_144);
or U960 (N_960,In_483,In_461);
nand U961 (N_961,In_17,In_223);
xnor U962 (N_962,In_444,In_175);
or U963 (N_963,In_53,In_445);
nand U964 (N_964,In_415,In_233);
nor U965 (N_965,In_249,In_328);
nor U966 (N_966,In_108,In_7);
xnor U967 (N_967,In_21,In_413);
nor U968 (N_968,In_251,In_372);
xnor U969 (N_969,In_395,In_16);
and U970 (N_970,In_483,In_19);
nand U971 (N_971,In_273,In_41);
and U972 (N_972,In_300,In_299);
and U973 (N_973,In_490,In_407);
xnor U974 (N_974,In_120,In_335);
xor U975 (N_975,In_113,In_14);
or U976 (N_976,In_482,In_241);
xnor U977 (N_977,In_443,In_17);
and U978 (N_978,In_466,In_100);
xor U979 (N_979,In_393,In_137);
and U980 (N_980,In_457,In_137);
and U981 (N_981,In_127,In_418);
or U982 (N_982,In_1,In_147);
xor U983 (N_983,In_250,In_366);
or U984 (N_984,In_244,In_354);
nor U985 (N_985,In_350,In_370);
nand U986 (N_986,In_123,In_183);
and U987 (N_987,In_287,In_134);
nand U988 (N_988,In_372,In_299);
xnor U989 (N_989,In_293,In_418);
and U990 (N_990,In_10,In_481);
nor U991 (N_991,In_452,In_389);
nor U992 (N_992,In_175,In_219);
nor U993 (N_993,In_239,In_336);
xnor U994 (N_994,In_490,In_212);
or U995 (N_995,In_378,In_411);
and U996 (N_996,In_129,In_437);
and U997 (N_997,In_376,In_155);
nor U998 (N_998,In_299,In_199);
or U999 (N_999,In_96,In_457);
xnor U1000 (N_1000,N_495,N_736);
nand U1001 (N_1001,N_774,N_571);
or U1002 (N_1002,N_458,N_218);
nor U1003 (N_1003,N_758,N_164);
xnor U1004 (N_1004,N_951,N_503);
or U1005 (N_1005,N_885,N_171);
and U1006 (N_1006,N_532,N_964);
nand U1007 (N_1007,N_611,N_589);
or U1008 (N_1008,N_80,N_876);
nand U1009 (N_1009,N_56,N_670);
xor U1010 (N_1010,N_497,N_804);
and U1011 (N_1011,N_788,N_903);
and U1012 (N_1012,N_666,N_916);
or U1013 (N_1013,N_309,N_721);
nor U1014 (N_1014,N_432,N_257);
nand U1015 (N_1015,N_368,N_239);
xnor U1016 (N_1016,N_592,N_905);
xnor U1017 (N_1017,N_699,N_891);
nor U1018 (N_1018,N_724,N_531);
or U1019 (N_1019,N_277,N_605);
nand U1020 (N_1020,N_601,N_476);
xor U1021 (N_1021,N_459,N_833);
or U1022 (N_1022,N_616,N_255);
and U1023 (N_1023,N_41,N_634);
xor U1024 (N_1024,N_513,N_940);
or U1025 (N_1025,N_379,N_273);
or U1026 (N_1026,N_682,N_490);
and U1027 (N_1027,N_930,N_545);
or U1028 (N_1028,N_895,N_477);
xor U1029 (N_1029,N_989,N_681);
nor U1030 (N_1030,N_92,N_374);
nand U1031 (N_1031,N_434,N_761);
or U1032 (N_1032,N_627,N_584);
xor U1033 (N_1033,N_506,N_159);
nand U1034 (N_1034,N_844,N_936);
xor U1035 (N_1035,N_677,N_34);
nor U1036 (N_1036,N_8,N_145);
or U1037 (N_1037,N_867,N_798);
or U1038 (N_1038,N_748,N_856);
nand U1039 (N_1039,N_829,N_566);
nand U1040 (N_1040,N_460,N_883);
nand U1041 (N_1041,N_600,N_962);
xor U1042 (N_1042,N_113,N_345);
and U1043 (N_1043,N_771,N_249);
nand U1044 (N_1044,N_69,N_384);
nand U1045 (N_1045,N_561,N_95);
xor U1046 (N_1046,N_609,N_737);
nor U1047 (N_1047,N_192,N_783);
or U1048 (N_1048,N_720,N_258);
nor U1049 (N_1049,N_117,N_908);
or U1050 (N_1050,N_24,N_728);
xnor U1051 (N_1051,N_517,N_295);
or U1052 (N_1052,N_94,N_990);
and U1053 (N_1053,N_684,N_168);
xor U1054 (N_1054,N_49,N_352);
nand U1055 (N_1055,N_158,N_410);
xnor U1056 (N_1056,N_195,N_147);
xor U1057 (N_1057,N_851,N_567);
and U1058 (N_1058,N_766,N_467);
nand U1059 (N_1059,N_418,N_734);
and U1060 (N_1060,N_902,N_57);
or U1061 (N_1061,N_583,N_852);
and U1062 (N_1062,N_603,N_128);
and U1063 (N_1063,N_144,N_645);
xnor U1064 (N_1064,N_123,N_698);
nand U1065 (N_1065,N_587,N_15);
xor U1066 (N_1066,N_875,N_568);
nor U1067 (N_1067,N_131,N_512);
or U1068 (N_1068,N_438,N_621);
or U1069 (N_1069,N_558,N_321);
and U1070 (N_1070,N_877,N_839);
nand U1071 (N_1071,N_719,N_780);
or U1072 (N_1072,N_840,N_188);
or U1073 (N_1073,N_140,N_620);
or U1074 (N_1074,N_918,N_400);
or U1075 (N_1075,N_527,N_61);
xnor U1076 (N_1076,N_830,N_557);
nand U1077 (N_1077,N_401,N_118);
xor U1078 (N_1078,N_360,N_661);
nand U1079 (N_1079,N_74,N_668);
nand U1080 (N_1080,N_626,N_900);
nor U1081 (N_1081,N_802,N_945);
xnor U1082 (N_1082,N_191,N_948);
nor U1083 (N_1083,N_484,N_493);
xor U1084 (N_1084,N_944,N_640);
nor U1085 (N_1085,N_283,N_546);
xnor U1086 (N_1086,N_970,N_959);
or U1087 (N_1087,N_664,N_404);
nor U1088 (N_1088,N_824,N_328);
and U1089 (N_1089,N_136,N_838);
xnor U1090 (N_1090,N_53,N_826);
nand U1091 (N_1091,N_955,N_949);
and U1092 (N_1092,N_845,N_542);
nand U1093 (N_1093,N_134,N_717);
or U1094 (N_1094,N_220,N_425);
nor U1095 (N_1095,N_86,N_831);
and U1096 (N_1096,N_124,N_373);
and U1097 (N_1097,N_262,N_937);
nor U1098 (N_1098,N_733,N_179);
xnor U1099 (N_1099,N_491,N_504);
nand U1100 (N_1100,N_577,N_770);
xor U1101 (N_1101,N_893,N_602);
and U1102 (N_1102,N_232,N_207);
and U1103 (N_1103,N_525,N_90);
or U1104 (N_1104,N_66,N_420);
xnor U1105 (N_1105,N_186,N_166);
nor U1106 (N_1106,N_597,N_173);
or U1107 (N_1107,N_246,N_11);
or U1108 (N_1108,N_977,N_644);
or U1109 (N_1109,N_399,N_789);
or U1110 (N_1110,N_863,N_254);
and U1111 (N_1111,N_496,N_860);
xor U1112 (N_1112,N_541,N_763);
xor U1113 (N_1113,N_806,N_339);
xnor U1114 (N_1114,N_377,N_746);
nand U1115 (N_1115,N_628,N_430);
nor U1116 (N_1116,N_884,N_827);
and U1117 (N_1117,N_242,N_1);
nor U1118 (N_1118,N_213,N_613);
nand U1119 (N_1119,N_755,N_472);
and U1120 (N_1120,N_350,N_271);
xnor U1121 (N_1121,N_966,N_741);
nand U1122 (N_1122,N_894,N_279);
nor U1123 (N_1123,N_22,N_904);
and U1124 (N_1124,N_615,N_501);
and U1125 (N_1125,N_396,N_642);
or U1126 (N_1126,N_554,N_729);
and U1127 (N_1127,N_853,N_198);
nand U1128 (N_1128,N_311,N_935);
nand U1129 (N_1129,N_578,N_610);
nor U1130 (N_1130,N_381,N_669);
nand U1131 (N_1131,N_227,N_530);
and U1132 (N_1132,N_565,N_727);
xnor U1133 (N_1133,N_992,N_837);
xor U1134 (N_1134,N_482,N_248);
or U1135 (N_1135,N_552,N_139);
and U1136 (N_1136,N_26,N_237);
nand U1137 (N_1137,N_285,N_890);
and U1138 (N_1138,N_362,N_375);
and U1139 (N_1139,N_222,N_141);
or U1140 (N_1140,N_658,N_45);
or U1141 (N_1141,N_920,N_585);
and U1142 (N_1142,N_292,N_97);
and U1143 (N_1143,N_161,N_330);
xor U1144 (N_1144,N_987,N_431);
and U1145 (N_1145,N_67,N_183);
nand U1146 (N_1146,N_991,N_533);
nor U1147 (N_1147,N_929,N_429);
xnor U1148 (N_1148,N_800,N_997);
or U1149 (N_1149,N_87,N_243);
or U1150 (N_1150,N_957,N_570);
nand U1151 (N_1151,N_986,N_457);
xnor U1152 (N_1152,N_214,N_960);
xor U1153 (N_1153,N_88,N_743);
or U1154 (N_1154,N_163,N_639);
and U1155 (N_1155,N_397,N_767);
and U1156 (N_1156,N_31,N_725);
or U1157 (N_1157,N_974,N_520);
nand U1158 (N_1158,N_849,N_581);
nand U1159 (N_1159,N_662,N_599);
nor U1160 (N_1160,N_760,N_641);
xor U1161 (N_1161,N_125,N_282);
nor U1162 (N_1162,N_363,N_126);
nand U1163 (N_1163,N_475,N_749);
and U1164 (N_1164,N_251,N_665);
and U1165 (N_1165,N_842,N_180);
or U1166 (N_1166,N_44,N_478);
nor U1167 (N_1167,N_96,N_809);
nand U1168 (N_1168,N_395,N_932);
and U1169 (N_1169,N_435,N_726);
or U1170 (N_1170,N_921,N_704);
nand U1171 (N_1171,N_33,N_596);
and U1172 (N_1172,N_209,N_101);
and U1173 (N_1173,N_151,N_83);
nor U1174 (N_1174,N_694,N_233);
xnor U1175 (N_1175,N_730,N_316);
or U1176 (N_1176,N_318,N_569);
nor U1177 (N_1177,N_102,N_127);
nand U1178 (N_1178,N_910,N_19);
or U1179 (N_1179,N_975,N_906);
xor U1180 (N_1180,N_494,N_693);
and U1181 (N_1181,N_518,N_836);
or U1182 (N_1182,N_408,N_288);
or U1183 (N_1183,N_414,N_355);
xnor U1184 (N_1184,N_388,N_701);
nand U1185 (N_1185,N_708,N_301);
or U1186 (N_1186,N_394,N_72);
and U1187 (N_1187,N_276,N_911);
or U1188 (N_1188,N_632,N_941);
nor U1189 (N_1189,N_857,N_866);
and U1190 (N_1190,N_331,N_286);
and U1191 (N_1191,N_17,N_290);
and U1192 (N_1192,N_865,N_73);
and U1193 (N_1193,N_712,N_353);
or U1194 (N_1194,N_441,N_190);
nand U1195 (N_1195,N_591,N_137);
or U1196 (N_1196,N_456,N_696);
xor U1197 (N_1197,N_415,N_750);
xor U1198 (N_1198,N_656,N_793);
xor U1199 (N_1199,N_272,N_998);
nand U1200 (N_1200,N_588,N_116);
or U1201 (N_1201,N_858,N_573);
xor U1202 (N_1202,N_773,N_357);
and U1203 (N_1203,N_98,N_341);
xnor U1204 (N_1204,N_796,N_108);
nand U1205 (N_1205,N_864,N_12);
nor U1206 (N_1206,N_466,N_489);
nand U1207 (N_1207,N_185,N_202);
nor U1208 (N_1208,N_488,N_419);
or U1209 (N_1209,N_580,N_46);
and U1210 (N_1210,N_486,N_203);
xnor U1211 (N_1211,N_535,N_818);
or U1212 (N_1212,N_556,N_988);
or U1213 (N_1213,N_953,N_236);
nand U1214 (N_1214,N_38,N_965);
nand U1215 (N_1215,N_71,N_739);
nor U1216 (N_1216,N_35,N_59);
nor U1217 (N_1217,N_536,N_336);
or U1218 (N_1218,N_607,N_91);
nand U1219 (N_1219,N_923,N_797);
and U1220 (N_1220,N_526,N_99);
nor U1221 (N_1221,N_688,N_174);
xnor U1222 (N_1222,N_176,N_927);
nand U1223 (N_1223,N_274,N_428);
and U1224 (N_1224,N_828,N_299);
nand U1225 (N_1225,N_332,N_383);
and U1226 (N_1226,N_514,N_454);
or U1227 (N_1227,N_700,N_560);
nand U1228 (N_1228,N_901,N_60);
nand U1229 (N_1229,N_643,N_846);
xor U1230 (N_1230,N_50,N_892);
xor U1231 (N_1231,N_424,N_452);
nand U1232 (N_1232,N_338,N_742);
nand U1233 (N_1233,N_317,N_82);
nand U1234 (N_1234,N_646,N_483);
nand U1235 (N_1235,N_64,N_740);
xnor U1236 (N_1236,N_914,N_834);
and U1237 (N_1237,N_764,N_691);
nand U1238 (N_1238,N_303,N_278);
nor U1239 (N_1239,N_954,N_300);
and U1240 (N_1240,N_722,N_4);
xor U1241 (N_1241,N_982,N_630);
xor U1242 (N_1242,N_551,N_337);
and U1243 (N_1243,N_680,N_356);
nor U1244 (N_1244,N_215,N_267);
or U1245 (N_1245,N_887,N_469);
and U1246 (N_1246,N_543,N_201);
nand U1247 (N_1247,N_983,N_412);
xor U1248 (N_1248,N_690,N_706);
xnor U1249 (N_1249,N_792,N_559);
xnor U1250 (N_1250,N_105,N_575);
xor U1251 (N_1251,N_859,N_847);
xor U1252 (N_1252,N_507,N_745);
nor U1253 (N_1253,N_405,N_407);
or U1254 (N_1254,N_385,N_651);
xnor U1255 (N_1255,N_816,N_9);
or U1256 (N_1256,N_241,N_463);
and U1257 (N_1257,N_178,N_505);
nand U1258 (N_1258,N_453,N_259);
nor U1259 (N_1259,N_121,N_473);
nor U1260 (N_1260,N_713,N_487);
xnor U1261 (N_1261,N_678,N_247);
or U1262 (N_1262,N_446,N_679);
or U1263 (N_1263,N_335,N_897);
or U1264 (N_1264,N_219,N_791);
nand U1265 (N_1265,N_814,N_122);
xor U1266 (N_1266,N_156,N_667);
xnor U1267 (N_1267,N_817,N_182);
nand U1268 (N_1268,N_305,N_206);
and U1269 (N_1269,N_62,N_112);
nor U1270 (N_1270,N_870,N_976);
xor U1271 (N_1271,N_735,N_2);
or U1272 (N_1272,N_996,N_785);
or U1273 (N_1273,N_302,N_969);
or U1274 (N_1274,N_75,N_896);
nor U1275 (N_1275,N_448,N_426);
and U1276 (N_1276,N_985,N_508);
or U1277 (N_1277,N_835,N_413);
and U1278 (N_1278,N_268,N_593);
nand U1279 (N_1279,N_820,N_617);
or U1280 (N_1280,N_406,N_703);
xor U1281 (N_1281,N_629,N_150);
or U1282 (N_1282,N_564,N_462);
and U1283 (N_1283,N_622,N_912);
and U1284 (N_1284,N_813,N_369);
nand U1285 (N_1285,N_440,N_398);
xor U1286 (N_1286,N_931,N_325);
nand U1287 (N_1287,N_114,N_380);
xor U1288 (N_1288,N_315,N_579);
nor U1289 (N_1289,N_909,N_153);
xor U1290 (N_1290,N_221,N_881);
xnor U1291 (N_1291,N_281,N_653);
and U1292 (N_1292,N_547,N_873);
and U1293 (N_1293,N_528,N_898);
nand U1294 (N_1294,N_880,N_657);
or U1295 (N_1295,N_275,N_784);
nor U1296 (N_1296,N_226,N_874);
or U1297 (N_1297,N_769,N_205);
nand U1298 (N_1298,N_386,N_808);
nor U1299 (N_1299,N_915,N_790);
nand U1300 (N_1300,N_324,N_138);
nor U1301 (N_1301,N_778,N_549);
nand U1302 (N_1302,N_815,N_170);
xor U1303 (N_1303,N_878,N_674);
and U1304 (N_1304,N_686,N_768);
or U1305 (N_1305,N_417,N_652);
and U1306 (N_1306,N_943,N_444);
nand U1307 (N_1307,N_42,N_794);
xnor U1308 (N_1308,N_157,N_821);
or U1309 (N_1309,N_200,N_421);
and U1310 (N_1310,N_994,N_172);
nand U1311 (N_1311,N_539,N_479);
and U1312 (N_1312,N_78,N_786);
or U1313 (N_1313,N_129,N_442);
and U1314 (N_1314,N_284,N_625);
xnor U1315 (N_1315,N_772,N_614);
xnor U1316 (N_1316,N_437,N_481);
and U1317 (N_1317,N_155,N_304);
xor U1318 (N_1318,N_582,N_624);
and U1319 (N_1319,N_20,N_346);
xnor U1320 (N_1320,N_294,N_744);
or U1321 (N_1321,N_54,N_225);
nor U1322 (N_1322,N_832,N_886);
xor U1323 (N_1323,N_208,N_608);
xnor U1324 (N_1324,N_104,N_216);
and U1325 (N_1325,N_590,N_563);
nor U1326 (N_1326,N_36,N_812);
or U1327 (N_1327,N_342,N_924);
xnor U1328 (N_1328,N_389,N_663);
nand U1329 (N_1329,N_650,N_862);
nand U1330 (N_1330,N_805,N_981);
or U1331 (N_1331,N_595,N_133);
and U1332 (N_1332,N_107,N_250);
and U1333 (N_1333,N_765,N_882);
nand U1334 (N_1334,N_572,N_963);
nand U1335 (N_1335,N_340,N_500);
or U1336 (N_1336,N_27,N_154);
or U1337 (N_1337,N_312,N_781);
or U1338 (N_1338,N_474,N_854);
or U1339 (N_1339,N_967,N_443);
or U1340 (N_1340,N_194,N_334);
or U1341 (N_1341,N_850,N_52);
nor U1342 (N_1342,N_197,N_55);
nor U1343 (N_1343,N_803,N_934);
xnor U1344 (N_1344,N_217,N_958);
nand U1345 (N_1345,N_320,N_752);
xnor U1346 (N_1346,N_30,N_451);
nand U1347 (N_1347,N_310,N_926);
and U1348 (N_1348,N_229,N_28);
and U1349 (N_1349,N_524,N_687);
or U1350 (N_1350,N_319,N_471);
nand U1351 (N_1351,N_499,N_636);
nor U1352 (N_1352,N_149,N_37);
xor U1353 (N_1353,N_939,N_747);
nand U1354 (N_1354,N_120,N_825);
and U1355 (N_1355,N_43,N_79);
and U1356 (N_1356,N_888,N_231);
nor U1357 (N_1357,N_58,N_868);
and U1358 (N_1358,N_439,N_106);
nor U1359 (N_1359,N_979,N_252);
and U1360 (N_1360,N_461,N_754);
nand U1361 (N_1361,N_184,N_757);
or U1362 (N_1362,N_177,N_409);
or U1363 (N_1363,N_638,N_390);
or U1364 (N_1364,N_907,N_972);
or U1365 (N_1365,N_210,N_899);
or U1366 (N_1366,N_296,N_775);
nor U1367 (N_1367,N_685,N_671);
nor U1368 (N_1368,N_841,N_348);
nor U1369 (N_1369,N_77,N_928);
nand U1370 (N_1370,N_598,N_152);
nand U1371 (N_1371,N_553,N_253);
nand U1372 (N_1372,N_287,N_879);
nor U1373 (N_1373,N_869,N_485);
and U1374 (N_1374,N_81,N_423);
nand U1375 (N_1375,N_995,N_63);
nand U1376 (N_1376,N_692,N_509);
and U1377 (N_1377,N_673,N_984);
nand U1378 (N_1378,N_25,N_498);
xor U1379 (N_1379,N_973,N_952);
nor U1380 (N_1380,N_689,N_40);
xnor U1381 (N_1381,N_978,N_606);
xor U1382 (N_1382,N_297,N_85);
or U1383 (N_1383,N_354,N_619);
or U1384 (N_1384,N_540,N_212);
or U1385 (N_1385,N_371,N_811);
nand U1386 (N_1386,N_807,N_445);
nor U1387 (N_1387,N_515,N_810);
or U1388 (N_1388,N_5,N_779);
nor U1389 (N_1389,N_801,N_110);
or U1390 (N_1390,N_672,N_387);
xor U1391 (N_1391,N_326,N_84);
nor U1392 (N_1392,N_534,N_544);
nor U1393 (N_1393,N_234,N_710);
and U1394 (N_1394,N_89,N_738);
xnor U1395 (N_1395,N_649,N_65);
nor U1396 (N_1396,N_366,N_705);
nor U1397 (N_1397,N_211,N_162);
nor U1398 (N_1398,N_942,N_871);
and U1399 (N_1399,N_364,N_165);
nor U1400 (N_1400,N_416,N_464);
nand U1401 (N_1401,N_100,N_917);
xnor U1402 (N_1402,N_47,N_576);
and U1403 (N_1403,N_29,N_269);
and U1404 (N_1404,N_470,N_130);
and U1405 (N_1405,N_822,N_391);
xor U1406 (N_1406,N_999,N_289);
or U1407 (N_1407,N_16,N_716);
xor U1408 (N_1408,N_313,N_298);
nor U1409 (N_1409,N_510,N_968);
nor U1410 (N_1410,N_68,N_925);
nand U1411 (N_1411,N_633,N_13);
nor U1412 (N_1412,N_612,N_635);
xnor U1413 (N_1413,N_648,N_922);
xor U1414 (N_1414,N_433,N_245);
nor U1415 (N_1415,N_683,N_93);
xor U1416 (N_1416,N_76,N_146);
xnor U1417 (N_1417,N_715,N_18);
or U1418 (N_1418,N_538,N_115);
and U1419 (N_1419,N_946,N_14);
xor U1420 (N_1420,N_148,N_956);
nor U1421 (N_1421,N_261,N_230);
xor U1422 (N_1422,N_266,N_280);
nor U1423 (N_1423,N_23,N_32);
xnor U1424 (N_1424,N_732,N_109);
nor U1425 (N_1425,N_731,N_293);
xnor U1426 (N_1426,N_502,N_586);
xor U1427 (N_1427,N_187,N_776);
nand U1428 (N_1428,N_919,N_529);
xor U1429 (N_1429,N_135,N_327);
nor U1430 (N_1430,N_223,N_160);
or U1431 (N_1431,N_333,N_306);
nor U1432 (N_1432,N_378,N_594);
nand U1433 (N_1433,N_235,N_132);
nor U1434 (N_1434,N_143,N_753);
nand U1435 (N_1435,N_971,N_181);
xor U1436 (N_1436,N_468,N_308);
and U1437 (N_1437,N_455,N_10);
nand U1438 (N_1438,N_6,N_711);
or U1439 (N_1439,N_376,N_933);
and U1440 (N_1440,N_695,N_392);
and U1441 (N_1441,N_861,N_167);
and U1442 (N_1442,N_823,N_659);
nor U1443 (N_1443,N_938,N_193);
and U1444 (N_1444,N_655,N_782);
xor U1445 (N_1445,N_950,N_993);
and U1446 (N_1446,N_411,N_343);
or U1447 (N_1447,N_367,N_307);
and U1448 (N_1448,N_361,N_169);
and U1449 (N_1449,N_228,N_522);
nor U1450 (N_1450,N_647,N_344);
and U1451 (N_1451,N_224,N_119);
nor U1452 (N_1452,N_372,N_359);
or U1453 (N_1453,N_855,N_51);
xnor U1454 (N_1454,N_48,N_323);
xnor U1455 (N_1455,N_0,N_365);
nand U1456 (N_1456,N_947,N_393);
or U1457 (N_1457,N_702,N_492);
nor U1458 (N_1458,N_175,N_263);
and U1459 (N_1459,N_604,N_3);
and U1460 (N_1460,N_872,N_260);
nor U1461 (N_1461,N_777,N_819);
xor U1462 (N_1462,N_21,N_618);
and U1463 (N_1463,N_189,N_382);
xnor U1464 (N_1464,N_322,N_521);
or U1465 (N_1465,N_291,N_799);
nand U1466 (N_1466,N_270,N_519);
nand U1467 (N_1467,N_631,N_111);
nand U1468 (N_1468,N_103,N_70);
xnor U1469 (N_1469,N_244,N_714);
and U1470 (N_1470,N_351,N_436);
nor U1471 (N_1471,N_759,N_913);
or U1472 (N_1472,N_265,N_349);
nand U1473 (N_1473,N_562,N_654);
nor U1474 (N_1474,N_718,N_196);
xnor U1475 (N_1475,N_422,N_675);
nor U1476 (N_1476,N_403,N_548);
nand U1477 (N_1477,N_795,N_848);
xor U1478 (N_1478,N_142,N_204);
and U1479 (N_1479,N_555,N_980);
and U1480 (N_1480,N_756,N_427);
xnor U1481 (N_1481,N_39,N_709);
nand U1482 (N_1482,N_537,N_402);
nand U1483 (N_1483,N_329,N_843);
nand U1484 (N_1484,N_370,N_314);
xor U1485 (N_1485,N_623,N_7);
xor U1486 (N_1486,N_358,N_762);
and U1487 (N_1487,N_511,N_465);
or U1488 (N_1488,N_961,N_723);
or U1489 (N_1489,N_240,N_707);
and U1490 (N_1490,N_676,N_480);
nand U1491 (N_1491,N_660,N_637);
nand U1492 (N_1492,N_199,N_264);
nand U1493 (N_1493,N_697,N_450);
or U1494 (N_1494,N_889,N_523);
and U1495 (N_1495,N_516,N_347);
nor U1496 (N_1496,N_238,N_449);
nor U1497 (N_1497,N_751,N_550);
and U1498 (N_1498,N_787,N_574);
nor U1499 (N_1499,N_256,N_447);
or U1500 (N_1500,N_610,N_552);
xor U1501 (N_1501,N_579,N_2);
xor U1502 (N_1502,N_328,N_921);
nor U1503 (N_1503,N_483,N_575);
nor U1504 (N_1504,N_13,N_384);
xor U1505 (N_1505,N_583,N_913);
and U1506 (N_1506,N_580,N_934);
or U1507 (N_1507,N_690,N_797);
nor U1508 (N_1508,N_678,N_450);
nor U1509 (N_1509,N_692,N_987);
and U1510 (N_1510,N_146,N_427);
or U1511 (N_1511,N_608,N_712);
xor U1512 (N_1512,N_633,N_380);
and U1513 (N_1513,N_938,N_509);
nand U1514 (N_1514,N_188,N_971);
xor U1515 (N_1515,N_509,N_762);
nand U1516 (N_1516,N_100,N_570);
and U1517 (N_1517,N_80,N_669);
or U1518 (N_1518,N_731,N_498);
xor U1519 (N_1519,N_182,N_883);
or U1520 (N_1520,N_754,N_364);
and U1521 (N_1521,N_293,N_381);
or U1522 (N_1522,N_664,N_952);
and U1523 (N_1523,N_186,N_576);
and U1524 (N_1524,N_26,N_148);
and U1525 (N_1525,N_174,N_179);
or U1526 (N_1526,N_451,N_73);
nand U1527 (N_1527,N_711,N_166);
xnor U1528 (N_1528,N_818,N_404);
and U1529 (N_1529,N_223,N_247);
nand U1530 (N_1530,N_938,N_847);
nand U1531 (N_1531,N_587,N_820);
nand U1532 (N_1532,N_92,N_421);
or U1533 (N_1533,N_982,N_513);
and U1534 (N_1534,N_625,N_866);
xor U1535 (N_1535,N_981,N_22);
xor U1536 (N_1536,N_239,N_874);
xnor U1537 (N_1537,N_171,N_496);
xor U1538 (N_1538,N_822,N_847);
or U1539 (N_1539,N_772,N_196);
xor U1540 (N_1540,N_936,N_379);
nand U1541 (N_1541,N_618,N_815);
or U1542 (N_1542,N_669,N_384);
nor U1543 (N_1543,N_171,N_839);
and U1544 (N_1544,N_50,N_878);
nand U1545 (N_1545,N_942,N_60);
nor U1546 (N_1546,N_912,N_988);
or U1547 (N_1547,N_419,N_225);
xor U1548 (N_1548,N_613,N_43);
xnor U1549 (N_1549,N_435,N_599);
nor U1550 (N_1550,N_577,N_978);
nor U1551 (N_1551,N_97,N_499);
xor U1552 (N_1552,N_300,N_915);
nand U1553 (N_1553,N_597,N_126);
nand U1554 (N_1554,N_526,N_967);
or U1555 (N_1555,N_39,N_412);
nand U1556 (N_1556,N_66,N_269);
xor U1557 (N_1557,N_39,N_241);
xnor U1558 (N_1558,N_976,N_299);
nor U1559 (N_1559,N_85,N_806);
or U1560 (N_1560,N_197,N_427);
and U1561 (N_1561,N_236,N_119);
xnor U1562 (N_1562,N_93,N_959);
nand U1563 (N_1563,N_316,N_212);
xor U1564 (N_1564,N_569,N_365);
or U1565 (N_1565,N_276,N_625);
nor U1566 (N_1566,N_154,N_462);
and U1567 (N_1567,N_621,N_222);
or U1568 (N_1568,N_764,N_965);
or U1569 (N_1569,N_631,N_644);
nor U1570 (N_1570,N_549,N_11);
and U1571 (N_1571,N_812,N_849);
and U1572 (N_1572,N_701,N_820);
or U1573 (N_1573,N_187,N_936);
or U1574 (N_1574,N_93,N_867);
xor U1575 (N_1575,N_697,N_734);
nand U1576 (N_1576,N_704,N_270);
and U1577 (N_1577,N_353,N_922);
nand U1578 (N_1578,N_567,N_369);
nor U1579 (N_1579,N_679,N_27);
nand U1580 (N_1580,N_696,N_298);
nor U1581 (N_1581,N_961,N_262);
and U1582 (N_1582,N_550,N_695);
xor U1583 (N_1583,N_0,N_50);
nor U1584 (N_1584,N_893,N_695);
nor U1585 (N_1585,N_114,N_204);
xor U1586 (N_1586,N_146,N_787);
or U1587 (N_1587,N_829,N_86);
and U1588 (N_1588,N_296,N_30);
and U1589 (N_1589,N_308,N_546);
nand U1590 (N_1590,N_487,N_74);
xor U1591 (N_1591,N_695,N_97);
nor U1592 (N_1592,N_612,N_252);
nand U1593 (N_1593,N_45,N_918);
nor U1594 (N_1594,N_821,N_623);
xor U1595 (N_1595,N_421,N_1);
and U1596 (N_1596,N_641,N_42);
or U1597 (N_1597,N_826,N_635);
and U1598 (N_1598,N_95,N_773);
nand U1599 (N_1599,N_18,N_904);
xor U1600 (N_1600,N_256,N_250);
and U1601 (N_1601,N_251,N_150);
nor U1602 (N_1602,N_31,N_782);
nand U1603 (N_1603,N_141,N_400);
xor U1604 (N_1604,N_139,N_842);
or U1605 (N_1605,N_844,N_442);
or U1606 (N_1606,N_510,N_27);
nor U1607 (N_1607,N_363,N_819);
nand U1608 (N_1608,N_321,N_548);
nor U1609 (N_1609,N_495,N_348);
and U1610 (N_1610,N_523,N_893);
nand U1611 (N_1611,N_387,N_29);
and U1612 (N_1612,N_19,N_545);
xnor U1613 (N_1613,N_657,N_345);
or U1614 (N_1614,N_518,N_478);
nand U1615 (N_1615,N_430,N_618);
or U1616 (N_1616,N_313,N_379);
nor U1617 (N_1617,N_768,N_186);
nor U1618 (N_1618,N_3,N_721);
xnor U1619 (N_1619,N_526,N_587);
or U1620 (N_1620,N_986,N_72);
nand U1621 (N_1621,N_363,N_477);
nand U1622 (N_1622,N_725,N_194);
or U1623 (N_1623,N_57,N_803);
nor U1624 (N_1624,N_462,N_108);
nand U1625 (N_1625,N_840,N_566);
nor U1626 (N_1626,N_112,N_174);
nand U1627 (N_1627,N_261,N_898);
and U1628 (N_1628,N_783,N_89);
nand U1629 (N_1629,N_486,N_817);
nand U1630 (N_1630,N_244,N_96);
xnor U1631 (N_1631,N_440,N_190);
nor U1632 (N_1632,N_724,N_120);
or U1633 (N_1633,N_515,N_559);
nor U1634 (N_1634,N_522,N_781);
xnor U1635 (N_1635,N_535,N_113);
and U1636 (N_1636,N_187,N_503);
nor U1637 (N_1637,N_395,N_54);
nor U1638 (N_1638,N_987,N_142);
nand U1639 (N_1639,N_623,N_234);
or U1640 (N_1640,N_495,N_173);
and U1641 (N_1641,N_606,N_930);
or U1642 (N_1642,N_509,N_145);
and U1643 (N_1643,N_279,N_620);
nor U1644 (N_1644,N_40,N_366);
and U1645 (N_1645,N_485,N_404);
nor U1646 (N_1646,N_152,N_440);
xnor U1647 (N_1647,N_373,N_238);
or U1648 (N_1648,N_685,N_629);
nand U1649 (N_1649,N_259,N_812);
and U1650 (N_1650,N_735,N_259);
nand U1651 (N_1651,N_333,N_537);
nand U1652 (N_1652,N_138,N_78);
nor U1653 (N_1653,N_13,N_586);
and U1654 (N_1654,N_187,N_569);
nor U1655 (N_1655,N_513,N_404);
and U1656 (N_1656,N_969,N_378);
nand U1657 (N_1657,N_802,N_271);
nand U1658 (N_1658,N_704,N_447);
nand U1659 (N_1659,N_338,N_918);
nand U1660 (N_1660,N_139,N_157);
and U1661 (N_1661,N_49,N_120);
nand U1662 (N_1662,N_202,N_959);
or U1663 (N_1663,N_75,N_32);
nor U1664 (N_1664,N_111,N_650);
or U1665 (N_1665,N_522,N_907);
nand U1666 (N_1666,N_612,N_86);
xor U1667 (N_1667,N_760,N_632);
xnor U1668 (N_1668,N_286,N_926);
or U1669 (N_1669,N_827,N_54);
nand U1670 (N_1670,N_381,N_646);
or U1671 (N_1671,N_138,N_39);
nand U1672 (N_1672,N_485,N_637);
and U1673 (N_1673,N_332,N_219);
or U1674 (N_1674,N_783,N_222);
or U1675 (N_1675,N_20,N_587);
nand U1676 (N_1676,N_280,N_102);
xnor U1677 (N_1677,N_551,N_126);
nand U1678 (N_1678,N_754,N_745);
nand U1679 (N_1679,N_884,N_283);
nand U1680 (N_1680,N_175,N_909);
xnor U1681 (N_1681,N_817,N_489);
or U1682 (N_1682,N_894,N_736);
or U1683 (N_1683,N_389,N_215);
and U1684 (N_1684,N_249,N_304);
and U1685 (N_1685,N_957,N_815);
and U1686 (N_1686,N_267,N_184);
xor U1687 (N_1687,N_347,N_436);
nor U1688 (N_1688,N_257,N_293);
nand U1689 (N_1689,N_924,N_632);
nand U1690 (N_1690,N_138,N_876);
nor U1691 (N_1691,N_801,N_61);
and U1692 (N_1692,N_708,N_299);
nor U1693 (N_1693,N_232,N_30);
nor U1694 (N_1694,N_723,N_410);
and U1695 (N_1695,N_42,N_928);
or U1696 (N_1696,N_125,N_151);
and U1697 (N_1697,N_683,N_988);
xnor U1698 (N_1698,N_241,N_439);
xor U1699 (N_1699,N_501,N_18);
nor U1700 (N_1700,N_200,N_970);
nand U1701 (N_1701,N_297,N_663);
nand U1702 (N_1702,N_845,N_951);
nor U1703 (N_1703,N_362,N_865);
xnor U1704 (N_1704,N_774,N_715);
and U1705 (N_1705,N_934,N_58);
or U1706 (N_1706,N_823,N_391);
or U1707 (N_1707,N_134,N_928);
nor U1708 (N_1708,N_645,N_553);
nor U1709 (N_1709,N_494,N_295);
nand U1710 (N_1710,N_826,N_581);
xnor U1711 (N_1711,N_240,N_658);
nand U1712 (N_1712,N_345,N_797);
xor U1713 (N_1713,N_419,N_640);
nor U1714 (N_1714,N_913,N_742);
and U1715 (N_1715,N_958,N_302);
nand U1716 (N_1716,N_468,N_298);
and U1717 (N_1717,N_984,N_148);
nor U1718 (N_1718,N_602,N_367);
nand U1719 (N_1719,N_717,N_188);
nor U1720 (N_1720,N_133,N_159);
nand U1721 (N_1721,N_923,N_281);
or U1722 (N_1722,N_209,N_896);
nand U1723 (N_1723,N_960,N_380);
nor U1724 (N_1724,N_843,N_140);
and U1725 (N_1725,N_584,N_527);
nor U1726 (N_1726,N_747,N_443);
and U1727 (N_1727,N_464,N_249);
and U1728 (N_1728,N_909,N_806);
xor U1729 (N_1729,N_546,N_745);
and U1730 (N_1730,N_833,N_162);
nor U1731 (N_1731,N_650,N_914);
and U1732 (N_1732,N_464,N_949);
nand U1733 (N_1733,N_440,N_28);
and U1734 (N_1734,N_368,N_397);
or U1735 (N_1735,N_631,N_832);
nor U1736 (N_1736,N_332,N_756);
nor U1737 (N_1737,N_174,N_927);
and U1738 (N_1738,N_715,N_698);
or U1739 (N_1739,N_343,N_423);
or U1740 (N_1740,N_140,N_785);
and U1741 (N_1741,N_122,N_936);
or U1742 (N_1742,N_74,N_876);
or U1743 (N_1743,N_947,N_664);
nand U1744 (N_1744,N_17,N_20);
nand U1745 (N_1745,N_113,N_692);
or U1746 (N_1746,N_22,N_535);
nand U1747 (N_1747,N_60,N_777);
xor U1748 (N_1748,N_173,N_371);
or U1749 (N_1749,N_958,N_879);
or U1750 (N_1750,N_815,N_921);
nand U1751 (N_1751,N_298,N_384);
nand U1752 (N_1752,N_87,N_527);
xor U1753 (N_1753,N_753,N_947);
or U1754 (N_1754,N_183,N_806);
and U1755 (N_1755,N_998,N_180);
or U1756 (N_1756,N_62,N_290);
xnor U1757 (N_1757,N_635,N_906);
nand U1758 (N_1758,N_481,N_462);
nand U1759 (N_1759,N_607,N_735);
and U1760 (N_1760,N_801,N_574);
nor U1761 (N_1761,N_348,N_837);
and U1762 (N_1762,N_27,N_702);
nor U1763 (N_1763,N_692,N_138);
xor U1764 (N_1764,N_53,N_240);
nand U1765 (N_1765,N_695,N_348);
or U1766 (N_1766,N_185,N_799);
nor U1767 (N_1767,N_605,N_589);
and U1768 (N_1768,N_886,N_468);
nand U1769 (N_1769,N_852,N_664);
and U1770 (N_1770,N_415,N_595);
xnor U1771 (N_1771,N_952,N_200);
xor U1772 (N_1772,N_118,N_965);
nor U1773 (N_1773,N_705,N_92);
and U1774 (N_1774,N_539,N_401);
or U1775 (N_1775,N_903,N_332);
nor U1776 (N_1776,N_385,N_675);
or U1777 (N_1777,N_279,N_84);
xor U1778 (N_1778,N_560,N_141);
nand U1779 (N_1779,N_78,N_882);
nand U1780 (N_1780,N_437,N_250);
and U1781 (N_1781,N_446,N_904);
nor U1782 (N_1782,N_908,N_102);
nand U1783 (N_1783,N_483,N_389);
nand U1784 (N_1784,N_897,N_46);
nor U1785 (N_1785,N_874,N_449);
xnor U1786 (N_1786,N_435,N_835);
nand U1787 (N_1787,N_802,N_640);
and U1788 (N_1788,N_571,N_2);
or U1789 (N_1789,N_512,N_41);
nor U1790 (N_1790,N_539,N_474);
nand U1791 (N_1791,N_112,N_848);
nand U1792 (N_1792,N_355,N_586);
nand U1793 (N_1793,N_204,N_418);
nor U1794 (N_1794,N_510,N_279);
xnor U1795 (N_1795,N_568,N_855);
nand U1796 (N_1796,N_647,N_436);
and U1797 (N_1797,N_859,N_910);
xor U1798 (N_1798,N_794,N_839);
or U1799 (N_1799,N_309,N_941);
nand U1800 (N_1800,N_747,N_212);
and U1801 (N_1801,N_937,N_669);
and U1802 (N_1802,N_589,N_245);
nor U1803 (N_1803,N_101,N_393);
or U1804 (N_1804,N_631,N_686);
nand U1805 (N_1805,N_190,N_963);
xor U1806 (N_1806,N_795,N_127);
and U1807 (N_1807,N_321,N_255);
nor U1808 (N_1808,N_725,N_79);
or U1809 (N_1809,N_327,N_447);
and U1810 (N_1810,N_899,N_879);
nand U1811 (N_1811,N_100,N_979);
or U1812 (N_1812,N_233,N_662);
nand U1813 (N_1813,N_347,N_317);
nand U1814 (N_1814,N_38,N_589);
nand U1815 (N_1815,N_439,N_445);
nand U1816 (N_1816,N_220,N_404);
or U1817 (N_1817,N_792,N_325);
nand U1818 (N_1818,N_959,N_972);
xor U1819 (N_1819,N_251,N_529);
nor U1820 (N_1820,N_514,N_199);
nand U1821 (N_1821,N_254,N_394);
nor U1822 (N_1822,N_402,N_243);
xnor U1823 (N_1823,N_57,N_752);
or U1824 (N_1824,N_819,N_263);
or U1825 (N_1825,N_482,N_570);
nor U1826 (N_1826,N_166,N_400);
or U1827 (N_1827,N_895,N_843);
nand U1828 (N_1828,N_338,N_824);
and U1829 (N_1829,N_775,N_908);
or U1830 (N_1830,N_583,N_882);
or U1831 (N_1831,N_547,N_199);
or U1832 (N_1832,N_346,N_311);
nor U1833 (N_1833,N_483,N_591);
nand U1834 (N_1834,N_755,N_25);
and U1835 (N_1835,N_883,N_238);
xor U1836 (N_1836,N_259,N_884);
xnor U1837 (N_1837,N_166,N_971);
nor U1838 (N_1838,N_366,N_860);
and U1839 (N_1839,N_414,N_679);
nor U1840 (N_1840,N_631,N_768);
xor U1841 (N_1841,N_395,N_946);
nand U1842 (N_1842,N_283,N_191);
or U1843 (N_1843,N_617,N_537);
nand U1844 (N_1844,N_479,N_167);
xnor U1845 (N_1845,N_939,N_190);
nand U1846 (N_1846,N_773,N_336);
xnor U1847 (N_1847,N_350,N_419);
and U1848 (N_1848,N_135,N_315);
and U1849 (N_1849,N_345,N_950);
and U1850 (N_1850,N_843,N_966);
xor U1851 (N_1851,N_571,N_196);
and U1852 (N_1852,N_350,N_314);
or U1853 (N_1853,N_713,N_796);
nor U1854 (N_1854,N_979,N_755);
nor U1855 (N_1855,N_455,N_959);
and U1856 (N_1856,N_549,N_968);
nand U1857 (N_1857,N_808,N_380);
and U1858 (N_1858,N_979,N_233);
xor U1859 (N_1859,N_716,N_524);
and U1860 (N_1860,N_968,N_908);
and U1861 (N_1861,N_128,N_19);
or U1862 (N_1862,N_538,N_219);
or U1863 (N_1863,N_158,N_572);
or U1864 (N_1864,N_521,N_535);
and U1865 (N_1865,N_351,N_350);
or U1866 (N_1866,N_750,N_343);
or U1867 (N_1867,N_385,N_149);
and U1868 (N_1868,N_74,N_390);
and U1869 (N_1869,N_760,N_947);
and U1870 (N_1870,N_221,N_549);
and U1871 (N_1871,N_721,N_636);
nand U1872 (N_1872,N_176,N_937);
xnor U1873 (N_1873,N_384,N_664);
xor U1874 (N_1874,N_425,N_390);
nand U1875 (N_1875,N_273,N_929);
nor U1876 (N_1876,N_885,N_344);
nand U1877 (N_1877,N_379,N_626);
or U1878 (N_1878,N_228,N_818);
or U1879 (N_1879,N_286,N_656);
nand U1880 (N_1880,N_767,N_679);
and U1881 (N_1881,N_502,N_279);
and U1882 (N_1882,N_294,N_678);
xnor U1883 (N_1883,N_770,N_776);
nor U1884 (N_1884,N_234,N_295);
nor U1885 (N_1885,N_477,N_64);
xor U1886 (N_1886,N_838,N_76);
nor U1887 (N_1887,N_944,N_135);
or U1888 (N_1888,N_84,N_330);
or U1889 (N_1889,N_805,N_722);
nand U1890 (N_1890,N_353,N_122);
nor U1891 (N_1891,N_97,N_802);
nand U1892 (N_1892,N_678,N_732);
nand U1893 (N_1893,N_918,N_654);
nand U1894 (N_1894,N_930,N_565);
nor U1895 (N_1895,N_879,N_272);
xor U1896 (N_1896,N_545,N_793);
or U1897 (N_1897,N_539,N_73);
or U1898 (N_1898,N_161,N_750);
and U1899 (N_1899,N_939,N_115);
or U1900 (N_1900,N_904,N_510);
nor U1901 (N_1901,N_223,N_320);
xor U1902 (N_1902,N_28,N_953);
nand U1903 (N_1903,N_564,N_305);
and U1904 (N_1904,N_842,N_602);
xnor U1905 (N_1905,N_45,N_617);
or U1906 (N_1906,N_460,N_786);
nor U1907 (N_1907,N_310,N_306);
and U1908 (N_1908,N_701,N_550);
nand U1909 (N_1909,N_658,N_884);
xor U1910 (N_1910,N_415,N_936);
xnor U1911 (N_1911,N_640,N_963);
xnor U1912 (N_1912,N_799,N_924);
nor U1913 (N_1913,N_178,N_257);
and U1914 (N_1914,N_669,N_70);
or U1915 (N_1915,N_992,N_54);
or U1916 (N_1916,N_375,N_310);
or U1917 (N_1917,N_798,N_546);
and U1918 (N_1918,N_708,N_856);
or U1919 (N_1919,N_553,N_876);
nand U1920 (N_1920,N_583,N_607);
nand U1921 (N_1921,N_872,N_309);
nor U1922 (N_1922,N_295,N_886);
xnor U1923 (N_1923,N_374,N_698);
nor U1924 (N_1924,N_541,N_419);
or U1925 (N_1925,N_652,N_725);
and U1926 (N_1926,N_743,N_516);
nand U1927 (N_1927,N_636,N_230);
nor U1928 (N_1928,N_882,N_347);
or U1929 (N_1929,N_348,N_674);
xor U1930 (N_1930,N_257,N_188);
xor U1931 (N_1931,N_656,N_230);
and U1932 (N_1932,N_360,N_677);
and U1933 (N_1933,N_910,N_294);
or U1934 (N_1934,N_562,N_387);
xnor U1935 (N_1935,N_669,N_37);
nor U1936 (N_1936,N_213,N_905);
xnor U1937 (N_1937,N_30,N_649);
nand U1938 (N_1938,N_2,N_438);
or U1939 (N_1939,N_74,N_679);
nand U1940 (N_1940,N_487,N_669);
or U1941 (N_1941,N_639,N_840);
or U1942 (N_1942,N_739,N_578);
nor U1943 (N_1943,N_615,N_786);
and U1944 (N_1944,N_102,N_612);
nand U1945 (N_1945,N_860,N_839);
and U1946 (N_1946,N_825,N_711);
or U1947 (N_1947,N_33,N_897);
xor U1948 (N_1948,N_150,N_709);
nand U1949 (N_1949,N_250,N_374);
or U1950 (N_1950,N_866,N_889);
xor U1951 (N_1951,N_615,N_209);
and U1952 (N_1952,N_682,N_70);
and U1953 (N_1953,N_426,N_133);
xor U1954 (N_1954,N_702,N_2);
nand U1955 (N_1955,N_225,N_499);
xor U1956 (N_1956,N_834,N_405);
xnor U1957 (N_1957,N_6,N_284);
or U1958 (N_1958,N_983,N_909);
xor U1959 (N_1959,N_954,N_447);
and U1960 (N_1960,N_86,N_660);
nor U1961 (N_1961,N_473,N_216);
nor U1962 (N_1962,N_390,N_534);
or U1963 (N_1963,N_380,N_66);
nor U1964 (N_1964,N_884,N_233);
nor U1965 (N_1965,N_823,N_541);
nand U1966 (N_1966,N_287,N_643);
nor U1967 (N_1967,N_984,N_797);
nor U1968 (N_1968,N_78,N_899);
or U1969 (N_1969,N_245,N_73);
or U1970 (N_1970,N_143,N_516);
xor U1971 (N_1971,N_652,N_280);
or U1972 (N_1972,N_332,N_556);
and U1973 (N_1973,N_544,N_514);
xor U1974 (N_1974,N_793,N_945);
xnor U1975 (N_1975,N_664,N_437);
and U1976 (N_1976,N_409,N_513);
or U1977 (N_1977,N_846,N_765);
nor U1978 (N_1978,N_605,N_340);
nand U1979 (N_1979,N_470,N_99);
nor U1980 (N_1980,N_80,N_792);
or U1981 (N_1981,N_891,N_963);
xor U1982 (N_1982,N_511,N_66);
xor U1983 (N_1983,N_549,N_817);
nor U1984 (N_1984,N_338,N_253);
or U1985 (N_1985,N_929,N_123);
or U1986 (N_1986,N_103,N_964);
nand U1987 (N_1987,N_107,N_745);
xor U1988 (N_1988,N_238,N_537);
and U1989 (N_1989,N_695,N_56);
nor U1990 (N_1990,N_949,N_401);
and U1991 (N_1991,N_720,N_468);
xnor U1992 (N_1992,N_312,N_161);
and U1993 (N_1993,N_871,N_859);
nand U1994 (N_1994,N_374,N_301);
and U1995 (N_1995,N_117,N_225);
xor U1996 (N_1996,N_10,N_327);
nor U1997 (N_1997,N_970,N_955);
nand U1998 (N_1998,N_150,N_504);
nor U1999 (N_1999,N_655,N_79);
or U2000 (N_2000,N_1549,N_1780);
nor U2001 (N_2001,N_1828,N_1504);
or U2002 (N_2002,N_1756,N_1318);
nand U2003 (N_2003,N_1604,N_1298);
or U2004 (N_2004,N_1147,N_1131);
nor U2005 (N_2005,N_1000,N_1190);
and U2006 (N_2006,N_1117,N_1309);
or U2007 (N_2007,N_1542,N_1195);
xor U2008 (N_2008,N_1682,N_1956);
nand U2009 (N_2009,N_1693,N_1483);
nor U2010 (N_2010,N_1789,N_1167);
nand U2011 (N_2011,N_1787,N_1754);
nand U2012 (N_2012,N_1784,N_1215);
nand U2013 (N_2013,N_1002,N_1364);
nand U2014 (N_2014,N_1750,N_1622);
and U2015 (N_2015,N_1181,N_1518);
or U2016 (N_2016,N_1731,N_1475);
nor U2017 (N_2017,N_1362,N_1858);
xnor U2018 (N_2018,N_1418,N_1101);
xnor U2019 (N_2019,N_1809,N_1659);
nor U2020 (N_2020,N_1871,N_1861);
and U2021 (N_2021,N_1714,N_1816);
xnor U2022 (N_2022,N_1407,N_1900);
nand U2023 (N_2023,N_1217,N_1284);
or U2024 (N_2024,N_1462,N_1010);
and U2025 (N_2025,N_1645,N_1069);
xor U2026 (N_2026,N_1235,N_1559);
nand U2027 (N_2027,N_1749,N_1239);
nand U2028 (N_2028,N_1737,N_1401);
xor U2029 (N_2029,N_1981,N_1951);
xnor U2030 (N_2030,N_1820,N_1599);
or U2031 (N_2031,N_1114,N_1478);
nor U2032 (N_2032,N_1908,N_1838);
and U2033 (N_2033,N_1579,N_1937);
xnor U2034 (N_2034,N_1484,N_1895);
nor U2035 (N_2035,N_1026,N_1493);
nor U2036 (N_2036,N_1589,N_1328);
xor U2037 (N_2037,N_1095,N_1991);
nor U2038 (N_2038,N_1297,N_1705);
nor U2039 (N_2039,N_1869,N_1548);
nor U2040 (N_2040,N_1607,N_1474);
nor U2041 (N_2041,N_1977,N_1431);
or U2042 (N_2042,N_1487,N_1072);
nor U2043 (N_2043,N_1471,N_1014);
nor U2044 (N_2044,N_1121,N_1827);
xor U2045 (N_2045,N_1893,N_1176);
and U2046 (N_2046,N_1930,N_1736);
or U2047 (N_2047,N_1551,N_1844);
nor U2048 (N_2048,N_1755,N_1430);
nor U2049 (N_2049,N_1161,N_1821);
xnor U2050 (N_2050,N_1106,N_1265);
xor U2051 (N_2051,N_1798,N_1142);
nand U2052 (N_2052,N_1843,N_1845);
nand U2053 (N_2053,N_1728,N_1360);
or U2054 (N_2054,N_1247,N_1839);
and U2055 (N_2055,N_1313,N_1251);
or U2056 (N_2056,N_1437,N_1453);
and U2057 (N_2057,N_1870,N_1996);
nor U2058 (N_2058,N_1301,N_1842);
nand U2059 (N_2059,N_1074,N_1440);
or U2060 (N_2060,N_1066,N_1635);
or U2061 (N_2061,N_1519,N_1145);
or U2062 (N_2062,N_1130,N_1802);
and U2063 (N_2063,N_1993,N_1379);
and U2064 (N_2064,N_1334,N_1073);
or U2065 (N_2065,N_1102,N_1079);
nor U2066 (N_2066,N_1968,N_1243);
nand U2067 (N_2067,N_1155,N_1425);
xor U2068 (N_2068,N_1322,N_1347);
and U2069 (N_2069,N_1323,N_1473);
or U2070 (N_2070,N_1357,N_1090);
and U2071 (N_2071,N_1086,N_1510);
nor U2072 (N_2072,N_1806,N_1982);
xnor U2073 (N_2073,N_1007,N_1184);
and U2074 (N_2074,N_1372,N_1275);
or U2075 (N_2075,N_1625,N_1605);
and U2076 (N_2076,N_1550,N_1189);
nor U2077 (N_2077,N_1495,N_1950);
nand U2078 (N_2078,N_1448,N_1533);
nor U2079 (N_2079,N_1303,N_1928);
and U2080 (N_2080,N_1777,N_1192);
or U2081 (N_2081,N_1132,N_1249);
nor U2082 (N_2082,N_1432,N_1915);
xnor U2083 (N_2083,N_1030,N_1733);
nand U2084 (N_2084,N_1637,N_1641);
and U2085 (N_2085,N_1391,N_1927);
nor U2086 (N_2086,N_1560,N_1967);
and U2087 (N_2087,N_1429,N_1214);
and U2088 (N_2088,N_1566,N_1517);
xnor U2089 (N_2089,N_1295,N_1596);
or U2090 (N_2090,N_1329,N_1123);
or U2091 (N_2091,N_1608,N_1253);
nand U2092 (N_2092,N_1224,N_1907);
nand U2093 (N_2093,N_1291,N_1396);
and U2094 (N_2094,N_1831,N_1266);
and U2095 (N_2095,N_1187,N_1149);
or U2096 (N_2096,N_1726,N_1655);
nor U2097 (N_2097,N_1819,N_1267);
xor U2098 (N_2098,N_1212,N_1242);
xnor U2099 (N_2099,N_1025,N_1120);
or U2100 (N_2100,N_1099,N_1640);
and U2101 (N_2101,N_1125,N_1051);
nand U2102 (N_2102,N_1032,N_1994);
or U2103 (N_2103,N_1972,N_1541);
or U2104 (N_2104,N_1618,N_1966);
or U2105 (N_2105,N_1415,N_1216);
nand U2106 (N_2106,N_1355,N_1445);
nor U2107 (N_2107,N_1709,N_1875);
and U2108 (N_2108,N_1642,N_1888);
and U2109 (N_2109,N_1741,N_1676);
and U2110 (N_2110,N_1801,N_1720);
nor U2111 (N_2111,N_1979,N_1384);
or U2112 (N_2112,N_1923,N_1077);
nand U2113 (N_2113,N_1552,N_1724);
nor U2114 (N_2114,N_1053,N_1345);
or U2115 (N_2115,N_1172,N_1068);
nand U2116 (N_2116,N_1496,N_1206);
nand U2117 (N_2117,N_1882,N_1006);
xnor U2118 (N_2118,N_1260,N_1924);
or U2119 (N_2119,N_1535,N_1444);
or U2120 (N_2120,N_1946,N_1490);
nand U2121 (N_2121,N_1286,N_1526);
or U2122 (N_2122,N_1038,N_1922);
nor U2123 (N_2123,N_1408,N_1082);
and U2124 (N_2124,N_1521,N_1417);
nor U2125 (N_2125,N_1998,N_1857);
nand U2126 (N_2126,N_1906,N_1853);
xor U2127 (N_2127,N_1188,N_1416);
and U2128 (N_2128,N_1442,N_1788);
xor U2129 (N_2129,N_1804,N_1454);
or U2130 (N_2130,N_1942,N_1494);
nand U2131 (N_2131,N_1520,N_1909);
xnor U2132 (N_2132,N_1547,N_1868);
nor U2133 (N_2133,N_1333,N_1449);
nand U2134 (N_2134,N_1234,N_1402);
xnor U2135 (N_2135,N_1472,N_1925);
and U2136 (N_2136,N_1228,N_1648);
and U2137 (N_2137,N_1610,N_1537);
or U2138 (N_2138,N_1557,N_1088);
or U2139 (N_2139,N_1151,N_1044);
or U2140 (N_2140,N_1764,N_1336);
nand U2141 (N_2141,N_1913,N_1603);
nand U2142 (N_2142,N_1245,N_1898);
and U2143 (N_2143,N_1227,N_1973);
and U2144 (N_2144,N_1037,N_1467);
xnor U2145 (N_2145,N_1230,N_1005);
xnor U2146 (N_2146,N_1264,N_1530);
nor U2147 (N_2147,N_1910,N_1631);
and U2148 (N_2148,N_1990,N_1770);
or U2149 (N_2149,N_1594,N_1085);
nand U2150 (N_2150,N_1374,N_1470);
or U2151 (N_2151,N_1835,N_1887);
nand U2152 (N_2152,N_1489,N_1897);
or U2153 (N_2153,N_1776,N_1400);
nand U2154 (N_2154,N_1775,N_1292);
and U2155 (N_2155,N_1896,N_1822);
xor U2156 (N_2156,N_1033,N_1282);
xor U2157 (N_2157,N_1795,N_1246);
xor U2158 (N_2158,N_1052,N_1342);
and U2159 (N_2159,N_1156,N_1287);
and U2160 (N_2160,N_1719,N_1562);
nand U2161 (N_2161,N_1883,N_1008);
nor U2162 (N_2162,N_1258,N_1715);
nor U2163 (N_2163,N_1685,N_1110);
nand U2164 (N_2164,N_1276,N_1237);
or U2165 (N_2165,N_1995,N_1867);
or U2166 (N_2166,N_1054,N_1522);
xnor U2167 (N_2167,N_1670,N_1353);
nor U2168 (N_2168,N_1461,N_1646);
and U2169 (N_2169,N_1294,N_1613);
or U2170 (N_2170,N_1210,N_1314);
and U2171 (N_2171,N_1615,N_1649);
and U2172 (N_2172,N_1945,N_1791);
and U2173 (N_2173,N_1892,N_1580);
nor U2174 (N_2174,N_1865,N_1527);
nand U2175 (N_2175,N_1019,N_1406);
or U2176 (N_2176,N_1177,N_1879);
nor U2177 (N_2177,N_1955,N_1654);
xor U2178 (N_2178,N_1499,N_1439);
or U2179 (N_2179,N_1338,N_1277);
or U2180 (N_2180,N_1988,N_1143);
nand U2181 (N_2181,N_1675,N_1056);
or U2182 (N_2182,N_1585,N_1890);
nor U2183 (N_2183,N_1766,N_1463);
and U2184 (N_2184,N_1790,N_1704);
and U2185 (N_2185,N_1860,N_1466);
or U2186 (N_2186,N_1129,N_1076);
or U2187 (N_2187,N_1969,N_1725);
xor U2188 (N_2188,N_1647,N_1539);
nor U2189 (N_2189,N_1039,N_1511);
nand U2190 (N_2190,N_1711,N_1751);
nor U2191 (N_2191,N_1092,N_1501);
nand U2192 (N_2192,N_1786,N_1901);
nand U2193 (N_2193,N_1986,N_1952);
or U2194 (N_2194,N_1723,N_1045);
xnor U2195 (N_2195,N_1359,N_1738);
and U2196 (N_2196,N_1279,N_1633);
nand U2197 (N_2197,N_1699,N_1023);
or U2198 (N_2198,N_1034,N_1285);
nor U2199 (N_2199,N_1220,N_1783);
or U2200 (N_2200,N_1639,N_1089);
xnor U2201 (N_2201,N_1450,N_1672);
xor U2202 (N_2202,N_1399,N_1435);
nor U2203 (N_2203,N_1523,N_1859);
nor U2204 (N_2204,N_1219,N_1381);
and U2205 (N_2205,N_1884,N_1962);
nand U2206 (N_2206,N_1398,N_1061);
and U2207 (N_2207,N_1757,N_1743);
nor U2208 (N_2208,N_1043,N_1954);
and U2209 (N_2209,N_1133,N_1146);
xor U2210 (N_2210,N_1834,N_1272);
and U2211 (N_2211,N_1252,N_1304);
or U2212 (N_2212,N_1614,N_1105);
and U2213 (N_2213,N_1710,N_1911);
nand U2214 (N_2214,N_1824,N_1638);
or U2215 (N_2215,N_1278,N_1346);
and U2216 (N_2216,N_1361,N_1348);
or U2217 (N_2217,N_1390,N_1446);
or U2218 (N_2218,N_1706,N_1096);
or U2219 (N_2219,N_1035,N_1624);
xor U2220 (N_2220,N_1274,N_1491);
nand U2221 (N_2221,N_1752,N_1593);
xnor U2222 (N_2222,N_1876,N_1104);
nor U2223 (N_2223,N_1931,N_1084);
or U2224 (N_2224,N_1627,N_1315);
and U2225 (N_2225,N_1582,N_1600);
xor U2226 (N_2226,N_1331,N_1564);
xor U2227 (N_2227,N_1358,N_1040);
xor U2228 (N_2228,N_1540,N_1047);
or U2229 (N_2229,N_1815,N_1576);
and U2230 (N_2230,N_1070,N_1921);
nor U2231 (N_2231,N_1847,N_1970);
xor U2232 (N_2232,N_1207,N_1311);
nand U2233 (N_2233,N_1457,N_1165);
or U2234 (N_2234,N_1332,N_1062);
and U2235 (N_2235,N_1350,N_1586);
nor U2236 (N_2236,N_1205,N_1094);
or U2237 (N_2237,N_1203,N_1632);
xnor U2238 (N_2238,N_1001,N_1846);
nor U2239 (N_2239,N_1735,N_1620);
xor U2240 (N_2240,N_1984,N_1310);
nor U2241 (N_2241,N_1296,N_1810);
or U2242 (N_2242,N_1367,N_1138);
nor U2243 (N_2243,N_1700,N_1083);
and U2244 (N_2244,N_1943,N_1273);
and U2245 (N_2245,N_1811,N_1833);
or U2246 (N_2246,N_1468,N_1373);
nor U2247 (N_2247,N_1257,N_1111);
nand U2248 (N_2248,N_1081,N_1936);
xor U2249 (N_2249,N_1889,N_1781);
nand U2250 (N_2250,N_1959,N_1060);
and U2251 (N_2251,N_1160,N_1744);
nor U2252 (N_2252,N_1651,N_1413);
or U2253 (N_2253,N_1914,N_1231);
xor U2254 (N_2254,N_1690,N_1388);
nor U2255 (N_2255,N_1201,N_1691);
or U2256 (N_2256,N_1729,N_1222);
or U2257 (N_2257,N_1689,N_1712);
xor U2258 (N_2258,N_1525,N_1335);
nand U2259 (N_2259,N_1570,N_1182);
nor U2260 (N_2260,N_1592,N_1912);
xnor U2261 (N_2261,N_1387,N_1029);
nor U2262 (N_2262,N_1629,N_1880);
xor U2263 (N_2263,N_1109,N_1563);
and U2264 (N_2264,N_1202,N_1856);
or U2265 (N_2265,N_1877,N_1515);
nand U2266 (N_2266,N_1103,N_1113);
nand U2267 (N_2267,N_1727,N_1899);
or U2268 (N_2268,N_1785,N_1339);
nor U2269 (N_2269,N_1696,N_1602);
nand U2270 (N_2270,N_1154,N_1141);
and U2271 (N_2271,N_1739,N_1978);
xor U2272 (N_2272,N_1989,N_1209);
xnor U2273 (N_2273,N_1905,N_1574);
or U2274 (N_2274,N_1740,N_1091);
and U2275 (N_2275,N_1263,N_1366);
or U2276 (N_2276,N_1657,N_1153);
or U2277 (N_2277,N_1852,N_1702);
or U2278 (N_2278,N_1866,N_1269);
nand U2279 (N_2279,N_1481,N_1538);
xnor U2280 (N_2280,N_1166,N_1926);
nand U2281 (N_2281,N_1581,N_1404);
nor U2282 (N_2282,N_1380,N_1953);
or U2283 (N_2283,N_1948,N_1512);
nor U2284 (N_2284,N_1464,N_1163);
or U2285 (N_2285,N_1768,N_1771);
nor U2286 (N_2286,N_1067,N_1665);
nand U2287 (N_2287,N_1941,N_1392);
nand U2288 (N_2288,N_1619,N_1573);
or U2289 (N_2289,N_1558,N_1306);
nand U2290 (N_2290,N_1722,N_1058);
nor U2291 (N_2291,N_1971,N_1634);
nor U2292 (N_2292,N_1862,N_1606);
nor U2293 (N_2293,N_1503,N_1137);
nor U2294 (N_2294,N_1410,N_1903);
and U2295 (N_2295,N_1456,N_1612);
nand U2296 (N_2296,N_1544,N_1807);
nand U2297 (N_2297,N_1352,N_1127);
xor U2298 (N_2298,N_1250,N_1716);
nor U2299 (N_2299,N_1830,N_1934);
nand U2300 (N_2300,N_1703,N_1695);
nand U2301 (N_2301,N_1904,N_1588);
nand U2302 (N_2302,N_1004,N_1280);
xnor U2303 (N_2303,N_1041,N_1148);
or U2304 (N_2304,N_1183,N_1204);
nand U2305 (N_2305,N_1003,N_1874);
xor U2306 (N_2306,N_1497,N_1112);
and U2307 (N_2307,N_1157,N_1759);
xor U2308 (N_2308,N_1351,N_1916);
xor U2309 (N_2309,N_1940,N_1508);
xnor U2310 (N_2310,N_1344,N_1221);
nand U2311 (N_2311,N_1377,N_1393);
xnor U2312 (N_2312,N_1590,N_1211);
or U2313 (N_2313,N_1383,N_1595);
nand U2314 (N_2314,N_1658,N_1832);
or U2315 (N_2315,N_1268,N_1196);
and U2316 (N_2316,N_1488,N_1370);
and U2317 (N_2317,N_1920,N_1150);
xnor U2318 (N_2318,N_1863,N_1836);
nand U2319 (N_2319,N_1546,N_1218);
nand U2320 (N_2320,N_1681,N_1507);
xor U2321 (N_2321,N_1017,N_1135);
or U2322 (N_2322,N_1529,N_1721);
xnor U2323 (N_2323,N_1375,N_1628);
and U2324 (N_2324,N_1479,N_1983);
nand U2325 (N_2325,N_1200,N_1194);
nor U2326 (N_2326,N_1568,N_1584);
nor U2327 (N_2327,N_1571,N_1403);
xnor U2328 (N_2328,N_1779,N_1116);
xor U2329 (N_2329,N_1611,N_1477);
nand U2330 (N_2330,N_1371,N_1963);
xor U2331 (N_2331,N_1609,N_1668);
and U2332 (N_2332,N_1742,N_1022);
or U2333 (N_2333,N_1554,N_1411);
or U2334 (N_2334,N_1307,N_1841);
nand U2335 (N_2335,N_1808,N_1575);
or U2336 (N_2336,N_1075,N_1687);
or U2337 (N_2337,N_1536,N_1319);
or U2338 (N_2338,N_1349,N_1763);
and U2339 (N_2339,N_1162,N_1621);
nor U2340 (N_2340,N_1389,N_1947);
nand U2341 (N_2341,N_1680,N_1509);
nor U2342 (N_2342,N_1917,N_1302);
or U2343 (N_2343,N_1918,N_1958);
nor U2344 (N_2344,N_1486,N_1837);
nor U2345 (N_2345,N_1233,N_1433);
xor U2346 (N_2346,N_1452,N_1236);
and U2347 (N_2347,N_1271,N_1572);
or U2348 (N_2348,N_1769,N_1792);
xor U2349 (N_2349,N_1248,N_1369);
or U2350 (N_2350,N_1164,N_1087);
xor U2351 (N_2351,N_1556,N_1059);
or U2352 (N_2352,N_1261,N_1814);
nand U2353 (N_2353,N_1476,N_1666);
or U2354 (N_2354,N_1255,N_1553);
nor U2355 (N_2355,N_1935,N_1762);
nand U2356 (N_2356,N_1223,N_1394);
nor U2357 (N_2357,N_1299,N_1420);
or U2358 (N_2358,N_1193,N_1321);
nor U2359 (N_2359,N_1027,N_1506);
or U2360 (N_2360,N_1823,N_1175);
nand U2361 (N_2361,N_1308,N_1532);
nor U2362 (N_2362,N_1938,N_1701);
nand U2363 (N_2363,N_1365,N_1505);
and U2364 (N_2364,N_1199,N_1050);
nand U2365 (N_2365,N_1097,N_1840);
and U2366 (N_2366,N_1140,N_1144);
nand U2367 (N_2367,N_1078,N_1797);
xnor U2368 (N_2368,N_1262,N_1326);
or U2369 (N_2369,N_1340,N_1290);
and U2370 (N_2370,N_1016,N_1692);
or U2371 (N_2371,N_1660,N_1885);
xor U2372 (N_2372,N_1385,N_1854);
nand U2373 (N_2373,N_1974,N_1965);
and U2374 (N_2374,N_1434,N_1734);
xor U2375 (N_2375,N_1849,N_1213);
or U2376 (N_2376,N_1598,N_1591);
or U2377 (N_2377,N_1485,N_1796);
or U2378 (N_2378,N_1949,N_1020);
and U2379 (N_2379,N_1569,N_1881);
xnor U2380 (N_2380,N_1674,N_1441);
xor U2381 (N_2381,N_1939,N_1305);
or U2382 (N_2382,N_1800,N_1327);
nand U2383 (N_2383,N_1760,N_1873);
and U2384 (N_2384,N_1409,N_1697);
xor U2385 (N_2385,N_1480,N_1065);
or U2386 (N_2386,N_1341,N_1492);
nor U2387 (N_2387,N_1708,N_1850);
and U2388 (N_2388,N_1980,N_1136);
nand U2389 (N_2389,N_1186,N_1232);
and U2390 (N_2390,N_1555,N_1872);
xnor U2391 (N_2391,N_1669,N_1288);
xnor U2392 (N_2392,N_1656,N_1688);
or U2393 (N_2393,N_1259,N_1878);
nor U2394 (N_2394,N_1363,N_1662);
nand U2395 (N_2395,N_1851,N_1225);
xnor U2396 (N_2396,N_1270,N_1829);
nor U2397 (N_2397,N_1601,N_1169);
xor U2398 (N_2398,N_1765,N_1782);
and U2399 (N_2399,N_1451,N_1644);
nor U2400 (N_2400,N_1577,N_1178);
xor U2401 (N_2401,N_1254,N_1894);
or U2402 (N_2402,N_1343,N_1864);
nand U2403 (N_2403,N_1185,N_1929);
or U2404 (N_2404,N_1009,N_1667);
or U2405 (N_2405,N_1122,N_1671);
nor U2406 (N_2406,N_1957,N_1049);
xnor U2407 (N_2407,N_1356,N_1747);
or U2408 (N_2408,N_1414,N_1805);
xor U2409 (N_2409,N_1482,N_1975);
or U2410 (N_2410,N_1197,N_1855);
and U2411 (N_2411,N_1997,N_1015);
and U2412 (N_2412,N_1534,N_1173);
nor U2413 (N_2413,N_1567,N_1686);
and U2414 (N_2414,N_1118,N_1528);
and U2415 (N_2415,N_1987,N_1745);
and U2416 (N_2416,N_1071,N_1198);
nor U2417 (N_2417,N_1337,N_1652);
and U2418 (N_2418,N_1767,N_1717);
or U2419 (N_2419,N_1678,N_1126);
and U2420 (N_2420,N_1458,N_1664);
or U2421 (N_2421,N_1500,N_1813);
nand U2422 (N_2422,N_1630,N_1502);
xnor U2423 (N_2423,N_1565,N_1064);
nand U2424 (N_2424,N_1436,N_1443);
nor U2425 (N_2425,N_1428,N_1524);
xnor U2426 (N_2426,N_1803,N_1158);
nand U2427 (N_2427,N_1730,N_1080);
nor U2428 (N_2428,N_1048,N_1324);
nand U2429 (N_2429,N_1180,N_1683);
nor U2430 (N_2430,N_1794,N_1932);
nand U2431 (N_2431,N_1698,N_1397);
or U2432 (N_2432,N_1650,N_1057);
nand U2433 (N_2433,N_1168,N_1818);
nand U2434 (N_2434,N_1694,N_1985);
or U2435 (N_2435,N_1159,N_1028);
nand U2436 (N_2436,N_1679,N_1382);
and U2437 (N_2437,N_1152,N_1663);
and U2438 (N_2438,N_1438,N_1677);
xnor U2439 (N_2439,N_1684,N_1423);
nand U2440 (N_2440,N_1317,N_1597);
nand U2441 (N_2441,N_1139,N_1626);
nand U2442 (N_2442,N_1902,N_1012);
xor U2443 (N_2443,N_1960,N_1093);
or U2444 (N_2444,N_1531,N_1999);
xor U2445 (N_2445,N_1812,N_1514);
nor U2446 (N_2446,N_1545,N_1108);
and U2447 (N_2447,N_1325,N_1773);
nor U2448 (N_2448,N_1386,N_1179);
xor U2449 (N_2449,N_1636,N_1459);
nand U2450 (N_2450,N_1241,N_1011);
nor U2451 (N_2451,N_1447,N_1419);
nand U2452 (N_2452,N_1405,N_1424);
xnor U2453 (N_2453,N_1718,N_1661);
nand U2454 (N_2454,N_1191,N_1761);
and U2455 (N_2455,N_1330,N_1376);
or U2456 (N_2456,N_1455,N_1238);
xnor U2457 (N_2457,N_1115,N_1244);
nand U2458 (N_2458,N_1226,N_1300);
and U2459 (N_2459,N_1281,N_1772);
xor U2460 (N_2460,N_1498,N_1170);
xor U2461 (N_2461,N_1976,N_1427);
nand U2462 (N_2462,N_1623,N_1320);
xor U2463 (N_2463,N_1107,N_1460);
nand U2464 (N_2464,N_1098,N_1748);
nor U2465 (N_2465,N_1289,N_1395);
nor U2466 (N_2466,N_1616,N_1793);
nor U2467 (N_2467,N_1774,N_1055);
nor U2468 (N_2468,N_1021,N_1799);
and U2469 (N_2469,N_1583,N_1673);
or U2470 (N_2470,N_1031,N_1992);
and U2471 (N_2471,N_1516,N_1426);
or U2472 (N_2472,N_1778,N_1513);
and U2473 (N_2473,N_1421,N_1293);
and U2474 (N_2474,N_1653,N_1171);
nor U2475 (N_2475,N_1378,N_1312);
nor U2476 (N_2476,N_1046,N_1208);
nor U2477 (N_2477,N_1024,N_1543);
and U2478 (N_2478,N_1964,N_1354);
xor U2479 (N_2479,N_1933,N_1758);
nor U2480 (N_2480,N_1817,N_1063);
or U2481 (N_2481,N_1919,N_1124);
xnor U2482 (N_2482,N_1746,N_1886);
or U2483 (N_2483,N_1412,N_1578);
or U2484 (N_2484,N_1961,N_1707);
xor U2485 (N_2485,N_1469,N_1617);
nor U2486 (N_2486,N_1256,N_1643);
and U2487 (N_2487,N_1018,N_1825);
or U2488 (N_2488,N_1732,N_1368);
and U2489 (N_2489,N_1134,N_1561);
or U2490 (N_2490,N_1465,N_1753);
and U2491 (N_2491,N_1240,N_1283);
xnor U2492 (N_2492,N_1036,N_1587);
nand U2493 (N_2493,N_1042,N_1848);
or U2494 (N_2494,N_1826,N_1174);
xnor U2495 (N_2495,N_1128,N_1119);
nor U2496 (N_2496,N_1013,N_1229);
and U2497 (N_2497,N_1316,N_1422);
nand U2498 (N_2498,N_1944,N_1713);
xnor U2499 (N_2499,N_1100,N_1891);
or U2500 (N_2500,N_1970,N_1400);
xor U2501 (N_2501,N_1912,N_1650);
nor U2502 (N_2502,N_1110,N_1583);
nor U2503 (N_2503,N_1812,N_1958);
nand U2504 (N_2504,N_1860,N_1894);
or U2505 (N_2505,N_1033,N_1241);
nor U2506 (N_2506,N_1433,N_1532);
or U2507 (N_2507,N_1626,N_1816);
xnor U2508 (N_2508,N_1245,N_1390);
xnor U2509 (N_2509,N_1855,N_1483);
xnor U2510 (N_2510,N_1490,N_1936);
nand U2511 (N_2511,N_1029,N_1187);
nor U2512 (N_2512,N_1589,N_1880);
nor U2513 (N_2513,N_1600,N_1088);
nor U2514 (N_2514,N_1879,N_1701);
or U2515 (N_2515,N_1656,N_1816);
nand U2516 (N_2516,N_1895,N_1822);
and U2517 (N_2517,N_1594,N_1111);
nor U2518 (N_2518,N_1191,N_1795);
and U2519 (N_2519,N_1275,N_1867);
and U2520 (N_2520,N_1403,N_1106);
nor U2521 (N_2521,N_1843,N_1872);
xnor U2522 (N_2522,N_1895,N_1354);
nand U2523 (N_2523,N_1223,N_1315);
nor U2524 (N_2524,N_1088,N_1572);
xnor U2525 (N_2525,N_1269,N_1591);
and U2526 (N_2526,N_1641,N_1111);
xnor U2527 (N_2527,N_1776,N_1594);
nor U2528 (N_2528,N_1401,N_1967);
and U2529 (N_2529,N_1657,N_1481);
nor U2530 (N_2530,N_1753,N_1257);
nor U2531 (N_2531,N_1081,N_1580);
and U2532 (N_2532,N_1142,N_1616);
xnor U2533 (N_2533,N_1117,N_1054);
xor U2534 (N_2534,N_1348,N_1631);
and U2535 (N_2535,N_1134,N_1630);
nor U2536 (N_2536,N_1300,N_1237);
or U2537 (N_2537,N_1341,N_1409);
nand U2538 (N_2538,N_1619,N_1885);
nor U2539 (N_2539,N_1315,N_1128);
or U2540 (N_2540,N_1165,N_1295);
xnor U2541 (N_2541,N_1387,N_1594);
or U2542 (N_2542,N_1480,N_1754);
xnor U2543 (N_2543,N_1538,N_1329);
nor U2544 (N_2544,N_1019,N_1674);
xnor U2545 (N_2545,N_1225,N_1812);
nand U2546 (N_2546,N_1043,N_1420);
xnor U2547 (N_2547,N_1876,N_1668);
xnor U2548 (N_2548,N_1108,N_1095);
or U2549 (N_2549,N_1359,N_1036);
or U2550 (N_2550,N_1040,N_1307);
nor U2551 (N_2551,N_1219,N_1489);
nand U2552 (N_2552,N_1019,N_1638);
or U2553 (N_2553,N_1915,N_1697);
nand U2554 (N_2554,N_1247,N_1689);
nand U2555 (N_2555,N_1468,N_1762);
or U2556 (N_2556,N_1925,N_1706);
or U2557 (N_2557,N_1963,N_1380);
and U2558 (N_2558,N_1021,N_1589);
xnor U2559 (N_2559,N_1583,N_1689);
or U2560 (N_2560,N_1679,N_1964);
nand U2561 (N_2561,N_1167,N_1696);
and U2562 (N_2562,N_1016,N_1488);
nor U2563 (N_2563,N_1841,N_1481);
and U2564 (N_2564,N_1644,N_1268);
and U2565 (N_2565,N_1793,N_1783);
nor U2566 (N_2566,N_1802,N_1257);
nor U2567 (N_2567,N_1537,N_1953);
nor U2568 (N_2568,N_1657,N_1664);
nor U2569 (N_2569,N_1540,N_1549);
and U2570 (N_2570,N_1982,N_1613);
xor U2571 (N_2571,N_1723,N_1801);
and U2572 (N_2572,N_1126,N_1564);
nor U2573 (N_2573,N_1696,N_1031);
xnor U2574 (N_2574,N_1197,N_1962);
xnor U2575 (N_2575,N_1162,N_1214);
or U2576 (N_2576,N_1011,N_1538);
or U2577 (N_2577,N_1606,N_1340);
or U2578 (N_2578,N_1263,N_1045);
nand U2579 (N_2579,N_1236,N_1597);
or U2580 (N_2580,N_1067,N_1405);
xnor U2581 (N_2581,N_1575,N_1943);
nand U2582 (N_2582,N_1449,N_1152);
and U2583 (N_2583,N_1522,N_1135);
and U2584 (N_2584,N_1631,N_1922);
nor U2585 (N_2585,N_1989,N_1921);
xor U2586 (N_2586,N_1491,N_1853);
and U2587 (N_2587,N_1189,N_1588);
and U2588 (N_2588,N_1794,N_1177);
and U2589 (N_2589,N_1081,N_1610);
or U2590 (N_2590,N_1476,N_1391);
or U2591 (N_2591,N_1018,N_1356);
xor U2592 (N_2592,N_1329,N_1466);
and U2593 (N_2593,N_1221,N_1797);
and U2594 (N_2594,N_1043,N_1717);
xor U2595 (N_2595,N_1955,N_1785);
nand U2596 (N_2596,N_1829,N_1537);
xor U2597 (N_2597,N_1772,N_1298);
nor U2598 (N_2598,N_1513,N_1184);
and U2599 (N_2599,N_1510,N_1679);
nand U2600 (N_2600,N_1585,N_1668);
nand U2601 (N_2601,N_1439,N_1161);
and U2602 (N_2602,N_1921,N_1077);
xor U2603 (N_2603,N_1247,N_1479);
nor U2604 (N_2604,N_1769,N_1488);
and U2605 (N_2605,N_1853,N_1113);
or U2606 (N_2606,N_1648,N_1296);
or U2607 (N_2607,N_1826,N_1791);
nand U2608 (N_2608,N_1217,N_1708);
or U2609 (N_2609,N_1774,N_1978);
nand U2610 (N_2610,N_1723,N_1288);
and U2611 (N_2611,N_1335,N_1871);
xnor U2612 (N_2612,N_1007,N_1751);
nor U2613 (N_2613,N_1735,N_1780);
nor U2614 (N_2614,N_1403,N_1648);
or U2615 (N_2615,N_1053,N_1329);
nand U2616 (N_2616,N_1431,N_1883);
or U2617 (N_2617,N_1566,N_1217);
nand U2618 (N_2618,N_1207,N_1775);
and U2619 (N_2619,N_1711,N_1803);
and U2620 (N_2620,N_1323,N_1748);
and U2621 (N_2621,N_1240,N_1749);
xnor U2622 (N_2622,N_1290,N_1450);
or U2623 (N_2623,N_1774,N_1225);
nand U2624 (N_2624,N_1060,N_1906);
or U2625 (N_2625,N_1305,N_1643);
and U2626 (N_2626,N_1894,N_1953);
nand U2627 (N_2627,N_1170,N_1019);
and U2628 (N_2628,N_1825,N_1342);
nor U2629 (N_2629,N_1673,N_1117);
or U2630 (N_2630,N_1182,N_1489);
xnor U2631 (N_2631,N_1590,N_1753);
or U2632 (N_2632,N_1045,N_1308);
nand U2633 (N_2633,N_1168,N_1444);
nor U2634 (N_2634,N_1477,N_1944);
nor U2635 (N_2635,N_1031,N_1968);
nand U2636 (N_2636,N_1609,N_1328);
nor U2637 (N_2637,N_1474,N_1914);
and U2638 (N_2638,N_1841,N_1730);
nor U2639 (N_2639,N_1593,N_1945);
nand U2640 (N_2640,N_1639,N_1574);
xor U2641 (N_2641,N_1569,N_1635);
or U2642 (N_2642,N_1431,N_1812);
and U2643 (N_2643,N_1450,N_1217);
and U2644 (N_2644,N_1985,N_1739);
and U2645 (N_2645,N_1665,N_1878);
nand U2646 (N_2646,N_1132,N_1785);
or U2647 (N_2647,N_1592,N_1593);
or U2648 (N_2648,N_1821,N_1704);
nor U2649 (N_2649,N_1323,N_1676);
xnor U2650 (N_2650,N_1453,N_1913);
nand U2651 (N_2651,N_1144,N_1005);
and U2652 (N_2652,N_1027,N_1264);
xnor U2653 (N_2653,N_1119,N_1656);
nor U2654 (N_2654,N_1604,N_1063);
nand U2655 (N_2655,N_1908,N_1186);
and U2656 (N_2656,N_1558,N_1216);
nand U2657 (N_2657,N_1597,N_1346);
nor U2658 (N_2658,N_1396,N_1448);
xor U2659 (N_2659,N_1946,N_1063);
xor U2660 (N_2660,N_1240,N_1515);
nor U2661 (N_2661,N_1252,N_1726);
nand U2662 (N_2662,N_1945,N_1738);
nand U2663 (N_2663,N_1755,N_1929);
or U2664 (N_2664,N_1632,N_1732);
xor U2665 (N_2665,N_1656,N_1366);
and U2666 (N_2666,N_1094,N_1244);
or U2667 (N_2667,N_1507,N_1344);
or U2668 (N_2668,N_1635,N_1602);
and U2669 (N_2669,N_1702,N_1598);
xor U2670 (N_2670,N_1682,N_1807);
or U2671 (N_2671,N_1226,N_1337);
or U2672 (N_2672,N_1390,N_1370);
and U2673 (N_2673,N_1258,N_1122);
nor U2674 (N_2674,N_1656,N_1585);
and U2675 (N_2675,N_1006,N_1357);
and U2676 (N_2676,N_1619,N_1638);
and U2677 (N_2677,N_1035,N_1547);
and U2678 (N_2678,N_1790,N_1392);
nor U2679 (N_2679,N_1524,N_1357);
and U2680 (N_2680,N_1096,N_1703);
nor U2681 (N_2681,N_1684,N_1249);
xnor U2682 (N_2682,N_1110,N_1813);
nor U2683 (N_2683,N_1035,N_1430);
or U2684 (N_2684,N_1849,N_1751);
and U2685 (N_2685,N_1364,N_1860);
and U2686 (N_2686,N_1724,N_1527);
nor U2687 (N_2687,N_1215,N_1690);
xnor U2688 (N_2688,N_1618,N_1678);
and U2689 (N_2689,N_1392,N_1428);
nor U2690 (N_2690,N_1339,N_1178);
xor U2691 (N_2691,N_1379,N_1633);
nand U2692 (N_2692,N_1999,N_1345);
or U2693 (N_2693,N_1375,N_1004);
and U2694 (N_2694,N_1737,N_1745);
xor U2695 (N_2695,N_1471,N_1819);
or U2696 (N_2696,N_1206,N_1514);
nand U2697 (N_2697,N_1896,N_1585);
or U2698 (N_2698,N_1341,N_1599);
nand U2699 (N_2699,N_1825,N_1425);
nand U2700 (N_2700,N_1208,N_1568);
and U2701 (N_2701,N_1952,N_1427);
and U2702 (N_2702,N_1651,N_1068);
or U2703 (N_2703,N_1034,N_1458);
nor U2704 (N_2704,N_1523,N_1702);
or U2705 (N_2705,N_1293,N_1164);
nand U2706 (N_2706,N_1473,N_1956);
and U2707 (N_2707,N_1695,N_1429);
nand U2708 (N_2708,N_1974,N_1443);
nand U2709 (N_2709,N_1663,N_1819);
nand U2710 (N_2710,N_1058,N_1419);
xnor U2711 (N_2711,N_1028,N_1921);
xnor U2712 (N_2712,N_1917,N_1935);
nand U2713 (N_2713,N_1859,N_1787);
or U2714 (N_2714,N_1885,N_1315);
xor U2715 (N_2715,N_1738,N_1948);
nand U2716 (N_2716,N_1839,N_1130);
and U2717 (N_2717,N_1476,N_1066);
nand U2718 (N_2718,N_1235,N_1830);
nor U2719 (N_2719,N_1638,N_1258);
or U2720 (N_2720,N_1154,N_1717);
and U2721 (N_2721,N_1162,N_1625);
and U2722 (N_2722,N_1283,N_1540);
nor U2723 (N_2723,N_1616,N_1960);
nor U2724 (N_2724,N_1539,N_1205);
nor U2725 (N_2725,N_1486,N_1751);
nand U2726 (N_2726,N_1026,N_1308);
or U2727 (N_2727,N_1562,N_1884);
or U2728 (N_2728,N_1657,N_1160);
xnor U2729 (N_2729,N_1009,N_1687);
nor U2730 (N_2730,N_1282,N_1074);
or U2731 (N_2731,N_1837,N_1634);
nand U2732 (N_2732,N_1686,N_1467);
xor U2733 (N_2733,N_1411,N_1356);
and U2734 (N_2734,N_1424,N_1876);
or U2735 (N_2735,N_1244,N_1981);
xor U2736 (N_2736,N_1846,N_1176);
nor U2737 (N_2737,N_1303,N_1350);
or U2738 (N_2738,N_1007,N_1426);
and U2739 (N_2739,N_1834,N_1179);
xor U2740 (N_2740,N_1933,N_1870);
or U2741 (N_2741,N_1507,N_1281);
nor U2742 (N_2742,N_1196,N_1524);
and U2743 (N_2743,N_1869,N_1774);
and U2744 (N_2744,N_1060,N_1191);
xor U2745 (N_2745,N_1447,N_1253);
or U2746 (N_2746,N_1006,N_1562);
nor U2747 (N_2747,N_1436,N_1463);
and U2748 (N_2748,N_1586,N_1305);
xnor U2749 (N_2749,N_1642,N_1338);
nand U2750 (N_2750,N_1000,N_1282);
nand U2751 (N_2751,N_1301,N_1503);
xor U2752 (N_2752,N_1471,N_1950);
xor U2753 (N_2753,N_1032,N_1601);
xnor U2754 (N_2754,N_1657,N_1752);
xnor U2755 (N_2755,N_1188,N_1454);
xor U2756 (N_2756,N_1260,N_1934);
xnor U2757 (N_2757,N_1606,N_1875);
nand U2758 (N_2758,N_1024,N_1642);
xnor U2759 (N_2759,N_1030,N_1439);
nor U2760 (N_2760,N_1355,N_1870);
nand U2761 (N_2761,N_1116,N_1993);
nand U2762 (N_2762,N_1994,N_1951);
nand U2763 (N_2763,N_1139,N_1787);
nor U2764 (N_2764,N_1651,N_1860);
xor U2765 (N_2765,N_1636,N_1591);
nand U2766 (N_2766,N_1594,N_1025);
or U2767 (N_2767,N_1038,N_1066);
nand U2768 (N_2768,N_1523,N_1627);
xor U2769 (N_2769,N_1066,N_1165);
and U2770 (N_2770,N_1829,N_1114);
and U2771 (N_2771,N_1897,N_1507);
and U2772 (N_2772,N_1735,N_1331);
nor U2773 (N_2773,N_1254,N_1710);
or U2774 (N_2774,N_1380,N_1458);
nand U2775 (N_2775,N_1723,N_1816);
nand U2776 (N_2776,N_1278,N_1628);
nand U2777 (N_2777,N_1945,N_1807);
xor U2778 (N_2778,N_1959,N_1034);
xor U2779 (N_2779,N_1023,N_1343);
and U2780 (N_2780,N_1133,N_1393);
nand U2781 (N_2781,N_1142,N_1351);
xnor U2782 (N_2782,N_1309,N_1308);
nand U2783 (N_2783,N_1599,N_1614);
or U2784 (N_2784,N_1387,N_1695);
nor U2785 (N_2785,N_1783,N_1116);
or U2786 (N_2786,N_1304,N_1446);
xor U2787 (N_2787,N_1778,N_1951);
nand U2788 (N_2788,N_1554,N_1339);
xnor U2789 (N_2789,N_1847,N_1514);
nor U2790 (N_2790,N_1140,N_1635);
or U2791 (N_2791,N_1857,N_1478);
and U2792 (N_2792,N_1179,N_1080);
xnor U2793 (N_2793,N_1235,N_1644);
nand U2794 (N_2794,N_1774,N_1748);
nand U2795 (N_2795,N_1986,N_1283);
and U2796 (N_2796,N_1788,N_1512);
or U2797 (N_2797,N_1596,N_1270);
and U2798 (N_2798,N_1744,N_1279);
nand U2799 (N_2799,N_1538,N_1769);
nand U2800 (N_2800,N_1221,N_1994);
xnor U2801 (N_2801,N_1437,N_1523);
xnor U2802 (N_2802,N_1734,N_1858);
nand U2803 (N_2803,N_1066,N_1649);
and U2804 (N_2804,N_1532,N_1205);
nor U2805 (N_2805,N_1351,N_1130);
nand U2806 (N_2806,N_1528,N_1231);
xnor U2807 (N_2807,N_1972,N_1159);
xnor U2808 (N_2808,N_1925,N_1211);
nor U2809 (N_2809,N_1680,N_1897);
and U2810 (N_2810,N_1580,N_1627);
nor U2811 (N_2811,N_1363,N_1139);
and U2812 (N_2812,N_1758,N_1852);
nand U2813 (N_2813,N_1865,N_1120);
nand U2814 (N_2814,N_1815,N_1232);
xor U2815 (N_2815,N_1373,N_1673);
and U2816 (N_2816,N_1374,N_1511);
or U2817 (N_2817,N_1165,N_1657);
and U2818 (N_2818,N_1892,N_1606);
nor U2819 (N_2819,N_1190,N_1266);
or U2820 (N_2820,N_1467,N_1877);
and U2821 (N_2821,N_1576,N_1296);
nand U2822 (N_2822,N_1020,N_1423);
or U2823 (N_2823,N_1886,N_1640);
nand U2824 (N_2824,N_1237,N_1651);
xor U2825 (N_2825,N_1506,N_1919);
xor U2826 (N_2826,N_1433,N_1093);
and U2827 (N_2827,N_1362,N_1231);
nand U2828 (N_2828,N_1292,N_1261);
and U2829 (N_2829,N_1900,N_1486);
and U2830 (N_2830,N_1580,N_1800);
and U2831 (N_2831,N_1477,N_1525);
xor U2832 (N_2832,N_1208,N_1364);
or U2833 (N_2833,N_1136,N_1126);
and U2834 (N_2834,N_1388,N_1458);
and U2835 (N_2835,N_1806,N_1280);
and U2836 (N_2836,N_1117,N_1160);
and U2837 (N_2837,N_1971,N_1294);
or U2838 (N_2838,N_1257,N_1491);
or U2839 (N_2839,N_1555,N_1128);
xor U2840 (N_2840,N_1729,N_1017);
and U2841 (N_2841,N_1796,N_1784);
nor U2842 (N_2842,N_1219,N_1163);
nor U2843 (N_2843,N_1948,N_1786);
nor U2844 (N_2844,N_1114,N_1697);
nor U2845 (N_2845,N_1819,N_1336);
xnor U2846 (N_2846,N_1934,N_1787);
or U2847 (N_2847,N_1627,N_1737);
nand U2848 (N_2848,N_1021,N_1612);
or U2849 (N_2849,N_1590,N_1234);
and U2850 (N_2850,N_1811,N_1789);
and U2851 (N_2851,N_1735,N_1877);
nand U2852 (N_2852,N_1912,N_1456);
nand U2853 (N_2853,N_1921,N_1428);
or U2854 (N_2854,N_1569,N_1564);
and U2855 (N_2855,N_1322,N_1233);
or U2856 (N_2856,N_1501,N_1338);
xnor U2857 (N_2857,N_1624,N_1236);
and U2858 (N_2858,N_1093,N_1241);
nor U2859 (N_2859,N_1965,N_1158);
xor U2860 (N_2860,N_1499,N_1423);
and U2861 (N_2861,N_1161,N_1056);
nor U2862 (N_2862,N_1506,N_1629);
nand U2863 (N_2863,N_1606,N_1900);
xnor U2864 (N_2864,N_1357,N_1970);
nand U2865 (N_2865,N_1148,N_1969);
or U2866 (N_2866,N_1988,N_1440);
nor U2867 (N_2867,N_1070,N_1700);
or U2868 (N_2868,N_1769,N_1395);
nor U2869 (N_2869,N_1674,N_1162);
xor U2870 (N_2870,N_1574,N_1454);
nand U2871 (N_2871,N_1670,N_1746);
or U2872 (N_2872,N_1412,N_1588);
or U2873 (N_2873,N_1447,N_1817);
and U2874 (N_2874,N_1032,N_1507);
nand U2875 (N_2875,N_1992,N_1491);
xor U2876 (N_2876,N_1179,N_1695);
and U2877 (N_2877,N_1372,N_1893);
and U2878 (N_2878,N_1510,N_1660);
or U2879 (N_2879,N_1760,N_1714);
nor U2880 (N_2880,N_1468,N_1957);
nand U2881 (N_2881,N_1716,N_1160);
and U2882 (N_2882,N_1424,N_1152);
or U2883 (N_2883,N_1522,N_1283);
and U2884 (N_2884,N_1883,N_1876);
and U2885 (N_2885,N_1847,N_1851);
nor U2886 (N_2886,N_1068,N_1202);
and U2887 (N_2887,N_1270,N_1954);
nor U2888 (N_2888,N_1950,N_1103);
nand U2889 (N_2889,N_1376,N_1258);
xnor U2890 (N_2890,N_1523,N_1451);
and U2891 (N_2891,N_1140,N_1205);
nand U2892 (N_2892,N_1514,N_1231);
and U2893 (N_2893,N_1483,N_1022);
nand U2894 (N_2894,N_1122,N_1369);
and U2895 (N_2895,N_1385,N_1309);
nor U2896 (N_2896,N_1397,N_1296);
or U2897 (N_2897,N_1026,N_1560);
xnor U2898 (N_2898,N_1125,N_1901);
nand U2899 (N_2899,N_1154,N_1595);
nand U2900 (N_2900,N_1061,N_1107);
nand U2901 (N_2901,N_1676,N_1794);
nand U2902 (N_2902,N_1331,N_1458);
nor U2903 (N_2903,N_1766,N_1332);
nand U2904 (N_2904,N_1251,N_1578);
xnor U2905 (N_2905,N_1350,N_1301);
and U2906 (N_2906,N_1149,N_1879);
nor U2907 (N_2907,N_1693,N_1992);
nor U2908 (N_2908,N_1505,N_1765);
and U2909 (N_2909,N_1314,N_1183);
xor U2910 (N_2910,N_1704,N_1525);
xnor U2911 (N_2911,N_1904,N_1229);
nand U2912 (N_2912,N_1477,N_1022);
nor U2913 (N_2913,N_1104,N_1536);
or U2914 (N_2914,N_1592,N_1338);
and U2915 (N_2915,N_1730,N_1839);
nor U2916 (N_2916,N_1436,N_1029);
xnor U2917 (N_2917,N_1565,N_1285);
nor U2918 (N_2918,N_1095,N_1625);
nand U2919 (N_2919,N_1578,N_1605);
nand U2920 (N_2920,N_1279,N_1322);
or U2921 (N_2921,N_1117,N_1919);
xor U2922 (N_2922,N_1585,N_1072);
and U2923 (N_2923,N_1455,N_1253);
nand U2924 (N_2924,N_1410,N_1996);
nor U2925 (N_2925,N_1884,N_1830);
or U2926 (N_2926,N_1556,N_1113);
and U2927 (N_2927,N_1037,N_1200);
or U2928 (N_2928,N_1121,N_1879);
nor U2929 (N_2929,N_1840,N_1286);
or U2930 (N_2930,N_1000,N_1449);
nand U2931 (N_2931,N_1233,N_1560);
or U2932 (N_2932,N_1920,N_1142);
or U2933 (N_2933,N_1318,N_1732);
nor U2934 (N_2934,N_1558,N_1627);
nor U2935 (N_2935,N_1175,N_1205);
or U2936 (N_2936,N_1978,N_1322);
nand U2937 (N_2937,N_1425,N_1555);
xnor U2938 (N_2938,N_1126,N_1177);
or U2939 (N_2939,N_1632,N_1689);
and U2940 (N_2940,N_1116,N_1303);
or U2941 (N_2941,N_1801,N_1882);
nor U2942 (N_2942,N_1816,N_1136);
nor U2943 (N_2943,N_1979,N_1482);
xnor U2944 (N_2944,N_1515,N_1960);
nand U2945 (N_2945,N_1030,N_1063);
xnor U2946 (N_2946,N_1606,N_1397);
nand U2947 (N_2947,N_1211,N_1213);
nor U2948 (N_2948,N_1671,N_1073);
or U2949 (N_2949,N_1836,N_1707);
and U2950 (N_2950,N_1548,N_1103);
xnor U2951 (N_2951,N_1193,N_1267);
or U2952 (N_2952,N_1773,N_1645);
nand U2953 (N_2953,N_1364,N_1514);
xor U2954 (N_2954,N_1650,N_1512);
xor U2955 (N_2955,N_1107,N_1486);
nor U2956 (N_2956,N_1311,N_1489);
or U2957 (N_2957,N_1181,N_1968);
and U2958 (N_2958,N_1258,N_1117);
nand U2959 (N_2959,N_1855,N_1773);
nor U2960 (N_2960,N_1447,N_1346);
xor U2961 (N_2961,N_1288,N_1161);
nor U2962 (N_2962,N_1034,N_1804);
and U2963 (N_2963,N_1228,N_1622);
xor U2964 (N_2964,N_1177,N_1728);
nor U2965 (N_2965,N_1018,N_1205);
or U2966 (N_2966,N_1573,N_1624);
xor U2967 (N_2967,N_1989,N_1680);
and U2968 (N_2968,N_1288,N_1910);
nand U2969 (N_2969,N_1289,N_1066);
or U2970 (N_2970,N_1318,N_1911);
xor U2971 (N_2971,N_1939,N_1220);
nor U2972 (N_2972,N_1536,N_1497);
nor U2973 (N_2973,N_1831,N_1784);
xnor U2974 (N_2974,N_1056,N_1314);
xor U2975 (N_2975,N_1228,N_1896);
nand U2976 (N_2976,N_1705,N_1357);
or U2977 (N_2977,N_1547,N_1929);
xor U2978 (N_2978,N_1037,N_1520);
nand U2979 (N_2979,N_1534,N_1866);
or U2980 (N_2980,N_1875,N_1581);
and U2981 (N_2981,N_1294,N_1608);
or U2982 (N_2982,N_1776,N_1840);
xnor U2983 (N_2983,N_1412,N_1195);
nand U2984 (N_2984,N_1434,N_1740);
or U2985 (N_2985,N_1803,N_1561);
and U2986 (N_2986,N_1489,N_1121);
nand U2987 (N_2987,N_1364,N_1901);
or U2988 (N_2988,N_1882,N_1211);
nand U2989 (N_2989,N_1759,N_1838);
nor U2990 (N_2990,N_1024,N_1195);
or U2991 (N_2991,N_1968,N_1079);
and U2992 (N_2992,N_1843,N_1588);
xor U2993 (N_2993,N_1132,N_1662);
and U2994 (N_2994,N_1871,N_1486);
nor U2995 (N_2995,N_1101,N_1823);
and U2996 (N_2996,N_1198,N_1140);
nand U2997 (N_2997,N_1722,N_1520);
and U2998 (N_2998,N_1550,N_1902);
nor U2999 (N_2999,N_1088,N_1265);
and UO_0 (O_0,N_2249,N_2967);
nor UO_1 (O_1,N_2140,N_2165);
nand UO_2 (O_2,N_2102,N_2812);
xnor UO_3 (O_3,N_2137,N_2283);
and UO_4 (O_4,N_2033,N_2459);
nand UO_5 (O_5,N_2418,N_2681);
or UO_6 (O_6,N_2118,N_2891);
nor UO_7 (O_7,N_2186,N_2245);
nand UO_8 (O_8,N_2021,N_2873);
nor UO_9 (O_9,N_2913,N_2398);
xor UO_10 (O_10,N_2668,N_2863);
or UO_11 (O_11,N_2430,N_2853);
and UO_12 (O_12,N_2049,N_2498);
nand UO_13 (O_13,N_2496,N_2910);
nand UO_14 (O_14,N_2030,N_2545);
nor UO_15 (O_15,N_2223,N_2592);
nand UO_16 (O_16,N_2674,N_2969);
and UO_17 (O_17,N_2754,N_2895);
nand UO_18 (O_18,N_2004,N_2002);
nor UO_19 (O_19,N_2390,N_2840);
or UO_20 (O_20,N_2847,N_2228);
nand UO_21 (O_21,N_2092,N_2145);
or UO_22 (O_22,N_2638,N_2098);
or UO_23 (O_23,N_2501,N_2193);
xor UO_24 (O_24,N_2904,N_2793);
or UO_25 (O_25,N_2234,N_2476);
xor UO_26 (O_26,N_2360,N_2747);
and UO_27 (O_27,N_2054,N_2426);
nand UO_28 (O_28,N_2125,N_2805);
nor UO_29 (O_29,N_2900,N_2475);
and UO_30 (O_30,N_2264,N_2888);
nor UO_31 (O_31,N_2774,N_2645);
xor UO_32 (O_32,N_2407,N_2865);
or UO_33 (O_33,N_2593,N_2875);
nor UO_34 (O_34,N_2235,N_2502);
and UO_35 (O_35,N_2979,N_2539);
or UO_36 (O_36,N_2351,N_2159);
xnor UO_37 (O_37,N_2604,N_2704);
nor UO_38 (O_38,N_2301,N_2141);
or UO_39 (O_39,N_2016,N_2014);
xnor UO_40 (O_40,N_2542,N_2233);
nand UO_41 (O_41,N_2968,N_2838);
or UO_42 (O_42,N_2737,N_2236);
nor UO_43 (O_43,N_2596,N_2981);
nor UO_44 (O_44,N_2254,N_2787);
or UO_45 (O_45,N_2685,N_2286);
or UO_46 (O_46,N_2522,N_2497);
and UO_47 (O_47,N_2210,N_2250);
nand UO_48 (O_48,N_2915,N_2640);
nand UO_49 (O_49,N_2688,N_2794);
nand UO_50 (O_50,N_2658,N_2636);
nor UO_51 (O_51,N_2296,N_2831);
and UO_52 (O_52,N_2661,N_2244);
nor UO_53 (O_53,N_2409,N_2833);
nor UO_54 (O_54,N_2791,N_2150);
and UO_55 (O_55,N_2386,N_2748);
or UO_56 (O_56,N_2918,N_2100);
xnor UO_57 (O_57,N_2288,N_2729);
nand UO_58 (O_58,N_2926,N_2275);
nand UO_59 (O_59,N_2733,N_2716);
xnor UO_60 (O_60,N_2346,N_2119);
and UO_61 (O_61,N_2023,N_2856);
xnor UO_62 (O_62,N_2877,N_2608);
and UO_63 (O_63,N_2491,N_2077);
or UO_64 (O_64,N_2870,N_2213);
and UO_65 (O_65,N_2835,N_2574);
nand UO_66 (O_66,N_2220,N_2515);
and UO_67 (O_67,N_2225,N_2821);
and UO_68 (O_68,N_2544,N_2701);
nand UO_69 (O_69,N_2783,N_2667);
and UO_70 (O_70,N_2956,N_2586);
or UO_71 (O_71,N_2813,N_2919);
nand UO_72 (O_72,N_2778,N_2078);
nor UO_73 (O_73,N_2690,N_2139);
or UO_74 (O_74,N_2735,N_2138);
and UO_75 (O_75,N_2019,N_2417);
or UO_76 (O_76,N_2192,N_2914);
or UO_77 (O_77,N_2975,N_2180);
and UO_78 (O_78,N_2982,N_2558);
nor UO_79 (O_79,N_2676,N_2441);
xor UO_80 (O_80,N_2583,N_2185);
and UO_81 (O_81,N_2200,N_2908);
nor UO_82 (O_82,N_2206,N_2530);
nand UO_83 (O_83,N_2601,N_2034);
and UO_84 (O_84,N_2897,N_2896);
and UO_85 (O_85,N_2719,N_2988);
or UO_86 (O_86,N_2340,N_2328);
nand UO_87 (O_87,N_2463,N_2284);
nand UO_88 (O_88,N_2932,N_2204);
or UO_89 (O_89,N_2788,N_2972);
nor UO_90 (O_90,N_2957,N_2955);
nand UO_91 (O_91,N_2770,N_2556);
and UO_92 (O_92,N_2759,N_2945);
nor UO_93 (O_93,N_2209,N_2026);
nor UO_94 (O_94,N_2304,N_2166);
and UO_95 (O_95,N_2557,N_2632);
xnor UO_96 (O_96,N_2858,N_2101);
nand UO_97 (O_97,N_2650,N_2769);
nand UO_98 (O_98,N_2256,N_2818);
nand UO_99 (O_99,N_2798,N_2698);
nor UO_100 (O_100,N_2610,N_2790);
and UO_101 (O_101,N_2299,N_2191);
and UO_102 (O_102,N_2440,N_2089);
and UO_103 (O_103,N_2480,N_2113);
and UO_104 (O_104,N_2776,N_2810);
nand UO_105 (O_105,N_2451,N_2103);
nor UO_106 (O_106,N_2452,N_2365);
or UO_107 (O_107,N_2073,N_2152);
nand UO_108 (O_108,N_2302,N_2285);
nor UO_109 (O_109,N_2190,N_2934);
xnor UO_110 (O_110,N_2987,N_2461);
nand UO_111 (O_111,N_2414,N_2611);
or UO_112 (O_112,N_2552,N_2907);
and UO_113 (O_113,N_2994,N_2857);
xnor UO_114 (O_114,N_2133,N_2282);
xnor UO_115 (O_115,N_2902,N_2991);
and UO_116 (O_116,N_2197,N_2731);
nand UO_117 (O_117,N_2664,N_2112);
nand UO_118 (O_118,N_2713,N_2757);
nand UO_119 (O_119,N_2621,N_2983);
and UO_120 (O_120,N_2773,N_2076);
nand UO_121 (O_121,N_2694,N_2024);
nand UO_122 (O_122,N_2511,N_2270);
xnor UO_123 (O_123,N_2356,N_2624);
xnor UO_124 (O_124,N_2447,N_2115);
nor UO_125 (O_125,N_2478,N_2564);
and UO_126 (O_126,N_2846,N_2408);
nor UO_127 (O_127,N_2040,N_2110);
or UO_128 (O_128,N_2022,N_2059);
xnor UO_129 (O_129,N_2927,N_2425);
xor UO_130 (O_130,N_2460,N_2384);
nor UO_131 (O_131,N_2550,N_2976);
nand UO_132 (O_132,N_2796,N_2037);
or UO_133 (O_133,N_2855,N_2208);
and UO_134 (O_134,N_2643,N_2240);
or UO_135 (O_135,N_2971,N_2699);
and UO_136 (O_136,N_2817,N_2600);
and UO_137 (O_137,N_2506,N_2553);
xnor UO_138 (O_138,N_2160,N_2682);
and UO_139 (O_139,N_2266,N_2175);
or UO_140 (O_140,N_2067,N_2294);
xnor UO_141 (O_141,N_2268,N_2939);
and UO_142 (O_142,N_2368,N_2135);
nor UO_143 (O_143,N_2859,N_2602);
xor UO_144 (O_144,N_2289,N_2909);
and UO_145 (O_145,N_2966,N_2074);
or UO_146 (O_146,N_2538,N_2349);
or UO_147 (O_147,N_2797,N_2011);
nor UO_148 (O_148,N_2095,N_2996);
xnor UO_149 (O_149,N_2094,N_2876);
or UO_150 (O_150,N_2861,N_2869);
xor UO_151 (O_151,N_2132,N_2973);
nor UO_152 (O_152,N_2534,N_2064);
xor UO_153 (O_153,N_2068,N_2819);
and UO_154 (O_154,N_2130,N_2168);
nand UO_155 (O_155,N_2952,N_2446);
or UO_156 (O_156,N_2305,N_2518);
nor UO_157 (O_157,N_2397,N_2670);
nor UO_158 (O_158,N_2255,N_2317);
nand UO_159 (O_159,N_2388,N_2320);
nand UO_160 (O_160,N_2663,N_2756);
or UO_161 (O_161,N_2815,N_2382);
xnor UO_162 (O_162,N_2651,N_2623);
nor UO_163 (O_163,N_2344,N_2237);
xnor UO_164 (O_164,N_2916,N_2111);
nand UO_165 (O_165,N_2614,N_2992);
or UO_166 (O_166,N_2563,N_2046);
xnor UO_167 (O_167,N_2482,N_2609);
or UO_168 (O_168,N_2196,N_2226);
xnor UO_169 (O_169,N_2779,N_2198);
nor UO_170 (O_170,N_2717,N_2371);
nand UO_171 (O_171,N_2726,N_2993);
or UO_172 (O_172,N_2619,N_2671);
nor UO_173 (O_173,N_2510,N_2874);
nor UO_174 (O_174,N_2436,N_2703);
nor UO_175 (O_175,N_2995,N_2848);
nor UO_176 (O_176,N_2679,N_2814);
nand UO_177 (O_177,N_2761,N_2649);
xnor UO_178 (O_178,N_2692,N_2470);
and UO_179 (O_179,N_2924,N_2310);
and UO_180 (O_180,N_2946,N_2325);
and UO_181 (O_181,N_2566,N_2540);
nor UO_182 (O_182,N_2584,N_2655);
xor UO_183 (O_183,N_2380,N_2706);
and UO_184 (O_184,N_2758,N_2507);
or UO_185 (O_185,N_2247,N_2312);
nor UO_186 (O_186,N_2938,N_2804);
nor UO_187 (O_187,N_2999,N_2803);
nand UO_188 (O_188,N_2599,N_2322);
xnor UO_189 (O_189,N_2777,N_2029);
nor UO_190 (O_190,N_2653,N_2811);
nand UO_191 (O_191,N_2280,N_2087);
or UO_192 (O_192,N_2048,N_2156);
and UO_193 (O_193,N_2309,N_2546);
nor UO_194 (O_194,N_2732,N_2837);
xnor UO_195 (O_195,N_2686,N_2764);
nor UO_196 (O_196,N_2224,N_2977);
nor UO_197 (O_197,N_2867,N_2271);
nand UO_198 (O_198,N_2017,N_2324);
or UO_199 (O_199,N_2830,N_2462);
nor UO_200 (O_200,N_2575,N_2943);
nor UO_201 (O_201,N_2164,N_2457);
nand UO_202 (O_202,N_2262,N_2474);
nor UO_203 (O_203,N_2001,N_2702);
or UO_204 (O_204,N_2389,N_2307);
nor UO_205 (O_205,N_2750,N_2172);
and UO_206 (O_206,N_2730,N_2646);
and UO_207 (O_207,N_2494,N_2598);
and UO_208 (O_208,N_2618,N_2473);
xor UO_209 (O_209,N_2925,N_2134);
nor UO_210 (O_210,N_2944,N_2625);
and UO_211 (O_211,N_2772,N_2121);
nor UO_212 (O_212,N_2431,N_2882);
or UO_213 (O_213,N_2472,N_2594);
nor UO_214 (O_214,N_2961,N_2079);
and UO_215 (O_215,N_2560,N_2525);
and UO_216 (O_216,N_2025,N_2062);
or UO_217 (O_217,N_2069,N_2050);
nor UO_218 (O_218,N_2744,N_2099);
and UO_219 (O_219,N_2573,N_2454);
xor UO_220 (O_220,N_2066,N_2845);
and UO_221 (O_221,N_2958,N_2199);
and UO_222 (O_222,N_2456,N_2438);
and UO_223 (O_223,N_2617,N_2905);
nand UO_224 (O_224,N_2147,N_2400);
nor UO_225 (O_225,N_2162,N_2490);
nand UO_226 (O_226,N_2263,N_2242);
nor UO_227 (O_227,N_2229,N_2535);
nor UO_228 (O_228,N_2372,N_2889);
nand UO_229 (O_229,N_2660,N_2736);
and UO_230 (O_230,N_2032,N_2331);
and UO_231 (O_231,N_2038,N_2136);
nand UO_232 (O_232,N_2509,N_2612);
xnor UO_233 (O_233,N_2767,N_2959);
and UO_234 (O_234,N_2687,N_2942);
or UO_235 (O_235,N_2370,N_2158);
xnor UO_236 (O_236,N_2261,N_2469);
and UO_237 (O_237,N_2170,N_2207);
xor UO_238 (O_238,N_2523,N_2217);
and UO_239 (O_239,N_2215,N_2551);
nor UO_240 (O_240,N_2559,N_2669);
xnor UO_241 (O_241,N_2738,N_2792);
nor UO_242 (O_242,N_2298,N_2708);
nor UO_243 (O_243,N_2595,N_2258);
and UO_244 (O_244,N_2639,N_2931);
nor UO_245 (O_245,N_2826,N_2657);
and UO_246 (O_246,N_2448,N_2107);
nor UO_247 (O_247,N_2072,N_2238);
and UO_248 (O_248,N_2720,N_2093);
nor UO_249 (O_249,N_2505,N_2316);
and UO_250 (O_250,N_2526,N_2176);
or UO_251 (O_251,N_2755,N_2589);
xor UO_252 (O_252,N_2230,N_2760);
nand UO_253 (O_253,N_2058,N_2297);
or UO_254 (O_254,N_2485,N_2013);
nor UO_255 (O_255,N_2082,N_2562);
nand UO_256 (O_256,N_2854,N_2892);
nor UO_257 (O_257,N_2424,N_2823);
nand UO_258 (O_258,N_2585,N_2742);
nor UO_259 (O_259,N_2007,N_2027);
nor UO_260 (O_260,N_2543,N_2203);
and UO_261 (O_261,N_2412,N_2303);
xor UO_262 (O_262,N_2520,N_2568);
and UO_263 (O_263,N_2597,N_2878);
xnor UO_264 (O_264,N_2061,N_2127);
nand UO_265 (O_265,N_2241,N_2403);
nor UO_266 (O_266,N_2329,N_2642);
or UO_267 (O_267,N_2850,N_2008);
and UO_268 (O_268,N_2691,N_2739);
or UO_269 (O_269,N_2375,N_2871);
nor UO_270 (O_270,N_2253,N_2091);
nand UO_271 (O_271,N_2930,N_2359);
nand UO_272 (O_272,N_2762,N_2071);
nor UO_273 (O_273,N_2807,N_2269);
nand UO_274 (O_274,N_2637,N_2039);
nand UO_275 (O_275,N_2277,N_2222);
or UO_276 (O_276,N_2827,N_2753);
nor UO_277 (O_277,N_2290,N_2377);
nor UO_278 (O_278,N_2334,N_2405);
or UO_279 (O_279,N_2746,N_2465);
xor UO_280 (O_280,N_2323,N_2784);
nor UO_281 (O_281,N_2893,N_2721);
nor UO_282 (O_282,N_2260,N_2672);
and UO_283 (O_283,N_2808,N_2012);
and UO_284 (O_284,N_2894,N_2665);
and UO_285 (O_285,N_2512,N_2142);
nand UO_286 (O_286,N_2627,N_2464);
or UO_287 (O_287,N_2257,N_2644);
nor UO_288 (O_288,N_2392,N_2697);
nand UO_289 (O_289,N_2188,N_2962);
nor UO_290 (O_290,N_2080,N_2187);
and UO_291 (O_291,N_2898,N_2728);
or UO_292 (O_292,N_2443,N_2194);
or UO_293 (O_293,N_2361,N_2528);
xnor UO_294 (O_294,N_2727,N_2911);
xnor UO_295 (O_295,N_2399,N_2547);
or UO_296 (O_296,N_2393,N_2343);
or UO_297 (O_297,N_2477,N_2824);
nor UO_298 (O_298,N_2481,N_2153);
nand UO_299 (O_299,N_2626,N_2899);
xnor UO_300 (O_300,N_2933,N_2886);
nor UO_301 (O_301,N_2381,N_2493);
xor UO_302 (O_302,N_2467,N_2834);
and UO_303 (O_303,N_2536,N_2173);
xnor UO_304 (O_304,N_2885,N_2364);
xnor UO_305 (O_305,N_2537,N_2345);
or UO_306 (O_306,N_2265,N_2555);
nand UO_307 (O_307,N_2171,N_2144);
and UO_308 (O_308,N_2503,N_2321);
and UO_309 (O_309,N_2274,N_2065);
nor UO_310 (O_310,N_2028,N_2785);
and UO_311 (O_311,N_2000,N_2648);
and UO_312 (O_312,N_2851,N_2581);
nor UO_313 (O_313,N_2775,N_2832);
and UO_314 (O_314,N_2211,N_2906);
and UO_315 (O_315,N_2281,N_2383);
or UO_316 (O_316,N_2378,N_2741);
and UO_317 (O_317,N_2852,N_2332);
or UO_318 (O_318,N_2395,N_2060);
or UO_319 (O_319,N_2953,N_2391);
or UO_320 (O_320,N_2567,N_2630);
and UO_321 (O_321,N_2096,N_2590);
nor UO_322 (O_322,N_2516,N_2531);
and UO_323 (O_323,N_2278,N_2572);
and UO_324 (O_324,N_2843,N_2117);
nor UO_325 (O_325,N_2734,N_2056);
or UO_326 (O_326,N_2579,N_2561);
and UO_327 (O_327,N_2689,N_2921);
and UO_328 (O_328,N_2009,N_2654);
and UO_329 (O_329,N_2723,N_2363);
nand UO_330 (O_330,N_2148,N_2327);
nor UO_331 (O_331,N_2471,N_2844);
nor UO_332 (O_332,N_2887,N_2554);
xor UO_333 (O_333,N_2202,N_2696);
nand UO_334 (O_334,N_2695,N_2251);
nand UO_335 (O_335,N_2890,N_2415);
xnor UO_336 (O_336,N_2177,N_2097);
nor UO_337 (O_337,N_2569,N_2300);
nand UO_338 (O_338,N_2293,N_2315);
nand UO_339 (O_339,N_2883,N_2864);
and UO_340 (O_340,N_2126,N_2923);
nor UO_341 (O_341,N_2880,N_2167);
nand UO_342 (O_342,N_2974,N_2718);
xnor UO_343 (O_343,N_2517,N_2053);
and UO_344 (O_344,N_2725,N_2429);
nand UO_345 (O_345,N_2740,N_2419);
and UO_346 (O_346,N_2155,N_2860);
xnor UO_347 (O_347,N_2114,N_2521);
and UO_348 (O_348,N_2951,N_2189);
nor UO_349 (O_349,N_2291,N_2036);
nand UO_350 (O_350,N_2181,N_2984);
nor UO_351 (O_351,N_2675,N_2105);
nor UO_352 (O_352,N_2453,N_2709);
and UO_353 (O_353,N_2184,N_2513);
and UO_354 (O_354,N_2435,N_2404);
or UO_355 (O_355,N_2295,N_2495);
and UO_356 (O_356,N_2629,N_2766);
nor UO_357 (O_357,N_2083,N_2163);
nand UO_358 (O_358,N_2620,N_2809);
or UO_359 (O_359,N_2673,N_2998);
and UO_360 (O_360,N_2929,N_2582);
nand UO_361 (O_361,N_2591,N_2680);
nor UO_362 (O_362,N_2862,N_2088);
nand UO_363 (O_363,N_2780,N_2527);
nor UO_364 (O_364,N_2635,N_2120);
or UO_365 (O_365,N_2311,N_2489);
and UO_366 (O_366,N_2086,N_2352);
or UO_367 (O_367,N_2326,N_2006);
nand UO_368 (O_368,N_2990,N_2122);
xnor UO_369 (O_369,N_2355,N_2276);
nand UO_370 (O_370,N_2109,N_2336);
or UO_371 (O_371,N_2178,N_2917);
nand UO_372 (O_372,N_2588,N_2500);
and UO_373 (O_373,N_2935,N_2123);
nor UO_374 (O_374,N_2106,N_2980);
or UO_375 (O_375,N_2928,N_2949);
xor UO_376 (O_376,N_2052,N_2337);
and UO_377 (O_377,N_2920,N_2499);
nand UO_378 (O_378,N_2442,N_2458);
nand UO_379 (O_379,N_2116,N_2428);
nor UO_380 (O_380,N_2248,N_2487);
and UO_381 (O_381,N_2912,N_2801);
or UO_382 (O_382,N_2950,N_2339);
xnor UO_383 (O_383,N_2411,N_2684);
or UO_384 (O_384,N_2259,N_2410);
xnor UO_385 (O_385,N_2580,N_2903);
xor UO_386 (O_386,N_2722,N_2745);
nor UO_387 (O_387,N_2450,N_2342);
xor UO_388 (O_388,N_2524,N_2444);
nand UO_389 (O_389,N_2752,N_2070);
nor UO_390 (O_390,N_2439,N_2347);
xor UO_391 (O_391,N_2149,N_2633);
and UO_392 (O_392,N_2587,N_2711);
nand UO_393 (O_393,N_2246,N_2104);
nand UO_394 (O_394,N_2267,N_2947);
and UO_395 (O_395,N_2353,N_2394);
and UO_396 (O_396,N_2018,N_2763);
nor UO_397 (O_397,N_2318,N_2806);
and UO_398 (O_398,N_2872,N_2603);
or UO_399 (O_399,N_2108,N_2182);
nor UO_400 (O_400,N_2940,N_2369);
and UO_401 (O_401,N_2964,N_2997);
or UO_402 (O_402,N_2252,N_2214);
xor UO_403 (O_403,N_2146,N_2292);
xnor UO_404 (O_404,N_2936,N_2357);
nor UO_405 (O_405,N_2789,N_2045);
and UO_406 (O_406,N_2514,N_2641);
nor UO_407 (O_407,N_2143,N_2035);
nor UO_408 (O_408,N_2492,N_2565);
and UO_409 (O_409,N_2948,N_2652);
and UO_410 (O_410,N_2751,N_2707);
nand UO_411 (O_411,N_2350,N_2705);
xnor UO_412 (O_412,N_2666,N_2047);
xnor UO_413 (O_413,N_2421,N_2010);
nand UO_414 (O_414,N_2548,N_2710);
or UO_415 (O_415,N_2423,N_2437);
and UO_416 (O_416,N_2479,N_2771);
xor UO_417 (O_417,N_2161,N_2578);
and UO_418 (O_418,N_2678,N_2020);
nand UO_419 (O_419,N_2434,N_2941);
or UO_420 (O_420,N_2628,N_2041);
nor UO_421 (O_421,N_2055,N_2432);
or UO_422 (O_422,N_2985,N_2571);
xnor UO_423 (O_423,N_2279,N_2455);
and UO_424 (O_424,N_2227,N_2715);
nor UO_425 (O_425,N_2549,N_2786);
and UO_426 (O_426,N_2273,N_2484);
xor UO_427 (O_427,N_2607,N_2802);
nor UO_428 (O_428,N_2151,N_2358);
xor UO_429 (O_429,N_2634,N_2179);
xor UO_430 (O_430,N_2057,N_2659);
or UO_431 (O_431,N_2243,N_2216);
and UO_432 (O_432,N_2605,N_2842);
xnor UO_433 (O_433,N_2348,N_2396);
or UO_434 (O_434,N_2768,N_2306);
or UO_435 (O_435,N_2828,N_2005);
or UO_436 (O_436,N_2700,N_2239);
nand UO_437 (O_437,N_2800,N_2376);
nor UO_438 (O_438,N_2385,N_2174);
or UO_439 (O_439,N_2965,N_2970);
nor UO_440 (O_440,N_2677,N_2205);
and UO_441 (O_441,N_2231,N_2195);
xor UO_442 (O_442,N_2799,N_2313);
nand UO_443 (O_443,N_2922,N_2272);
nand UO_444 (O_444,N_2362,N_2615);
and UO_445 (O_445,N_2577,N_2820);
xor UO_446 (O_446,N_2221,N_2308);
and UO_447 (O_447,N_2051,N_2401);
and UO_448 (O_448,N_2433,N_2081);
xor UO_449 (O_449,N_2402,N_2374);
xnor UO_450 (O_450,N_2154,N_2314);
and UO_451 (O_451,N_2884,N_2468);
or UO_452 (O_452,N_2075,N_2712);
and UO_453 (O_453,N_2631,N_2367);
nor UO_454 (O_454,N_2341,N_2816);
nand UO_455 (O_455,N_2849,N_2466);
nor UO_456 (O_456,N_2606,N_2338);
or UO_457 (O_457,N_2131,N_2868);
nor UO_458 (O_458,N_2781,N_2084);
xnor UO_459 (O_459,N_2085,N_2330);
or UO_460 (O_460,N_2218,N_2124);
nand UO_461 (O_461,N_2042,N_2866);
xnor UO_462 (O_462,N_2379,N_2157);
and UO_463 (O_463,N_2129,N_2519);
nor UO_464 (O_464,N_2570,N_2406);
xnor UO_465 (O_465,N_2044,N_2782);
and UO_466 (O_466,N_2413,N_2795);
and UO_467 (O_467,N_2647,N_2743);
and UO_468 (O_468,N_2825,N_2765);
nor UO_469 (O_469,N_2839,N_2219);
xor UO_470 (O_470,N_2881,N_2201);
or UO_471 (O_471,N_2532,N_2387);
or UO_472 (O_472,N_2989,N_2613);
and UO_473 (O_473,N_2829,N_2529);
and UO_474 (O_474,N_2822,N_2879);
nand UO_475 (O_475,N_2841,N_2616);
nand UO_476 (O_476,N_2128,N_2576);
nand UO_477 (O_477,N_2749,N_2483);
nand UO_478 (O_478,N_2937,N_2486);
nand UO_479 (O_479,N_2978,N_2954);
xor UO_480 (O_480,N_2986,N_2335);
nor UO_481 (O_481,N_2043,N_2090);
or UO_482 (O_482,N_2427,N_2504);
or UO_483 (O_483,N_2366,N_2488);
nand UO_484 (O_484,N_2354,N_2508);
or UO_485 (O_485,N_2319,N_2003);
xor UO_486 (O_486,N_2063,N_2836);
nor UO_487 (O_487,N_2212,N_2287);
and UO_488 (O_488,N_2373,N_2232);
and UO_489 (O_489,N_2169,N_2724);
and UO_490 (O_490,N_2015,N_2333);
nor UO_491 (O_491,N_2901,N_2533);
nand UO_492 (O_492,N_2449,N_2445);
nor UO_493 (O_493,N_2963,N_2693);
nor UO_494 (O_494,N_2183,N_2714);
nand UO_495 (O_495,N_2422,N_2541);
nor UO_496 (O_496,N_2420,N_2031);
or UO_497 (O_497,N_2416,N_2960);
xor UO_498 (O_498,N_2662,N_2683);
nand UO_499 (O_499,N_2622,N_2656);
endmodule