module basic_750_5000_1000_50_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_656,In_431);
xor U1 (N_1,In_627,In_718);
nor U2 (N_2,In_318,In_104);
nand U3 (N_3,In_412,In_187);
nor U4 (N_4,In_630,In_554);
nor U5 (N_5,In_542,In_138);
nand U6 (N_6,In_529,In_15);
and U7 (N_7,In_163,In_514);
and U8 (N_8,In_18,In_705);
nor U9 (N_9,In_308,In_592);
xor U10 (N_10,In_657,In_22);
or U11 (N_11,In_570,In_80);
xnor U12 (N_12,In_414,In_694);
and U13 (N_13,In_714,In_648);
nand U14 (N_14,In_75,In_443);
or U15 (N_15,In_739,In_241);
nand U16 (N_16,In_321,In_229);
xor U17 (N_17,In_166,In_237);
nand U18 (N_18,In_181,In_496);
nor U19 (N_19,In_84,In_268);
nor U20 (N_20,In_704,In_549);
xor U21 (N_21,In_30,In_196);
or U22 (N_22,In_48,In_668);
xor U23 (N_23,In_628,In_482);
and U24 (N_24,In_429,In_493);
or U25 (N_25,In_355,In_591);
nand U26 (N_26,In_349,In_449);
nand U27 (N_27,In_444,In_541);
or U28 (N_28,In_586,In_117);
and U29 (N_29,In_233,In_525);
nand U30 (N_30,In_463,In_157);
or U31 (N_31,In_269,In_722);
or U32 (N_32,In_122,In_40);
or U33 (N_33,In_597,In_401);
xor U34 (N_34,In_235,In_400);
or U35 (N_35,In_97,In_361);
xnor U36 (N_36,In_475,In_394);
or U37 (N_37,In_484,In_527);
or U38 (N_38,In_497,In_596);
xor U39 (N_39,In_639,In_370);
xor U40 (N_40,In_43,In_650);
nor U41 (N_41,In_425,In_142);
nor U42 (N_42,In_430,In_141);
and U43 (N_43,In_432,In_248);
nand U44 (N_44,In_252,In_522);
or U45 (N_45,In_28,In_683);
nand U46 (N_46,In_659,In_682);
or U47 (N_47,In_615,In_297);
and U48 (N_48,In_69,In_508);
and U49 (N_49,In_93,In_372);
nand U50 (N_50,In_144,In_102);
xor U51 (N_51,In_261,In_510);
nand U52 (N_52,In_366,In_505);
or U53 (N_53,In_538,In_222);
nor U54 (N_54,In_500,In_553);
xnor U55 (N_55,In_31,In_346);
and U56 (N_56,In_253,In_576);
nand U57 (N_57,In_748,In_292);
and U58 (N_58,In_531,In_2);
nand U59 (N_59,In_495,In_384);
xnor U60 (N_60,In_691,In_634);
nor U61 (N_61,In_280,In_464);
nand U62 (N_62,In_119,In_378);
and U63 (N_63,In_127,In_621);
nor U64 (N_64,In_582,In_109);
and U65 (N_65,In_351,In_546);
nor U66 (N_66,In_534,In_439);
or U67 (N_67,In_338,In_712);
xor U68 (N_68,In_204,In_289);
xnor U69 (N_69,In_502,In_517);
and U70 (N_70,In_695,In_25);
and U71 (N_71,In_573,In_279);
nand U72 (N_72,In_106,In_152);
nand U73 (N_73,In_640,In_353);
xnor U74 (N_74,In_710,In_636);
nand U75 (N_75,In_588,In_348);
and U76 (N_76,In_317,In_281);
or U77 (N_77,In_260,In_337);
and U78 (N_78,In_175,In_479);
or U79 (N_79,In_651,In_571);
and U80 (N_80,In_96,In_134);
or U81 (N_81,In_539,In_188);
nor U82 (N_82,In_516,In_403);
or U83 (N_83,In_442,In_396);
or U84 (N_84,In_87,In_364);
nor U85 (N_85,In_202,In_362);
or U86 (N_86,In_558,In_247);
nor U87 (N_87,In_208,In_44);
nand U88 (N_88,In_115,In_267);
and U89 (N_89,In_226,In_619);
or U90 (N_90,In_397,In_552);
or U91 (N_91,In_580,In_740);
nand U92 (N_92,In_262,In_441);
nand U93 (N_93,In_209,In_72);
or U94 (N_94,In_437,In_277);
and U95 (N_95,In_551,In_713);
nor U96 (N_96,In_193,In_221);
nor U97 (N_97,In_41,In_742);
xor U98 (N_98,In_257,In_436);
nor U99 (N_99,In_426,In_136);
xor U100 (N_100,In_333,In_14);
xnor U101 (N_101,In_575,In_38);
nor U102 (N_102,In_206,In_164);
or U103 (N_103,In_697,In_563);
nor U104 (N_104,N_70,In_418);
and U105 (N_105,In_368,N_55);
nand U106 (N_106,N_35,N_51);
nor U107 (N_107,In_327,In_145);
nand U108 (N_108,In_335,In_275);
nand U109 (N_109,In_377,In_13);
xnor U110 (N_110,In_34,In_466);
and U111 (N_111,In_227,In_734);
xor U112 (N_112,In_618,In_322);
nor U113 (N_113,In_357,In_238);
nand U114 (N_114,In_10,In_339);
nand U115 (N_115,In_11,N_34);
xor U116 (N_116,In_33,In_293);
xnor U117 (N_117,In_744,In_32);
xnor U118 (N_118,In_191,In_453);
nor U119 (N_119,In_633,N_50);
nand U120 (N_120,In_27,In_194);
nand U121 (N_121,In_341,In_201);
xnor U122 (N_122,In_644,In_290);
and U123 (N_123,In_524,In_46);
and U124 (N_124,In_399,In_314);
nand U125 (N_125,N_30,In_489);
xnor U126 (N_126,In_245,In_8);
nand U127 (N_127,In_310,In_477);
or U128 (N_128,In_455,In_729);
nand U129 (N_129,In_60,In_133);
and U130 (N_130,In_675,In_79);
nor U131 (N_131,In_231,In_647);
nand U132 (N_132,In_66,In_398);
and U133 (N_133,In_78,In_402);
or U134 (N_134,In_182,In_203);
nand U135 (N_135,In_3,In_161);
nor U136 (N_136,N_99,N_38);
nor U137 (N_137,In_513,N_62);
nand U138 (N_138,N_29,In_602);
nor U139 (N_139,In_108,In_409);
or U140 (N_140,In_299,In_424);
and U141 (N_141,In_550,In_715);
and U142 (N_142,In_120,In_471);
or U143 (N_143,In_135,In_146);
xor U144 (N_144,In_730,In_434);
nand U145 (N_145,In_249,In_548);
or U146 (N_146,In_666,In_311);
nand U147 (N_147,In_47,In_223);
nor U148 (N_148,In_411,In_385);
nor U149 (N_149,In_143,In_658);
nand U150 (N_150,In_101,N_74);
xor U151 (N_151,In_124,N_57);
and U152 (N_152,In_719,In_218);
and U153 (N_153,In_153,In_460);
nor U154 (N_154,In_59,In_367);
or U155 (N_155,In_745,In_693);
nand U156 (N_156,In_200,In_230);
nor U157 (N_157,N_37,In_587);
nand U158 (N_158,In_701,In_741);
and U159 (N_159,N_83,In_149);
nor U160 (N_160,In_568,In_645);
nor U161 (N_161,In_100,In_506);
and U162 (N_162,N_9,In_560);
xnor U163 (N_163,N_7,In_649);
nand U164 (N_164,N_10,In_688);
or U165 (N_165,In_50,In_625);
nand U166 (N_166,In_438,In_601);
nor U167 (N_167,In_64,In_94);
nand U168 (N_168,In_51,N_45);
and U169 (N_169,In_259,In_356);
xor U170 (N_170,N_20,In_354);
and U171 (N_171,In_26,In_263);
nor U172 (N_172,In_670,In_234);
and U173 (N_173,N_40,In_557);
nand U174 (N_174,In_16,In_726);
nand U175 (N_175,In_749,In_156);
nand U176 (N_176,In_604,In_244);
nand U177 (N_177,In_129,In_663);
or U178 (N_178,In_501,In_448);
nor U179 (N_179,In_700,In_386);
or U180 (N_180,N_82,In_83);
xnor U181 (N_181,N_96,N_31);
nor U182 (N_182,In_283,In_265);
nand U183 (N_183,N_81,N_86);
and U184 (N_184,In_415,In_99);
or U185 (N_185,In_336,In_696);
or U186 (N_186,In_536,In_264);
nor U187 (N_187,In_492,In_105);
and U188 (N_188,In_476,In_637);
nor U189 (N_189,In_215,N_71);
nor U190 (N_190,N_60,In_556);
and U191 (N_191,In_147,In_232);
and U192 (N_192,In_139,In_90);
nor U193 (N_193,In_148,In_130);
xor U194 (N_194,In_583,N_84);
and U195 (N_195,N_72,In_428);
and U196 (N_196,In_315,In_211);
or U197 (N_197,In_172,In_302);
xnor U198 (N_198,In_114,N_75);
xnor U199 (N_199,N_98,N_42);
or U200 (N_200,In_427,In_388);
and U201 (N_201,In_251,In_521);
or U202 (N_202,N_47,N_6);
xnor U203 (N_203,N_92,In_155);
nand U204 (N_204,In_635,N_172);
or U205 (N_205,N_149,In_422);
nand U206 (N_206,In_89,In_612);
and U207 (N_207,N_25,In_125);
xnor U208 (N_208,In_532,In_594);
nor U209 (N_209,In_599,In_490);
or U210 (N_210,N_129,In_217);
and U211 (N_211,In_140,In_363);
nor U212 (N_212,N_16,In_390);
xnor U213 (N_213,In_486,In_53);
nand U214 (N_214,In_35,N_1);
xnor U215 (N_215,N_122,N_39);
and U216 (N_216,In_451,In_344);
or U217 (N_217,In_555,N_27);
and U218 (N_218,In_733,N_137);
xor U219 (N_219,In_373,In_665);
nor U220 (N_220,In_55,In_509);
xor U221 (N_221,In_503,In_306);
nand U222 (N_222,N_178,In_176);
or U223 (N_223,In_669,N_180);
nand U224 (N_224,N_186,N_170);
or U225 (N_225,In_562,In_52);
nand U226 (N_226,In_325,N_93);
or U227 (N_227,In_608,In_126);
nand U228 (N_228,N_28,N_103);
and U229 (N_229,N_53,In_512);
nor U230 (N_230,In_36,In_76);
xor U231 (N_231,N_118,In_408);
nor U232 (N_232,In_447,In_452);
nand U233 (N_233,In_242,In_585);
nor U234 (N_234,In_676,N_156);
nor U235 (N_235,In_199,In_481);
or U236 (N_236,In_123,N_18);
nand U237 (N_237,N_148,N_36);
xor U238 (N_238,In_685,N_65);
nor U239 (N_239,N_67,In_56);
and U240 (N_240,In_724,In_620);
or U241 (N_241,In_407,In_5);
nor U242 (N_242,N_79,In_326);
nand U243 (N_243,In_660,N_183);
nor U244 (N_244,In_622,N_187);
xnor U245 (N_245,N_163,In_699);
or U246 (N_246,In_276,In_567);
xor U247 (N_247,N_134,In_406);
or U248 (N_248,In_365,N_115);
nand U249 (N_249,In_708,N_164);
nand U250 (N_250,In_111,N_44);
and U251 (N_251,In_116,In_731);
nor U252 (N_252,N_123,N_193);
nor U253 (N_253,N_26,In_375);
xnor U254 (N_254,N_117,In_716);
or U255 (N_255,In_255,N_77);
or U256 (N_256,In_530,N_155);
or U257 (N_257,In_154,In_271);
nor U258 (N_258,In_137,In_369);
and U259 (N_259,In_273,In_379);
nor U260 (N_260,N_4,In_473);
nand U261 (N_261,In_65,In_494);
xor U262 (N_262,N_197,In_721);
nand U263 (N_263,In_632,In_313);
or U264 (N_264,N_141,In_616);
nand U265 (N_265,In_684,N_56);
nor U266 (N_266,In_345,In_171);
nand U267 (N_267,N_23,In_667);
xor U268 (N_268,N_24,N_184);
xnor U269 (N_269,N_21,In_340);
and U270 (N_270,In_646,In_746);
or U271 (N_271,In_7,In_214);
nor U272 (N_272,In_186,In_499);
and U273 (N_273,N_12,In_631);
xor U274 (N_274,In_23,N_135);
xnor U275 (N_275,In_81,In_461);
or U276 (N_276,N_119,N_124);
xor U277 (N_277,N_32,In_416);
nand U278 (N_278,In_711,In_526);
nand U279 (N_279,In_160,In_605);
nor U280 (N_280,In_507,N_150);
nor U281 (N_281,N_152,In_284);
or U282 (N_282,N_132,In_286);
xnor U283 (N_283,N_173,N_109);
xnor U284 (N_284,N_159,In_57);
or U285 (N_285,In_296,In_282);
nor U286 (N_286,N_113,In_165);
or U287 (N_287,N_61,In_572);
xor U288 (N_288,In_421,In_528);
nor U289 (N_289,N_89,N_140);
nor U290 (N_290,In_566,In_70);
nor U291 (N_291,N_46,In_504);
nor U292 (N_292,N_154,N_151);
xnor U293 (N_293,N_13,In_167);
xnor U294 (N_294,In_62,In_178);
or U295 (N_295,In_545,N_106);
and U296 (N_296,In_488,In_598);
xor U297 (N_297,In_653,In_19);
nand U298 (N_298,In_158,In_435);
or U299 (N_299,N_69,In_458);
nand U300 (N_300,N_213,N_284);
nand U301 (N_301,In_274,In_298);
nand U302 (N_302,N_203,N_139);
nor U303 (N_303,N_282,In_417);
and U304 (N_304,In_638,In_564);
and U305 (N_305,N_285,In_450);
and U306 (N_306,In_626,N_259);
or U307 (N_307,In_595,In_641);
nand U308 (N_308,N_162,N_297);
or U309 (N_309,In_547,In_332);
nand U310 (N_310,In_1,N_97);
or U311 (N_311,N_226,N_52);
and U312 (N_312,In_291,N_271);
nor U313 (N_313,N_225,In_391);
and U314 (N_314,N_205,N_209);
nor U315 (N_315,In_270,In_679);
and U316 (N_316,In_86,In_459);
or U317 (N_317,In_12,In_629);
or U318 (N_318,In_523,In_623);
or U319 (N_319,In_617,In_183);
or U320 (N_320,N_239,N_232);
nor U321 (N_321,In_518,In_686);
nand U322 (N_322,In_383,In_128);
or U323 (N_323,In_216,N_112);
xnor U324 (N_324,N_107,In_39);
nor U325 (N_325,In_738,In_9);
xnor U326 (N_326,In_743,In_423);
nor U327 (N_327,In_358,In_577);
xnor U328 (N_328,N_78,N_263);
xnor U329 (N_329,N_298,N_66);
nand U330 (N_330,N_276,In_454);
nor U331 (N_331,N_176,N_182);
nor U332 (N_332,In_170,In_574);
xor U333 (N_333,In_520,In_457);
nor U334 (N_334,N_288,N_17);
or U335 (N_335,N_270,N_102);
and U336 (N_336,N_269,In_288);
nor U337 (N_337,In_687,N_181);
nor U338 (N_338,N_262,In_74);
xor U339 (N_339,In_278,N_90);
nand U340 (N_340,In_258,In_17);
or U341 (N_341,N_299,N_255);
and U342 (N_342,In_533,N_231);
xnor U343 (N_343,In_413,N_188);
or U344 (N_344,N_174,In_329);
or U345 (N_345,N_33,N_260);
xor U346 (N_346,N_167,In_614);
xor U347 (N_347,In_150,N_22);
and U348 (N_348,In_680,N_126);
and U349 (N_349,In_540,In_728);
nor U350 (N_350,In_462,In_88);
and U351 (N_351,In_295,In_184);
and U352 (N_352,N_100,N_206);
or U353 (N_353,N_168,N_292);
xnor U354 (N_354,In_236,In_698);
or U355 (N_355,In_467,N_41);
nor U356 (N_356,N_281,N_295);
xnor U357 (N_357,N_216,N_198);
or U358 (N_358,In_6,In_590);
nor U359 (N_359,N_287,In_674);
xnor U360 (N_360,In_323,In_350);
and U361 (N_361,In_535,In_82);
nand U362 (N_362,In_690,In_611);
xor U363 (N_363,N_220,N_114);
nor U364 (N_364,In_440,N_166);
or U365 (N_365,N_8,N_202);
nor U366 (N_366,In_581,In_519);
nand U367 (N_367,N_131,In_543);
and U368 (N_368,N_95,N_235);
or U369 (N_369,In_132,In_382);
and U370 (N_370,In_256,N_64);
nand U371 (N_371,N_175,N_251);
xor U372 (N_372,In_266,In_703);
or U373 (N_373,In_707,In_747);
or U374 (N_374,N_294,N_48);
nor U375 (N_375,In_254,N_63);
nand U376 (N_376,N_91,In_374);
xor U377 (N_377,N_219,N_19);
nand U378 (N_378,N_236,In_228);
xnor U379 (N_379,N_240,N_212);
or U380 (N_380,N_179,N_234);
nand U381 (N_381,N_49,N_241);
or U382 (N_382,N_272,N_215);
nor U383 (N_383,In_446,N_254);
and U384 (N_384,In_624,In_304);
nand U385 (N_385,In_73,In_29);
and U386 (N_386,In_515,N_111);
and U387 (N_387,In_285,N_116);
nand U388 (N_388,In_118,In_702);
nor U389 (N_389,In_607,N_273);
or U390 (N_390,In_192,In_312);
and U391 (N_391,N_143,In_359);
and U392 (N_392,In_643,In_709);
nor U393 (N_393,In_190,In_381);
or U394 (N_394,In_664,N_125);
xor U395 (N_395,N_199,In_606);
and U396 (N_396,In_672,In_21);
or U397 (N_397,N_138,In_389);
xor U398 (N_398,In_307,N_153);
nand U399 (N_399,N_160,N_246);
xnor U400 (N_400,N_320,In_376);
or U401 (N_401,N_247,In_420);
or U402 (N_402,N_108,In_207);
and U403 (N_403,In_294,N_300);
nand U404 (N_404,In_405,In_24);
or U405 (N_405,N_303,N_275);
nand U406 (N_406,N_353,In_395);
nand U407 (N_407,In_37,In_272);
nor U408 (N_408,In_578,In_661);
xnor U409 (N_409,N_369,N_323);
nand U410 (N_410,In_305,In_303);
nor U411 (N_411,N_265,In_95);
or U412 (N_412,N_194,In_565);
xor U413 (N_413,N_238,N_195);
nand U414 (N_414,In_85,In_92);
nor U415 (N_415,N_296,In_469);
nand U416 (N_416,In_246,N_157);
nor U417 (N_417,In_67,N_110);
or U418 (N_418,N_347,In_107);
nand U419 (N_419,N_261,N_346);
xor U420 (N_420,N_395,N_85);
or U421 (N_421,N_351,N_366);
and U422 (N_422,N_319,N_316);
nand U423 (N_423,N_229,N_3);
nor U424 (N_424,N_377,In_58);
and U425 (N_425,N_189,N_383);
nand U426 (N_426,In_706,N_222);
and U427 (N_427,N_399,N_248);
or U428 (N_428,N_249,In_681);
nand U429 (N_429,In_652,N_348);
and U430 (N_430,N_54,N_308);
xor U431 (N_431,In_677,In_225);
nand U432 (N_432,N_237,N_15);
nand U433 (N_433,N_207,N_368);
nor U434 (N_434,N_358,N_144);
xnor U435 (N_435,N_146,In_54);
and U436 (N_436,N_59,In_655);
and U437 (N_437,In_404,In_559);
nand U438 (N_438,N_228,In_342);
nor U439 (N_439,N_338,N_252);
and U440 (N_440,N_11,N_253);
and U441 (N_441,N_210,In_243);
nor U442 (N_442,In_671,N_373);
or U443 (N_443,In_309,In_723);
nor U444 (N_444,In_732,In_180);
or U445 (N_445,In_613,In_393);
or U446 (N_446,In_603,In_673);
nand U447 (N_447,In_220,In_205);
nand U448 (N_448,In_380,N_268);
or U449 (N_449,In_174,N_387);
nor U450 (N_450,In_537,N_283);
nand U451 (N_451,N_136,N_43);
xor U452 (N_452,N_190,N_76);
or U453 (N_453,N_333,In_360);
xnor U454 (N_454,N_344,N_214);
nand U455 (N_455,In_433,N_312);
nor U456 (N_456,In_470,In_20);
nor U457 (N_457,In_737,N_177);
xnor U458 (N_458,In_113,In_419);
nand U459 (N_459,N_267,N_349);
nand U460 (N_460,In_593,N_318);
nor U461 (N_461,N_289,N_374);
or U462 (N_462,N_329,In_544);
and U463 (N_463,N_356,N_58);
nand U464 (N_464,In_131,N_257);
nor U465 (N_465,In_456,N_359);
and U466 (N_466,N_342,N_200);
and U467 (N_467,N_304,N_2);
or U468 (N_468,N_171,In_168);
and U469 (N_469,N_0,In_121);
or U470 (N_470,In_487,In_330);
nor U471 (N_471,N_165,N_310);
or U472 (N_472,In_727,In_725);
or U473 (N_473,In_103,In_98);
nor U474 (N_474,In_169,N_365);
nor U475 (N_475,N_302,N_360);
xnor U476 (N_476,N_233,In_343);
and U477 (N_477,N_361,In_720);
nor U478 (N_478,N_397,N_370);
xnor U479 (N_479,N_381,N_80);
nor U480 (N_480,In_480,In_589);
xnor U481 (N_481,In_213,In_42);
xor U482 (N_482,In_445,N_309);
nor U483 (N_483,In_112,N_391);
or U484 (N_484,In_316,N_5);
xnor U485 (N_485,In_347,In_210);
xor U486 (N_486,N_73,In_179);
nand U487 (N_487,In_162,N_317);
xnor U488 (N_488,N_277,N_307);
xnor U489 (N_489,N_293,N_392);
and U490 (N_490,In_91,N_336);
xor U491 (N_491,In_662,N_221);
nand U492 (N_492,In_195,In_642);
nand U493 (N_493,In_600,N_389);
nand U494 (N_494,N_322,N_311);
nand U495 (N_495,N_133,N_379);
and U496 (N_496,In_224,N_121);
nor U497 (N_497,In_324,N_334);
or U498 (N_498,N_280,N_345);
nand U499 (N_499,N_208,N_367);
nor U500 (N_500,N_321,N_378);
xor U501 (N_501,In_177,N_414);
and U502 (N_502,N_423,N_415);
nor U503 (N_503,N_279,N_352);
xor U504 (N_504,In_579,N_455);
nor U505 (N_505,N_402,N_362);
nor U506 (N_506,N_404,N_419);
and U507 (N_507,N_488,N_459);
xor U508 (N_508,N_453,N_436);
and U509 (N_509,N_492,N_439);
or U510 (N_510,N_357,N_473);
xnor U511 (N_511,N_313,N_274);
nor U512 (N_512,N_458,N_230);
nand U513 (N_513,N_490,N_485);
xor U514 (N_514,In_485,In_474);
nor U515 (N_515,N_305,N_472);
and U516 (N_516,N_448,In_483);
nand U517 (N_517,In_219,N_486);
nand U518 (N_518,N_371,N_421);
nor U519 (N_519,N_407,In_240);
or U520 (N_520,N_426,N_196);
nor U521 (N_521,N_433,In_410);
nor U522 (N_522,N_393,N_211);
or U523 (N_523,N_330,N_244);
and U524 (N_524,N_364,N_68);
nand U525 (N_525,N_372,In_173);
and U526 (N_526,N_406,In_678);
or U527 (N_527,N_417,N_243);
xor U528 (N_528,N_185,In_472);
nand U529 (N_529,N_491,In_392);
xnor U530 (N_530,N_382,N_290);
xor U531 (N_531,N_14,N_227);
or U532 (N_532,In_735,N_420);
nor U533 (N_533,N_324,N_245);
nand U534 (N_534,N_489,In_498);
and U535 (N_535,In_151,N_158);
nand U536 (N_536,N_350,In_717);
and U537 (N_537,N_256,N_388);
nor U538 (N_538,In_569,N_478);
nand U539 (N_539,N_306,N_428);
or U540 (N_540,N_384,In_0);
or U541 (N_541,N_449,N_401);
or U542 (N_542,N_474,In_45);
nand U543 (N_543,N_468,N_408);
and U544 (N_544,In_239,N_94);
xnor U545 (N_545,In_561,N_441);
or U546 (N_546,N_482,N_412);
or U547 (N_547,N_437,N_130);
or U548 (N_548,In_212,In_68);
nand U549 (N_549,N_467,N_494);
nand U550 (N_550,In_300,N_444);
or U551 (N_551,N_440,N_487);
or U552 (N_552,In_250,In_328);
nand U553 (N_553,N_435,N_331);
and U554 (N_554,N_355,N_461);
xnor U555 (N_555,In_287,N_427);
nor U556 (N_556,N_496,N_454);
xnor U557 (N_557,N_477,N_470);
and U558 (N_558,N_396,N_484);
or U559 (N_559,N_405,N_169);
nand U560 (N_560,In_189,In_689);
nor U561 (N_561,In_49,In_4);
or U562 (N_562,N_264,N_464);
nor U563 (N_563,N_327,N_218);
nor U564 (N_564,N_340,N_410);
and U565 (N_565,In_159,N_498);
nand U566 (N_566,N_466,N_335);
xnor U567 (N_567,N_456,N_339);
and U568 (N_568,N_201,In_736);
and U569 (N_569,N_483,N_495);
and U570 (N_570,N_398,N_104);
nand U571 (N_571,N_325,N_416);
and U572 (N_572,N_314,N_462);
or U573 (N_573,N_88,N_409);
and U574 (N_574,N_443,N_403);
nor U575 (N_575,In_468,N_223);
or U576 (N_576,N_434,N_127);
xnor U577 (N_577,N_442,N_192);
and U578 (N_578,N_147,N_278);
nand U579 (N_579,In_110,In_491);
or U580 (N_580,N_204,N_445);
and U581 (N_581,N_286,N_469);
nor U582 (N_582,N_394,In_584);
xor U583 (N_583,N_424,In_610);
nand U584 (N_584,N_386,N_142);
nor U585 (N_585,N_217,N_250);
xnor U586 (N_586,N_326,N_258);
nand U587 (N_587,N_120,N_380);
and U588 (N_588,N_431,N_497);
nand U589 (N_589,N_224,In_478);
and U590 (N_590,In_71,N_479);
nand U591 (N_591,N_438,N_413);
xnor U592 (N_592,In_654,N_457);
nor U593 (N_593,N_128,N_465);
nand U594 (N_594,In_320,N_145);
nand U595 (N_595,N_463,N_446);
xnor U596 (N_596,N_101,N_432);
xnor U597 (N_597,In_334,N_450);
nand U598 (N_598,In_371,N_363);
xnor U599 (N_599,N_161,In_319);
xor U600 (N_600,In_609,N_525);
and U601 (N_601,In_511,In_692);
xor U602 (N_602,N_522,N_460);
nor U603 (N_603,N_588,N_545);
xor U604 (N_604,N_581,N_390);
or U605 (N_605,N_537,N_481);
or U606 (N_606,N_531,In_198);
nand U607 (N_607,N_575,N_541);
or U608 (N_608,In_63,N_564);
xnor U609 (N_609,N_480,N_563);
and U610 (N_610,N_505,N_514);
xnor U611 (N_611,N_573,N_337);
nor U612 (N_612,N_506,N_570);
xor U613 (N_613,N_552,N_593);
nand U614 (N_614,N_315,N_341);
nand U615 (N_615,N_569,In_465);
or U616 (N_616,N_551,N_536);
and U617 (N_617,N_567,N_538);
and U618 (N_618,N_429,N_447);
nand U619 (N_619,N_475,N_568);
xor U620 (N_620,In_77,N_559);
xnor U621 (N_621,N_580,N_534);
nand U622 (N_622,N_560,N_430);
nor U623 (N_623,N_515,N_594);
xnor U624 (N_624,N_596,N_558);
nand U625 (N_625,N_291,N_599);
xnor U626 (N_626,N_526,N_520);
or U627 (N_627,N_543,N_418);
or U628 (N_628,N_385,In_61);
nor U629 (N_629,N_519,N_535);
nand U630 (N_630,N_509,In_301);
xor U631 (N_631,N_577,N_562);
xnor U632 (N_632,N_571,N_533);
nand U633 (N_633,N_493,In_197);
or U634 (N_634,N_583,N_516);
nand U635 (N_635,N_502,N_343);
and U636 (N_636,N_511,N_266);
nor U637 (N_637,N_504,N_574);
and U638 (N_638,N_422,N_555);
nor U639 (N_639,N_576,N_532);
nor U640 (N_640,N_523,N_510);
xnor U641 (N_641,N_354,In_185);
nor U642 (N_642,N_507,N_530);
and U643 (N_643,N_549,N_452);
and U644 (N_644,N_579,N_553);
nor U645 (N_645,N_595,N_554);
nand U646 (N_646,N_550,N_513);
nor U647 (N_647,N_556,N_425);
xnor U648 (N_648,N_561,N_546);
nand U649 (N_649,N_566,N_565);
nor U650 (N_650,N_527,N_521);
and U651 (N_651,N_517,N_585);
nand U652 (N_652,N_587,N_592);
or U653 (N_653,N_590,N_528);
or U654 (N_654,N_524,N_301);
nor U655 (N_655,N_589,N_508);
nand U656 (N_656,N_548,N_191);
or U657 (N_657,N_501,In_352);
nor U658 (N_658,N_544,N_332);
xor U659 (N_659,N_578,N_411);
and U660 (N_660,N_376,N_512);
nand U661 (N_661,N_582,N_542);
or U662 (N_662,N_584,In_331);
nand U663 (N_663,N_591,N_529);
xor U664 (N_664,N_503,N_500);
nor U665 (N_665,N_499,N_539);
nand U666 (N_666,N_547,N_598);
nand U667 (N_667,N_375,N_586);
xnor U668 (N_668,In_387,N_328);
nand U669 (N_669,N_105,N_451);
or U670 (N_670,N_518,N_540);
xnor U671 (N_671,N_471,N_87);
and U672 (N_672,N_572,N_476);
and U673 (N_673,N_597,N_400);
xnor U674 (N_674,N_242,N_557);
nor U675 (N_675,N_588,N_503);
nor U676 (N_676,N_593,N_567);
nor U677 (N_677,N_594,N_242);
nand U678 (N_678,N_589,N_571);
or U679 (N_679,N_527,N_341);
xnor U680 (N_680,N_425,N_516);
nand U681 (N_681,N_301,In_61);
nor U682 (N_682,N_594,N_551);
nor U683 (N_683,N_572,N_536);
nand U684 (N_684,N_585,N_592);
nor U685 (N_685,N_521,N_514);
and U686 (N_686,N_572,N_341);
or U687 (N_687,N_546,N_530);
and U688 (N_688,N_594,N_568);
nand U689 (N_689,N_475,N_541);
and U690 (N_690,N_507,N_547);
nand U691 (N_691,N_525,N_587);
xor U692 (N_692,N_566,N_516);
nand U693 (N_693,N_515,N_505);
nand U694 (N_694,N_519,N_542);
nor U695 (N_695,N_447,N_547);
xnor U696 (N_696,N_291,N_343);
nor U697 (N_697,N_354,N_594);
nand U698 (N_698,N_578,In_331);
xor U699 (N_699,N_592,N_597);
or U700 (N_700,N_622,N_686);
or U701 (N_701,N_627,N_677);
and U702 (N_702,N_668,N_632);
nand U703 (N_703,N_660,N_682);
xor U704 (N_704,N_626,N_631);
nand U705 (N_705,N_689,N_678);
or U706 (N_706,N_623,N_643);
nor U707 (N_707,N_697,N_640);
nand U708 (N_708,N_685,N_629);
or U709 (N_709,N_617,N_634);
or U710 (N_710,N_679,N_610);
and U711 (N_711,N_644,N_699);
nand U712 (N_712,N_606,N_664);
or U713 (N_713,N_661,N_618);
nor U714 (N_714,N_654,N_601);
and U715 (N_715,N_615,N_662);
nor U716 (N_716,N_674,N_665);
or U717 (N_717,N_655,N_688);
nand U718 (N_718,N_695,N_624);
or U719 (N_719,N_619,N_628);
or U720 (N_720,N_646,N_648);
or U721 (N_721,N_651,N_671);
nor U722 (N_722,N_639,N_692);
nor U723 (N_723,N_659,N_611);
nand U724 (N_724,N_653,N_636);
nor U725 (N_725,N_667,N_652);
or U726 (N_726,N_683,N_684);
xnor U727 (N_727,N_608,N_620);
xnor U728 (N_728,N_600,N_672);
or U729 (N_729,N_616,N_604);
nand U730 (N_730,N_613,N_656);
nand U731 (N_731,N_669,N_630);
and U732 (N_732,N_657,N_649);
or U733 (N_733,N_658,N_625);
nand U734 (N_734,N_666,N_609);
and U735 (N_735,N_621,N_693);
and U736 (N_736,N_663,N_633);
and U737 (N_737,N_675,N_676);
xor U738 (N_738,N_614,N_687);
nor U739 (N_739,N_612,N_603);
nand U740 (N_740,N_650,N_670);
xnor U741 (N_741,N_637,N_647);
nor U742 (N_742,N_602,N_694);
or U743 (N_743,N_691,N_681);
nand U744 (N_744,N_605,N_642);
or U745 (N_745,N_645,N_673);
nor U746 (N_746,N_698,N_696);
or U747 (N_747,N_638,N_690);
xnor U748 (N_748,N_680,N_641);
xnor U749 (N_749,N_635,N_607);
nand U750 (N_750,N_697,N_656);
or U751 (N_751,N_672,N_642);
nor U752 (N_752,N_695,N_656);
nor U753 (N_753,N_662,N_672);
nor U754 (N_754,N_643,N_652);
and U755 (N_755,N_665,N_613);
or U756 (N_756,N_636,N_658);
xor U757 (N_757,N_632,N_620);
nand U758 (N_758,N_615,N_613);
xor U759 (N_759,N_603,N_627);
xor U760 (N_760,N_669,N_696);
xnor U761 (N_761,N_654,N_699);
and U762 (N_762,N_623,N_670);
nor U763 (N_763,N_628,N_604);
nor U764 (N_764,N_661,N_628);
nor U765 (N_765,N_636,N_695);
xnor U766 (N_766,N_659,N_684);
nor U767 (N_767,N_694,N_618);
xor U768 (N_768,N_661,N_604);
nor U769 (N_769,N_627,N_672);
nor U770 (N_770,N_641,N_615);
nand U771 (N_771,N_611,N_609);
nor U772 (N_772,N_606,N_696);
or U773 (N_773,N_620,N_616);
xnor U774 (N_774,N_681,N_674);
and U775 (N_775,N_658,N_698);
nor U776 (N_776,N_629,N_694);
and U777 (N_777,N_612,N_668);
or U778 (N_778,N_682,N_650);
and U779 (N_779,N_603,N_672);
or U780 (N_780,N_635,N_620);
nor U781 (N_781,N_611,N_657);
or U782 (N_782,N_678,N_693);
nand U783 (N_783,N_688,N_613);
and U784 (N_784,N_611,N_631);
and U785 (N_785,N_607,N_684);
xnor U786 (N_786,N_674,N_686);
and U787 (N_787,N_632,N_614);
nor U788 (N_788,N_673,N_661);
nand U789 (N_789,N_609,N_645);
nor U790 (N_790,N_614,N_631);
nand U791 (N_791,N_653,N_662);
and U792 (N_792,N_649,N_664);
nor U793 (N_793,N_629,N_697);
nor U794 (N_794,N_613,N_676);
nand U795 (N_795,N_642,N_621);
nor U796 (N_796,N_643,N_680);
and U797 (N_797,N_671,N_665);
and U798 (N_798,N_664,N_659);
xor U799 (N_799,N_617,N_602);
nor U800 (N_800,N_707,N_724);
xor U801 (N_801,N_711,N_720);
and U802 (N_802,N_727,N_781);
nand U803 (N_803,N_732,N_700);
and U804 (N_804,N_706,N_744);
xor U805 (N_805,N_758,N_779);
and U806 (N_806,N_729,N_756);
xnor U807 (N_807,N_731,N_703);
xnor U808 (N_808,N_785,N_760);
and U809 (N_809,N_735,N_768);
and U810 (N_810,N_784,N_789);
xnor U811 (N_811,N_728,N_723);
nand U812 (N_812,N_701,N_775);
nor U813 (N_813,N_786,N_733);
xor U814 (N_814,N_738,N_797);
xnor U815 (N_815,N_763,N_777);
nor U816 (N_816,N_765,N_726);
xnor U817 (N_817,N_766,N_799);
nor U818 (N_818,N_746,N_709);
and U819 (N_819,N_773,N_712);
nand U820 (N_820,N_741,N_754);
and U821 (N_821,N_740,N_750);
xnor U822 (N_822,N_755,N_713);
nand U823 (N_823,N_788,N_761);
nor U824 (N_824,N_708,N_734);
nand U825 (N_825,N_783,N_798);
nor U826 (N_826,N_771,N_796);
xor U827 (N_827,N_751,N_717);
xnor U828 (N_828,N_743,N_742);
nor U829 (N_829,N_792,N_759);
xnor U830 (N_830,N_791,N_721);
or U831 (N_831,N_714,N_718);
nand U832 (N_832,N_794,N_767);
nor U833 (N_833,N_782,N_764);
xnor U834 (N_834,N_745,N_749);
nand U835 (N_835,N_736,N_705);
nand U836 (N_836,N_772,N_722);
or U837 (N_837,N_780,N_715);
nand U838 (N_838,N_716,N_702);
and U839 (N_839,N_757,N_704);
or U840 (N_840,N_769,N_710);
nand U841 (N_841,N_795,N_752);
xor U842 (N_842,N_739,N_787);
and U843 (N_843,N_719,N_776);
nor U844 (N_844,N_774,N_730);
nand U845 (N_845,N_793,N_790);
xor U846 (N_846,N_753,N_748);
nor U847 (N_847,N_770,N_762);
and U848 (N_848,N_778,N_725);
xnor U849 (N_849,N_747,N_737);
nor U850 (N_850,N_785,N_745);
and U851 (N_851,N_700,N_727);
nor U852 (N_852,N_764,N_778);
and U853 (N_853,N_763,N_796);
nand U854 (N_854,N_721,N_742);
and U855 (N_855,N_739,N_798);
nand U856 (N_856,N_711,N_736);
nor U857 (N_857,N_716,N_730);
nand U858 (N_858,N_785,N_766);
and U859 (N_859,N_759,N_723);
nand U860 (N_860,N_728,N_739);
or U861 (N_861,N_707,N_730);
or U862 (N_862,N_716,N_768);
nor U863 (N_863,N_770,N_748);
and U864 (N_864,N_711,N_722);
and U865 (N_865,N_776,N_743);
and U866 (N_866,N_797,N_768);
nor U867 (N_867,N_741,N_758);
nor U868 (N_868,N_756,N_711);
or U869 (N_869,N_714,N_746);
nand U870 (N_870,N_740,N_747);
xnor U871 (N_871,N_758,N_707);
nand U872 (N_872,N_713,N_798);
nor U873 (N_873,N_704,N_762);
or U874 (N_874,N_756,N_704);
xnor U875 (N_875,N_730,N_732);
and U876 (N_876,N_778,N_775);
or U877 (N_877,N_795,N_797);
nor U878 (N_878,N_742,N_723);
nor U879 (N_879,N_760,N_787);
or U880 (N_880,N_749,N_707);
nand U881 (N_881,N_756,N_735);
nand U882 (N_882,N_715,N_746);
and U883 (N_883,N_729,N_771);
nor U884 (N_884,N_716,N_763);
nand U885 (N_885,N_792,N_725);
nand U886 (N_886,N_714,N_787);
nand U887 (N_887,N_768,N_778);
or U888 (N_888,N_736,N_714);
or U889 (N_889,N_725,N_740);
and U890 (N_890,N_741,N_747);
and U891 (N_891,N_743,N_730);
nor U892 (N_892,N_788,N_757);
xor U893 (N_893,N_756,N_730);
and U894 (N_894,N_767,N_789);
nand U895 (N_895,N_715,N_709);
nand U896 (N_896,N_790,N_748);
nor U897 (N_897,N_742,N_726);
xor U898 (N_898,N_775,N_777);
xnor U899 (N_899,N_769,N_757);
nand U900 (N_900,N_893,N_807);
nand U901 (N_901,N_874,N_882);
xnor U902 (N_902,N_838,N_822);
or U903 (N_903,N_891,N_832);
nand U904 (N_904,N_870,N_894);
and U905 (N_905,N_873,N_829);
nand U906 (N_906,N_876,N_869);
xor U907 (N_907,N_821,N_812);
and U908 (N_908,N_826,N_802);
xor U909 (N_909,N_849,N_806);
nor U910 (N_910,N_872,N_848);
nor U911 (N_911,N_845,N_879);
nor U912 (N_912,N_881,N_840);
nor U913 (N_913,N_864,N_871);
or U914 (N_914,N_813,N_839);
or U915 (N_915,N_854,N_837);
xnor U916 (N_916,N_867,N_842);
xnor U917 (N_917,N_835,N_805);
nor U918 (N_918,N_863,N_841);
nand U919 (N_919,N_819,N_852);
and U920 (N_920,N_817,N_823);
nand U921 (N_921,N_833,N_804);
or U922 (N_922,N_898,N_855);
nand U923 (N_923,N_814,N_801);
xor U924 (N_924,N_883,N_824);
or U925 (N_925,N_857,N_808);
nand U926 (N_926,N_811,N_856);
nand U927 (N_927,N_830,N_853);
or U928 (N_928,N_896,N_892);
nor U929 (N_929,N_800,N_899);
or U930 (N_930,N_831,N_834);
and U931 (N_931,N_816,N_858);
or U932 (N_932,N_868,N_884);
nor U933 (N_933,N_820,N_846);
and U934 (N_934,N_862,N_803);
xor U935 (N_935,N_861,N_825);
xnor U936 (N_936,N_827,N_860);
nand U937 (N_937,N_815,N_818);
nand U938 (N_938,N_836,N_859);
and U939 (N_939,N_844,N_897);
or U940 (N_940,N_875,N_889);
xnor U941 (N_941,N_895,N_885);
nand U942 (N_942,N_810,N_843);
or U943 (N_943,N_887,N_847);
xnor U944 (N_944,N_866,N_888);
nor U945 (N_945,N_865,N_851);
nor U946 (N_946,N_809,N_886);
nor U947 (N_947,N_880,N_890);
and U948 (N_948,N_877,N_878);
nor U949 (N_949,N_828,N_850);
and U950 (N_950,N_861,N_873);
xnor U951 (N_951,N_810,N_817);
or U952 (N_952,N_807,N_881);
and U953 (N_953,N_812,N_873);
and U954 (N_954,N_800,N_898);
nand U955 (N_955,N_879,N_858);
or U956 (N_956,N_859,N_863);
and U957 (N_957,N_840,N_890);
xnor U958 (N_958,N_827,N_805);
nor U959 (N_959,N_805,N_868);
nand U960 (N_960,N_887,N_807);
and U961 (N_961,N_842,N_868);
nand U962 (N_962,N_845,N_858);
nand U963 (N_963,N_881,N_876);
nor U964 (N_964,N_807,N_876);
nor U965 (N_965,N_800,N_837);
or U966 (N_966,N_886,N_841);
and U967 (N_967,N_820,N_826);
or U968 (N_968,N_804,N_818);
xor U969 (N_969,N_837,N_887);
nor U970 (N_970,N_885,N_858);
nor U971 (N_971,N_861,N_806);
xor U972 (N_972,N_843,N_825);
xor U973 (N_973,N_865,N_875);
nor U974 (N_974,N_824,N_872);
nor U975 (N_975,N_806,N_862);
xor U976 (N_976,N_847,N_822);
xnor U977 (N_977,N_807,N_875);
or U978 (N_978,N_858,N_871);
nor U979 (N_979,N_892,N_841);
xor U980 (N_980,N_846,N_866);
and U981 (N_981,N_879,N_899);
nor U982 (N_982,N_837,N_862);
nand U983 (N_983,N_802,N_818);
nand U984 (N_984,N_870,N_850);
and U985 (N_985,N_800,N_834);
and U986 (N_986,N_800,N_897);
nand U987 (N_987,N_884,N_855);
or U988 (N_988,N_863,N_886);
nor U989 (N_989,N_839,N_846);
xnor U990 (N_990,N_868,N_888);
nand U991 (N_991,N_859,N_885);
nand U992 (N_992,N_854,N_856);
nor U993 (N_993,N_885,N_824);
xor U994 (N_994,N_892,N_837);
nand U995 (N_995,N_822,N_882);
nand U996 (N_996,N_887,N_872);
and U997 (N_997,N_854,N_863);
nand U998 (N_998,N_825,N_819);
nor U999 (N_999,N_838,N_848);
xor U1000 (N_1000,N_973,N_993);
and U1001 (N_1001,N_976,N_962);
xor U1002 (N_1002,N_991,N_915);
and U1003 (N_1003,N_907,N_909);
or U1004 (N_1004,N_922,N_918);
or U1005 (N_1005,N_964,N_956);
xor U1006 (N_1006,N_946,N_903);
nand U1007 (N_1007,N_969,N_932);
xnor U1008 (N_1008,N_949,N_986);
and U1009 (N_1009,N_957,N_951);
nor U1010 (N_1010,N_975,N_988);
xnor U1011 (N_1011,N_917,N_960);
nand U1012 (N_1012,N_929,N_919);
nor U1013 (N_1013,N_979,N_965);
and U1014 (N_1014,N_924,N_998);
nor U1015 (N_1015,N_931,N_980);
or U1016 (N_1016,N_985,N_952);
nand U1017 (N_1017,N_983,N_926);
nand U1018 (N_1018,N_984,N_982);
nand U1019 (N_1019,N_959,N_941);
and U1020 (N_1020,N_910,N_923);
nor U1021 (N_1021,N_999,N_987);
nor U1022 (N_1022,N_958,N_936);
or U1023 (N_1023,N_934,N_968);
nor U1024 (N_1024,N_977,N_928);
and U1025 (N_1025,N_990,N_927);
or U1026 (N_1026,N_908,N_955);
and U1027 (N_1027,N_971,N_916);
xor U1028 (N_1028,N_981,N_950);
or U1029 (N_1029,N_992,N_914);
or U1030 (N_1030,N_948,N_944);
or U1031 (N_1031,N_940,N_904);
nand U1032 (N_1032,N_933,N_995);
xor U1033 (N_1033,N_989,N_930);
nor U1034 (N_1034,N_913,N_911);
nand U1035 (N_1035,N_994,N_978);
nor U1036 (N_1036,N_942,N_902);
nor U1037 (N_1037,N_974,N_953);
nand U1038 (N_1038,N_920,N_901);
nor U1039 (N_1039,N_947,N_935);
nand U1040 (N_1040,N_961,N_906);
nand U1041 (N_1041,N_945,N_966);
and U1042 (N_1042,N_905,N_925);
and U1043 (N_1043,N_939,N_970);
and U1044 (N_1044,N_943,N_937);
and U1045 (N_1045,N_954,N_997);
xnor U1046 (N_1046,N_921,N_963);
xor U1047 (N_1047,N_912,N_996);
and U1048 (N_1048,N_938,N_900);
and U1049 (N_1049,N_967,N_972);
or U1050 (N_1050,N_904,N_953);
nor U1051 (N_1051,N_907,N_968);
and U1052 (N_1052,N_920,N_951);
nand U1053 (N_1053,N_970,N_944);
xnor U1054 (N_1054,N_917,N_952);
or U1055 (N_1055,N_930,N_954);
nor U1056 (N_1056,N_921,N_994);
xor U1057 (N_1057,N_972,N_926);
and U1058 (N_1058,N_913,N_955);
or U1059 (N_1059,N_954,N_938);
or U1060 (N_1060,N_986,N_923);
and U1061 (N_1061,N_981,N_953);
and U1062 (N_1062,N_928,N_907);
and U1063 (N_1063,N_938,N_997);
or U1064 (N_1064,N_975,N_964);
xor U1065 (N_1065,N_971,N_965);
or U1066 (N_1066,N_998,N_967);
xor U1067 (N_1067,N_998,N_994);
nor U1068 (N_1068,N_930,N_983);
or U1069 (N_1069,N_997,N_983);
xnor U1070 (N_1070,N_968,N_984);
nand U1071 (N_1071,N_918,N_980);
nand U1072 (N_1072,N_984,N_981);
xor U1073 (N_1073,N_958,N_995);
xnor U1074 (N_1074,N_910,N_956);
and U1075 (N_1075,N_975,N_972);
nand U1076 (N_1076,N_955,N_965);
and U1077 (N_1077,N_947,N_930);
nand U1078 (N_1078,N_966,N_923);
nor U1079 (N_1079,N_947,N_949);
xor U1080 (N_1080,N_901,N_985);
nand U1081 (N_1081,N_990,N_973);
and U1082 (N_1082,N_926,N_942);
and U1083 (N_1083,N_982,N_900);
xor U1084 (N_1084,N_960,N_954);
and U1085 (N_1085,N_997,N_936);
nand U1086 (N_1086,N_981,N_961);
or U1087 (N_1087,N_972,N_927);
and U1088 (N_1088,N_993,N_992);
nand U1089 (N_1089,N_952,N_910);
or U1090 (N_1090,N_924,N_985);
or U1091 (N_1091,N_926,N_936);
or U1092 (N_1092,N_946,N_944);
nand U1093 (N_1093,N_919,N_915);
or U1094 (N_1094,N_983,N_939);
or U1095 (N_1095,N_971,N_967);
nor U1096 (N_1096,N_981,N_940);
or U1097 (N_1097,N_950,N_987);
nor U1098 (N_1098,N_953,N_920);
or U1099 (N_1099,N_983,N_987);
or U1100 (N_1100,N_1096,N_1066);
nor U1101 (N_1101,N_1026,N_1071);
nand U1102 (N_1102,N_1088,N_1091);
nor U1103 (N_1103,N_1075,N_1014);
nand U1104 (N_1104,N_1092,N_1017);
and U1105 (N_1105,N_1064,N_1070);
nand U1106 (N_1106,N_1034,N_1004);
nor U1107 (N_1107,N_1047,N_1054);
and U1108 (N_1108,N_1036,N_1097);
and U1109 (N_1109,N_1023,N_1062);
nor U1110 (N_1110,N_1039,N_1061);
nand U1111 (N_1111,N_1051,N_1006);
or U1112 (N_1112,N_1024,N_1065);
nor U1113 (N_1113,N_1030,N_1005);
xor U1114 (N_1114,N_1019,N_1059);
or U1115 (N_1115,N_1077,N_1080);
nand U1116 (N_1116,N_1067,N_1044);
nor U1117 (N_1117,N_1037,N_1053);
nand U1118 (N_1118,N_1015,N_1057);
nand U1119 (N_1119,N_1007,N_1031);
nor U1120 (N_1120,N_1073,N_1018);
xor U1121 (N_1121,N_1011,N_1008);
and U1122 (N_1122,N_1090,N_1046);
nor U1123 (N_1123,N_1093,N_1033);
nand U1124 (N_1124,N_1068,N_1016);
and U1125 (N_1125,N_1048,N_1042);
or U1126 (N_1126,N_1003,N_1086);
nand U1127 (N_1127,N_1083,N_1098);
xor U1128 (N_1128,N_1052,N_1069);
xor U1129 (N_1129,N_1040,N_1022);
nor U1130 (N_1130,N_1058,N_1087);
xor U1131 (N_1131,N_1095,N_1060);
and U1132 (N_1132,N_1082,N_1000);
nor U1133 (N_1133,N_1041,N_1055);
nor U1134 (N_1134,N_1038,N_1078);
or U1135 (N_1135,N_1063,N_1089);
nand U1136 (N_1136,N_1084,N_1076);
or U1137 (N_1137,N_1085,N_1021);
xnor U1138 (N_1138,N_1009,N_1079);
or U1139 (N_1139,N_1043,N_1081);
and U1140 (N_1140,N_1074,N_1072);
nor U1141 (N_1141,N_1002,N_1050);
xor U1142 (N_1142,N_1099,N_1025);
and U1143 (N_1143,N_1028,N_1045);
nand U1144 (N_1144,N_1094,N_1035);
or U1145 (N_1145,N_1049,N_1010);
and U1146 (N_1146,N_1012,N_1001);
or U1147 (N_1147,N_1056,N_1020);
xor U1148 (N_1148,N_1013,N_1032);
and U1149 (N_1149,N_1029,N_1027);
and U1150 (N_1150,N_1091,N_1060);
nand U1151 (N_1151,N_1065,N_1052);
or U1152 (N_1152,N_1078,N_1072);
or U1153 (N_1153,N_1091,N_1053);
xnor U1154 (N_1154,N_1059,N_1033);
and U1155 (N_1155,N_1044,N_1063);
nand U1156 (N_1156,N_1061,N_1046);
and U1157 (N_1157,N_1007,N_1035);
nand U1158 (N_1158,N_1084,N_1025);
or U1159 (N_1159,N_1049,N_1016);
and U1160 (N_1160,N_1094,N_1098);
or U1161 (N_1161,N_1047,N_1078);
nand U1162 (N_1162,N_1044,N_1068);
nand U1163 (N_1163,N_1063,N_1080);
and U1164 (N_1164,N_1062,N_1058);
or U1165 (N_1165,N_1033,N_1019);
xor U1166 (N_1166,N_1051,N_1097);
nor U1167 (N_1167,N_1084,N_1028);
and U1168 (N_1168,N_1001,N_1032);
nor U1169 (N_1169,N_1060,N_1093);
and U1170 (N_1170,N_1095,N_1008);
xnor U1171 (N_1171,N_1025,N_1064);
xor U1172 (N_1172,N_1009,N_1084);
or U1173 (N_1173,N_1075,N_1077);
and U1174 (N_1174,N_1044,N_1041);
nor U1175 (N_1175,N_1047,N_1015);
nand U1176 (N_1176,N_1035,N_1027);
or U1177 (N_1177,N_1054,N_1023);
nand U1178 (N_1178,N_1050,N_1007);
and U1179 (N_1179,N_1001,N_1078);
nor U1180 (N_1180,N_1046,N_1064);
or U1181 (N_1181,N_1093,N_1065);
or U1182 (N_1182,N_1014,N_1003);
or U1183 (N_1183,N_1078,N_1083);
and U1184 (N_1184,N_1092,N_1057);
or U1185 (N_1185,N_1017,N_1032);
and U1186 (N_1186,N_1048,N_1018);
xnor U1187 (N_1187,N_1085,N_1039);
nor U1188 (N_1188,N_1064,N_1097);
xnor U1189 (N_1189,N_1052,N_1083);
nor U1190 (N_1190,N_1097,N_1053);
or U1191 (N_1191,N_1096,N_1013);
and U1192 (N_1192,N_1053,N_1060);
nor U1193 (N_1193,N_1056,N_1078);
xor U1194 (N_1194,N_1045,N_1092);
and U1195 (N_1195,N_1094,N_1005);
and U1196 (N_1196,N_1069,N_1041);
or U1197 (N_1197,N_1060,N_1081);
or U1198 (N_1198,N_1015,N_1050);
and U1199 (N_1199,N_1089,N_1072);
or U1200 (N_1200,N_1120,N_1159);
nor U1201 (N_1201,N_1101,N_1174);
and U1202 (N_1202,N_1123,N_1199);
nor U1203 (N_1203,N_1129,N_1157);
and U1204 (N_1204,N_1190,N_1164);
and U1205 (N_1205,N_1156,N_1127);
and U1206 (N_1206,N_1138,N_1134);
or U1207 (N_1207,N_1109,N_1185);
or U1208 (N_1208,N_1105,N_1113);
nor U1209 (N_1209,N_1178,N_1128);
nor U1210 (N_1210,N_1132,N_1151);
or U1211 (N_1211,N_1126,N_1144);
xnor U1212 (N_1212,N_1106,N_1116);
or U1213 (N_1213,N_1167,N_1114);
and U1214 (N_1214,N_1158,N_1107);
nand U1215 (N_1215,N_1170,N_1194);
nand U1216 (N_1216,N_1110,N_1141);
and U1217 (N_1217,N_1111,N_1108);
or U1218 (N_1218,N_1118,N_1176);
or U1219 (N_1219,N_1161,N_1188);
and U1220 (N_1220,N_1184,N_1149);
nand U1221 (N_1221,N_1104,N_1122);
and U1222 (N_1222,N_1154,N_1179);
xor U1223 (N_1223,N_1183,N_1115);
nor U1224 (N_1224,N_1139,N_1177);
and U1225 (N_1225,N_1192,N_1195);
nand U1226 (N_1226,N_1135,N_1133);
nand U1227 (N_1227,N_1163,N_1100);
xnor U1228 (N_1228,N_1166,N_1143);
nor U1229 (N_1229,N_1119,N_1112);
nand U1230 (N_1230,N_1169,N_1180);
or U1231 (N_1231,N_1137,N_1162);
nor U1232 (N_1232,N_1160,N_1136);
nand U1233 (N_1233,N_1124,N_1173);
and U1234 (N_1234,N_1196,N_1148);
xnor U1235 (N_1235,N_1172,N_1103);
or U1236 (N_1236,N_1165,N_1131);
nor U1237 (N_1237,N_1146,N_1125);
nor U1238 (N_1238,N_1191,N_1198);
or U1239 (N_1239,N_1168,N_1140);
or U1240 (N_1240,N_1153,N_1152);
xor U1241 (N_1241,N_1155,N_1117);
nor U1242 (N_1242,N_1121,N_1193);
nand U1243 (N_1243,N_1145,N_1181);
nor U1244 (N_1244,N_1197,N_1182);
nor U1245 (N_1245,N_1147,N_1187);
nand U1246 (N_1246,N_1102,N_1186);
and U1247 (N_1247,N_1171,N_1189);
xnor U1248 (N_1248,N_1130,N_1175);
or U1249 (N_1249,N_1150,N_1142);
nand U1250 (N_1250,N_1184,N_1182);
nand U1251 (N_1251,N_1185,N_1181);
xnor U1252 (N_1252,N_1131,N_1120);
and U1253 (N_1253,N_1124,N_1180);
and U1254 (N_1254,N_1135,N_1134);
xnor U1255 (N_1255,N_1161,N_1197);
nor U1256 (N_1256,N_1156,N_1114);
nand U1257 (N_1257,N_1105,N_1187);
and U1258 (N_1258,N_1168,N_1179);
xnor U1259 (N_1259,N_1136,N_1150);
or U1260 (N_1260,N_1139,N_1114);
xor U1261 (N_1261,N_1116,N_1144);
or U1262 (N_1262,N_1185,N_1179);
xor U1263 (N_1263,N_1147,N_1124);
xnor U1264 (N_1264,N_1135,N_1173);
or U1265 (N_1265,N_1181,N_1174);
xor U1266 (N_1266,N_1121,N_1147);
nor U1267 (N_1267,N_1155,N_1101);
or U1268 (N_1268,N_1123,N_1153);
or U1269 (N_1269,N_1166,N_1163);
nor U1270 (N_1270,N_1195,N_1177);
nor U1271 (N_1271,N_1121,N_1133);
nor U1272 (N_1272,N_1135,N_1191);
or U1273 (N_1273,N_1157,N_1181);
or U1274 (N_1274,N_1199,N_1180);
nand U1275 (N_1275,N_1101,N_1106);
xor U1276 (N_1276,N_1155,N_1162);
xnor U1277 (N_1277,N_1160,N_1149);
nand U1278 (N_1278,N_1123,N_1152);
nor U1279 (N_1279,N_1119,N_1153);
or U1280 (N_1280,N_1141,N_1100);
nor U1281 (N_1281,N_1145,N_1136);
xnor U1282 (N_1282,N_1152,N_1189);
and U1283 (N_1283,N_1120,N_1163);
xnor U1284 (N_1284,N_1185,N_1100);
xnor U1285 (N_1285,N_1138,N_1195);
nand U1286 (N_1286,N_1198,N_1180);
or U1287 (N_1287,N_1135,N_1139);
nand U1288 (N_1288,N_1146,N_1160);
nor U1289 (N_1289,N_1138,N_1130);
xor U1290 (N_1290,N_1164,N_1185);
xor U1291 (N_1291,N_1192,N_1199);
nand U1292 (N_1292,N_1102,N_1116);
or U1293 (N_1293,N_1100,N_1152);
nor U1294 (N_1294,N_1106,N_1109);
or U1295 (N_1295,N_1143,N_1133);
xor U1296 (N_1296,N_1112,N_1177);
xor U1297 (N_1297,N_1152,N_1144);
xor U1298 (N_1298,N_1143,N_1165);
and U1299 (N_1299,N_1106,N_1199);
nand U1300 (N_1300,N_1244,N_1254);
and U1301 (N_1301,N_1212,N_1231);
xor U1302 (N_1302,N_1207,N_1203);
or U1303 (N_1303,N_1288,N_1242);
or U1304 (N_1304,N_1278,N_1273);
and U1305 (N_1305,N_1299,N_1260);
nand U1306 (N_1306,N_1239,N_1255);
and U1307 (N_1307,N_1274,N_1248);
nand U1308 (N_1308,N_1293,N_1219);
and U1309 (N_1309,N_1232,N_1262);
nand U1310 (N_1310,N_1227,N_1202);
xor U1311 (N_1311,N_1281,N_1291);
and U1312 (N_1312,N_1211,N_1250);
nor U1313 (N_1313,N_1275,N_1265);
and U1314 (N_1314,N_1208,N_1253);
nand U1315 (N_1315,N_1261,N_1240);
nor U1316 (N_1316,N_1276,N_1285);
or U1317 (N_1317,N_1286,N_1216);
nand U1318 (N_1318,N_1201,N_1230);
nand U1319 (N_1319,N_1225,N_1247);
or U1320 (N_1320,N_1218,N_1249);
xnor U1321 (N_1321,N_1271,N_1295);
and U1322 (N_1322,N_1277,N_1263);
nand U1323 (N_1323,N_1214,N_1257);
or U1324 (N_1324,N_1259,N_1283);
and U1325 (N_1325,N_1205,N_1289);
xor U1326 (N_1326,N_1223,N_1251);
nor U1327 (N_1327,N_1252,N_1292);
xnor U1328 (N_1328,N_1282,N_1279);
xor U1329 (N_1329,N_1264,N_1204);
nor U1330 (N_1330,N_1243,N_1296);
nor U1331 (N_1331,N_1297,N_1210);
nand U1332 (N_1332,N_1268,N_1267);
xnor U1333 (N_1333,N_1270,N_1234);
and U1334 (N_1334,N_1258,N_1235);
and U1335 (N_1335,N_1272,N_1284);
xor U1336 (N_1336,N_1221,N_1266);
nand U1337 (N_1337,N_1245,N_1220);
and U1338 (N_1338,N_1206,N_1269);
nor U1339 (N_1339,N_1298,N_1217);
or U1340 (N_1340,N_1241,N_1236);
nor U1341 (N_1341,N_1228,N_1224);
xor U1342 (N_1342,N_1226,N_1213);
xor U1343 (N_1343,N_1294,N_1222);
nor U1344 (N_1344,N_1256,N_1209);
or U1345 (N_1345,N_1200,N_1237);
or U1346 (N_1346,N_1229,N_1233);
nor U1347 (N_1347,N_1290,N_1287);
nor U1348 (N_1348,N_1238,N_1280);
nor U1349 (N_1349,N_1215,N_1246);
nand U1350 (N_1350,N_1257,N_1284);
xnor U1351 (N_1351,N_1271,N_1231);
nand U1352 (N_1352,N_1206,N_1233);
nor U1353 (N_1353,N_1201,N_1221);
nand U1354 (N_1354,N_1262,N_1200);
xor U1355 (N_1355,N_1298,N_1215);
and U1356 (N_1356,N_1243,N_1266);
xnor U1357 (N_1357,N_1231,N_1215);
and U1358 (N_1358,N_1290,N_1234);
and U1359 (N_1359,N_1265,N_1231);
nand U1360 (N_1360,N_1269,N_1227);
xor U1361 (N_1361,N_1248,N_1246);
nor U1362 (N_1362,N_1263,N_1243);
or U1363 (N_1363,N_1276,N_1256);
or U1364 (N_1364,N_1283,N_1231);
nor U1365 (N_1365,N_1257,N_1283);
and U1366 (N_1366,N_1228,N_1203);
nor U1367 (N_1367,N_1274,N_1225);
nand U1368 (N_1368,N_1208,N_1236);
xor U1369 (N_1369,N_1225,N_1241);
and U1370 (N_1370,N_1262,N_1246);
nor U1371 (N_1371,N_1275,N_1289);
nor U1372 (N_1372,N_1235,N_1204);
nand U1373 (N_1373,N_1250,N_1281);
nand U1374 (N_1374,N_1251,N_1283);
xor U1375 (N_1375,N_1203,N_1264);
nand U1376 (N_1376,N_1297,N_1265);
and U1377 (N_1377,N_1253,N_1215);
xor U1378 (N_1378,N_1267,N_1296);
or U1379 (N_1379,N_1249,N_1251);
and U1380 (N_1380,N_1283,N_1268);
nand U1381 (N_1381,N_1210,N_1257);
xor U1382 (N_1382,N_1298,N_1274);
or U1383 (N_1383,N_1283,N_1227);
nand U1384 (N_1384,N_1286,N_1293);
xor U1385 (N_1385,N_1227,N_1200);
nand U1386 (N_1386,N_1216,N_1227);
and U1387 (N_1387,N_1202,N_1262);
nor U1388 (N_1388,N_1245,N_1292);
xnor U1389 (N_1389,N_1251,N_1271);
and U1390 (N_1390,N_1259,N_1278);
and U1391 (N_1391,N_1227,N_1250);
nor U1392 (N_1392,N_1278,N_1294);
or U1393 (N_1393,N_1294,N_1244);
or U1394 (N_1394,N_1213,N_1237);
xnor U1395 (N_1395,N_1286,N_1229);
or U1396 (N_1396,N_1292,N_1281);
or U1397 (N_1397,N_1238,N_1251);
and U1398 (N_1398,N_1224,N_1208);
or U1399 (N_1399,N_1206,N_1219);
or U1400 (N_1400,N_1317,N_1395);
nand U1401 (N_1401,N_1349,N_1301);
nor U1402 (N_1402,N_1351,N_1309);
nand U1403 (N_1403,N_1371,N_1383);
nor U1404 (N_1404,N_1394,N_1393);
xor U1405 (N_1405,N_1300,N_1318);
and U1406 (N_1406,N_1359,N_1397);
nand U1407 (N_1407,N_1319,N_1335);
xnor U1408 (N_1408,N_1315,N_1381);
nor U1409 (N_1409,N_1326,N_1337);
or U1410 (N_1410,N_1306,N_1396);
and U1411 (N_1411,N_1348,N_1332);
and U1412 (N_1412,N_1331,N_1361);
nor U1413 (N_1413,N_1388,N_1343);
nor U1414 (N_1414,N_1305,N_1314);
xnor U1415 (N_1415,N_1312,N_1342);
nand U1416 (N_1416,N_1344,N_1323);
xor U1417 (N_1417,N_1313,N_1320);
xnor U1418 (N_1418,N_1324,N_1368);
or U1419 (N_1419,N_1322,N_1329);
nor U1420 (N_1420,N_1378,N_1307);
or U1421 (N_1421,N_1303,N_1357);
nor U1422 (N_1422,N_1386,N_1310);
and U1423 (N_1423,N_1377,N_1390);
xor U1424 (N_1424,N_1362,N_1352);
xnor U1425 (N_1425,N_1355,N_1384);
xnor U1426 (N_1426,N_1380,N_1321);
or U1427 (N_1427,N_1366,N_1360);
xnor U1428 (N_1428,N_1374,N_1365);
xnor U1429 (N_1429,N_1304,N_1347);
nand U1430 (N_1430,N_1379,N_1325);
or U1431 (N_1431,N_1302,N_1385);
xor U1432 (N_1432,N_1399,N_1370);
nor U1433 (N_1433,N_1330,N_1369);
nor U1434 (N_1434,N_1389,N_1363);
or U1435 (N_1435,N_1345,N_1350);
nand U1436 (N_1436,N_1336,N_1376);
or U1437 (N_1437,N_1316,N_1356);
and U1438 (N_1438,N_1334,N_1308);
or U1439 (N_1439,N_1339,N_1353);
nor U1440 (N_1440,N_1382,N_1333);
xor U1441 (N_1441,N_1328,N_1364);
and U1442 (N_1442,N_1367,N_1392);
xnor U1443 (N_1443,N_1372,N_1338);
and U1444 (N_1444,N_1311,N_1340);
or U1445 (N_1445,N_1346,N_1354);
or U1446 (N_1446,N_1341,N_1398);
nor U1447 (N_1447,N_1358,N_1387);
or U1448 (N_1448,N_1373,N_1391);
xor U1449 (N_1449,N_1375,N_1327);
xnor U1450 (N_1450,N_1363,N_1310);
and U1451 (N_1451,N_1320,N_1311);
nand U1452 (N_1452,N_1354,N_1301);
and U1453 (N_1453,N_1386,N_1356);
or U1454 (N_1454,N_1337,N_1343);
nor U1455 (N_1455,N_1382,N_1390);
xor U1456 (N_1456,N_1312,N_1368);
nor U1457 (N_1457,N_1352,N_1320);
or U1458 (N_1458,N_1314,N_1346);
and U1459 (N_1459,N_1393,N_1370);
nand U1460 (N_1460,N_1366,N_1313);
or U1461 (N_1461,N_1331,N_1334);
or U1462 (N_1462,N_1323,N_1312);
and U1463 (N_1463,N_1312,N_1348);
and U1464 (N_1464,N_1320,N_1369);
and U1465 (N_1465,N_1300,N_1364);
or U1466 (N_1466,N_1347,N_1395);
nor U1467 (N_1467,N_1330,N_1301);
or U1468 (N_1468,N_1302,N_1368);
or U1469 (N_1469,N_1307,N_1395);
xor U1470 (N_1470,N_1392,N_1361);
nor U1471 (N_1471,N_1335,N_1313);
xor U1472 (N_1472,N_1393,N_1372);
and U1473 (N_1473,N_1366,N_1330);
or U1474 (N_1474,N_1358,N_1309);
or U1475 (N_1475,N_1327,N_1318);
nor U1476 (N_1476,N_1365,N_1379);
nand U1477 (N_1477,N_1354,N_1343);
nor U1478 (N_1478,N_1302,N_1327);
nand U1479 (N_1479,N_1384,N_1320);
or U1480 (N_1480,N_1388,N_1342);
and U1481 (N_1481,N_1368,N_1387);
nor U1482 (N_1482,N_1375,N_1312);
nor U1483 (N_1483,N_1315,N_1399);
nor U1484 (N_1484,N_1342,N_1311);
nand U1485 (N_1485,N_1368,N_1362);
or U1486 (N_1486,N_1349,N_1317);
and U1487 (N_1487,N_1323,N_1314);
or U1488 (N_1488,N_1353,N_1391);
xnor U1489 (N_1489,N_1307,N_1360);
and U1490 (N_1490,N_1369,N_1385);
nor U1491 (N_1491,N_1361,N_1301);
or U1492 (N_1492,N_1354,N_1371);
nand U1493 (N_1493,N_1348,N_1399);
nand U1494 (N_1494,N_1374,N_1350);
nor U1495 (N_1495,N_1360,N_1378);
xor U1496 (N_1496,N_1369,N_1349);
nor U1497 (N_1497,N_1374,N_1379);
and U1498 (N_1498,N_1359,N_1330);
nand U1499 (N_1499,N_1301,N_1316);
or U1500 (N_1500,N_1471,N_1420);
nor U1501 (N_1501,N_1449,N_1466);
xor U1502 (N_1502,N_1477,N_1422);
xnor U1503 (N_1503,N_1464,N_1454);
nand U1504 (N_1504,N_1491,N_1472);
xnor U1505 (N_1505,N_1485,N_1415);
and U1506 (N_1506,N_1460,N_1438);
nor U1507 (N_1507,N_1493,N_1469);
nand U1508 (N_1508,N_1497,N_1408);
nand U1509 (N_1509,N_1459,N_1429);
nand U1510 (N_1510,N_1479,N_1487);
nand U1511 (N_1511,N_1489,N_1437);
xor U1512 (N_1512,N_1423,N_1416);
and U1513 (N_1513,N_1412,N_1448);
nand U1514 (N_1514,N_1401,N_1457);
xor U1515 (N_1515,N_1427,N_1417);
nand U1516 (N_1516,N_1446,N_1425);
or U1517 (N_1517,N_1419,N_1495);
nand U1518 (N_1518,N_1400,N_1490);
nor U1519 (N_1519,N_1467,N_1444);
and U1520 (N_1520,N_1436,N_1439);
and U1521 (N_1521,N_1405,N_1410);
and U1522 (N_1522,N_1481,N_1453);
nand U1523 (N_1523,N_1480,N_1432);
xnor U1524 (N_1524,N_1431,N_1406);
or U1525 (N_1525,N_1465,N_1474);
nor U1526 (N_1526,N_1450,N_1463);
xor U1527 (N_1527,N_1407,N_1430);
nand U1528 (N_1528,N_1426,N_1435);
nand U1529 (N_1529,N_1482,N_1413);
and U1530 (N_1530,N_1462,N_1496);
xor U1531 (N_1531,N_1486,N_1452);
nor U1532 (N_1532,N_1440,N_1494);
nor U1533 (N_1533,N_1473,N_1458);
nor U1534 (N_1534,N_1483,N_1456);
nor U1535 (N_1535,N_1421,N_1475);
nand U1536 (N_1536,N_1403,N_1411);
nor U1537 (N_1537,N_1484,N_1409);
or U1538 (N_1538,N_1476,N_1434);
nor U1539 (N_1539,N_1404,N_1447);
nand U1540 (N_1540,N_1414,N_1492);
or U1541 (N_1541,N_1468,N_1455);
nor U1542 (N_1542,N_1418,N_1402);
or U1543 (N_1543,N_1424,N_1478);
nor U1544 (N_1544,N_1445,N_1498);
xnor U1545 (N_1545,N_1443,N_1433);
or U1546 (N_1546,N_1470,N_1461);
xnor U1547 (N_1547,N_1442,N_1441);
and U1548 (N_1548,N_1488,N_1428);
nand U1549 (N_1549,N_1499,N_1451);
and U1550 (N_1550,N_1427,N_1434);
nand U1551 (N_1551,N_1485,N_1489);
nand U1552 (N_1552,N_1448,N_1453);
xor U1553 (N_1553,N_1406,N_1427);
nand U1554 (N_1554,N_1433,N_1493);
xor U1555 (N_1555,N_1443,N_1498);
xnor U1556 (N_1556,N_1459,N_1406);
nor U1557 (N_1557,N_1428,N_1402);
or U1558 (N_1558,N_1452,N_1455);
xor U1559 (N_1559,N_1427,N_1418);
nor U1560 (N_1560,N_1469,N_1425);
xnor U1561 (N_1561,N_1442,N_1494);
xnor U1562 (N_1562,N_1494,N_1413);
nand U1563 (N_1563,N_1445,N_1411);
xor U1564 (N_1564,N_1462,N_1477);
and U1565 (N_1565,N_1457,N_1460);
xor U1566 (N_1566,N_1458,N_1442);
nor U1567 (N_1567,N_1446,N_1427);
and U1568 (N_1568,N_1416,N_1466);
nand U1569 (N_1569,N_1441,N_1458);
nor U1570 (N_1570,N_1417,N_1413);
xor U1571 (N_1571,N_1414,N_1410);
nor U1572 (N_1572,N_1420,N_1483);
and U1573 (N_1573,N_1418,N_1432);
xnor U1574 (N_1574,N_1417,N_1432);
xor U1575 (N_1575,N_1489,N_1440);
or U1576 (N_1576,N_1415,N_1469);
nand U1577 (N_1577,N_1488,N_1401);
nand U1578 (N_1578,N_1433,N_1402);
nand U1579 (N_1579,N_1497,N_1492);
nor U1580 (N_1580,N_1420,N_1489);
xor U1581 (N_1581,N_1422,N_1407);
and U1582 (N_1582,N_1442,N_1498);
nand U1583 (N_1583,N_1493,N_1418);
or U1584 (N_1584,N_1477,N_1409);
nor U1585 (N_1585,N_1433,N_1474);
and U1586 (N_1586,N_1426,N_1484);
xnor U1587 (N_1587,N_1426,N_1481);
and U1588 (N_1588,N_1498,N_1404);
or U1589 (N_1589,N_1405,N_1420);
nor U1590 (N_1590,N_1439,N_1412);
nor U1591 (N_1591,N_1466,N_1422);
and U1592 (N_1592,N_1450,N_1452);
nand U1593 (N_1593,N_1480,N_1476);
nor U1594 (N_1594,N_1497,N_1417);
xnor U1595 (N_1595,N_1427,N_1423);
xor U1596 (N_1596,N_1477,N_1450);
nor U1597 (N_1597,N_1416,N_1442);
nor U1598 (N_1598,N_1484,N_1487);
and U1599 (N_1599,N_1431,N_1439);
nand U1600 (N_1600,N_1552,N_1530);
or U1601 (N_1601,N_1523,N_1564);
nand U1602 (N_1602,N_1582,N_1593);
or U1603 (N_1603,N_1576,N_1540);
xor U1604 (N_1604,N_1544,N_1585);
xor U1605 (N_1605,N_1589,N_1597);
nand U1606 (N_1606,N_1577,N_1569);
xor U1607 (N_1607,N_1584,N_1524);
nand U1608 (N_1608,N_1547,N_1556);
xnor U1609 (N_1609,N_1574,N_1551);
nor U1610 (N_1610,N_1555,N_1545);
and U1611 (N_1611,N_1517,N_1565);
nor U1612 (N_1612,N_1522,N_1503);
and U1613 (N_1613,N_1508,N_1521);
nor U1614 (N_1614,N_1578,N_1587);
and U1615 (N_1615,N_1543,N_1553);
or U1616 (N_1616,N_1583,N_1533);
or U1617 (N_1617,N_1535,N_1562);
and U1618 (N_1618,N_1526,N_1572);
nand U1619 (N_1619,N_1595,N_1502);
nor U1620 (N_1620,N_1550,N_1531);
and U1621 (N_1621,N_1575,N_1558);
nor U1622 (N_1622,N_1512,N_1501);
or U1623 (N_1623,N_1528,N_1504);
or U1624 (N_1624,N_1596,N_1588);
and U1625 (N_1625,N_1559,N_1500);
or U1626 (N_1626,N_1586,N_1527);
xor U1627 (N_1627,N_1554,N_1509);
or U1628 (N_1628,N_1541,N_1506);
nor U1629 (N_1629,N_1516,N_1599);
or U1630 (N_1630,N_1520,N_1567);
nor U1631 (N_1631,N_1537,N_1581);
xnor U1632 (N_1632,N_1557,N_1592);
and U1633 (N_1633,N_1525,N_1519);
xor U1634 (N_1634,N_1542,N_1536);
nand U1635 (N_1635,N_1511,N_1573);
or U1636 (N_1636,N_1566,N_1539);
and U1637 (N_1637,N_1532,N_1548);
nor U1638 (N_1638,N_1518,N_1549);
nand U1639 (N_1639,N_1594,N_1515);
nor U1640 (N_1640,N_1598,N_1560);
nor U1641 (N_1641,N_1538,N_1510);
xnor U1642 (N_1642,N_1563,N_1579);
nand U1643 (N_1643,N_1580,N_1570);
nor U1644 (N_1644,N_1571,N_1561);
or U1645 (N_1645,N_1529,N_1534);
or U1646 (N_1646,N_1590,N_1514);
nor U1647 (N_1647,N_1546,N_1568);
nor U1648 (N_1648,N_1507,N_1513);
nand U1649 (N_1649,N_1505,N_1591);
and U1650 (N_1650,N_1544,N_1512);
or U1651 (N_1651,N_1547,N_1523);
nand U1652 (N_1652,N_1561,N_1554);
and U1653 (N_1653,N_1553,N_1589);
nor U1654 (N_1654,N_1520,N_1508);
nand U1655 (N_1655,N_1543,N_1517);
or U1656 (N_1656,N_1558,N_1561);
or U1657 (N_1657,N_1512,N_1511);
or U1658 (N_1658,N_1513,N_1525);
xor U1659 (N_1659,N_1521,N_1530);
nor U1660 (N_1660,N_1585,N_1573);
nand U1661 (N_1661,N_1509,N_1572);
nand U1662 (N_1662,N_1517,N_1501);
or U1663 (N_1663,N_1525,N_1591);
nand U1664 (N_1664,N_1531,N_1567);
nand U1665 (N_1665,N_1594,N_1567);
xor U1666 (N_1666,N_1535,N_1571);
nor U1667 (N_1667,N_1576,N_1584);
xnor U1668 (N_1668,N_1521,N_1582);
nand U1669 (N_1669,N_1519,N_1512);
nor U1670 (N_1670,N_1576,N_1529);
xnor U1671 (N_1671,N_1595,N_1503);
xnor U1672 (N_1672,N_1563,N_1512);
xor U1673 (N_1673,N_1533,N_1546);
nand U1674 (N_1674,N_1582,N_1530);
xor U1675 (N_1675,N_1539,N_1580);
nor U1676 (N_1676,N_1558,N_1519);
nor U1677 (N_1677,N_1548,N_1599);
and U1678 (N_1678,N_1506,N_1578);
nor U1679 (N_1679,N_1546,N_1520);
or U1680 (N_1680,N_1590,N_1506);
and U1681 (N_1681,N_1564,N_1583);
nor U1682 (N_1682,N_1540,N_1575);
xor U1683 (N_1683,N_1532,N_1580);
nand U1684 (N_1684,N_1545,N_1588);
and U1685 (N_1685,N_1560,N_1529);
xor U1686 (N_1686,N_1529,N_1502);
nor U1687 (N_1687,N_1551,N_1564);
xor U1688 (N_1688,N_1589,N_1581);
xnor U1689 (N_1689,N_1594,N_1536);
nand U1690 (N_1690,N_1553,N_1561);
or U1691 (N_1691,N_1508,N_1516);
xor U1692 (N_1692,N_1598,N_1520);
nor U1693 (N_1693,N_1584,N_1571);
xor U1694 (N_1694,N_1598,N_1537);
and U1695 (N_1695,N_1549,N_1531);
nor U1696 (N_1696,N_1580,N_1508);
xor U1697 (N_1697,N_1509,N_1505);
and U1698 (N_1698,N_1544,N_1554);
xor U1699 (N_1699,N_1579,N_1540);
nor U1700 (N_1700,N_1673,N_1658);
xnor U1701 (N_1701,N_1644,N_1623);
or U1702 (N_1702,N_1633,N_1693);
nor U1703 (N_1703,N_1687,N_1683);
nor U1704 (N_1704,N_1694,N_1605);
or U1705 (N_1705,N_1625,N_1608);
xor U1706 (N_1706,N_1612,N_1651);
nor U1707 (N_1707,N_1606,N_1661);
or U1708 (N_1708,N_1632,N_1672);
or U1709 (N_1709,N_1689,N_1637);
and U1710 (N_1710,N_1682,N_1648);
or U1711 (N_1711,N_1669,N_1696);
nand U1712 (N_1712,N_1653,N_1602);
nor U1713 (N_1713,N_1667,N_1601);
xor U1714 (N_1714,N_1628,N_1626);
and U1715 (N_1715,N_1665,N_1692);
xor U1716 (N_1716,N_1611,N_1620);
and U1717 (N_1717,N_1685,N_1629);
and U1718 (N_1718,N_1691,N_1610);
or U1719 (N_1719,N_1674,N_1695);
nor U1720 (N_1720,N_1668,N_1614);
nand U1721 (N_1721,N_1646,N_1636);
xnor U1722 (N_1722,N_1662,N_1624);
and U1723 (N_1723,N_1638,N_1698);
or U1724 (N_1724,N_1655,N_1634);
xor U1725 (N_1725,N_1681,N_1675);
xor U1726 (N_1726,N_1643,N_1642);
nor U1727 (N_1727,N_1603,N_1676);
xnor U1728 (N_1728,N_1615,N_1607);
or U1729 (N_1729,N_1641,N_1619);
or U1730 (N_1730,N_1635,N_1617);
nand U1731 (N_1731,N_1616,N_1664);
xnor U1732 (N_1732,N_1627,N_1659);
and U1733 (N_1733,N_1671,N_1686);
or U1734 (N_1734,N_1657,N_1690);
and U1735 (N_1735,N_1656,N_1600);
nor U1736 (N_1736,N_1679,N_1652);
nand U1737 (N_1737,N_1618,N_1666);
xor U1738 (N_1738,N_1640,N_1630);
xnor U1739 (N_1739,N_1649,N_1678);
nand U1740 (N_1740,N_1677,N_1670);
xnor U1741 (N_1741,N_1645,N_1684);
nand U1742 (N_1742,N_1697,N_1639);
nand U1743 (N_1743,N_1647,N_1622);
nand U1744 (N_1744,N_1663,N_1650);
nand U1745 (N_1745,N_1680,N_1613);
nor U1746 (N_1746,N_1631,N_1699);
xor U1747 (N_1747,N_1688,N_1654);
and U1748 (N_1748,N_1604,N_1660);
or U1749 (N_1749,N_1621,N_1609);
or U1750 (N_1750,N_1648,N_1605);
or U1751 (N_1751,N_1623,N_1608);
nand U1752 (N_1752,N_1619,N_1600);
xnor U1753 (N_1753,N_1626,N_1653);
nor U1754 (N_1754,N_1641,N_1620);
or U1755 (N_1755,N_1696,N_1601);
or U1756 (N_1756,N_1627,N_1692);
and U1757 (N_1757,N_1661,N_1612);
and U1758 (N_1758,N_1622,N_1678);
nor U1759 (N_1759,N_1672,N_1656);
xor U1760 (N_1760,N_1680,N_1699);
xor U1761 (N_1761,N_1694,N_1676);
and U1762 (N_1762,N_1639,N_1631);
and U1763 (N_1763,N_1668,N_1656);
nor U1764 (N_1764,N_1693,N_1665);
or U1765 (N_1765,N_1667,N_1619);
nand U1766 (N_1766,N_1639,N_1686);
nor U1767 (N_1767,N_1611,N_1647);
and U1768 (N_1768,N_1643,N_1621);
and U1769 (N_1769,N_1659,N_1652);
nand U1770 (N_1770,N_1662,N_1626);
and U1771 (N_1771,N_1686,N_1681);
and U1772 (N_1772,N_1685,N_1657);
or U1773 (N_1773,N_1666,N_1611);
or U1774 (N_1774,N_1625,N_1631);
and U1775 (N_1775,N_1655,N_1670);
nand U1776 (N_1776,N_1671,N_1625);
or U1777 (N_1777,N_1642,N_1651);
nor U1778 (N_1778,N_1609,N_1651);
xnor U1779 (N_1779,N_1694,N_1647);
or U1780 (N_1780,N_1699,N_1687);
nor U1781 (N_1781,N_1692,N_1689);
nor U1782 (N_1782,N_1661,N_1699);
nor U1783 (N_1783,N_1637,N_1636);
nand U1784 (N_1784,N_1698,N_1648);
xor U1785 (N_1785,N_1685,N_1681);
nand U1786 (N_1786,N_1677,N_1621);
nand U1787 (N_1787,N_1665,N_1609);
nor U1788 (N_1788,N_1613,N_1628);
nand U1789 (N_1789,N_1657,N_1689);
or U1790 (N_1790,N_1696,N_1621);
nor U1791 (N_1791,N_1659,N_1688);
nor U1792 (N_1792,N_1691,N_1679);
or U1793 (N_1793,N_1633,N_1613);
or U1794 (N_1794,N_1623,N_1654);
and U1795 (N_1795,N_1651,N_1671);
or U1796 (N_1796,N_1661,N_1695);
or U1797 (N_1797,N_1619,N_1605);
nand U1798 (N_1798,N_1621,N_1637);
and U1799 (N_1799,N_1650,N_1659);
and U1800 (N_1800,N_1765,N_1777);
nand U1801 (N_1801,N_1762,N_1701);
nand U1802 (N_1802,N_1791,N_1704);
xnor U1803 (N_1803,N_1730,N_1718);
and U1804 (N_1804,N_1731,N_1737);
nand U1805 (N_1805,N_1763,N_1776);
xor U1806 (N_1806,N_1768,N_1735);
or U1807 (N_1807,N_1790,N_1781);
nand U1808 (N_1808,N_1753,N_1795);
nor U1809 (N_1809,N_1706,N_1734);
or U1810 (N_1810,N_1727,N_1717);
and U1811 (N_1811,N_1711,N_1750);
xnor U1812 (N_1812,N_1720,N_1788);
xor U1813 (N_1813,N_1738,N_1769);
or U1814 (N_1814,N_1756,N_1798);
and U1815 (N_1815,N_1779,N_1721);
and U1816 (N_1816,N_1749,N_1758);
xnor U1817 (N_1817,N_1725,N_1771);
nand U1818 (N_1818,N_1782,N_1732);
and U1819 (N_1819,N_1783,N_1702);
nand U1820 (N_1820,N_1722,N_1740);
or U1821 (N_1821,N_1736,N_1719);
nor U1822 (N_1822,N_1743,N_1709);
nand U1823 (N_1823,N_1767,N_1770);
nor U1824 (N_1824,N_1705,N_1744);
nor U1825 (N_1825,N_1733,N_1774);
xnor U1826 (N_1826,N_1755,N_1761);
nand U1827 (N_1827,N_1726,N_1741);
nor U1828 (N_1828,N_1728,N_1729);
or U1829 (N_1829,N_1759,N_1789);
xor U1830 (N_1830,N_1739,N_1714);
xnor U1831 (N_1831,N_1793,N_1724);
nand U1832 (N_1832,N_1766,N_1778);
nand U1833 (N_1833,N_1723,N_1713);
xor U1834 (N_1834,N_1715,N_1797);
and U1835 (N_1835,N_1785,N_1712);
and U1836 (N_1836,N_1752,N_1775);
xor U1837 (N_1837,N_1747,N_1700);
and U1838 (N_1838,N_1764,N_1742);
and U1839 (N_1839,N_1772,N_1787);
or U1840 (N_1840,N_1794,N_1708);
xnor U1841 (N_1841,N_1754,N_1707);
nor U1842 (N_1842,N_1703,N_1773);
nand U1843 (N_1843,N_1760,N_1786);
and U1844 (N_1844,N_1799,N_1757);
nand U1845 (N_1845,N_1745,N_1784);
nand U1846 (N_1846,N_1748,N_1746);
xnor U1847 (N_1847,N_1780,N_1710);
or U1848 (N_1848,N_1792,N_1796);
xor U1849 (N_1849,N_1751,N_1716);
or U1850 (N_1850,N_1716,N_1795);
and U1851 (N_1851,N_1725,N_1744);
or U1852 (N_1852,N_1709,N_1739);
nand U1853 (N_1853,N_1745,N_1765);
nand U1854 (N_1854,N_1722,N_1777);
xnor U1855 (N_1855,N_1731,N_1795);
nor U1856 (N_1856,N_1726,N_1751);
and U1857 (N_1857,N_1731,N_1766);
nor U1858 (N_1858,N_1789,N_1780);
and U1859 (N_1859,N_1789,N_1705);
and U1860 (N_1860,N_1725,N_1782);
nand U1861 (N_1861,N_1776,N_1787);
xor U1862 (N_1862,N_1723,N_1778);
xnor U1863 (N_1863,N_1778,N_1724);
and U1864 (N_1864,N_1799,N_1750);
or U1865 (N_1865,N_1706,N_1761);
or U1866 (N_1866,N_1728,N_1741);
and U1867 (N_1867,N_1793,N_1713);
nor U1868 (N_1868,N_1764,N_1728);
xnor U1869 (N_1869,N_1767,N_1797);
nand U1870 (N_1870,N_1791,N_1798);
nand U1871 (N_1871,N_1766,N_1746);
nand U1872 (N_1872,N_1798,N_1729);
xnor U1873 (N_1873,N_1704,N_1799);
nor U1874 (N_1874,N_1756,N_1791);
xor U1875 (N_1875,N_1758,N_1798);
nand U1876 (N_1876,N_1739,N_1778);
nor U1877 (N_1877,N_1735,N_1791);
or U1878 (N_1878,N_1714,N_1747);
and U1879 (N_1879,N_1777,N_1755);
or U1880 (N_1880,N_1720,N_1713);
or U1881 (N_1881,N_1733,N_1793);
or U1882 (N_1882,N_1736,N_1746);
nor U1883 (N_1883,N_1779,N_1791);
or U1884 (N_1884,N_1770,N_1781);
nor U1885 (N_1885,N_1768,N_1731);
or U1886 (N_1886,N_1745,N_1727);
nand U1887 (N_1887,N_1763,N_1755);
nand U1888 (N_1888,N_1713,N_1750);
xor U1889 (N_1889,N_1722,N_1799);
nand U1890 (N_1890,N_1773,N_1799);
xnor U1891 (N_1891,N_1731,N_1735);
or U1892 (N_1892,N_1775,N_1776);
xnor U1893 (N_1893,N_1793,N_1778);
and U1894 (N_1894,N_1730,N_1754);
xnor U1895 (N_1895,N_1732,N_1717);
or U1896 (N_1896,N_1762,N_1706);
nor U1897 (N_1897,N_1706,N_1763);
or U1898 (N_1898,N_1799,N_1751);
or U1899 (N_1899,N_1726,N_1758);
nor U1900 (N_1900,N_1896,N_1867);
nor U1901 (N_1901,N_1888,N_1873);
or U1902 (N_1902,N_1875,N_1828);
xnor U1903 (N_1903,N_1874,N_1881);
nand U1904 (N_1904,N_1857,N_1883);
or U1905 (N_1905,N_1818,N_1865);
nor U1906 (N_1906,N_1822,N_1880);
or U1907 (N_1907,N_1861,N_1829);
nor U1908 (N_1908,N_1887,N_1878);
or U1909 (N_1909,N_1834,N_1837);
nand U1910 (N_1910,N_1877,N_1846);
or U1911 (N_1911,N_1882,N_1805);
nor U1912 (N_1912,N_1842,N_1830);
nand U1913 (N_1913,N_1847,N_1819);
nor U1914 (N_1914,N_1870,N_1827);
xor U1915 (N_1915,N_1849,N_1871);
nand U1916 (N_1916,N_1848,N_1862);
or U1917 (N_1917,N_1840,N_1854);
nor U1918 (N_1918,N_1872,N_1839);
nand U1919 (N_1919,N_1864,N_1809);
xor U1920 (N_1920,N_1802,N_1841);
nand U1921 (N_1921,N_1823,N_1815);
and U1922 (N_1922,N_1812,N_1838);
nand U1923 (N_1923,N_1866,N_1821);
and U1924 (N_1924,N_1850,N_1894);
nor U1925 (N_1925,N_1852,N_1863);
nor U1926 (N_1926,N_1843,N_1803);
nor U1927 (N_1927,N_1895,N_1826);
nor U1928 (N_1928,N_1885,N_1801);
and U1929 (N_1929,N_1889,N_1820);
xnor U1930 (N_1930,N_1898,N_1876);
and U1931 (N_1931,N_1879,N_1853);
and U1932 (N_1932,N_1897,N_1891);
or U1933 (N_1933,N_1808,N_1859);
nor U1934 (N_1934,N_1884,N_1858);
nor U1935 (N_1935,N_1899,N_1817);
xnor U1936 (N_1936,N_1835,N_1831);
or U1937 (N_1937,N_1845,N_1890);
xor U1938 (N_1938,N_1836,N_1832);
or U1939 (N_1939,N_1806,N_1855);
nor U1940 (N_1940,N_1868,N_1869);
nor U1941 (N_1941,N_1810,N_1814);
or U1942 (N_1942,N_1800,N_1811);
and U1943 (N_1943,N_1844,N_1833);
nor U1944 (N_1944,N_1893,N_1804);
or U1945 (N_1945,N_1824,N_1856);
xor U1946 (N_1946,N_1825,N_1892);
and U1947 (N_1947,N_1807,N_1886);
and U1948 (N_1948,N_1816,N_1813);
nand U1949 (N_1949,N_1851,N_1860);
nor U1950 (N_1950,N_1893,N_1860);
or U1951 (N_1951,N_1852,N_1886);
nor U1952 (N_1952,N_1874,N_1891);
xnor U1953 (N_1953,N_1819,N_1845);
or U1954 (N_1954,N_1858,N_1890);
nand U1955 (N_1955,N_1809,N_1881);
and U1956 (N_1956,N_1869,N_1873);
nand U1957 (N_1957,N_1883,N_1807);
or U1958 (N_1958,N_1879,N_1869);
nand U1959 (N_1959,N_1802,N_1871);
and U1960 (N_1960,N_1808,N_1873);
or U1961 (N_1961,N_1885,N_1858);
nand U1962 (N_1962,N_1870,N_1879);
or U1963 (N_1963,N_1898,N_1828);
xnor U1964 (N_1964,N_1885,N_1884);
or U1965 (N_1965,N_1825,N_1885);
or U1966 (N_1966,N_1840,N_1849);
nor U1967 (N_1967,N_1840,N_1824);
nor U1968 (N_1968,N_1859,N_1836);
nor U1969 (N_1969,N_1851,N_1826);
nor U1970 (N_1970,N_1846,N_1807);
nor U1971 (N_1971,N_1803,N_1808);
xor U1972 (N_1972,N_1865,N_1880);
or U1973 (N_1973,N_1889,N_1886);
nor U1974 (N_1974,N_1826,N_1805);
or U1975 (N_1975,N_1881,N_1806);
nor U1976 (N_1976,N_1894,N_1819);
and U1977 (N_1977,N_1839,N_1848);
or U1978 (N_1978,N_1876,N_1812);
and U1979 (N_1979,N_1865,N_1892);
xnor U1980 (N_1980,N_1855,N_1842);
or U1981 (N_1981,N_1847,N_1872);
or U1982 (N_1982,N_1801,N_1870);
or U1983 (N_1983,N_1809,N_1866);
or U1984 (N_1984,N_1861,N_1812);
and U1985 (N_1985,N_1841,N_1819);
and U1986 (N_1986,N_1894,N_1831);
xnor U1987 (N_1987,N_1814,N_1884);
or U1988 (N_1988,N_1808,N_1810);
nand U1989 (N_1989,N_1883,N_1845);
nor U1990 (N_1990,N_1821,N_1858);
nand U1991 (N_1991,N_1844,N_1850);
nand U1992 (N_1992,N_1897,N_1893);
or U1993 (N_1993,N_1890,N_1877);
xor U1994 (N_1994,N_1805,N_1895);
nand U1995 (N_1995,N_1801,N_1835);
nand U1996 (N_1996,N_1829,N_1811);
nor U1997 (N_1997,N_1801,N_1828);
nor U1998 (N_1998,N_1879,N_1820);
xnor U1999 (N_1999,N_1828,N_1859);
xor U2000 (N_2000,N_1996,N_1933);
nor U2001 (N_2001,N_1975,N_1925);
nor U2002 (N_2002,N_1923,N_1972);
nand U2003 (N_2003,N_1980,N_1977);
xor U2004 (N_2004,N_1930,N_1954);
nand U2005 (N_2005,N_1911,N_1901);
and U2006 (N_2006,N_1963,N_1953);
or U2007 (N_2007,N_1982,N_1920);
xor U2008 (N_2008,N_1931,N_1917);
xnor U2009 (N_2009,N_1956,N_1987);
nor U2010 (N_2010,N_1902,N_1976);
xnor U2011 (N_2011,N_1909,N_1943);
nor U2012 (N_2012,N_1929,N_1948);
and U2013 (N_2013,N_1922,N_1952);
nor U2014 (N_2014,N_1918,N_1973);
nor U2015 (N_2015,N_1986,N_1958);
nor U2016 (N_2016,N_1966,N_1955);
nand U2017 (N_2017,N_1993,N_1944);
or U2018 (N_2018,N_1984,N_1971);
nand U2019 (N_2019,N_1978,N_1936);
and U2020 (N_2020,N_1928,N_1935);
and U2021 (N_2021,N_1919,N_1916);
nand U2022 (N_2022,N_1969,N_1912);
or U2023 (N_2023,N_1999,N_1974);
xnor U2024 (N_2024,N_1979,N_1932);
and U2025 (N_2025,N_1908,N_1939);
or U2026 (N_2026,N_1940,N_1970);
nand U2027 (N_2027,N_1937,N_1959);
and U2028 (N_2028,N_1949,N_1983);
nand U2029 (N_2029,N_1957,N_1941);
nor U2030 (N_2030,N_1900,N_1921);
nand U2031 (N_2031,N_1924,N_1915);
nand U2032 (N_2032,N_1934,N_1903);
nand U2033 (N_2033,N_1995,N_1905);
nor U2034 (N_2034,N_1907,N_1960);
or U2035 (N_2035,N_1994,N_1904);
nor U2036 (N_2036,N_1989,N_1990);
xor U2037 (N_2037,N_1967,N_1914);
or U2038 (N_2038,N_1992,N_1950);
nand U2039 (N_2039,N_1927,N_1910);
nor U2040 (N_2040,N_1962,N_1985);
nand U2041 (N_2041,N_1965,N_1938);
and U2042 (N_2042,N_1951,N_1998);
xor U2043 (N_2043,N_1947,N_1961);
nand U2044 (N_2044,N_1926,N_1968);
xnor U2045 (N_2045,N_1946,N_1981);
or U2046 (N_2046,N_1988,N_1942);
and U2047 (N_2047,N_1945,N_1997);
xor U2048 (N_2048,N_1964,N_1991);
xnor U2049 (N_2049,N_1906,N_1913);
nor U2050 (N_2050,N_1989,N_1934);
nor U2051 (N_2051,N_1979,N_1934);
and U2052 (N_2052,N_1998,N_1947);
or U2053 (N_2053,N_1907,N_1913);
nand U2054 (N_2054,N_1917,N_1910);
nor U2055 (N_2055,N_1941,N_1946);
or U2056 (N_2056,N_1922,N_1918);
xnor U2057 (N_2057,N_1956,N_1992);
and U2058 (N_2058,N_1929,N_1917);
xnor U2059 (N_2059,N_1933,N_1903);
and U2060 (N_2060,N_1934,N_1993);
and U2061 (N_2061,N_1972,N_1999);
and U2062 (N_2062,N_1980,N_1927);
nand U2063 (N_2063,N_1942,N_1933);
xnor U2064 (N_2064,N_1939,N_1917);
xor U2065 (N_2065,N_1931,N_1969);
xnor U2066 (N_2066,N_1942,N_1966);
nor U2067 (N_2067,N_1933,N_1987);
nor U2068 (N_2068,N_1930,N_1972);
and U2069 (N_2069,N_1967,N_1911);
and U2070 (N_2070,N_1997,N_1907);
nand U2071 (N_2071,N_1932,N_1965);
nand U2072 (N_2072,N_1961,N_1995);
or U2073 (N_2073,N_1966,N_1960);
nand U2074 (N_2074,N_1925,N_1952);
nor U2075 (N_2075,N_1952,N_1911);
nand U2076 (N_2076,N_1900,N_1969);
nor U2077 (N_2077,N_1977,N_1918);
nand U2078 (N_2078,N_1934,N_1988);
nor U2079 (N_2079,N_1983,N_1925);
xnor U2080 (N_2080,N_1988,N_1952);
xor U2081 (N_2081,N_1978,N_1998);
or U2082 (N_2082,N_1959,N_1970);
and U2083 (N_2083,N_1963,N_1984);
nand U2084 (N_2084,N_1904,N_1989);
or U2085 (N_2085,N_1990,N_1943);
and U2086 (N_2086,N_1935,N_1946);
nand U2087 (N_2087,N_1971,N_1993);
and U2088 (N_2088,N_1994,N_1937);
and U2089 (N_2089,N_1979,N_1904);
xor U2090 (N_2090,N_1908,N_1998);
nor U2091 (N_2091,N_1909,N_1900);
or U2092 (N_2092,N_1996,N_1940);
nor U2093 (N_2093,N_1943,N_1910);
and U2094 (N_2094,N_1910,N_1922);
xnor U2095 (N_2095,N_1961,N_1942);
xnor U2096 (N_2096,N_1992,N_1919);
xor U2097 (N_2097,N_1995,N_1955);
and U2098 (N_2098,N_1914,N_1940);
and U2099 (N_2099,N_1980,N_1938);
or U2100 (N_2100,N_2025,N_2094);
nand U2101 (N_2101,N_2042,N_2016);
or U2102 (N_2102,N_2075,N_2019);
nor U2103 (N_2103,N_2039,N_2077);
or U2104 (N_2104,N_2031,N_2046);
xnor U2105 (N_2105,N_2068,N_2084);
or U2106 (N_2106,N_2056,N_2035);
xor U2107 (N_2107,N_2028,N_2010);
or U2108 (N_2108,N_2003,N_2061);
xnor U2109 (N_2109,N_2098,N_2005);
and U2110 (N_2110,N_2032,N_2026);
nand U2111 (N_2111,N_2022,N_2096);
and U2112 (N_2112,N_2011,N_2050);
and U2113 (N_2113,N_2023,N_2013);
and U2114 (N_2114,N_2087,N_2059);
and U2115 (N_2115,N_2034,N_2091);
or U2116 (N_2116,N_2044,N_2021);
or U2117 (N_2117,N_2012,N_2043);
nand U2118 (N_2118,N_2008,N_2063);
nand U2119 (N_2119,N_2048,N_2051);
xnor U2120 (N_2120,N_2020,N_2000);
nor U2121 (N_2121,N_2041,N_2076);
nor U2122 (N_2122,N_2073,N_2055);
nand U2123 (N_2123,N_2058,N_2083);
or U2124 (N_2124,N_2018,N_2017);
xnor U2125 (N_2125,N_2082,N_2064);
xnor U2126 (N_2126,N_2053,N_2081);
nor U2127 (N_2127,N_2089,N_2072);
and U2128 (N_2128,N_2071,N_2024);
xnor U2129 (N_2129,N_2065,N_2070);
or U2130 (N_2130,N_2054,N_2027);
nand U2131 (N_2131,N_2066,N_2038);
nor U2132 (N_2132,N_2045,N_2015);
xor U2133 (N_2133,N_2036,N_2060);
and U2134 (N_2134,N_2079,N_2002);
nor U2135 (N_2135,N_2086,N_2097);
xor U2136 (N_2136,N_2092,N_2052);
and U2137 (N_2137,N_2069,N_2007);
nor U2138 (N_2138,N_2099,N_2014);
nand U2139 (N_2139,N_2009,N_2047);
or U2140 (N_2140,N_2078,N_2033);
nor U2141 (N_2141,N_2030,N_2095);
or U2142 (N_2142,N_2057,N_2001);
xnor U2143 (N_2143,N_2088,N_2029);
and U2144 (N_2144,N_2090,N_2006);
xor U2145 (N_2145,N_2067,N_2004);
nor U2146 (N_2146,N_2080,N_2037);
and U2147 (N_2147,N_2085,N_2062);
nor U2148 (N_2148,N_2049,N_2040);
or U2149 (N_2149,N_2093,N_2074);
or U2150 (N_2150,N_2088,N_2082);
or U2151 (N_2151,N_2003,N_2077);
nand U2152 (N_2152,N_2093,N_2028);
nand U2153 (N_2153,N_2058,N_2054);
nand U2154 (N_2154,N_2093,N_2051);
nor U2155 (N_2155,N_2043,N_2098);
or U2156 (N_2156,N_2053,N_2056);
or U2157 (N_2157,N_2087,N_2074);
xnor U2158 (N_2158,N_2086,N_2036);
nand U2159 (N_2159,N_2025,N_2092);
nand U2160 (N_2160,N_2072,N_2081);
and U2161 (N_2161,N_2024,N_2026);
or U2162 (N_2162,N_2067,N_2077);
nor U2163 (N_2163,N_2076,N_2089);
xor U2164 (N_2164,N_2097,N_2077);
nand U2165 (N_2165,N_2082,N_2018);
nor U2166 (N_2166,N_2057,N_2059);
and U2167 (N_2167,N_2082,N_2008);
and U2168 (N_2168,N_2072,N_2065);
or U2169 (N_2169,N_2080,N_2017);
and U2170 (N_2170,N_2048,N_2003);
nand U2171 (N_2171,N_2066,N_2096);
nor U2172 (N_2172,N_2052,N_2002);
xor U2173 (N_2173,N_2048,N_2085);
or U2174 (N_2174,N_2030,N_2023);
or U2175 (N_2175,N_2098,N_2042);
nand U2176 (N_2176,N_2006,N_2017);
xnor U2177 (N_2177,N_2031,N_2038);
nand U2178 (N_2178,N_2096,N_2056);
and U2179 (N_2179,N_2014,N_2084);
nand U2180 (N_2180,N_2009,N_2074);
and U2181 (N_2181,N_2046,N_2089);
nand U2182 (N_2182,N_2065,N_2016);
or U2183 (N_2183,N_2012,N_2064);
and U2184 (N_2184,N_2011,N_2018);
nor U2185 (N_2185,N_2098,N_2044);
nor U2186 (N_2186,N_2038,N_2051);
nor U2187 (N_2187,N_2006,N_2040);
nor U2188 (N_2188,N_2020,N_2034);
or U2189 (N_2189,N_2017,N_2041);
and U2190 (N_2190,N_2004,N_2062);
nor U2191 (N_2191,N_2035,N_2037);
and U2192 (N_2192,N_2035,N_2081);
nand U2193 (N_2193,N_2001,N_2095);
and U2194 (N_2194,N_2084,N_2000);
nand U2195 (N_2195,N_2063,N_2058);
nand U2196 (N_2196,N_2049,N_2077);
and U2197 (N_2197,N_2046,N_2024);
or U2198 (N_2198,N_2006,N_2080);
nand U2199 (N_2199,N_2062,N_2082);
xnor U2200 (N_2200,N_2127,N_2136);
nor U2201 (N_2201,N_2125,N_2179);
xor U2202 (N_2202,N_2191,N_2123);
nand U2203 (N_2203,N_2151,N_2103);
or U2204 (N_2204,N_2180,N_2117);
nor U2205 (N_2205,N_2157,N_2143);
nand U2206 (N_2206,N_2167,N_2153);
nor U2207 (N_2207,N_2197,N_2134);
xor U2208 (N_2208,N_2158,N_2121);
nor U2209 (N_2209,N_2198,N_2181);
xor U2210 (N_2210,N_2138,N_2106);
xor U2211 (N_2211,N_2186,N_2164);
xnor U2212 (N_2212,N_2182,N_2128);
or U2213 (N_2213,N_2101,N_2170);
xor U2214 (N_2214,N_2183,N_2160);
nand U2215 (N_2215,N_2144,N_2131);
xor U2216 (N_2216,N_2173,N_2176);
and U2217 (N_2217,N_2130,N_2199);
nand U2218 (N_2218,N_2169,N_2110);
xnor U2219 (N_2219,N_2135,N_2140);
or U2220 (N_2220,N_2190,N_2116);
xor U2221 (N_2221,N_2146,N_2113);
or U2222 (N_2222,N_2120,N_2174);
and U2223 (N_2223,N_2165,N_2119);
nand U2224 (N_2224,N_2133,N_2109);
or U2225 (N_2225,N_2188,N_2102);
or U2226 (N_2226,N_2155,N_2184);
or U2227 (N_2227,N_2172,N_2129);
and U2228 (N_2228,N_2168,N_2150);
and U2229 (N_2229,N_2145,N_2141);
xnor U2230 (N_2230,N_2139,N_2104);
and U2231 (N_2231,N_2162,N_2166);
xnor U2232 (N_2232,N_2159,N_2189);
xor U2233 (N_2233,N_2161,N_2122);
nand U2234 (N_2234,N_2111,N_2156);
or U2235 (N_2235,N_2107,N_2149);
nor U2236 (N_2236,N_2195,N_2147);
nor U2237 (N_2237,N_2126,N_2187);
nand U2238 (N_2238,N_2142,N_2114);
or U2239 (N_2239,N_2178,N_2124);
and U2240 (N_2240,N_2154,N_2192);
or U2241 (N_2241,N_2108,N_2196);
xor U2242 (N_2242,N_2194,N_2112);
or U2243 (N_2243,N_2137,N_2171);
or U2244 (N_2244,N_2177,N_2152);
and U2245 (N_2245,N_2175,N_2132);
xnor U2246 (N_2246,N_2148,N_2115);
and U2247 (N_2247,N_2185,N_2163);
and U2248 (N_2248,N_2193,N_2118);
nor U2249 (N_2249,N_2100,N_2105);
nor U2250 (N_2250,N_2194,N_2102);
nor U2251 (N_2251,N_2149,N_2162);
nand U2252 (N_2252,N_2190,N_2112);
and U2253 (N_2253,N_2198,N_2189);
and U2254 (N_2254,N_2198,N_2186);
xor U2255 (N_2255,N_2158,N_2199);
nand U2256 (N_2256,N_2198,N_2162);
and U2257 (N_2257,N_2181,N_2115);
or U2258 (N_2258,N_2179,N_2163);
nand U2259 (N_2259,N_2158,N_2191);
nor U2260 (N_2260,N_2185,N_2180);
or U2261 (N_2261,N_2162,N_2161);
xnor U2262 (N_2262,N_2123,N_2147);
nand U2263 (N_2263,N_2138,N_2108);
xnor U2264 (N_2264,N_2116,N_2145);
xnor U2265 (N_2265,N_2189,N_2126);
nor U2266 (N_2266,N_2179,N_2169);
nor U2267 (N_2267,N_2145,N_2126);
nand U2268 (N_2268,N_2199,N_2136);
xnor U2269 (N_2269,N_2188,N_2195);
and U2270 (N_2270,N_2135,N_2178);
and U2271 (N_2271,N_2113,N_2180);
and U2272 (N_2272,N_2107,N_2165);
or U2273 (N_2273,N_2114,N_2178);
and U2274 (N_2274,N_2150,N_2154);
nor U2275 (N_2275,N_2154,N_2136);
nand U2276 (N_2276,N_2110,N_2142);
nor U2277 (N_2277,N_2113,N_2108);
nor U2278 (N_2278,N_2145,N_2112);
and U2279 (N_2279,N_2117,N_2108);
nand U2280 (N_2280,N_2109,N_2132);
nand U2281 (N_2281,N_2127,N_2163);
xnor U2282 (N_2282,N_2118,N_2101);
or U2283 (N_2283,N_2103,N_2155);
nand U2284 (N_2284,N_2191,N_2173);
and U2285 (N_2285,N_2126,N_2128);
or U2286 (N_2286,N_2139,N_2127);
xor U2287 (N_2287,N_2143,N_2151);
or U2288 (N_2288,N_2103,N_2193);
or U2289 (N_2289,N_2112,N_2106);
and U2290 (N_2290,N_2126,N_2112);
nor U2291 (N_2291,N_2187,N_2120);
and U2292 (N_2292,N_2116,N_2127);
xnor U2293 (N_2293,N_2127,N_2134);
or U2294 (N_2294,N_2165,N_2152);
nor U2295 (N_2295,N_2114,N_2148);
xor U2296 (N_2296,N_2180,N_2148);
and U2297 (N_2297,N_2161,N_2151);
nor U2298 (N_2298,N_2158,N_2103);
and U2299 (N_2299,N_2134,N_2155);
or U2300 (N_2300,N_2250,N_2264);
nand U2301 (N_2301,N_2292,N_2259);
and U2302 (N_2302,N_2215,N_2296);
nor U2303 (N_2303,N_2251,N_2217);
or U2304 (N_2304,N_2254,N_2267);
xor U2305 (N_2305,N_2223,N_2270);
xnor U2306 (N_2306,N_2239,N_2234);
nor U2307 (N_2307,N_2258,N_2276);
nor U2308 (N_2308,N_2257,N_2238);
and U2309 (N_2309,N_2289,N_2214);
nand U2310 (N_2310,N_2260,N_2218);
nor U2311 (N_2311,N_2288,N_2242);
and U2312 (N_2312,N_2237,N_2284);
nand U2313 (N_2313,N_2248,N_2207);
xor U2314 (N_2314,N_2221,N_2219);
and U2315 (N_2315,N_2295,N_2256);
or U2316 (N_2316,N_2282,N_2266);
nand U2317 (N_2317,N_2236,N_2233);
nor U2318 (N_2318,N_2241,N_2231);
and U2319 (N_2319,N_2232,N_2261);
or U2320 (N_2320,N_2208,N_2212);
xor U2321 (N_2321,N_2286,N_2263);
nand U2322 (N_2322,N_2272,N_2287);
nor U2323 (N_2323,N_2255,N_2229);
or U2324 (N_2324,N_2243,N_2280);
nor U2325 (N_2325,N_2275,N_2235);
or U2326 (N_2326,N_2273,N_2293);
or U2327 (N_2327,N_2277,N_2216);
nand U2328 (N_2328,N_2203,N_2291);
nand U2329 (N_2329,N_2226,N_2262);
xnor U2330 (N_2330,N_2247,N_2202);
nor U2331 (N_2331,N_2298,N_2227);
nand U2332 (N_2332,N_2265,N_2244);
or U2333 (N_2333,N_2299,N_2274);
or U2334 (N_2334,N_2211,N_2201);
or U2335 (N_2335,N_2253,N_2240);
and U2336 (N_2336,N_2246,N_2297);
nand U2337 (N_2337,N_2213,N_2220);
nor U2338 (N_2338,N_2224,N_2205);
nor U2339 (N_2339,N_2294,N_2279);
and U2340 (N_2340,N_2271,N_2245);
or U2341 (N_2341,N_2206,N_2252);
or U2342 (N_2342,N_2249,N_2269);
nand U2343 (N_2343,N_2285,N_2281);
nor U2344 (N_2344,N_2230,N_2268);
or U2345 (N_2345,N_2200,N_2210);
xor U2346 (N_2346,N_2209,N_2290);
and U2347 (N_2347,N_2204,N_2222);
and U2348 (N_2348,N_2228,N_2225);
and U2349 (N_2349,N_2278,N_2283);
nand U2350 (N_2350,N_2218,N_2262);
and U2351 (N_2351,N_2253,N_2236);
nor U2352 (N_2352,N_2299,N_2257);
xnor U2353 (N_2353,N_2233,N_2246);
xor U2354 (N_2354,N_2214,N_2283);
nor U2355 (N_2355,N_2243,N_2249);
or U2356 (N_2356,N_2270,N_2293);
nor U2357 (N_2357,N_2223,N_2217);
nand U2358 (N_2358,N_2234,N_2214);
xnor U2359 (N_2359,N_2219,N_2282);
or U2360 (N_2360,N_2212,N_2266);
nand U2361 (N_2361,N_2239,N_2274);
xnor U2362 (N_2362,N_2289,N_2228);
xor U2363 (N_2363,N_2258,N_2283);
and U2364 (N_2364,N_2264,N_2211);
and U2365 (N_2365,N_2228,N_2216);
xnor U2366 (N_2366,N_2209,N_2274);
and U2367 (N_2367,N_2204,N_2254);
or U2368 (N_2368,N_2281,N_2276);
nor U2369 (N_2369,N_2276,N_2236);
xnor U2370 (N_2370,N_2267,N_2289);
and U2371 (N_2371,N_2262,N_2203);
xor U2372 (N_2372,N_2279,N_2202);
nor U2373 (N_2373,N_2260,N_2204);
or U2374 (N_2374,N_2219,N_2245);
nor U2375 (N_2375,N_2231,N_2213);
and U2376 (N_2376,N_2245,N_2243);
nor U2377 (N_2377,N_2270,N_2203);
nor U2378 (N_2378,N_2273,N_2251);
and U2379 (N_2379,N_2224,N_2252);
nand U2380 (N_2380,N_2206,N_2222);
nor U2381 (N_2381,N_2233,N_2296);
xnor U2382 (N_2382,N_2268,N_2254);
xnor U2383 (N_2383,N_2203,N_2298);
nand U2384 (N_2384,N_2250,N_2239);
nand U2385 (N_2385,N_2263,N_2215);
or U2386 (N_2386,N_2269,N_2205);
nand U2387 (N_2387,N_2269,N_2204);
nand U2388 (N_2388,N_2213,N_2221);
and U2389 (N_2389,N_2286,N_2208);
xor U2390 (N_2390,N_2241,N_2294);
nand U2391 (N_2391,N_2252,N_2235);
and U2392 (N_2392,N_2299,N_2239);
and U2393 (N_2393,N_2225,N_2215);
and U2394 (N_2394,N_2237,N_2290);
nor U2395 (N_2395,N_2255,N_2295);
or U2396 (N_2396,N_2272,N_2258);
or U2397 (N_2397,N_2288,N_2228);
nand U2398 (N_2398,N_2297,N_2276);
or U2399 (N_2399,N_2205,N_2287);
nand U2400 (N_2400,N_2351,N_2337);
and U2401 (N_2401,N_2387,N_2322);
or U2402 (N_2402,N_2384,N_2316);
nand U2403 (N_2403,N_2325,N_2308);
and U2404 (N_2404,N_2362,N_2341);
nand U2405 (N_2405,N_2335,N_2302);
and U2406 (N_2406,N_2339,N_2324);
nand U2407 (N_2407,N_2357,N_2328);
nor U2408 (N_2408,N_2393,N_2307);
nand U2409 (N_2409,N_2379,N_2381);
and U2410 (N_2410,N_2336,N_2354);
nor U2411 (N_2411,N_2358,N_2313);
nand U2412 (N_2412,N_2368,N_2378);
nor U2413 (N_2413,N_2303,N_2323);
nor U2414 (N_2414,N_2320,N_2388);
and U2415 (N_2415,N_2329,N_2355);
xnor U2416 (N_2416,N_2349,N_2359);
nor U2417 (N_2417,N_2318,N_2314);
or U2418 (N_2418,N_2300,N_2334);
xor U2419 (N_2419,N_2363,N_2306);
and U2420 (N_2420,N_2309,N_2389);
and U2421 (N_2421,N_2312,N_2360);
or U2422 (N_2422,N_2304,N_2352);
nand U2423 (N_2423,N_2348,N_2390);
nand U2424 (N_2424,N_2305,N_2376);
xnor U2425 (N_2425,N_2373,N_2398);
nand U2426 (N_2426,N_2311,N_2331);
or U2427 (N_2427,N_2338,N_2394);
nand U2428 (N_2428,N_2332,N_2371);
nand U2429 (N_2429,N_2391,N_2392);
nor U2430 (N_2430,N_2365,N_2374);
and U2431 (N_2431,N_2345,N_2369);
and U2432 (N_2432,N_2340,N_2367);
xnor U2433 (N_2433,N_2397,N_2364);
and U2434 (N_2434,N_2386,N_2385);
xor U2435 (N_2435,N_2350,N_2356);
or U2436 (N_2436,N_2321,N_2383);
xor U2437 (N_2437,N_2344,N_2333);
and U2438 (N_2438,N_2315,N_2380);
xor U2439 (N_2439,N_2372,N_2370);
nand U2440 (N_2440,N_2377,N_2346);
xor U2441 (N_2441,N_2319,N_2366);
or U2442 (N_2442,N_2396,N_2327);
xnor U2443 (N_2443,N_2353,N_2361);
or U2444 (N_2444,N_2347,N_2382);
and U2445 (N_2445,N_2399,N_2317);
and U2446 (N_2446,N_2395,N_2330);
or U2447 (N_2447,N_2343,N_2342);
and U2448 (N_2448,N_2375,N_2310);
nor U2449 (N_2449,N_2301,N_2326);
or U2450 (N_2450,N_2312,N_2348);
and U2451 (N_2451,N_2396,N_2392);
nor U2452 (N_2452,N_2355,N_2320);
xnor U2453 (N_2453,N_2311,N_2310);
nor U2454 (N_2454,N_2321,N_2304);
nand U2455 (N_2455,N_2366,N_2346);
nand U2456 (N_2456,N_2376,N_2374);
and U2457 (N_2457,N_2328,N_2344);
xor U2458 (N_2458,N_2343,N_2390);
nand U2459 (N_2459,N_2388,N_2377);
nor U2460 (N_2460,N_2386,N_2355);
nand U2461 (N_2461,N_2378,N_2327);
xor U2462 (N_2462,N_2393,N_2324);
and U2463 (N_2463,N_2395,N_2300);
xor U2464 (N_2464,N_2316,N_2325);
and U2465 (N_2465,N_2380,N_2361);
xor U2466 (N_2466,N_2302,N_2377);
nand U2467 (N_2467,N_2316,N_2370);
nor U2468 (N_2468,N_2384,N_2394);
nand U2469 (N_2469,N_2313,N_2352);
or U2470 (N_2470,N_2344,N_2340);
nand U2471 (N_2471,N_2342,N_2399);
and U2472 (N_2472,N_2367,N_2371);
nor U2473 (N_2473,N_2318,N_2363);
xnor U2474 (N_2474,N_2384,N_2303);
xnor U2475 (N_2475,N_2326,N_2325);
nor U2476 (N_2476,N_2386,N_2362);
or U2477 (N_2477,N_2376,N_2383);
and U2478 (N_2478,N_2384,N_2330);
nand U2479 (N_2479,N_2370,N_2357);
xnor U2480 (N_2480,N_2372,N_2317);
xnor U2481 (N_2481,N_2358,N_2386);
or U2482 (N_2482,N_2363,N_2371);
nand U2483 (N_2483,N_2380,N_2357);
and U2484 (N_2484,N_2320,N_2364);
nand U2485 (N_2485,N_2373,N_2304);
xor U2486 (N_2486,N_2358,N_2307);
or U2487 (N_2487,N_2383,N_2386);
nand U2488 (N_2488,N_2367,N_2323);
xor U2489 (N_2489,N_2321,N_2343);
nor U2490 (N_2490,N_2323,N_2313);
and U2491 (N_2491,N_2359,N_2369);
or U2492 (N_2492,N_2385,N_2325);
or U2493 (N_2493,N_2350,N_2360);
xor U2494 (N_2494,N_2320,N_2310);
nand U2495 (N_2495,N_2368,N_2334);
and U2496 (N_2496,N_2358,N_2355);
or U2497 (N_2497,N_2311,N_2385);
xnor U2498 (N_2498,N_2362,N_2339);
xor U2499 (N_2499,N_2368,N_2355);
or U2500 (N_2500,N_2452,N_2421);
nor U2501 (N_2501,N_2417,N_2498);
nor U2502 (N_2502,N_2454,N_2418);
or U2503 (N_2503,N_2485,N_2478);
xor U2504 (N_2504,N_2446,N_2451);
xor U2505 (N_2505,N_2455,N_2470);
nor U2506 (N_2506,N_2490,N_2435);
and U2507 (N_2507,N_2484,N_2458);
or U2508 (N_2508,N_2469,N_2493);
nor U2509 (N_2509,N_2433,N_2434);
nor U2510 (N_2510,N_2431,N_2477);
xnor U2511 (N_2511,N_2487,N_2447);
xnor U2512 (N_2512,N_2456,N_2440);
and U2513 (N_2513,N_2411,N_2423);
or U2514 (N_2514,N_2492,N_2460);
nor U2515 (N_2515,N_2481,N_2467);
or U2516 (N_2516,N_2429,N_2413);
nand U2517 (N_2517,N_2461,N_2479);
or U2518 (N_2518,N_2437,N_2459);
or U2519 (N_2519,N_2466,N_2400);
nor U2520 (N_2520,N_2457,N_2499);
nand U2521 (N_2521,N_2444,N_2428);
or U2522 (N_2522,N_2401,N_2419);
and U2523 (N_2523,N_2473,N_2409);
and U2524 (N_2524,N_2441,N_2443);
and U2525 (N_2525,N_2416,N_2450);
or U2526 (N_2526,N_2474,N_2449);
and U2527 (N_2527,N_2489,N_2425);
xnor U2528 (N_2528,N_2415,N_2476);
xnor U2529 (N_2529,N_2480,N_2436);
and U2530 (N_2530,N_2406,N_2439);
nor U2531 (N_2531,N_2472,N_2463);
xor U2532 (N_2532,N_2404,N_2488);
nor U2533 (N_2533,N_2427,N_2465);
nor U2534 (N_2534,N_2442,N_2412);
nor U2535 (N_2535,N_2420,N_2486);
nor U2536 (N_2536,N_2453,N_2438);
xor U2537 (N_2537,N_2424,N_2482);
and U2538 (N_2538,N_2405,N_2414);
nand U2539 (N_2539,N_2491,N_2475);
nand U2540 (N_2540,N_2448,N_2410);
xor U2541 (N_2541,N_2496,N_2497);
or U2542 (N_2542,N_2462,N_2471);
nor U2543 (N_2543,N_2426,N_2445);
nor U2544 (N_2544,N_2464,N_2402);
xnor U2545 (N_2545,N_2483,N_2408);
nand U2546 (N_2546,N_2422,N_2407);
xor U2547 (N_2547,N_2430,N_2495);
nor U2548 (N_2548,N_2403,N_2468);
nor U2549 (N_2549,N_2432,N_2494);
or U2550 (N_2550,N_2452,N_2410);
nor U2551 (N_2551,N_2462,N_2416);
or U2552 (N_2552,N_2425,N_2439);
nor U2553 (N_2553,N_2420,N_2478);
nand U2554 (N_2554,N_2444,N_2409);
nand U2555 (N_2555,N_2403,N_2458);
xor U2556 (N_2556,N_2442,N_2425);
nand U2557 (N_2557,N_2421,N_2436);
nor U2558 (N_2558,N_2477,N_2486);
or U2559 (N_2559,N_2404,N_2405);
nand U2560 (N_2560,N_2435,N_2485);
nor U2561 (N_2561,N_2439,N_2473);
and U2562 (N_2562,N_2470,N_2463);
nor U2563 (N_2563,N_2431,N_2455);
xor U2564 (N_2564,N_2419,N_2452);
and U2565 (N_2565,N_2435,N_2477);
or U2566 (N_2566,N_2400,N_2476);
xor U2567 (N_2567,N_2436,N_2437);
nor U2568 (N_2568,N_2468,N_2435);
nand U2569 (N_2569,N_2497,N_2412);
nor U2570 (N_2570,N_2408,N_2411);
or U2571 (N_2571,N_2477,N_2428);
nand U2572 (N_2572,N_2485,N_2443);
nor U2573 (N_2573,N_2474,N_2460);
xnor U2574 (N_2574,N_2443,N_2439);
or U2575 (N_2575,N_2466,N_2487);
nand U2576 (N_2576,N_2414,N_2418);
or U2577 (N_2577,N_2431,N_2414);
nor U2578 (N_2578,N_2487,N_2442);
xnor U2579 (N_2579,N_2440,N_2415);
nor U2580 (N_2580,N_2417,N_2449);
xnor U2581 (N_2581,N_2412,N_2443);
and U2582 (N_2582,N_2411,N_2428);
and U2583 (N_2583,N_2488,N_2487);
xor U2584 (N_2584,N_2448,N_2420);
and U2585 (N_2585,N_2434,N_2430);
nand U2586 (N_2586,N_2442,N_2406);
and U2587 (N_2587,N_2487,N_2425);
xnor U2588 (N_2588,N_2406,N_2444);
or U2589 (N_2589,N_2478,N_2467);
and U2590 (N_2590,N_2428,N_2410);
nor U2591 (N_2591,N_2418,N_2432);
nor U2592 (N_2592,N_2403,N_2441);
xor U2593 (N_2593,N_2433,N_2487);
nor U2594 (N_2594,N_2403,N_2475);
nor U2595 (N_2595,N_2465,N_2434);
xnor U2596 (N_2596,N_2467,N_2494);
nand U2597 (N_2597,N_2414,N_2432);
nand U2598 (N_2598,N_2405,N_2422);
xnor U2599 (N_2599,N_2461,N_2454);
and U2600 (N_2600,N_2518,N_2519);
xor U2601 (N_2601,N_2586,N_2505);
nand U2602 (N_2602,N_2566,N_2559);
or U2603 (N_2603,N_2544,N_2510);
xor U2604 (N_2604,N_2571,N_2537);
nand U2605 (N_2605,N_2500,N_2582);
nand U2606 (N_2606,N_2554,N_2520);
or U2607 (N_2607,N_2540,N_2546);
or U2608 (N_2608,N_2541,N_2576);
and U2609 (N_2609,N_2543,N_2588);
nor U2610 (N_2610,N_2532,N_2577);
xnor U2611 (N_2611,N_2530,N_2511);
or U2612 (N_2612,N_2597,N_2527);
nand U2613 (N_2613,N_2592,N_2512);
nand U2614 (N_2614,N_2517,N_2563);
xnor U2615 (N_2615,N_2545,N_2552);
and U2616 (N_2616,N_2598,N_2504);
nand U2617 (N_2617,N_2523,N_2565);
nand U2618 (N_2618,N_2580,N_2596);
or U2619 (N_2619,N_2553,N_2595);
nand U2620 (N_2620,N_2549,N_2562);
or U2621 (N_2621,N_2568,N_2539);
nand U2622 (N_2622,N_2521,N_2534);
xor U2623 (N_2623,N_2567,N_2579);
nor U2624 (N_2624,N_2536,N_2593);
nand U2625 (N_2625,N_2525,N_2501);
nand U2626 (N_2626,N_2550,N_2535);
and U2627 (N_2627,N_2594,N_2533);
nor U2628 (N_2628,N_2526,N_2529);
xnor U2629 (N_2629,N_2589,N_2502);
nor U2630 (N_2630,N_2514,N_2584);
xor U2631 (N_2631,N_2538,N_2547);
and U2632 (N_2632,N_2561,N_2564);
and U2633 (N_2633,N_2513,N_2555);
xor U2634 (N_2634,N_2542,N_2516);
nand U2635 (N_2635,N_2581,N_2509);
xor U2636 (N_2636,N_2508,N_2556);
nand U2637 (N_2637,N_2551,N_2587);
xnor U2638 (N_2638,N_2548,N_2531);
xor U2639 (N_2639,N_2583,N_2578);
nand U2640 (N_2640,N_2574,N_2503);
or U2641 (N_2641,N_2522,N_2528);
and U2642 (N_2642,N_2573,N_2590);
or U2643 (N_2643,N_2524,N_2507);
nand U2644 (N_2644,N_2591,N_2575);
and U2645 (N_2645,N_2585,N_2569);
or U2646 (N_2646,N_2599,N_2558);
nand U2647 (N_2647,N_2506,N_2515);
and U2648 (N_2648,N_2572,N_2560);
xnor U2649 (N_2649,N_2557,N_2570);
or U2650 (N_2650,N_2543,N_2592);
and U2651 (N_2651,N_2513,N_2518);
nor U2652 (N_2652,N_2565,N_2597);
nand U2653 (N_2653,N_2594,N_2599);
nand U2654 (N_2654,N_2537,N_2522);
or U2655 (N_2655,N_2559,N_2504);
and U2656 (N_2656,N_2516,N_2587);
nor U2657 (N_2657,N_2584,N_2583);
or U2658 (N_2658,N_2592,N_2596);
and U2659 (N_2659,N_2570,N_2571);
nand U2660 (N_2660,N_2529,N_2573);
or U2661 (N_2661,N_2595,N_2524);
nand U2662 (N_2662,N_2566,N_2580);
nand U2663 (N_2663,N_2594,N_2573);
xor U2664 (N_2664,N_2524,N_2570);
nor U2665 (N_2665,N_2577,N_2514);
and U2666 (N_2666,N_2574,N_2506);
or U2667 (N_2667,N_2584,N_2596);
or U2668 (N_2668,N_2529,N_2527);
nand U2669 (N_2669,N_2562,N_2582);
and U2670 (N_2670,N_2532,N_2534);
nor U2671 (N_2671,N_2504,N_2595);
and U2672 (N_2672,N_2569,N_2556);
nor U2673 (N_2673,N_2593,N_2533);
xnor U2674 (N_2674,N_2574,N_2510);
and U2675 (N_2675,N_2558,N_2517);
nand U2676 (N_2676,N_2585,N_2595);
or U2677 (N_2677,N_2569,N_2586);
xor U2678 (N_2678,N_2578,N_2537);
nand U2679 (N_2679,N_2593,N_2590);
or U2680 (N_2680,N_2583,N_2562);
and U2681 (N_2681,N_2594,N_2544);
xnor U2682 (N_2682,N_2576,N_2590);
nand U2683 (N_2683,N_2507,N_2589);
nor U2684 (N_2684,N_2568,N_2579);
and U2685 (N_2685,N_2524,N_2541);
or U2686 (N_2686,N_2508,N_2553);
and U2687 (N_2687,N_2569,N_2527);
nand U2688 (N_2688,N_2520,N_2502);
nand U2689 (N_2689,N_2545,N_2599);
or U2690 (N_2690,N_2595,N_2565);
and U2691 (N_2691,N_2530,N_2554);
xor U2692 (N_2692,N_2550,N_2501);
and U2693 (N_2693,N_2599,N_2568);
and U2694 (N_2694,N_2503,N_2544);
or U2695 (N_2695,N_2575,N_2515);
and U2696 (N_2696,N_2574,N_2532);
and U2697 (N_2697,N_2574,N_2521);
nor U2698 (N_2698,N_2515,N_2512);
nor U2699 (N_2699,N_2507,N_2586);
xor U2700 (N_2700,N_2620,N_2698);
and U2701 (N_2701,N_2697,N_2672);
xor U2702 (N_2702,N_2693,N_2627);
nand U2703 (N_2703,N_2609,N_2632);
or U2704 (N_2704,N_2699,N_2610);
and U2705 (N_2705,N_2624,N_2664);
and U2706 (N_2706,N_2602,N_2611);
nor U2707 (N_2707,N_2630,N_2660);
nor U2708 (N_2708,N_2638,N_2669);
nor U2709 (N_2709,N_2604,N_2651);
xor U2710 (N_2710,N_2637,N_2652);
xnor U2711 (N_2711,N_2655,N_2617);
nand U2712 (N_2712,N_2646,N_2645);
nand U2713 (N_2713,N_2670,N_2626);
xor U2714 (N_2714,N_2603,N_2692);
nand U2715 (N_2715,N_2668,N_2654);
and U2716 (N_2716,N_2607,N_2673);
or U2717 (N_2717,N_2621,N_2648);
xnor U2718 (N_2718,N_2663,N_2633);
xnor U2719 (N_2719,N_2671,N_2696);
or U2720 (N_2720,N_2639,N_2691);
and U2721 (N_2721,N_2682,N_2619);
and U2722 (N_2722,N_2600,N_2684);
xnor U2723 (N_2723,N_2658,N_2659);
nand U2724 (N_2724,N_2680,N_2675);
nor U2725 (N_2725,N_2613,N_2674);
or U2726 (N_2726,N_2641,N_2631);
xor U2727 (N_2727,N_2685,N_2643);
and U2728 (N_2728,N_2618,N_2678);
nor U2729 (N_2729,N_2647,N_2616);
nand U2730 (N_2730,N_2628,N_2653);
nand U2731 (N_2731,N_2612,N_2683);
or U2732 (N_2732,N_2677,N_2676);
and U2733 (N_2733,N_2667,N_2642);
nor U2734 (N_2734,N_2636,N_2649);
and U2735 (N_2735,N_2615,N_2686);
and U2736 (N_2736,N_2614,N_2608);
nand U2737 (N_2737,N_2656,N_2629);
nand U2738 (N_2738,N_2635,N_2640);
xor U2739 (N_2739,N_2666,N_2625);
or U2740 (N_2740,N_2644,N_2634);
xnor U2741 (N_2741,N_2662,N_2657);
nand U2742 (N_2742,N_2623,N_2679);
nor U2743 (N_2743,N_2689,N_2690);
and U2744 (N_2744,N_2622,N_2694);
nor U2745 (N_2745,N_2688,N_2605);
or U2746 (N_2746,N_2650,N_2601);
xnor U2747 (N_2747,N_2695,N_2661);
nor U2748 (N_2748,N_2606,N_2687);
and U2749 (N_2749,N_2681,N_2665);
and U2750 (N_2750,N_2679,N_2689);
and U2751 (N_2751,N_2687,N_2682);
nand U2752 (N_2752,N_2682,N_2612);
nand U2753 (N_2753,N_2672,N_2614);
xor U2754 (N_2754,N_2640,N_2664);
nor U2755 (N_2755,N_2649,N_2642);
nor U2756 (N_2756,N_2673,N_2626);
xor U2757 (N_2757,N_2665,N_2637);
or U2758 (N_2758,N_2676,N_2616);
xor U2759 (N_2759,N_2605,N_2633);
xnor U2760 (N_2760,N_2656,N_2664);
xor U2761 (N_2761,N_2689,N_2697);
nand U2762 (N_2762,N_2631,N_2636);
nand U2763 (N_2763,N_2635,N_2692);
xor U2764 (N_2764,N_2666,N_2622);
xnor U2765 (N_2765,N_2681,N_2613);
or U2766 (N_2766,N_2692,N_2636);
xnor U2767 (N_2767,N_2602,N_2694);
or U2768 (N_2768,N_2604,N_2659);
nor U2769 (N_2769,N_2683,N_2626);
nor U2770 (N_2770,N_2668,N_2681);
or U2771 (N_2771,N_2676,N_2615);
nor U2772 (N_2772,N_2652,N_2673);
and U2773 (N_2773,N_2626,N_2657);
nand U2774 (N_2774,N_2686,N_2632);
xnor U2775 (N_2775,N_2634,N_2667);
and U2776 (N_2776,N_2689,N_2674);
xnor U2777 (N_2777,N_2665,N_2657);
or U2778 (N_2778,N_2649,N_2651);
nor U2779 (N_2779,N_2681,N_2653);
nand U2780 (N_2780,N_2698,N_2668);
and U2781 (N_2781,N_2629,N_2631);
xor U2782 (N_2782,N_2602,N_2632);
nand U2783 (N_2783,N_2626,N_2611);
nor U2784 (N_2784,N_2640,N_2694);
nor U2785 (N_2785,N_2684,N_2634);
xnor U2786 (N_2786,N_2664,N_2620);
and U2787 (N_2787,N_2698,N_2650);
xnor U2788 (N_2788,N_2636,N_2619);
or U2789 (N_2789,N_2612,N_2604);
nand U2790 (N_2790,N_2657,N_2638);
nand U2791 (N_2791,N_2676,N_2696);
and U2792 (N_2792,N_2602,N_2687);
or U2793 (N_2793,N_2671,N_2607);
nand U2794 (N_2794,N_2694,N_2652);
xnor U2795 (N_2795,N_2698,N_2674);
xor U2796 (N_2796,N_2677,N_2672);
and U2797 (N_2797,N_2666,N_2698);
nand U2798 (N_2798,N_2647,N_2684);
nand U2799 (N_2799,N_2686,N_2638);
xor U2800 (N_2800,N_2727,N_2725);
xor U2801 (N_2801,N_2752,N_2726);
nor U2802 (N_2802,N_2724,N_2731);
or U2803 (N_2803,N_2775,N_2771);
xor U2804 (N_2804,N_2721,N_2760);
and U2805 (N_2805,N_2705,N_2782);
xor U2806 (N_2806,N_2745,N_2794);
nand U2807 (N_2807,N_2715,N_2722);
or U2808 (N_2808,N_2763,N_2723);
xor U2809 (N_2809,N_2714,N_2700);
and U2810 (N_2810,N_2785,N_2786);
nand U2811 (N_2811,N_2748,N_2730);
nand U2812 (N_2812,N_2793,N_2750);
or U2813 (N_2813,N_2741,N_2767);
and U2814 (N_2814,N_2756,N_2779);
and U2815 (N_2815,N_2704,N_2766);
and U2816 (N_2816,N_2747,N_2762);
nor U2817 (N_2817,N_2773,N_2784);
or U2818 (N_2818,N_2729,N_2795);
or U2819 (N_2819,N_2751,N_2736);
nor U2820 (N_2820,N_2708,N_2753);
xor U2821 (N_2821,N_2706,N_2798);
or U2822 (N_2822,N_2709,N_2716);
nor U2823 (N_2823,N_2769,N_2710);
and U2824 (N_2824,N_2718,N_2799);
xnor U2825 (N_2825,N_2738,N_2743);
nand U2826 (N_2826,N_2765,N_2761);
nand U2827 (N_2827,N_2789,N_2717);
or U2828 (N_2828,N_2713,N_2787);
nor U2829 (N_2829,N_2788,N_2758);
or U2830 (N_2830,N_2792,N_2732);
or U2831 (N_2831,N_2720,N_2757);
nor U2832 (N_2832,N_2764,N_2755);
xor U2833 (N_2833,N_2791,N_2781);
xnor U2834 (N_2834,N_2719,N_2707);
or U2835 (N_2835,N_2749,N_2701);
nand U2836 (N_2836,N_2790,N_2735);
nor U2837 (N_2837,N_2740,N_2733);
or U2838 (N_2838,N_2739,N_2754);
nand U2839 (N_2839,N_2744,N_2742);
and U2840 (N_2840,N_2776,N_2734);
xor U2841 (N_2841,N_2777,N_2774);
and U2842 (N_2842,N_2712,N_2711);
nand U2843 (N_2843,N_2778,N_2772);
xnor U2844 (N_2844,N_2796,N_2797);
nor U2845 (N_2845,N_2768,N_2737);
nand U2846 (N_2846,N_2703,N_2780);
or U2847 (N_2847,N_2702,N_2770);
nor U2848 (N_2848,N_2783,N_2746);
xnor U2849 (N_2849,N_2759,N_2728);
nand U2850 (N_2850,N_2799,N_2778);
xnor U2851 (N_2851,N_2728,N_2778);
or U2852 (N_2852,N_2743,N_2713);
and U2853 (N_2853,N_2761,N_2703);
or U2854 (N_2854,N_2774,N_2789);
nor U2855 (N_2855,N_2786,N_2797);
nand U2856 (N_2856,N_2797,N_2779);
nand U2857 (N_2857,N_2777,N_2715);
xor U2858 (N_2858,N_2705,N_2797);
nand U2859 (N_2859,N_2725,N_2708);
xor U2860 (N_2860,N_2779,N_2706);
nor U2861 (N_2861,N_2701,N_2752);
or U2862 (N_2862,N_2776,N_2715);
xnor U2863 (N_2863,N_2743,N_2715);
or U2864 (N_2864,N_2783,N_2756);
and U2865 (N_2865,N_2737,N_2750);
xor U2866 (N_2866,N_2737,N_2742);
nand U2867 (N_2867,N_2724,N_2765);
and U2868 (N_2868,N_2792,N_2778);
nor U2869 (N_2869,N_2780,N_2761);
nor U2870 (N_2870,N_2727,N_2726);
nand U2871 (N_2871,N_2762,N_2786);
nor U2872 (N_2872,N_2742,N_2711);
nand U2873 (N_2873,N_2745,N_2786);
or U2874 (N_2874,N_2723,N_2785);
xor U2875 (N_2875,N_2719,N_2745);
or U2876 (N_2876,N_2749,N_2714);
xor U2877 (N_2877,N_2762,N_2740);
nand U2878 (N_2878,N_2757,N_2755);
xnor U2879 (N_2879,N_2738,N_2715);
nand U2880 (N_2880,N_2793,N_2799);
nor U2881 (N_2881,N_2724,N_2773);
and U2882 (N_2882,N_2711,N_2787);
nor U2883 (N_2883,N_2757,N_2744);
and U2884 (N_2884,N_2763,N_2730);
nor U2885 (N_2885,N_2780,N_2763);
and U2886 (N_2886,N_2709,N_2700);
nor U2887 (N_2887,N_2700,N_2750);
and U2888 (N_2888,N_2792,N_2700);
nand U2889 (N_2889,N_2742,N_2779);
xnor U2890 (N_2890,N_2708,N_2775);
or U2891 (N_2891,N_2765,N_2784);
and U2892 (N_2892,N_2785,N_2705);
nor U2893 (N_2893,N_2713,N_2757);
and U2894 (N_2894,N_2781,N_2749);
or U2895 (N_2895,N_2796,N_2728);
xnor U2896 (N_2896,N_2781,N_2779);
nor U2897 (N_2897,N_2757,N_2705);
and U2898 (N_2898,N_2777,N_2741);
nor U2899 (N_2899,N_2790,N_2786);
nand U2900 (N_2900,N_2880,N_2891);
xnor U2901 (N_2901,N_2849,N_2872);
and U2902 (N_2902,N_2877,N_2894);
nand U2903 (N_2903,N_2855,N_2806);
nand U2904 (N_2904,N_2848,N_2852);
and U2905 (N_2905,N_2838,N_2842);
and U2906 (N_2906,N_2828,N_2865);
nor U2907 (N_2907,N_2885,N_2809);
and U2908 (N_2908,N_2823,N_2890);
and U2909 (N_2909,N_2854,N_2857);
xor U2910 (N_2910,N_2878,N_2863);
nand U2911 (N_2911,N_2811,N_2864);
xnor U2912 (N_2912,N_2861,N_2888);
xnor U2913 (N_2913,N_2841,N_2802);
or U2914 (N_2914,N_2850,N_2843);
nand U2915 (N_2915,N_2886,N_2853);
and U2916 (N_2916,N_2858,N_2898);
nand U2917 (N_2917,N_2830,N_2889);
nor U2918 (N_2918,N_2873,N_2800);
nand U2919 (N_2919,N_2803,N_2836);
xnor U2920 (N_2920,N_2810,N_2897);
xnor U2921 (N_2921,N_2815,N_2851);
nand U2922 (N_2922,N_2881,N_2859);
and U2923 (N_2923,N_2825,N_2821);
nor U2924 (N_2924,N_2847,N_2867);
and U2925 (N_2925,N_2899,N_2808);
and U2926 (N_2926,N_2871,N_2822);
xnor U2927 (N_2927,N_2845,N_2870);
nand U2928 (N_2928,N_2837,N_2805);
nor U2929 (N_2929,N_2835,N_2820);
or U2930 (N_2930,N_2844,N_2829);
nand U2931 (N_2931,N_2807,N_2812);
nand U2932 (N_2932,N_2868,N_2869);
xor U2933 (N_2933,N_2883,N_2801);
and U2934 (N_2934,N_2892,N_2846);
nor U2935 (N_2935,N_2896,N_2879);
xor U2936 (N_2936,N_2826,N_2832);
nor U2937 (N_2937,N_2819,N_2817);
nand U2938 (N_2938,N_2834,N_2875);
or U2939 (N_2939,N_2804,N_2818);
or U2940 (N_2940,N_2814,N_2831);
nand U2941 (N_2941,N_2876,N_2893);
nand U2942 (N_2942,N_2839,N_2884);
xnor U2943 (N_2943,N_2862,N_2874);
and U2944 (N_2944,N_2833,N_2887);
nor U2945 (N_2945,N_2816,N_2860);
and U2946 (N_2946,N_2840,N_2813);
or U2947 (N_2947,N_2856,N_2827);
nor U2948 (N_2948,N_2882,N_2824);
nor U2949 (N_2949,N_2895,N_2866);
or U2950 (N_2950,N_2820,N_2816);
nand U2951 (N_2951,N_2840,N_2841);
xor U2952 (N_2952,N_2802,N_2886);
or U2953 (N_2953,N_2826,N_2857);
nand U2954 (N_2954,N_2846,N_2810);
or U2955 (N_2955,N_2881,N_2897);
or U2956 (N_2956,N_2818,N_2858);
xor U2957 (N_2957,N_2853,N_2877);
and U2958 (N_2958,N_2879,N_2818);
nor U2959 (N_2959,N_2864,N_2836);
nand U2960 (N_2960,N_2849,N_2895);
and U2961 (N_2961,N_2812,N_2875);
and U2962 (N_2962,N_2868,N_2838);
or U2963 (N_2963,N_2836,N_2823);
or U2964 (N_2964,N_2806,N_2892);
and U2965 (N_2965,N_2889,N_2803);
nor U2966 (N_2966,N_2888,N_2871);
nor U2967 (N_2967,N_2891,N_2853);
and U2968 (N_2968,N_2881,N_2853);
nor U2969 (N_2969,N_2847,N_2872);
xor U2970 (N_2970,N_2895,N_2825);
and U2971 (N_2971,N_2890,N_2852);
xor U2972 (N_2972,N_2863,N_2803);
and U2973 (N_2973,N_2854,N_2888);
and U2974 (N_2974,N_2849,N_2893);
or U2975 (N_2975,N_2859,N_2829);
nand U2976 (N_2976,N_2835,N_2858);
nor U2977 (N_2977,N_2836,N_2879);
nand U2978 (N_2978,N_2825,N_2896);
nand U2979 (N_2979,N_2847,N_2881);
nand U2980 (N_2980,N_2854,N_2847);
nand U2981 (N_2981,N_2882,N_2885);
or U2982 (N_2982,N_2801,N_2874);
nand U2983 (N_2983,N_2802,N_2850);
nor U2984 (N_2984,N_2856,N_2881);
xor U2985 (N_2985,N_2874,N_2827);
or U2986 (N_2986,N_2870,N_2890);
or U2987 (N_2987,N_2802,N_2860);
xor U2988 (N_2988,N_2831,N_2811);
xor U2989 (N_2989,N_2878,N_2802);
nand U2990 (N_2990,N_2862,N_2831);
and U2991 (N_2991,N_2805,N_2820);
and U2992 (N_2992,N_2847,N_2862);
nor U2993 (N_2993,N_2813,N_2880);
and U2994 (N_2994,N_2851,N_2873);
and U2995 (N_2995,N_2813,N_2891);
xnor U2996 (N_2996,N_2823,N_2824);
nand U2997 (N_2997,N_2867,N_2857);
nor U2998 (N_2998,N_2882,N_2846);
xor U2999 (N_2999,N_2886,N_2855);
or U3000 (N_3000,N_2977,N_2994);
xnor U3001 (N_3001,N_2959,N_2922);
nor U3002 (N_3002,N_2976,N_2903);
nand U3003 (N_3003,N_2940,N_2954);
xnor U3004 (N_3004,N_2929,N_2999);
and U3005 (N_3005,N_2909,N_2943);
nand U3006 (N_3006,N_2955,N_2914);
and U3007 (N_3007,N_2950,N_2931);
and U3008 (N_3008,N_2962,N_2949);
or U3009 (N_3009,N_2987,N_2968);
nor U3010 (N_3010,N_2919,N_2956);
or U3011 (N_3011,N_2989,N_2918);
or U3012 (N_3012,N_2985,N_2921);
and U3013 (N_3013,N_2912,N_2917);
nand U3014 (N_3014,N_2951,N_2941);
nor U3015 (N_3015,N_2953,N_2998);
or U3016 (N_3016,N_2983,N_2945);
nor U3017 (N_3017,N_2933,N_2986);
nor U3018 (N_3018,N_2904,N_2958);
and U3019 (N_3019,N_2936,N_2997);
or U3020 (N_3020,N_2974,N_2916);
nand U3021 (N_3021,N_2978,N_2973);
nand U3022 (N_3022,N_2971,N_2923);
nor U3023 (N_3023,N_2930,N_2902);
nand U3024 (N_3024,N_2993,N_2970);
nor U3025 (N_3025,N_2915,N_2960);
xnor U3026 (N_3026,N_2907,N_2935);
or U3027 (N_3027,N_2957,N_2996);
or U3028 (N_3028,N_2961,N_2972);
nand U3029 (N_3029,N_2995,N_2984);
nand U3030 (N_3030,N_2980,N_2900);
and U3031 (N_3031,N_2992,N_2947);
nor U3032 (N_3032,N_2913,N_2939);
nand U3033 (N_3033,N_2966,N_2952);
nand U3034 (N_3034,N_2926,N_2908);
nor U3035 (N_3035,N_2990,N_2901);
or U3036 (N_3036,N_2948,N_2911);
or U3037 (N_3037,N_2924,N_2925);
nand U3038 (N_3038,N_2944,N_2982);
xnor U3039 (N_3039,N_2934,N_2938);
nor U3040 (N_3040,N_2928,N_2975);
or U3041 (N_3041,N_2981,N_2991);
and U3042 (N_3042,N_2969,N_2920);
xnor U3043 (N_3043,N_2942,N_2937);
nor U3044 (N_3044,N_2910,N_2932);
nor U3045 (N_3045,N_2963,N_2979);
nand U3046 (N_3046,N_2946,N_2905);
and U3047 (N_3047,N_2965,N_2988);
nor U3048 (N_3048,N_2967,N_2927);
nand U3049 (N_3049,N_2906,N_2964);
nand U3050 (N_3050,N_2904,N_2980);
or U3051 (N_3051,N_2991,N_2957);
or U3052 (N_3052,N_2964,N_2998);
and U3053 (N_3053,N_2925,N_2981);
nor U3054 (N_3054,N_2956,N_2988);
and U3055 (N_3055,N_2966,N_2907);
or U3056 (N_3056,N_2923,N_2912);
xor U3057 (N_3057,N_2976,N_2964);
xor U3058 (N_3058,N_2979,N_2994);
or U3059 (N_3059,N_2935,N_2981);
nand U3060 (N_3060,N_2964,N_2937);
nand U3061 (N_3061,N_2953,N_2959);
nand U3062 (N_3062,N_2909,N_2948);
or U3063 (N_3063,N_2990,N_2908);
nor U3064 (N_3064,N_2979,N_2967);
or U3065 (N_3065,N_2976,N_2913);
or U3066 (N_3066,N_2975,N_2989);
xor U3067 (N_3067,N_2929,N_2954);
nand U3068 (N_3068,N_2955,N_2976);
nand U3069 (N_3069,N_2920,N_2946);
nor U3070 (N_3070,N_2921,N_2906);
nor U3071 (N_3071,N_2970,N_2910);
and U3072 (N_3072,N_2918,N_2986);
nor U3073 (N_3073,N_2918,N_2947);
or U3074 (N_3074,N_2983,N_2912);
and U3075 (N_3075,N_2939,N_2911);
nand U3076 (N_3076,N_2916,N_2964);
nand U3077 (N_3077,N_2907,N_2929);
xor U3078 (N_3078,N_2971,N_2929);
or U3079 (N_3079,N_2988,N_2911);
or U3080 (N_3080,N_2906,N_2988);
or U3081 (N_3081,N_2931,N_2994);
xnor U3082 (N_3082,N_2942,N_2928);
xnor U3083 (N_3083,N_2962,N_2969);
or U3084 (N_3084,N_2980,N_2901);
xor U3085 (N_3085,N_2938,N_2959);
nand U3086 (N_3086,N_2954,N_2960);
nand U3087 (N_3087,N_2909,N_2976);
or U3088 (N_3088,N_2981,N_2977);
or U3089 (N_3089,N_2962,N_2937);
xor U3090 (N_3090,N_2919,N_2987);
or U3091 (N_3091,N_2900,N_2967);
nor U3092 (N_3092,N_2947,N_2932);
nor U3093 (N_3093,N_2963,N_2987);
xor U3094 (N_3094,N_2938,N_2975);
xor U3095 (N_3095,N_2965,N_2921);
nor U3096 (N_3096,N_2997,N_2983);
nand U3097 (N_3097,N_2949,N_2945);
nand U3098 (N_3098,N_2935,N_2976);
nor U3099 (N_3099,N_2910,N_2936);
xor U3100 (N_3100,N_3063,N_3048);
nor U3101 (N_3101,N_3024,N_3042);
xor U3102 (N_3102,N_3074,N_3045);
nor U3103 (N_3103,N_3060,N_3083);
or U3104 (N_3104,N_3058,N_3002);
xor U3105 (N_3105,N_3034,N_3015);
and U3106 (N_3106,N_3062,N_3089);
nand U3107 (N_3107,N_3037,N_3043);
xnor U3108 (N_3108,N_3029,N_3028);
nand U3109 (N_3109,N_3084,N_3082);
nand U3110 (N_3110,N_3080,N_3038);
or U3111 (N_3111,N_3092,N_3033);
or U3112 (N_3112,N_3039,N_3016);
or U3113 (N_3113,N_3066,N_3085);
or U3114 (N_3114,N_3075,N_3098);
xnor U3115 (N_3115,N_3049,N_3050);
or U3116 (N_3116,N_3069,N_3055);
xor U3117 (N_3117,N_3065,N_3009);
xnor U3118 (N_3118,N_3046,N_3001);
and U3119 (N_3119,N_3088,N_3004);
nand U3120 (N_3120,N_3000,N_3020);
or U3121 (N_3121,N_3078,N_3032);
xnor U3122 (N_3122,N_3041,N_3012);
or U3123 (N_3123,N_3067,N_3056);
nor U3124 (N_3124,N_3054,N_3070);
nand U3125 (N_3125,N_3052,N_3094);
or U3126 (N_3126,N_3003,N_3047);
xnor U3127 (N_3127,N_3036,N_3071);
xnor U3128 (N_3128,N_3030,N_3097);
nor U3129 (N_3129,N_3095,N_3079);
nor U3130 (N_3130,N_3076,N_3096);
or U3131 (N_3131,N_3011,N_3059);
or U3132 (N_3132,N_3057,N_3086);
nand U3133 (N_3133,N_3014,N_3051);
and U3134 (N_3134,N_3090,N_3099);
xor U3135 (N_3135,N_3025,N_3087);
xor U3136 (N_3136,N_3026,N_3093);
and U3137 (N_3137,N_3040,N_3064);
nor U3138 (N_3138,N_3077,N_3018);
nand U3139 (N_3139,N_3010,N_3006);
nor U3140 (N_3140,N_3044,N_3023);
or U3141 (N_3141,N_3073,N_3053);
nand U3142 (N_3142,N_3007,N_3027);
xnor U3143 (N_3143,N_3021,N_3017);
and U3144 (N_3144,N_3019,N_3035);
nor U3145 (N_3145,N_3013,N_3008);
xor U3146 (N_3146,N_3072,N_3022);
nand U3147 (N_3147,N_3031,N_3068);
xor U3148 (N_3148,N_3061,N_3005);
xnor U3149 (N_3149,N_3091,N_3081);
or U3150 (N_3150,N_3047,N_3059);
xnor U3151 (N_3151,N_3098,N_3071);
or U3152 (N_3152,N_3034,N_3026);
nand U3153 (N_3153,N_3023,N_3078);
or U3154 (N_3154,N_3060,N_3024);
nand U3155 (N_3155,N_3050,N_3075);
or U3156 (N_3156,N_3086,N_3085);
and U3157 (N_3157,N_3053,N_3029);
and U3158 (N_3158,N_3019,N_3022);
xor U3159 (N_3159,N_3017,N_3029);
and U3160 (N_3160,N_3039,N_3049);
nand U3161 (N_3161,N_3037,N_3036);
xnor U3162 (N_3162,N_3029,N_3024);
or U3163 (N_3163,N_3068,N_3040);
xor U3164 (N_3164,N_3098,N_3019);
or U3165 (N_3165,N_3010,N_3008);
nand U3166 (N_3166,N_3085,N_3071);
xor U3167 (N_3167,N_3047,N_3032);
and U3168 (N_3168,N_3076,N_3064);
and U3169 (N_3169,N_3049,N_3038);
and U3170 (N_3170,N_3004,N_3000);
xor U3171 (N_3171,N_3093,N_3000);
xor U3172 (N_3172,N_3005,N_3065);
nor U3173 (N_3173,N_3001,N_3042);
nand U3174 (N_3174,N_3004,N_3038);
or U3175 (N_3175,N_3067,N_3078);
and U3176 (N_3176,N_3090,N_3083);
or U3177 (N_3177,N_3001,N_3029);
nand U3178 (N_3178,N_3045,N_3095);
xor U3179 (N_3179,N_3014,N_3037);
nand U3180 (N_3180,N_3037,N_3052);
xor U3181 (N_3181,N_3089,N_3030);
nor U3182 (N_3182,N_3098,N_3016);
nor U3183 (N_3183,N_3089,N_3050);
and U3184 (N_3184,N_3036,N_3089);
nor U3185 (N_3185,N_3053,N_3014);
and U3186 (N_3186,N_3021,N_3099);
xnor U3187 (N_3187,N_3017,N_3074);
xor U3188 (N_3188,N_3029,N_3003);
or U3189 (N_3189,N_3010,N_3045);
nor U3190 (N_3190,N_3052,N_3025);
nand U3191 (N_3191,N_3025,N_3017);
or U3192 (N_3192,N_3034,N_3009);
or U3193 (N_3193,N_3081,N_3049);
nor U3194 (N_3194,N_3032,N_3094);
nor U3195 (N_3195,N_3015,N_3090);
or U3196 (N_3196,N_3067,N_3036);
nand U3197 (N_3197,N_3099,N_3014);
nand U3198 (N_3198,N_3078,N_3072);
nand U3199 (N_3199,N_3033,N_3038);
nor U3200 (N_3200,N_3157,N_3190);
or U3201 (N_3201,N_3120,N_3177);
and U3202 (N_3202,N_3173,N_3174);
or U3203 (N_3203,N_3102,N_3176);
nor U3204 (N_3204,N_3113,N_3140);
nor U3205 (N_3205,N_3128,N_3108);
xnor U3206 (N_3206,N_3165,N_3171);
or U3207 (N_3207,N_3194,N_3111);
or U3208 (N_3208,N_3135,N_3163);
nor U3209 (N_3209,N_3196,N_3147);
and U3210 (N_3210,N_3179,N_3175);
or U3211 (N_3211,N_3151,N_3188);
nor U3212 (N_3212,N_3185,N_3106);
nor U3213 (N_3213,N_3160,N_3118);
xor U3214 (N_3214,N_3178,N_3105);
nand U3215 (N_3215,N_3117,N_3167);
and U3216 (N_3216,N_3191,N_3141);
or U3217 (N_3217,N_3198,N_3158);
nor U3218 (N_3218,N_3187,N_3149);
and U3219 (N_3219,N_3148,N_3101);
and U3220 (N_3220,N_3142,N_3162);
and U3221 (N_3221,N_3136,N_3123);
and U3222 (N_3222,N_3130,N_3166);
nor U3223 (N_3223,N_3183,N_3100);
nand U3224 (N_3224,N_3180,N_3115);
nor U3225 (N_3225,N_3193,N_3181);
nand U3226 (N_3226,N_3137,N_3138);
or U3227 (N_3227,N_3146,N_3164);
and U3228 (N_3228,N_3172,N_3168);
or U3229 (N_3229,N_3131,N_3150);
xor U3230 (N_3230,N_3152,N_3169);
xnor U3231 (N_3231,N_3134,N_3116);
nor U3232 (N_3232,N_3155,N_3195);
nand U3233 (N_3233,N_3119,N_3109);
or U3234 (N_3234,N_3121,N_3125);
and U3235 (N_3235,N_3114,N_3143);
and U3236 (N_3236,N_3126,N_3144);
and U3237 (N_3237,N_3199,N_3139);
xnor U3238 (N_3238,N_3156,N_3154);
and U3239 (N_3239,N_3170,N_3184);
nor U3240 (N_3240,N_3129,N_3133);
nor U3241 (N_3241,N_3127,N_3104);
nor U3242 (N_3242,N_3124,N_3132);
nand U3243 (N_3243,N_3153,N_3145);
xor U3244 (N_3244,N_3103,N_3161);
nor U3245 (N_3245,N_3107,N_3182);
and U3246 (N_3246,N_3192,N_3159);
or U3247 (N_3247,N_3110,N_3197);
or U3248 (N_3248,N_3189,N_3122);
and U3249 (N_3249,N_3112,N_3186);
nor U3250 (N_3250,N_3197,N_3138);
xnor U3251 (N_3251,N_3172,N_3120);
or U3252 (N_3252,N_3151,N_3116);
xor U3253 (N_3253,N_3153,N_3196);
or U3254 (N_3254,N_3151,N_3170);
nor U3255 (N_3255,N_3100,N_3154);
nand U3256 (N_3256,N_3116,N_3148);
nand U3257 (N_3257,N_3191,N_3110);
nor U3258 (N_3258,N_3192,N_3145);
nor U3259 (N_3259,N_3137,N_3114);
xor U3260 (N_3260,N_3121,N_3141);
nand U3261 (N_3261,N_3148,N_3110);
or U3262 (N_3262,N_3197,N_3121);
and U3263 (N_3263,N_3145,N_3144);
nor U3264 (N_3264,N_3158,N_3127);
nor U3265 (N_3265,N_3110,N_3133);
and U3266 (N_3266,N_3134,N_3122);
nor U3267 (N_3267,N_3132,N_3178);
nand U3268 (N_3268,N_3141,N_3175);
and U3269 (N_3269,N_3191,N_3190);
nor U3270 (N_3270,N_3158,N_3191);
or U3271 (N_3271,N_3128,N_3176);
nand U3272 (N_3272,N_3113,N_3158);
nand U3273 (N_3273,N_3187,N_3119);
nand U3274 (N_3274,N_3158,N_3182);
nand U3275 (N_3275,N_3118,N_3164);
nor U3276 (N_3276,N_3128,N_3123);
nor U3277 (N_3277,N_3128,N_3133);
nand U3278 (N_3278,N_3154,N_3134);
nor U3279 (N_3279,N_3147,N_3198);
or U3280 (N_3280,N_3101,N_3105);
nor U3281 (N_3281,N_3183,N_3146);
and U3282 (N_3282,N_3150,N_3151);
nor U3283 (N_3283,N_3157,N_3142);
nand U3284 (N_3284,N_3140,N_3127);
or U3285 (N_3285,N_3109,N_3192);
or U3286 (N_3286,N_3145,N_3193);
nand U3287 (N_3287,N_3164,N_3130);
and U3288 (N_3288,N_3142,N_3117);
nand U3289 (N_3289,N_3171,N_3129);
and U3290 (N_3290,N_3171,N_3158);
nor U3291 (N_3291,N_3163,N_3175);
or U3292 (N_3292,N_3134,N_3135);
nand U3293 (N_3293,N_3181,N_3108);
xnor U3294 (N_3294,N_3177,N_3161);
and U3295 (N_3295,N_3162,N_3105);
or U3296 (N_3296,N_3112,N_3151);
or U3297 (N_3297,N_3101,N_3186);
nand U3298 (N_3298,N_3180,N_3162);
or U3299 (N_3299,N_3135,N_3115);
and U3300 (N_3300,N_3213,N_3249);
and U3301 (N_3301,N_3237,N_3238);
xnor U3302 (N_3302,N_3206,N_3285);
nand U3303 (N_3303,N_3227,N_3258);
and U3304 (N_3304,N_3261,N_3226);
nand U3305 (N_3305,N_3280,N_3231);
and U3306 (N_3306,N_3208,N_3256);
xor U3307 (N_3307,N_3266,N_3251);
xnor U3308 (N_3308,N_3236,N_3215);
nor U3309 (N_3309,N_3201,N_3287);
and U3310 (N_3310,N_3264,N_3297);
nor U3311 (N_3311,N_3254,N_3232);
xnor U3312 (N_3312,N_3291,N_3265);
and U3313 (N_3313,N_3222,N_3205);
nand U3314 (N_3314,N_3293,N_3294);
and U3315 (N_3315,N_3217,N_3246);
nand U3316 (N_3316,N_3239,N_3211);
nand U3317 (N_3317,N_3275,N_3292);
xor U3318 (N_3318,N_3240,N_3225);
and U3319 (N_3319,N_3224,N_3270);
xor U3320 (N_3320,N_3219,N_3267);
nor U3321 (N_3321,N_3210,N_3262);
xnor U3322 (N_3322,N_3273,N_3269);
or U3323 (N_3323,N_3242,N_3260);
and U3324 (N_3324,N_3200,N_3271);
nor U3325 (N_3325,N_3279,N_3255);
xor U3326 (N_3326,N_3290,N_3278);
and U3327 (N_3327,N_3281,N_3207);
nor U3328 (N_3328,N_3268,N_3299);
nor U3329 (N_3329,N_3272,N_3289);
and U3330 (N_3330,N_3230,N_3220);
xnor U3331 (N_3331,N_3202,N_3204);
or U3332 (N_3332,N_3248,N_3223);
nor U3333 (N_3333,N_3245,N_3298);
nand U3334 (N_3334,N_3241,N_3296);
and U3335 (N_3335,N_3234,N_3276);
or U3336 (N_3336,N_3274,N_3253);
nand U3337 (N_3337,N_3284,N_3235);
and U3338 (N_3338,N_3209,N_3286);
and U3339 (N_3339,N_3252,N_3250);
or U3340 (N_3340,N_3212,N_3228);
or U3341 (N_3341,N_3283,N_3244);
and U3342 (N_3342,N_3259,N_3257);
nand U3343 (N_3343,N_3214,N_3247);
xnor U3344 (N_3344,N_3295,N_3282);
xor U3345 (N_3345,N_3277,N_3218);
nor U3346 (N_3346,N_3203,N_3263);
nand U3347 (N_3347,N_3216,N_3229);
nor U3348 (N_3348,N_3288,N_3243);
or U3349 (N_3349,N_3233,N_3221);
nand U3350 (N_3350,N_3243,N_3234);
xor U3351 (N_3351,N_3201,N_3271);
nand U3352 (N_3352,N_3251,N_3250);
nand U3353 (N_3353,N_3219,N_3282);
or U3354 (N_3354,N_3228,N_3288);
nand U3355 (N_3355,N_3233,N_3218);
and U3356 (N_3356,N_3223,N_3221);
or U3357 (N_3357,N_3239,N_3226);
nand U3358 (N_3358,N_3236,N_3254);
or U3359 (N_3359,N_3240,N_3202);
or U3360 (N_3360,N_3231,N_3268);
or U3361 (N_3361,N_3298,N_3226);
xnor U3362 (N_3362,N_3201,N_3258);
and U3363 (N_3363,N_3290,N_3268);
nand U3364 (N_3364,N_3205,N_3249);
or U3365 (N_3365,N_3201,N_3222);
nand U3366 (N_3366,N_3265,N_3237);
xnor U3367 (N_3367,N_3253,N_3239);
nor U3368 (N_3368,N_3222,N_3281);
or U3369 (N_3369,N_3205,N_3261);
xor U3370 (N_3370,N_3240,N_3285);
xor U3371 (N_3371,N_3213,N_3200);
nor U3372 (N_3372,N_3285,N_3297);
nand U3373 (N_3373,N_3243,N_3263);
nand U3374 (N_3374,N_3251,N_3221);
nand U3375 (N_3375,N_3270,N_3292);
nor U3376 (N_3376,N_3262,N_3212);
nor U3377 (N_3377,N_3271,N_3204);
or U3378 (N_3378,N_3217,N_3237);
nor U3379 (N_3379,N_3233,N_3273);
nor U3380 (N_3380,N_3298,N_3240);
and U3381 (N_3381,N_3212,N_3284);
xor U3382 (N_3382,N_3224,N_3298);
nand U3383 (N_3383,N_3283,N_3260);
nor U3384 (N_3384,N_3296,N_3245);
nor U3385 (N_3385,N_3262,N_3284);
nand U3386 (N_3386,N_3202,N_3297);
or U3387 (N_3387,N_3233,N_3268);
and U3388 (N_3388,N_3228,N_3201);
nand U3389 (N_3389,N_3283,N_3275);
nor U3390 (N_3390,N_3275,N_3296);
xor U3391 (N_3391,N_3229,N_3250);
xor U3392 (N_3392,N_3295,N_3229);
and U3393 (N_3393,N_3273,N_3222);
and U3394 (N_3394,N_3259,N_3293);
nand U3395 (N_3395,N_3265,N_3292);
and U3396 (N_3396,N_3232,N_3218);
xnor U3397 (N_3397,N_3259,N_3220);
xor U3398 (N_3398,N_3220,N_3245);
nor U3399 (N_3399,N_3235,N_3287);
nor U3400 (N_3400,N_3396,N_3326);
nand U3401 (N_3401,N_3327,N_3355);
and U3402 (N_3402,N_3351,N_3390);
or U3403 (N_3403,N_3392,N_3307);
and U3404 (N_3404,N_3338,N_3369);
and U3405 (N_3405,N_3331,N_3315);
and U3406 (N_3406,N_3343,N_3388);
xnor U3407 (N_3407,N_3342,N_3382);
nand U3408 (N_3408,N_3375,N_3321);
xnor U3409 (N_3409,N_3362,N_3312);
or U3410 (N_3410,N_3376,N_3350);
and U3411 (N_3411,N_3360,N_3314);
nor U3412 (N_3412,N_3336,N_3325);
xor U3413 (N_3413,N_3364,N_3308);
nor U3414 (N_3414,N_3399,N_3334);
and U3415 (N_3415,N_3311,N_3368);
and U3416 (N_3416,N_3389,N_3394);
nor U3417 (N_3417,N_3391,N_3377);
xor U3418 (N_3418,N_3347,N_3352);
or U3419 (N_3419,N_3383,N_3319);
nand U3420 (N_3420,N_3341,N_3387);
xor U3421 (N_3421,N_3353,N_3324);
xor U3422 (N_3422,N_3304,N_3397);
or U3423 (N_3423,N_3313,N_3358);
and U3424 (N_3424,N_3303,N_3379);
and U3425 (N_3425,N_3398,N_3345);
or U3426 (N_3426,N_3320,N_3395);
and U3427 (N_3427,N_3354,N_3370);
xnor U3428 (N_3428,N_3349,N_3317);
and U3429 (N_3429,N_3359,N_3384);
nand U3430 (N_3430,N_3310,N_3372);
or U3431 (N_3431,N_3339,N_3357);
and U3432 (N_3432,N_3301,N_3309);
or U3433 (N_3433,N_3361,N_3374);
xnor U3434 (N_3434,N_3335,N_3340);
nor U3435 (N_3435,N_3305,N_3316);
or U3436 (N_3436,N_3323,N_3330);
xor U3437 (N_3437,N_3322,N_3328);
xor U3438 (N_3438,N_3329,N_3306);
xor U3439 (N_3439,N_3385,N_3356);
nand U3440 (N_3440,N_3302,N_3344);
nand U3441 (N_3441,N_3371,N_3365);
or U3442 (N_3442,N_3332,N_3393);
and U3443 (N_3443,N_3348,N_3386);
and U3444 (N_3444,N_3367,N_3373);
nor U3445 (N_3445,N_3346,N_3337);
nand U3446 (N_3446,N_3378,N_3380);
xor U3447 (N_3447,N_3363,N_3366);
or U3448 (N_3448,N_3381,N_3333);
nand U3449 (N_3449,N_3318,N_3300);
xor U3450 (N_3450,N_3385,N_3333);
and U3451 (N_3451,N_3312,N_3332);
or U3452 (N_3452,N_3372,N_3311);
and U3453 (N_3453,N_3356,N_3317);
xor U3454 (N_3454,N_3303,N_3320);
and U3455 (N_3455,N_3356,N_3364);
and U3456 (N_3456,N_3382,N_3304);
xnor U3457 (N_3457,N_3326,N_3315);
nand U3458 (N_3458,N_3335,N_3374);
nand U3459 (N_3459,N_3362,N_3302);
nor U3460 (N_3460,N_3364,N_3318);
and U3461 (N_3461,N_3361,N_3347);
and U3462 (N_3462,N_3372,N_3303);
nor U3463 (N_3463,N_3313,N_3351);
and U3464 (N_3464,N_3372,N_3351);
nor U3465 (N_3465,N_3373,N_3362);
xnor U3466 (N_3466,N_3310,N_3301);
xnor U3467 (N_3467,N_3343,N_3359);
or U3468 (N_3468,N_3338,N_3398);
or U3469 (N_3469,N_3300,N_3393);
nor U3470 (N_3470,N_3387,N_3361);
xor U3471 (N_3471,N_3360,N_3333);
nand U3472 (N_3472,N_3349,N_3320);
nand U3473 (N_3473,N_3312,N_3338);
nand U3474 (N_3474,N_3301,N_3328);
and U3475 (N_3475,N_3365,N_3368);
and U3476 (N_3476,N_3368,N_3326);
nor U3477 (N_3477,N_3308,N_3366);
and U3478 (N_3478,N_3356,N_3334);
or U3479 (N_3479,N_3306,N_3308);
or U3480 (N_3480,N_3324,N_3393);
or U3481 (N_3481,N_3376,N_3305);
and U3482 (N_3482,N_3364,N_3387);
or U3483 (N_3483,N_3363,N_3339);
nor U3484 (N_3484,N_3303,N_3312);
nand U3485 (N_3485,N_3385,N_3350);
and U3486 (N_3486,N_3370,N_3337);
and U3487 (N_3487,N_3342,N_3368);
nand U3488 (N_3488,N_3397,N_3300);
xor U3489 (N_3489,N_3347,N_3364);
nand U3490 (N_3490,N_3323,N_3394);
or U3491 (N_3491,N_3328,N_3308);
and U3492 (N_3492,N_3363,N_3364);
xor U3493 (N_3493,N_3357,N_3307);
and U3494 (N_3494,N_3327,N_3302);
xnor U3495 (N_3495,N_3327,N_3373);
or U3496 (N_3496,N_3379,N_3386);
nor U3497 (N_3497,N_3313,N_3317);
nor U3498 (N_3498,N_3304,N_3317);
xor U3499 (N_3499,N_3346,N_3327);
or U3500 (N_3500,N_3441,N_3415);
nand U3501 (N_3501,N_3435,N_3452);
and U3502 (N_3502,N_3455,N_3430);
xnor U3503 (N_3503,N_3480,N_3461);
nor U3504 (N_3504,N_3424,N_3498);
xnor U3505 (N_3505,N_3405,N_3477);
nand U3506 (N_3506,N_3484,N_3466);
or U3507 (N_3507,N_3453,N_3436);
nor U3508 (N_3508,N_3489,N_3412);
nor U3509 (N_3509,N_3403,N_3492);
xnor U3510 (N_3510,N_3422,N_3414);
nand U3511 (N_3511,N_3458,N_3467);
xor U3512 (N_3512,N_3486,N_3409);
and U3513 (N_3513,N_3476,N_3407);
nand U3514 (N_3514,N_3497,N_3428);
nand U3515 (N_3515,N_3410,N_3438);
nor U3516 (N_3516,N_3434,N_3446);
nor U3517 (N_3517,N_3419,N_3493);
or U3518 (N_3518,N_3468,N_3481);
nor U3519 (N_3519,N_3456,N_3423);
nor U3520 (N_3520,N_3447,N_3479);
and U3521 (N_3521,N_3426,N_3443);
or U3522 (N_3522,N_3487,N_3444);
or U3523 (N_3523,N_3491,N_3404);
and U3524 (N_3524,N_3400,N_3442);
nor U3525 (N_3525,N_3402,N_3496);
xnor U3526 (N_3526,N_3420,N_3413);
and U3527 (N_3527,N_3460,N_3482);
nor U3528 (N_3528,N_3457,N_3464);
nor U3529 (N_3529,N_3408,N_3440);
nand U3530 (N_3530,N_3499,N_3472);
or U3531 (N_3531,N_3478,N_3425);
nand U3532 (N_3532,N_3485,N_3473);
xor U3533 (N_3533,N_3469,N_3475);
and U3534 (N_3534,N_3437,N_3421);
xnor U3535 (N_3535,N_3454,N_3406);
or U3536 (N_3536,N_3427,N_3448);
xor U3537 (N_3537,N_3432,N_3445);
and U3538 (N_3538,N_3488,N_3439);
or U3539 (N_3539,N_3494,N_3462);
xnor U3540 (N_3540,N_3433,N_3465);
or U3541 (N_3541,N_3417,N_3463);
or U3542 (N_3542,N_3401,N_3490);
and U3543 (N_3543,N_3431,N_3471);
xnor U3544 (N_3544,N_3459,N_3474);
nor U3545 (N_3545,N_3495,N_3418);
or U3546 (N_3546,N_3429,N_3411);
nand U3547 (N_3547,N_3470,N_3483);
nor U3548 (N_3548,N_3451,N_3416);
or U3549 (N_3549,N_3449,N_3450);
xnor U3550 (N_3550,N_3406,N_3413);
nor U3551 (N_3551,N_3472,N_3465);
and U3552 (N_3552,N_3485,N_3467);
xnor U3553 (N_3553,N_3437,N_3448);
xor U3554 (N_3554,N_3409,N_3428);
and U3555 (N_3555,N_3490,N_3474);
nand U3556 (N_3556,N_3480,N_3468);
and U3557 (N_3557,N_3474,N_3495);
or U3558 (N_3558,N_3443,N_3422);
nand U3559 (N_3559,N_3453,N_3465);
nor U3560 (N_3560,N_3495,N_3411);
xor U3561 (N_3561,N_3469,N_3472);
or U3562 (N_3562,N_3442,N_3407);
nor U3563 (N_3563,N_3411,N_3444);
or U3564 (N_3564,N_3478,N_3448);
or U3565 (N_3565,N_3443,N_3447);
and U3566 (N_3566,N_3430,N_3467);
xor U3567 (N_3567,N_3423,N_3438);
nor U3568 (N_3568,N_3441,N_3432);
and U3569 (N_3569,N_3448,N_3454);
xnor U3570 (N_3570,N_3475,N_3427);
or U3571 (N_3571,N_3428,N_3498);
nand U3572 (N_3572,N_3497,N_3494);
and U3573 (N_3573,N_3418,N_3413);
nand U3574 (N_3574,N_3499,N_3437);
nand U3575 (N_3575,N_3440,N_3422);
or U3576 (N_3576,N_3401,N_3479);
and U3577 (N_3577,N_3472,N_3464);
nor U3578 (N_3578,N_3414,N_3452);
xor U3579 (N_3579,N_3403,N_3443);
xor U3580 (N_3580,N_3462,N_3410);
nor U3581 (N_3581,N_3479,N_3429);
and U3582 (N_3582,N_3462,N_3450);
nand U3583 (N_3583,N_3497,N_3463);
nand U3584 (N_3584,N_3468,N_3400);
or U3585 (N_3585,N_3496,N_3412);
or U3586 (N_3586,N_3450,N_3479);
or U3587 (N_3587,N_3499,N_3415);
and U3588 (N_3588,N_3421,N_3477);
xnor U3589 (N_3589,N_3429,N_3469);
nor U3590 (N_3590,N_3473,N_3468);
xor U3591 (N_3591,N_3424,N_3407);
and U3592 (N_3592,N_3465,N_3456);
nand U3593 (N_3593,N_3457,N_3482);
or U3594 (N_3594,N_3419,N_3428);
nand U3595 (N_3595,N_3497,N_3417);
nand U3596 (N_3596,N_3434,N_3420);
and U3597 (N_3597,N_3443,N_3445);
nor U3598 (N_3598,N_3420,N_3458);
or U3599 (N_3599,N_3444,N_3407);
or U3600 (N_3600,N_3545,N_3598);
nor U3601 (N_3601,N_3546,N_3507);
nor U3602 (N_3602,N_3528,N_3511);
xor U3603 (N_3603,N_3566,N_3573);
and U3604 (N_3604,N_3559,N_3542);
xnor U3605 (N_3605,N_3529,N_3592);
nor U3606 (N_3606,N_3583,N_3538);
nor U3607 (N_3607,N_3543,N_3510);
and U3608 (N_3608,N_3569,N_3568);
nor U3609 (N_3609,N_3547,N_3557);
nor U3610 (N_3610,N_3537,N_3512);
or U3611 (N_3611,N_3595,N_3500);
nor U3612 (N_3612,N_3553,N_3562);
nand U3613 (N_3613,N_3558,N_3524);
nand U3614 (N_3614,N_3530,N_3513);
xnor U3615 (N_3615,N_3575,N_3589);
nand U3616 (N_3616,N_3597,N_3514);
or U3617 (N_3617,N_3580,N_3596);
nor U3618 (N_3618,N_3518,N_3591);
nor U3619 (N_3619,N_3521,N_3556);
xor U3620 (N_3620,N_3523,N_3535);
nand U3621 (N_3621,N_3506,N_3549);
nor U3622 (N_3622,N_3544,N_3577);
nand U3623 (N_3623,N_3515,N_3552);
nor U3624 (N_3624,N_3576,N_3534);
xnor U3625 (N_3625,N_3555,N_3578);
nand U3626 (N_3626,N_3581,N_3531);
xor U3627 (N_3627,N_3590,N_3551);
xor U3628 (N_3628,N_3522,N_3582);
xnor U3629 (N_3629,N_3584,N_3571);
xnor U3630 (N_3630,N_3599,N_3563);
or U3631 (N_3631,N_3548,N_3560);
or U3632 (N_3632,N_3501,N_3564);
nand U3633 (N_3633,N_3503,N_3502);
and U3634 (N_3634,N_3532,N_3554);
nor U3635 (N_3635,N_3588,N_3526);
and U3636 (N_3636,N_3593,N_3505);
nand U3637 (N_3637,N_3572,N_3541);
or U3638 (N_3638,N_3587,N_3536);
nand U3639 (N_3639,N_3540,N_3520);
nand U3640 (N_3640,N_3570,N_3509);
nand U3641 (N_3641,N_3527,N_3508);
or U3642 (N_3642,N_3517,N_3585);
and U3643 (N_3643,N_3525,N_3565);
xnor U3644 (N_3644,N_3594,N_3574);
and U3645 (N_3645,N_3504,N_3567);
or U3646 (N_3646,N_3579,N_3516);
xor U3647 (N_3647,N_3561,N_3533);
nand U3648 (N_3648,N_3586,N_3539);
or U3649 (N_3649,N_3550,N_3519);
xor U3650 (N_3650,N_3580,N_3519);
or U3651 (N_3651,N_3578,N_3540);
nor U3652 (N_3652,N_3553,N_3504);
nor U3653 (N_3653,N_3552,N_3586);
nand U3654 (N_3654,N_3569,N_3549);
nand U3655 (N_3655,N_3551,N_3595);
and U3656 (N_3656,N_3541,N_3565);
and U3657 (N_3657,N_3530,N_3536);
nand U3658 (N_3658,N_3574,N_3592);
nor U3659 (N_3659,N_3556,N_3502);
nor U3660 (N_3660,N_3523,N_3582);
or U3661 (N_3661,N_3559,N_3586);
nand U3662 (N_3662,N_3599,N_3543);
xnor U3663 (N_3663,N_3509,N_3577);
nor U3664 (N_3664,N_3548,N_3568);
and U3665 (N_3665,N_3542,N_3568);
nand U3666 (N_3666,N_3504,N_3559);
nor U3667 (N_3667,N_3517,N_3575);
xor U3668 (N_3668,N_3585,N_3588);
nor U3669 (N_3669,N_3580,N_3529);
xor U3670 (N_3670,N_3524,N_3537);
nand U3671 (N_3671,N_3579,N_3534);
xor U3672 (N_3672,N_3532,N_3590);
and U3673 (N_3673,N_3545,N_3516);
or U3674 (N_3674,N_3522,N_3512);
and U3675 (N_3675,N_3503,N_3555);
or U3676 (N_3676,N_3576,N_3515);
and U3677 (N_3677,N_3539,N_3578);
nor U3678 (N_3678,N_3592,N_3554);
nor U3679 (N_3679,N_3583,N_3503);
nor U3680 (N_3680,N_3510,N_3572);
or U3681 (N_3681,N_3575,N_3569);
or U3682 (N_3682,N_3564,N_3506);
and U3683 (N_3683,N_3560,N_3530);
nor U3684 (N_3684,N_3527,N_3551);
nand U3685 (N_3685,N_3517,N_3580);
and U3686 (N_3686,N_3585,N_3596);
or U3687 (N_3687,N_3567,N_3530);
nand U3688 (N_3688,N_3538,N_3525);
and U3689 (N_3689,N_3553,N_3510);
nand U3690 (N_3690,N_3512,N_3596);
nand U3691 (N_3691,N_3599,N_3520);
nand U3692 (N_3692,N_3546,N_3584);
or U3693 (N_3693,N_3586,N_3538);
or U3694 (N_3694,N_3550,N_3557);
xor U3695 (N_3695,N_3571,N_3560);
or U3696 (N_3696,N_3508,N_3531);
nand U3697 (N_3697,N_3583,N_3586);
or U3698 (N_3698,N_3544,N_3572);
and U3699 (N_3699,N_3593,N_3566);
nor U3700 (N_3700,N_3641,N_3647);
nand U3701 (N_3701,N_3636,N_3642);
or U3702 (N_3702,N_3610,N_3666);
xor U3703 (N_3703,N_3605,N_3688);
nand U3704 (N_3704,N_3644,N_3696);
or U3705 (N_3705,N_3691,N_3604);
nand U3706 (N_3706,N_3640,N_3614);
nor U3707 (N_3707,N_3628,N_3646);
or U3708 (N_3708,N_3654,N_3602);
or U3709 (N_3709,N_3649,N_3618);
and U3710 (N_3710,N_3657,N_3612);
or U3711 (N_3711,N_3625,N_3693);
nand U3712 (N_3712,N_3624,N_3650);
xor U3713 (N_3713,N_3661,N_3664);
nand U3714 (N_3714,N_3615,N_3631);
or U3715 (N_3715,N_3665,N_3684);
and U3716 (N_3716,N_3619,N_3643);
or U3717 (N_3717,N_3689,N_3659);
nand U3718 (N_3718,N_3697,N_3621);
and U3719 (N_3719,N_3626,N_3681);
xnor U3720 (N_3720,N_3634,N_3671);
nor U3721 (N_3721,N_3668,N_3632);
xor U3722 (N_3722,N_3695,N_3682);
and U3723 (N_3723,N_3603,N_3670);
xnor U3724 (N_3724,N_3690,N_3679);
nor U3725 (N_3725,N_3635,N_3660);
xnor U3726 (N_3726,N_3617,N_3645);
xor U3727 (N_3727,N_3629,N_3637);
or U3728 (N_3728,N_3627,N_3620);
nor U3729 (N_3729,N_3663,N_3675);
nand U3730 (N_3730,N_3655,N_3658);
xnor U3731 (N_3731,N_3662,N_3601);
nand U3732 (N_3732,N_3648,N_3672);
xnor U3733 (N_3733,N_3623,N_3611);
xor U3734 (N_3734,N_3609,N_3669);
xor U3735 (N_3735,N_3673,N_3613);
xor U3736 (N_3736,N_3638,N_3699);
nor U3737 (N_3737,N_3694,N_3677);
nand U3738 (N_3738,N_3608,N_3698);
and U3739 (N_3739,N_3687,N_3651);
nand U3740 (N_3740,N_3616,N_3674);
xnor U3741 (N_3741,N_3683,N_3656);
and U3742 (N_3742,N_3678,N_3630);
and U3743 (N_3743,N_3633,N_3686);
nand U3744 (N_3744,N_3676,N_3653);
nor U3745 (N_3745,N_3600,N_3680);
or U3746 (N_3746,N_3692,N_3652);
nand U3747 (N_3747,N_3607,N_3606);
nor U3748 (N_3748,N_3667,N_3622);
nor U3749 (N_3749,N_3685,N_3639);
nand U3750 (N_3750,N_3600,N_3648);
and U3751 (N_3751,N_3661,N_3631);
nand U3752 (N_3752,N_3669,N_3670);
nand U3753 (N_3753,N_3682,N_3665);
nor U3754 (N_3754,N_3624,N_3627);
and U3755 (N_3755,N_3609,N_3684);
and U3756 (N_3756,N_3619,N_3604);
and U3757 (N_3757,N_3620,N_3619);
and U3758 (N_3758,N_3649,N_3662);
nor U3759 (N_3759,N_3616,N_3631);
nor U3760 (N_3760,N_3630,N_3615);
or U3761 (N_3761,N_3669,N_3685);
nor U3762 (N_3762,N_3605,N_3666);
nor U3763 (N_3763,N_3643,N_3682);
and U3764 (N_3764,N_3694,N_3672);
nor U3765 (N_3765,N_3654,N_3628);
and U3766 (N_3766,N_3681,N_3661);
nand U3767 (N_3767,N_3625,N_3659);
xnor U3768 (N_3768,N_3694,N_3625);
or U3769 (N_3769,N_3657,N_3652);
nor U3770 (N_3770,N_3654,N_3604);
nor U3771 (N_3771,N_3631,N_3663);
xor U3772 (N_3772,N_3684,N_3637);
or U3773 (N_3773,N_3615,N_3611);
and U3774 (N_3774,N_3622,N_3651);
xor U3775 (N_3775,N_3621,N_3602);
xor U3776 (N_3776,N_3675,N_3632);
nor U3777 (N_3777,N_3631,N_3695);
or U3778 (N_3778,N_3686,N_3606);
nor U3779 (N_3779,N_3649,N_3677);
and U3780 (N_3780,N_3653,N_3639);
and U3781 (N_3781,N_3678,N_3665);
and U3782 (N_3782,N_3634,N_3653);
or U3783 (N_3783,N_3604,N_3626);
or U3784 (N_3784,N_3681,N_3656);
or U3785 (N_3785,N_3678,N_3623);
nand U3786 (N_3786,N_3631,N_3693);
nor U3787 (N_3787,N_3668,N_3620);
xnor U3788 (N_3788,N_3639,N_3679);
or U3789 (N_3789,N_3632,N_3646);
and U3790 (N_3790,N_3684,N_3691);
nor U3791 (N_3791,N_3660,N_3661);
nand U3792 (N_3792,N_3685,N_3637);
and U3793 (N_3793,N_3629,N_3663);
nand U3794 (N_3794,N_3696,N_3685);
or U3795 (N_3795,N_3673,N_3612);
or U3796 (N_3796,N_3602,N_3639);
xnor U3797 (N_3797,N_3688,N_3656);
and U3798 (N_3798,N_3641,N_3639);
xnor U3799 (N_3799,N_3630,N_3694);
xor U3800 (N_3800,N_3707,N_3733);
xnor U3801 (N_3801,N_3741,N_3795);
xor U3802 (N_3802,N_3713,N_3780);
or U3803 (N_3803,N_3727,N_3710);
nand U3804 (N_3804,N_3749,N_3769);
nor U3805 (N_3805,N_3785,N_3717);
and U3806 (N_3806,N_3737,N_3793);
xnor U3807 (N_3807,N_3789,N_3778);
and U3808 (N_3808,N_3792,N_3768);
nor U3809 (N_3809,N_3734,N_3758);
or U3810 (N_3810,N_3746,N_3744);
nand U3811 (N_3811,N_3714,N_3740);
or U3812 (N_3812,N_3797,N_3757);
or U3813 (N_3813,N_3738,N_3700);
and U3814 (N_3814,N_3777,N_3796);
and U3815 (N_3815,N_3799,N_3763);
xnor U3816 (N_3816,N_3794,N_3776);
and U3817 (N_3817,N_3748,N_3730);
xnor U3818 (N_3818,N_3701,N_3742);
or U3819 (N_3819,N_3703,N_3761);
and U3820 (N_3820,N_3772,N_3722);
xnor U3821 (N_3821,N_3736,N_3715);
nand U3822 (N_3822,N_3729,N_3702);
nor U3823 (N_3823,N_3716,N_3764);
xnor U3824 (N_3824,N_3782,N_3739);
xnor U3825 (N_3825,N_3786,N_3723);
or U3826 (N_3826,N_3732,N_3765);
nor U3827 (N_3827,N_3783,N_3760);
xnor U3828 (N_3828,N_3728,N_3753);
nand U3829 (N_3829,N_3773,N_3718);
xnor U3830 (N_3830,N_3770,N_3712);
nand U3831 (N_3831,N_3775,N_3750);
nor U3832 (N_3832,N_3705,N_3709);
nand U3833 (N_3833,N_3711,N_3754);
nor U3834 (N_3834,N_3731,N_3706);
nor U3835 (N_3835,N_3798,N_3791);
and U3836 (N_3836,N_3762,N_3755);
nor U3837 (N_3837,N_3719,N_3790);
xor U3838 (N_3838,N_3704,N_3788);
nor U3839 (N_3839,N_3751,N_3726);
xnor U3840 (N_3840,N_3759,N_3784);
or U3841 (N_3841,N_3743,N_3779);
xnor U3842 (N_3842,N_3745,N_3767);
and U3843 (N_3843,N_3766,N_3708);
and U3844 (N_3844,N_3774,N_3735);
nor U3845 (N_3845,N_3721,N_3752);
or U3846 (N_3846,N_3724,N_3787);
and U3847 (N_3847,N_3781,N_3747);
and U3848 (N_3848,N_3725,N_3756);
or U3849 (N_3849,N_3771,N_3720);
nor U3850 (N_3850,N_3778,N_3706);
nand U3851 (N_3851,N_3756,N_3763);
nand U3852 (N_3852,N_3767,N_3706);
or U3853 (N_3853,N_3795,N_3765);
nor U3854 (N_3854,N_3728,N_3726);
nor U3855 (N_3855,N_3766,N_3751);
and U3856 (N_3856,N_3755,N_3757);
or U3857 (N_3857,N_3723,N_3765);
nor U3858 (N_3858,N_3786,N_3718);
and U3859 (N_3859,N_3783,N_3719);
nand U3860 (N_3860,N_3734,N_3766);
xor U3861 (N_3861,N_3789,N_3752);
or U3862 (N_3862,N_3712,N_3710);
nand U3863 (N_3863,N_3763,N_3732);
nor U3864 (N_3864,N_3746,N_3713);
nor U3865 (N_3865,N_3753,N_3759);
nor U3866 (N_3866,N_3740,N_3751);
or U3867 (N_3867,N_3732,N_3719);
and U3868 (N_3868,N_3753,N_3730);
and U3869 (N_3869,N_3754,N_3790);
xor U3870 (N_3870,N_3795,N_3756);
and U3871 (N_3871,N_3730,N_3704);
xnor U3872 (N_3872,N_3731,N_3738);
and U3873 (N_3873,N_3730,N_3710);
or U3874 (N_3874,N_3708,N_3740);
xnor U3875 (N_3875,N_3746,N_3755);
nand U3876 (N_3876,N_3760,N_3788);
xnor U3877 (N_3877,N_3702,N_3765);
nor U3878 (N_3878,N_3730,N_3760);
and U3879 (N_3879,N_3746,N_3712);
nand U3880 (N_3880,N_3733,N_3790);
xnor U3881 (N_3881,N_3760,N_3776);
nand U3882 (N_3882,N_3706,N_3740);
or U3883 (N_3883,N_3759,N_3732);
nor U3884 (N_3884,N_3720,N_3733);
nand U3885 (N_3885,N_3773,N_3733);
xnor U3886 (N_3886,N_3721,N_3763);
or U3887 (N_3887,N_3794,N_3700);
xor U3888 (N_3888,N_3710,N_3793);
or U3889 (N_3889,N_3726,N_3779);
nand U3890 (N_3890,N_3774,N_3738);
nand U3891 (N_3891,N_3739,N_3737);
xor U3892 (N_3892,N_3747,N_3767);
nand U3893 (N_3893,N_3780,N_3775);
and U3894 (N_3894,N_3705,N_3751);
xnor U3895 (N_3895,N_3745,N_3731);
xor U3896 (N_3896,N_3728,N_3720);
nor U3897 (N_3897,N_3701,N_3750);
or U3898 (N_3898,N_3756,N_3711);
and U3899 (N_3899,N_3788,N_3774);
nand U3900 (N_3900,N_3882,N_3896);
or U3901 (N_3901,N_3835,N_3866);
xor U3902 (N_3902,N_3815,N_3893);
or U3903 (N_3903,N_3862,N_3821);
xor U3904 (N_3904,N_3875,N_3861);
nand U3905 (N_3905,N_3845,N_3826);
or U3906 (N_3906,N_3880,N_3856);
or U3907 (N_3907,N_3859,N_3819);
or U3908 (N_3908,N_3841,N_3812);
or U3909 (N_3909,N_3889,N_3803);
and U3910 (N_3910,N_3843,N_3873);
nand U3911 (N_3911,N_3886,N_3885);
xor U3912 (N_3912,N_3813,N_3838);
nor U3913 (N_3913,N_3850,N_3876);
nand U3914 (N_3914,N_3809,N_3808);
nand U3915 (N_3915,N_3833,N_3810);
nor U3916 (N_3916,N_3837,N_3872);
nand U3917 (N_3917,N_3820,N_3802);
nand U3918 (N_3918,N_3839,N_3848);
nor U3919 (N_3919,N_3867,N_3818);
nor U3920 (N_3920,N_3864,N_3868);
nor U3921 (N_3921,N_3888,N_3877);
nor U3922 (N_3922,N_3842,N_3807);
and U3923 (N_3923,N_3863,N_3897);
xnor U3924 (N_3924,N_3849,N_3806);
and U3925 (N_3925,N_3816,N_3891);
nor U3926 (N_3926,N_3895,N_3881);
nand U3927 (N_3927,N_3854,N_3894);
nand U3928 (N_3928,N_3829,N_3857);
or U3929 (N_3929,N_3871,N_3814);
or U3930 (N_3930,N_3822,N_3878);
or U3931 (N_3931,N_3805,N_3832);
nor U3932 (N_3932,N_3858,N_3887);
or U3933 (N_3933,N_3827,N_3898);
nand U3934 (N_3934,N_3824,N_3870);
xor U3935 (N_3935,N_3836,N_3847);
and U3936 (N_3936,N_3840,N_3800);
and U3937 (N_3937,N_3801,N_3869);
xnor U3938 (N_3938,N_3865,N_3890);
nand U3939 (N_3939,N_3817,N_3834);
nor U3940 (N_3940,N_3855,N_3899);
nor U3941 (N_3941,N_3828,N_3884);
nand U3942 (N_3942,N_3830,N_3811);
or U3943 (N_3943,N_3879,N_3852);
and U3944 (N_3944,N_3851,N_3892);
nand U3945 (N_3945,N_3831,N_3846);
or U3946 (N_3946,N_3883,N_3825);
nor U3947 (N_3947,N_3853,N_3823);
and U3948 (N_3948,N_3874,N_3804);
or U3949 (N_3949,N_3844,N_3860);
xor U3950 (N_3950,N_3800,N_3823);
or U3951 (N_3951,N_3898,N_3869);
and U3952 (N_3952,N_3859,N_3805);
nand U3953 (N_3953,N_3866,N_3818);
xnor U3954 (N_3954,N_3807,N_3860);
or U3955 (N_3955,N_3848,N_3890);
xnor U3956 (N_3956,N_3818,N_3846);
and U3957 (N_3957,N_3822,N_3870);
xnor U3958 (N_3958,N_3861,N_3883);
nor U3959 (N_3959,N_3866,N_3847);
nor U3960 (N_3960,N_3829,N_3889);
nand U3961 (N_3961,N_3833,N_3865);
or U3962 (N_3962,N_3824,N_3839);
or U3963 (N_3963,N_3851,N_3878);
and U3964 (N_3964,N_3870,N_3835);
xor U3965 (N_3965,N_3845,N_3898);
nand U3966 (N_3966,N_3814,N_3850);
xnor U3967 (N_3967,N_3801,N_3852);
xor U3968 (N_3968,N_3865,N_3878);
and U3969 (N_3969,N_3819,N_3872);
and U3970 (N_3970,N_3811,N_3848);
xnor U3971 (N_3971,N_3803,N_3816);
or U3972 (N_3972,N_3859,N_3841);
and U3973 (N_3973,N_3835,N_3838);
nor U3974 (N_3974,N_3822,N_3833);
xnor U3975 (N_3975,N_3827,N_3899);
or U3976 (N_3976,N_3896,N_3820);
nor U3977 (N_3977,N_3820,N_3876);
xnor U3978 (N_3978,N_3899,N_3856);
and U3979 (N_3979,N_3857,N_3881);
nor U3980 (N_3980,N_3821,N_3838);
nand U3981 (N_3981,N_3808,N_3857);
nand U3982 (N_3982,N_3883,N_3878);
and U3983 (N_3983,N_3852,N_3825);
xnor U3984 (N_3984,N_3898,N_3886);
or U3985 (N_3985,N_3819,N_3852);
nand U3986 (N_3986,N_3811,N_3834);
nand U3987 (N_3987,N_3805,N_3867);
nand U3988 (N_3988,N_3838,N_3884);
nand U3989 (N_3989,N_3884,N_3840);
or U3990 (N_3990,N_3848,N_3819);
xor U3991 (N_3991,N_3890,N_3862);
or U3992 (N_3992,N_3880,N_3887);
nand U3993 (N_3993,N_3894,N_3863);
xnor U3994 (N_3994,N_3831,N_3849);
nand U3995 (N_3995,N_3842,N_3857);
nor U3996 (N_3996,N_3809,N_3853);
and U3997 (N_3997,N_3804,N_3864);
nor U3998 (N_3998,N_3800,N_3882);
nand U3999 (N_3999,N_3832,N_3817);
nor U4000 (N_4000,N_3918,N_3953);
nand U4001 (N_4001,N_3923,N_3908);
nor U4002 (N_4002,N_3983,N_3999);
nor U4003 (N_4003,N_3945,N_3914);
nor U4004 (N_4004,N_3912,N_3966);
and U4005 (N_4005,N_3915,N_3933);
nor U4006 (N_4006,N_3967,N_3954);
nor U4007 (N_4007,N_3971,N_3920);
and U4008 (N_4008,N_3955,N_3994);
or U4009 (N_4009,N_3903,N_3993);
nor U4010 (N_4010,N_3924,N_3905);
and U4011 (N_4011,N_3981,N_3942);
nor U4012 (N_4012,N_3950,N_3921);
nand U4013 (N_4013,N_3960,N_3986);
and U4014 (N_4014,N_3909,N_3929);
nor U4015 (N_4015,N_3944,N_3963);
or U4016 (N_4016,N_3925,N_3926);
or U4017 (N_4017,N_3906,N_3941);
nand U4018 (N_4018,N_3968,N_3943);
or U4019 (N_4019,N_3985,N_3965);
nand U4020 (N_4020,N_3989,N_3947);
nor U4021 (N_4021,N_3922,N_3916);
nor U4022 (N_4022,N_3919,N_3928);
and U4023 (N_4023,N_3984,N_3964);
nor U4024 (N_4024,N_3932,N_3998);
nand U4025 (N_4025,N_3996,N_3902);
or U4026 (N_4026,N_3973,N_3992);
and U4027 (N_4027,N_3982,N_3957);
nor U4028 (N_4028,N_3951,N_3961);
nor U4029 (N_4029,N_3976,N_3904);
or U4030 (N_4030,N_3978,N_3938);
xnor U4031 (N_4031,N_3969,N_3979);
nand U4032 (N_4032,N_3975,N_3949);
nand U4033 (N_4033,N_3956,N_3972);
xor U4034 (N_4034,N_3974,N_3997);
or U4035 (N_4035,N_3901,N_3913);
nand U4036 (N_4036,N_3940,N_3952);
nand U4037 (N_4037,N_3911,N_3930);
nor U4038 (N_4038,N_3980,N_3939);
and U4039 (N_4039,N_3987,N_3995);
nor U4040 (N_4040,N_3990,N_3936);
xnor U4041 (N_4041,N_3931,N_3958);
xnor U4042 (N_4042,N_3907,N_3937);
or U4043 (N_4043,N_3948,N_3977);
or U4044 (N_4044,N_3900,N_3935);
or U4045 (N_4045,N_3988,N_3934);
and U4046 (N_4046,N_3970,N_3991);
nor U4047 (N_4047,N_3910,N_3917);
or U4048 (N_4048,N_3959,N_3962);
nand U4049 (N_4049,N_3927,N_3946);
or U4050 (N_4050,N_3901,N_3959);
nand U4051 (N_4051,N_3927,N_3902);
or U4052 (N_4052,N_3942,N_3999);
or U4053 (N_4053,N_3945,N_3996);
or U4054 (N_4054,N_3931,N_3941);
or U4055 (N_4055,N_3991,N_3998);
or U4056 (N_4056,N_3901,N_3997);
and U4057 (N_4057,N_3939,N_3976);
nand U4058 (N_4058,N_3929,N_3982);
xor U4059 (N_4059,N_3969,N_3964);
nand U4060 (N_4060,N_3910,N_3991);
nor U4061 (N_4061,N_3987,N_3965);
or U4062 (N_4062,N_3929,N_3930);
and U4063 (N_4063,N_3937,N_3913);
nor U4064 (N_4064,N_3918,N_3997);
or U4065 (N_4065,N_3968,N_3948);
or U4066 (N_4066,N_3958,N_3909);
xor U4067 (N_4067,N_3967,N_3976);
or U4068 (N_4068,N_3983,N_3927);
xor U4069 (N_4069,N_3987,N_3980);
nand U4070 (N_4070,N_3983,N_3903);
and U4071 (N_4071,N_3930,N_3980);
and U4072 (N_4072,N_3928,N_3930);
and U4073 (N_4073,N_3951,N_3932);
xnor U4074 (N_4074,N_3937,N_3939);
xor U4075 (N_4075,N_3911,N_3977);
or U4076 (N_4076,N_3970,N_3969);
and U4077 (N_4077,N_3941,N_3943);
or U4078 (N_4078,N_3965,N_3980);
xor U4079 (N_4079,N_3934,N_3994);
xnor U4080 (N_4080,N_3920,N_3949);
or U4081 (N_4081,N_3989,N_3936);
and U4082 (N_4082,N_3949,N_3931);
or U4083 (N_4083,N_3920,N_3988);
and U4084 (N_4084,N_3907,N_3929);
or U4085 (N_4085,N_3958,N_3924);
and U4086 (N_4086,N_3995,N_3915);
and U4087 (N_4087,N_3969,N_3908);
or U4088 (N_4088,N_3944,N_3959);
or U4089 (N_4089,N_3943,N_3922);
nand U4090 (N_4090,N_3969,N_3921);
nand U4091 (N_4091,N_3941,N_3998);
and U4092 (N_4092,N_3986,N_3998);
nor U4093 (N_4093,N_3975,N_3920);
xnor U4094 (N_4094,N_3952,N_3989);
xor U4095 (N_4095,N_3933,N_3942);
xnor U4096 (N_4096,N_3955,N_3986);
nand U4097 (N_4097,N_3903,N_3974);
nand U4098 (N_4098,N_3930,N_3967);
or U4099 (N_4099,N_3987,N_3914);
xor U4100 (N_4100,N_4072,N_4022);
nor U4101 (N_4101,N_4068,N_4060);
and U4102 (N_4102,N_4049,N_4025);
nand U4103 (N_4103,N_4077,N_4043);
nand U4104 (N_4104,N_4075,N_4092);
or U4105 (N_4105,N_4094,N_4061);
or U4106 (N_4106,N_4058,N_4093);
and U4107 (N_4107,N_4003,N_4037);
and U4108 (N_4108,N_4021,N_4083);
and U4109 (N_4109,N_4034,N_4045);
nand U4110 (N_4110,N_4063,N_4005);
xnor U4111 (N_4111,N_4010,N_4029);
or U4112 (N_4112,N_4059,N_4056);
xor U4113 (N_4113,N_4054,N_4076);
or U4114 (N_4114,N_4028,N_4085);
nand U4115 (N_4115,N_4013,N_4008);
or U4116 (N_4116,N_4053,N_4002);
or U4117 (N_4117,N_4070,N_4023);
xor U4118 (N_4118,N_4071,N_4065);
and U4119 (N_4119,N_4016,N_4082);
and U4120 (N_4120,N_4007,N_4015);
and U4121 (N_4121,N_4036,N_4064);
nor U4122 (N_4122,N_4051,N_4011);
or U4123 (N_4123,N_4035,N_4097);
nor U4124 (N_4124,N_4088,N_4026);
or U4125 (N_4125,N_4087,N_4039);
and U4126 (N_4126,N_4030,N_4084);
nand U4127 (N_4127,N_4078,N_4024);
and U4128 (N_4128,N_4032,N_4086);
or U4129 (N_4129,N_4006,N_4090);
nand U4130 (N_4130,N_4091,N_4089);
and U4131 (N_4131,N_4000,N_4027);
xor U4132 (N_4132,N_4062,N_4066);
nor U4133 (N_4133,N_4057,N_4052);
nand U4134 (N_4134,N_4009,N_4038);
nand U4135 (N_4135,N_4042,N_4017);
and U4136 (N_4136,N_4046,N_4096);
xor U4137 (N_4137,N_4014,N_4074);
xnor U4138 (N_4138,N_4099,N_4012);
xnor U4139 (N_4139,N_4004,N_4081);
and U4140 (N_4140,N_4019,N_4020);
xor U4141 (N_4141,N_4098,N_4044);
or U4142 (N_4142,N_4001,N_4080);
nand U4143 (N_4143,N_4050,N_4079);
or U4144 (N_4144,N_4095,N_4055);
xnor U4145 (N_4145,N_4040,N_4048);
nor U4146 (N_4146,N_4069,N_4018);
or U4147 (N_4147,N_4073,N_4067);
xor U4148 (N_4148,N_4041,N_4047);
or U4149 (N_4149,N_4031,N_4033);
and U4150 (N_4150,N_4029,N_4056);
and U4151 (N_4151,N_4060,N_4091);
xor U4152 (N_4152,N_4033,N_4001);
or U4153 (N_4153,N_4005,N_4074);
or U4154 (N_4154,N_4013,N_4042);
xor U4155 (N_4155,N_4017,N_4006);
xnor U4156 (N_4156,N_4057,N_4078);
or U4157 (N_4157,N_4061,N_4028);
or U4158 (N_4158,N_4093,N_4089);
or U4159 (N_4159,N_4075,N_4027);
nor U4160 (N_4160,N_4031,N_4023);
or U4161 (N_4161,N_4012,N_4055);
nand U4162 (N_4162,N_4034,N_4044);
nor U4163 (N_4163,N_4049,N_4044);
or U4164 (N_4164,N_4059,N_4072);
nand U4165 (N_4165,N_4075,N_4046);
nand U4166 (N_4166,N_4086,N_4049);
nand U4167 (N_4167,N_4077,N_4070);
nor U4168 (N_4168,N_4025,N_4062);
nor U4169 (N_4169,N_4027,N_4042);
nand U4170 (N_4170,N_4062,N_4046);
xnor U4171 (N_4171,N_4075,N_4070);
nor U4172 (N_4172,N_4040,N_4023);
and U4173 (N_4173,N_4094,N_4084);
xnor U4174 (N_4174,N_4089,N_4098);
and U4175 (N_4175,N_4056,N_4063);
nand U4176 (N_4176,N_4014,N_4024);
nor U4177 (N_4177,N_4001,N_4004);
xor U4178 (N_4178,N_4010,N_4055);
nor U4179 (N_4179,N_4011,N_4061);
and U4180 (N_4180,N_4029,N_4061);
nor U4181 (N_4181,N_4094,N_4000);
nor U4182 (N_4182,N_4039,N_4081);
and U4183 (N_4183,N_4025,N_4013);
nand U4184 (N_4184,N_4075,N_4072);
nand U4185 (N_4185,N_4054,N_4006);
nor U4186 (N_4186,N_4075,N_4001);
xor U4187 (N_4187,N_4002,N_4039);
nor U4188 (N_4188,N_4061,N_4004);
nor U4189 (N_4189,N_4067,N_4024);
or U4190 (N_4190,N_4078,N_4097);
xnor U4191 (N_4191,N_4044,N_4022);
or U4192 (N_4192,N_4027,N_4039);
or U4193 (N_4193,N_4080,N_4062);
or U4194 (N_4194,N_4039,N_4021);
nor U4195 (N_4195,N_4060,N_4070);
xor U4196 (N_4196,N_4086,N_4047);
or U4197 (N_4197,N_4056,N_4028);
or U4198 (N_4198,N_4084,N_4003);
or U4199 (N_4199,N_4080,N_4055);
nand U4200 (N_4200,N_4105,N_4166);
xor U4201 (N_4201,N_4167,N_4102);
xor U4202 (N_4202,N_4162,N_4160);
xnor U4203 (N_4203,N_4116,N_4173);
nor U4204 (N_4204,N_4178,N_4161);
nand U4205 (N_4205,N_4182,N_4188);
xor U4206 (N_4206,N_4148,N_4126);
and U4207 (N_4207,N_4129,N_4135);
nand U4208 (N_4208,N_4111,N_4122);
or U4209 (N_4209,N_4133,N_4156);
or U4210 (N_4210,N_4170,N_4165);
nor U4211 (N_4211,N_4198,N_4128);
and U4212 (N_4212,N_4120,N_4138);
xor U4213 (N_4213,N_4186,N_4121);
nand U4214 (N_4214,N_4113,N_4172);
nor U4215 (N_4215,N_4143,N_4100);
nand U4216 (N_4216,N_4181,N_4191);
nor U4217 (N_4217,N_4108,N_4192);
nor U4218 (N_4218,N_4180,N_4136);
xnor U4219 (N_4219,N_4104,N_4157);
nor U4220 (N_4220,N_4183,N_4154);
nor U4221 (N_4221,N_4125,N_4123);
xor U4222 (N_4222,N_4149,N_4164);
nor U4223 (N_4223,N_4152,N_4185);
nor U4224 (N_4224,N_4151,N_4114);
nand U4225 (N_4225,N_4144,N_4124);
xor U4226 (N_4226,N_4117,N_4190);
nor U4227 (N_4227,N_4134,N_4140);
or U4228 (N_4228,N_4194,N_4137);
nor U4229 (N_4229,N_4103,N_4175);
nor U4230 (N_4230,N_4101,N_4141);
and U4231 (N_4231,N_4118,N_4150);
or U4232 (N_4232,N_4176,N_4130);
and U4233 (N_4233,N_4158,N_4184);
xnor U4234 (N_4234,N_4127,N_4187);
xnor U4235 (N_4235,N_4168,N_4107);
or U4236 (N_4236,N_4145,N_4112);
and U4237 (N_4237,N_4147,N_4110);
xnor U4238 (N_4238,N_4179,N_4109);
and U4239 (N_4239,N_4115,N_4153);
or U4240 (N_4240,N_4196,N_4177);
and U4241 (N_4241,N_4132,N_4169);
xnor U4242 (N_4242,N_4146,N_4171);
nor U4243 (N_4243,N_4163,N_4174);
and U4244 (N_4244,N_4106,N_4131);
or U4245 (N_4245,N_4195,N_4142);
nand U4246 (N_4246,N_4155,N_4139);
or U4247 (N_4247,N_4193,N_4159);
and U4248 (N_4248,N_4199,N_4189);
nor U4249 (N_4249,N_4119,N_4197);
and U4250 (N_4250,N_4170,N_4159);
and U4251 (N_4251,N_4153,N_4191);
nor U4252 (N_4252,N_4133,N_4106);
xnor U4253 (N_4253,N_4110,N_4172);
nand U4254 (N_4254,N_4186,N_4173);
or U4255 (N_4255,N_4177,N_4149);
or U4256 (N_4256,N_4195,N_4138);
and U4257 (N_4257,N_4189,N_4146);
nand U4258 (N_4258,N_4194,N_4183);
nor U4259 (N_4259,N_4113,N_4131);
nand U4260 (N_4260,N_4135,N_4193);
xnor U4261 (N_4261,N_4179,N_4166);
nor U4262 (N_4262,N_4127,N_4192);
nand U4263 (N_4263,N_4143,N_4151);
and U4264 (N_4264,N_4105,N_4136);
and U4265 (N_4265,N_4150,N_4132);
nor U4266 (N_4266,N_4104,N_4150);
xor U4267 (N_4267,N_4125,N_4178);
nor U4268 (N_4268,N_4112,N_4176);
or U4269 (N_4269,N_4100,N_4102);
nand U4270 (N_4270,N_4151,N_4146);
nor U4271 (N_4271,N_4145,N_4142);
or U4272 (N_4272,N_4116,N_4117);
or U4273 (N_4273,N_4107,N_4173);
nor U4274 (N_4274,N_4159,N_4116);
or U4275 (N_4275,N_4166,N_4132);
nand U4276 (N_4276,N_4137,N_4127);
or U4277 (N_4277,N_4177,N_4184);
and U4278 (N_4278,N_4110,N_4157);
nor U4279 (N_4279,N_4186,N_4192);
and U4280 (N_4280,N_4169,N_4170);
xnor U4281 (N_4281,N_4185,N_4194);
nor U4282 (N_4282,N_4129,N_4150);
nand U4283 (N_4283,N_4141,N_4127);
nor U4284 (N_4284,N_4174,N_4161);
nor U4285 (N_4285,N_4124,N_4199);
nor U4286 (N_4286,N_4118,N_4134);
nor U4287 (N_4287,N_4157,N_4173);
nand U4288 (N_4288,N_4196,N_4132);
or U4289 (N_4289,N_4151,N_4171);
xor U4290 (N_4290,N_4189,N_4156);
or U4291 (N_4291,N_4106,N_4195);
xnor U4292 (N_4292,N_4164,N_4112);
nand U4293 (N_4293,N_4114,N_4129);
and U4294 (N_4294,N_4187,N_4128);
or U4295 (N_4295,N_4112,N_4159);
nand U4296 (N_4296,N_4146,N_4124);
or U4297 (N_4297,N_4155,N_4118);
nor U4298 (N_4298,N_4104,N_4158);
or U4299 (N_4299,N_4101,N_4130);
or U4300 (N_4300,N_4288,N_4277);
xor U4301 (N_4301,N_4233,N_4252);
and U4302 (N_4302,N_4287,N_4265);
xnor U4303 (N_4303,N_4215,N_4225);
nand U4304 (N_4304,N_4208,N_4238);
or U4305 (N_4305,N_4244,N_4294);
xor U4306 (N_4306,N_4247,N_4211);
xor U4307 (N_4307,N_4201,N_4284);
nand U4308 (N_4308,N_4228,N_4281);
nor U4309 (N_4309,N_4236,N_4246);
xnor U4310 (N_4310,N_4261,N_4266);
xnor U4311 (N_4311,N_4235,N_4275);
xnor U4312 (N_4312,N_4285,N_4292);
nor U4313 (N_4313,N_4242,N_4226);
and U4314 (N_4314,N_4276,N_4218);
xnor U4315 (N_4315,N_4249,N_4258);
and U4316 (N_4316,N_4248,N_4210);
or U4317 (N_4317,N_4202,N_4282);
or U4318 (N_4318,N_4262,N_4256);
nor U4319 (N_4319,N_4203,N_4255);
and U4320 (N_4320,N_4296,N_4254);
and U4321 (N_4321,N_4273,N_4293);
nor U4322 (N_4322,N_4278,N_4237);
nand U4323 (N_4323,N_4253,N_4269);
nor U4324 (N_4324,N_4232,N_4243);
nand U4325 (N_4325,N_4299,N_4268);
and U4326 (N_4326,N_4209,N_4272);
xnor U4327 (N_4327,N_4222,N_4224);
and U4328 (N_4328,N_4200,N_4206);
xor U4329 (N_4329,N_4290,N_4229);
and U4330 (N_4330,N_4220,N_4295);
or U4331 (N_4331,N_4217,N_4257);
or U4332 (N_4332,N_4214,N_4298);
xnor U4333 (N_4333,N_4259,N_4283);
and U4334 (N_4334,N_4223,N_4207);
and U4335 (N_4335,N_4274,N_4216);
xor U4336 (N_4336,N_4212,N_4264);
or U4337 (N_4337,N_4250,N_4297);
and U4338 (N_4338,N_4289,N_4270);
nor U4339 (N_4339,N_4219,N_4251);
nand U4340 (N_4340,N_4241,N_4234);
or U4341 (N_4341,N_4240,N_4205);
and U4342 (N_4342,N_4260,N_4227);
or U4343 (N_4343,N_4231,N_4279);
nor U4344 (N_4344,N_4271,N_4245);
and U4345 (N_4345,N_4204,N_4280);
nor U4346 (N_4346,N_4213,N_4267);
xnor U4347 (N_4347,N_4221,N_4291);
nor U4348 (N_4348,N_4230,N_4239);
nand U4349 (N_4349,N_4263,N_4286);
nor U4350 (N_4350,N_4205,N_4221);
xor U4351 (N_4351,N_4220,N_4211);
or U4352 (N_4352,N_4232,N_4276);
or U4353 (N_4353,N_4280,N_4220);
xor U4354 (N_4354,N_4286,N_4289);
nor U4355 (N_4355,N_4256,N_4261);
nand U4356 (N_4356,N_4259,N_4241);
nand U4357 (N_4357,N_4224,N_4254);
or U4358 (N_4358,N_4258,N_4269);
nand U4359 (N_4359,N_4272,N_4236);
nand U4360 (N_4360,N_4291,N_4240);
or U4361 (N_4361,N_4202,N_4278);
nor U4362 (N_4362,N_4296,N_4206);
nor U4363 (N_4363,N_4282,N_4238);
nand U4364 (N_4364,N_4231,N_4286);
xnor U4365 (N_4365,N_4252,N_4204);
xor U4366 (N_4366,N_4233,N_4261);
and U4367 (N_4367,N_4216,N_4277);
or U4368 (N_4368,N_4290,N_4285);
and U4369 (N_4369,N_4239,N_4223);
xnor U4370 (N_4370,N_4251,N_4275);
nor U4371 (N_4371,N_4288,N_4235);
nand U4372 (N_4372,N_4200,N_4262);
nand U4373 (N_4373,N_4277,N_4282);
xnor U4374 (N_4374,N_4292,N_4208);
nand U4375 (N_4375,N_4233,N_4237);
nand U4376 (N_4376,N_4222,N_4258);
xor U4377 (N_4377,N_4280,N_4244);
xnor U4378 (N_4378,N_4299,N_4218);
and U4379 (N_4379,N_4231,N_4215);
nand U4380 (N_4380,N_4282,N_4208);
xor U4381 (N_4381,N_4206,N_4246);
nor U4382 (N_4382,N_4231,N_4213);
or U4383 (N_4383,N_4230,N_4235);
xor U4384 (N_4384,N_4208,N_4245);
xor U4385 (N_4385,N_4232,N_4214);
nand U4386 (N_4386,N_4257,N_4232);
xor U4387 (N_4387,N_4200,N_4238);
and U4388 (N_4388,N_4273,N_4256);
or U4389 (N_4389,N_4249,N_4231);
and U4390 (N_4390,N_4252,N_4247);
or U4391 (N_4391,N_4215,N_4263);
nor U4392 (N_4392,N_4297,N_4227);
nor U4393 (N_4393,N_4279,N_4263);
nor U4394 (N_4394,N_4229,N_4224);
and U4395 (N_4395,N_4226,N_4290);
xnor U4396 (N_4396,N_4270,N_4278);
or U4397 (N_4397,N_4257,N_4262);
nor U4398 (N_4398,N_4228,N_4288);
or U4399 (N_4399,N_4231,N_4219);
nor U4400 (N_4400,N_4343,N_4333);
nor U4401 (N_4401,N_4351,N_4308);
and U4402 (N_4402,N_4356,N_4344);
xor U4403 (N_4403,N_4352,N_4332);
nor U4404 (N_4404,N_4391,N_4335);
xnor U4405 (N_4405,N_4366,N_4377);
and U4406 (N_4406,N_4342,N_4311);
xor U4407 (N_4407,N_4367,N_4358);
and U4408 (N_4408,N_4390,N_4399);
nand U4409 (N_4409,N_4318,N_4387);
or U4410 (N_4410,N_4393,N_4378);
or U4411 (N_4411,N_4386,N_4381);
xor U4412 (N_4412,N_4310,N_4364);
nor U4413 (N_4413,N_4327,N_4306);
xor U4414 (N_4414,N_4350,N_4374);
nor U4415 (N_4415,N_4355,N_4368);
or U4416 (N_4416,N_4330,N_4321);
xnor U4417 (N_4417,N_4360,N_4315);
or U4418 (N_4418,N_4380,N_4357);
and U4419 (N_4419,N_4392,N_4307);
nor U4420 (N_4420,N_4340,N_4371);
nand U4421 (N_4421,N_4336,N_4362);
nand U4422 (N_4422,N_4398,N_4396);
and U4423 (N_4423,N_4313,N_4388);
nand U4424 (N_4424,N_4383,N_4379);
nand U4425 (N_4425,N_4361,N_4394);
and U4426 (N_4426,N_4322,N_4317);
nor U4427 (N_4427,N_4348,N_4305);
nand U4428 (N_4428,N_4373,N_4359);
nand U4429 (N_4429,N_4363,N_4303);
and U4430 (N_4430,N_4353,N_4384);
nor U4431 (N_4431,N_4375,N_4389);
nand U4432 (N_4432,N_4300,N_4304);
and U4433 (N_4433,N_4382,N_4397);
or U4434 (N_4434,N_4334,N_4329);
or U4435 (N_4435,N_4339,N_4370);
and U4436 (N_4436,N_4309,N_4345);
or U4437 (N_4437,N_4346,N_4316);
and U4438 (N_4438,N_4324,N_4320);
and U4439 (N_4439,N_4347,N_4301);
or U4440 (N_4440,N_4372,N_4319);
xor U4441 (N_4441,N_4365,N_4326);
or U4442 (N_4442,N_4328,N_4338);
or U4443 (N_4443,N_4395,N_4376);
nor U4444 (N_4444,N_4312,N_4323);
or U4445 (N_4445,N_4325,N_4385);
nand U4446 (N_4446,N_4337,N_4354);
and U4447 (N_4447,N_4314,N_4349);
xor U4448 (N_4448,N_4331,N_4369);
xor U4449 (N_4449,N_4302,N_4341);
or U4450 (N_4450,N_4365,N_4352);
nor U4451 (N_4451,N_4320,N_4327);
xnor U4452 (N_4452,N_4327,N_4328);
nor U4453 (N_4453,N_4303,N_4315);
or U4454 (N_4454,N_4318,N_4388);
and U4455 (N_4455,N_4389,N_4382);
xnor U4456 (N_4456,N_4399,N_4349);
and U4457 (N_4457,N_4329,N_4388);
and U4458 (N_4458,N_4316,N_4379);
and U4459 (N_4459,N_4334,N_4344);
and U4460 (N_4460,N_4357,N_4373);
and U4461 (N_4461,N_4353,N_4301);
xnor U4462 (N_4462,N_4392,N_4322);
nor U4463 (N_4463,N_4307,N_4354);
xor U4464 (N_4464,N_4326,N_4332);
or U4465 (N_4465,N_4314,N_4326);
nor U4466 (N_4466,N_4343,N_4389);
and U4467 (N_4467,N_4354,N_4355);
nor U4468 (N_4468,N_4300,N_4382);
xnor U4469 (N_4469,N_4342,N_4344);
xor U4470 (N_4470,N_4323,N_4316);
nand U4471 (N_4471,N_4370,N_4324);
and U4472 (N_4472,N_4322,N_4371);
and U4473 (N_4473,N_4327,N_4301);
and U4474 (N_4474,N_4317,N_4301);
and U4475 (N_4475,N_4396,N_4363);
nor U4476 (N_4476,N_4390,N_4301);
or U4477 (N_4477,N_4346,N_4399);
nor U4478 (N_4478,N_4347,N_4361);
or U4479 (N_4479,N_4330,N_4332);
nor U4480 (N_4480,N_4341,N_4309);
xnor U4481 (N_4481,N_4341,N_4330);
or U4482 (N_4482,N_4389,N_4309);
xor U4483 (N_4483,N_4344,N_4321);
nor U4484 (N_4484,N_4340,N_4367);
or U4485 (N_4485,N_4328,N_4352);
or U4486 (N_4486,N_4362,N_4387);
and U4487 (N_4487,N_4340,N_4307);
nor U4488 (N_4488,N_4354,N_4397);
nor U4489 (N_4489,N_4306,N_4304);
and U4490 (N_4490,N_4395,N_4324);
xor U4491 (N_4491,N_4373,N_4321);
and U4492 (N_4492,N_4347,N_4333);
nand U4493 (N_4493,N_4338,N_4346);
xnor U4494 (N_4494,N_4353,N_4316);
nor U4495 (N_4495,N_4393,N_4381);
xor U4496 (N_4496,N_4346,N_4328);
nand U4497 (N_4497,N_4374,N_4330);
xnor U4498 (N_4498,N_4379,N_4378);
or U4499 (N_4499,N_4332,N_4307);
or U4500 (N_4500,N_4457,N_4437);
and U4501 (N_4501,N_4491,N_4439);
xnor U4502 (N_4502,N_4468,N_4464);
nand U4503 (N_4503,N_4443,N_4486);
xor U4504 (N_4504,N_4481,N_4467);
xnor U4505 (N_4505,N_4466,N_4415);
or U4506 (N_4506,N_4490,N_4450);
and U4507 (N_4507,N_4444,N_4478);
or U4508 (N_4508,N_4483,N_4494);
nor U4509 (N_4509,N_4452,N_4487);
nand U4510 (N_4510,N_4488,N_4469);
and U4511 (N_4511,N_4414,N_4477);
nor U4512 (N_4512,N_4470,N_4479);
nor U4513 (N_4513,N_4407,N_4465);
nand U4514 (N_4514,N_4424,N_4423);
nand U4515 (N_4515,N_4411,N_4434);
nor U4516 (N_4516,N_4475,N_4417);
xnor U4517 (N_4517,N_4436,N_4440);
nor U4518 (N_4518,N_4449,N_4410);
nand U4519 (N_4519,N_4427,N_4442);
nor U4520 (N_4520,N_4463,N_4460);
nand U4521 (N_4521,N_4422,N_4435);
or U4522 (N_4522,N_4433,N_4413);
and U4523 (N_4523,N_4462,N_4472);
or U4524 (N_4524,N_4471,N_4459);
xnor U4525 (N_4525,N_4429,N_4425);
nor U4526 (N_4526,N_4493,N_4484);
xnor U4527 (N_4527,N_4441,N_4453);
xnor U4528 (N_4528,N_4418,N_4431);
xnor U4529 (N_4529,N_4445,N_4421);
nor U4530 (N_4530,N_4455,N_4498);
and U4531 (N_4531,N_4448,N_4426);
or U4532 (N_4532,N_4480,N_4495);
or U4533 (N_4533,N_4416,N_4405);
nor U4534 (N_4534,N_4447,N_4430);
nor U4535 (N_4535,N_4499,N_4482);
nor U4536 (N_4536,N_4404,N_4432);
nand U4537 (N_4537,N_4461,N_4428);
nor U4538 (N_4538,N_4446,N_4401);
nand U4539 (N_4539,N_4496,N_4403);
or U4540 (N_4540,N_4419,N_4458);
or U4541 (N_4541,N_4451,N_4408);
or U4542 (N_4542,N_4412,N_4420);
nand U4543 (N_4543,N_4456,N_4400);
xor U4544 (N_4544,N_4438,N_4489);
nand U4545 (N_4545,N_4473,N_4409);
or U4546 (N_4546,N_4454,N_4485);
or U4547 (N_4547,N_4406,N_4492);
xnor U4548 (N_4548,N_4497,N_4474);
nor U4549 (N_4549,N_4476,N_4402);
nor U4550 (N_4550,N_4488,N_4423);
or U4551 (N_4551,N_4466,N_4402);
nand U4552 (N_4552,N_4427,N_4430);
or U4553 (N_4553,N_4426,N_4479);
and U4554 (N_4554,N_4486,N_4490);
nand U4555 (N_4555,N_4420,N_4463);
nand U4556 (N_4556,N_4402,N_4429);
nand U4557 (N_4557,N_4455,N_4444);
xor U4558 (N_4558,N_4402,N_4461);
and U4559 (N_4559,N_4479,N_4415);
or U4560 (N_4560,N_4452,N_4443);
xor U4561 (N_4561,N_4412,N_4492);
xor U4562 (N_4562,N_4494,N_4422);
nor U4563 (N_4563,N_4499,N_4474);
and U4564 (N_4564,N_4472,N_4419);
nand U4565 (N_4565,N_4462,N_4498);
xor U4566 (N_4566,N_4459,N_4449);
nand U4567 (N_4567,N_4430,N_4404);
or U4568 (N_4568,N_4475,N_4486);
or U4569 (N_4569,N_4495,N_4452);
xnor U4570 (N_4570,N_4466,N_4484);
or U4571 (N_4571,N_4439,N_4455);
nand U4572 (N_4572,N_4468,N_4452);
and U4573 (N_4573,N_4447,N_4469);
or U4574 (N_4574,N_4430,N_4436);
or U4575 (N_4575,N_4473,N_4444);
xnor U4576 (N_4576,N_4406,N_4494);
nand U4577 (N_4577,N_4404,N_4409);
or U4578 (N_4578,N_4498,N_4482);
nor U4579 (N_4579,N_4429,N_4496);
nand U4580 (N_4580,N_4433,N_4415);
or U4581 (N_4581,N_4460,N_4455);
nand U4582 (N_4582,N_4440,N_4434);
or U4583 (N_4583,N_4431,N_4466);
or U4584 (N_4584,N_4436,N_4444);
nand U4585 (N_4585,N_4437,N_4466);
nand U4586 (N_4586,N_4455,N_4448);
nor U4587 (N_4587,N_4404,N_4462);
xor U4588 (N_4588,N_4470,N_4473);
nor U4589 (N_4589,N_4439,N_4402);
or U4590 (N_4590,N_4446,N_4474);
or U4591 (N_4591,N_4493,N_4495);
xor U4592 (N_4592,N_4491,N_4432);
nor U4593 (N_4593,N_4445,N_4473);
nand U4594 (N_4594,N_4400,N_4483);
nand U4595 (N_4595,N_4426,N_4457);
nand U4596 (N_4596,N_4410,N_4472);
nor U4597 (N_4597,N_4472,N_4411);
nor U4598 (N_4598,N_4463,N_4467);
nor U4599 (N_4599,N_4459,N_4403);
nand U4600 (N_4600,N_4597,N_4560);
nand U4601 (N_4601,N_4535,N_4562);
or U4602 (N_4602,N_4534,N_4513);
xor U4603 (N_4603,N_4577,N_4553);
and U4604 (N_4604,N_4551,N_4502);
nand U4605 (N_4605,N_4547,N_4532);
nor U4606 (N_4606,N_4517,N_4536);
or U4607 (N_4607,N_4518,N_4509);
nor U4608 (N_4608,N_4521,N_4545);
nor U4609 (N_4609,N_4539,N_4530);
xor U4610 (N_4610,N_4572,N_4564);
and U4611 (N_4611,N_4510,N_4507);
xnor U4612 (N_4612,N_4574,N_4592);
nor U4613 (N_4613,N_4582,N_4581);
nor U4614 (N_4614,N_4526,N_4541);
nand U4615 (N_4615,N_4566,N_4549);
nor U4616 (N_4616,N_4515,N_4593);
and U4617 (N_4617,N_4568,N_4580);
nand U4618 (N_4618,N_4500,N_4542);
and U4619 (N_4619,N_4557,N_4588);
or U4620 (N_4620,N_4563,N_4514);
xor U4621 (N_4621,N_4561,N_4573);
nand U4622 (N_4622,N_4578,N_4525);
nor U4623 (N_4623,N_4567,N_4585);
and U4624 (N_4624,N_4558,N_4505);
nor U4625 (N_4625,N_4544,N_4516);
xnor U4626 (N_4626,N_4520,N_4524);
and U4627 (N_4627,N_4501,N_4599);
nand U4628 (N_4628,N_4537,N_4576);
nand U4629 (N_4629,N_4552,N_4579);
or U4630 (N_4630,N_4506,N_4559);
nor U4631 (N_4631,N_4598,N_4508);
or U4632 (N_4632,N_4519,N_4569);
nand U4633 (N_4633,N_4543,N_4546);
xnor U4634 (N_4634,N_4531,N_4538);
and U4635 (N_4635,N_4586,N_4528);
or U4636 (N_4636,N_4589,N_4504);
nor U4637 (N_4637,N_4596,N_4584);
and U4638 (N_4638,N_4548,N_4522);
and U4639 (N_4639,N_4511,N_4575);
or U4640 (N_4640,N_4503,N_4571);
xor U4641 (N_4641,N_4550,N_4529);
nor U4642 (N_4642,N_4590,N_4587);
nor U4643 (N_4643,N_4512,N_4565);
xor U4644 (N_4644,N_4591,N_4594);
xnor U4645 (N_4645,N_4595,N_4554);
or U4646 (N_4646,N_4540,N_4527);
nand U4647 (N_4647,N_4555,N_4556);
nand U4648 (N_4648,N_4523,N_4533);
xor U4649 (N_4649,N_4570,N_4583);
xor U4650 (N_4650,N_4540,N_4557);
or U4651 (N_4651,N_4500,N_4507);
xnor U4652 (N_4652,N_4539,N_4513);
xor U4653 (N_4653,N_4524,N_4578);
nor U4654 (N_4654,N_4561,N_4519);
nor U4655 (N_4655,N_4532,N_4586);
or U4656 (N_4656,N_4569,N_4552);
or U4657 (N_4657,N_4578,N_4521);
nor U4658 (N_4658,N_4585,N_4514);
nor U4659 (N_4659,N_4583,N_4512);
or U4660 (N_4660,N_4535,N_4501);
nand U4661 (N_4661,N_4575,N_4570);
nor U4662 (N_4662,N_4501,N_4589);
and U4663 (N_4663,N_4533,N_4510);
xnor U4664 (N_4664,N_4531,N_4590);
or U4665 (N_4665,N_4553,N_4568);
or U4666 (N_4666,N_4573,N_4574);
nor U4667 (N_4667,N_4570,N_4597);
or U4668 (N_4668,N_4536,N_4569);
nand U4669 (N_4669,N_4504,N_4500);
nor U4670 (N_4670,N_4567,N_4572);
xor U4671 (N_4671,N_4588,N_4561);
xor U4672 (N_4672,N_4508,N_4533);
or U4673 (N_4673,N_4528,N_4513);
or U4674 (N_4674,N_4512,N_4568);
or U4675 (N_4675,N_4590,N_4565);
and U4676 (N_4676,N_4578,N_4590);
nand U4677 (N_4677,N_4525,N_4536);
and U4678 (N_4678,N_4577,N_4575);
or U4679 (N_4679,N_4506,N_4507);
nand U4680 (N_4680,N_4557,N_4525);
and U4681 (N_4681,N_4593,N_4518);
nor U4682 (N_4682,N_4577,N_4532);
nor U4683 (N_4683,N_4579,N_4507);
nand U4684 (N_4684,N_4510,N_4536);
and U4685 (N_4685,N_4569,N_4540);
or U4686 (N_4686,N_4573,N_4537);
and U4687 (N_4687,N_4533,N_4559);
xor U4688 (N_4688,N_4531,N_4581);
nor U4689 (N_4689,N_4562,N_4588);
and U4690 (N_4690,N_4526,N_4590);
nand U4691 (N_4691,N_4550,N_4544);
or U4692 (N_4692,N_4597,N_4545);
xnor U4693 (N_4693,N_4543,N_4510);
nor U4694 (N_4694,N_4505,N_4521);
nand U4695 (N_4695,N_4505,N_4589);
nand U4696 (N_4696,N_4510,N_4517);
and U4697 (N_4697,N_4584,N_4587);
nor U4698 (N_4698,N_4589,N_4537);
nor U4699 (N_4699,N_4573,N_4591);
or U4700 (N_4700,N_4632,N_4654);
nand U4701 (N_4701,N_4622,N_4604);
nand U4702 (N_4702,N_4665,N_4680);
nor U4703 (N_4703,N_4698,N_4645);
and U4704 (N_4704,N_4615,N_4638);
xnor U4705 (N_4705,N_4686,N_4695);
nor U4706 (N_4706,N_4652,N_4666);
or U4707 (N_4707,N_4625,N_4685);
nor U4708 (N_4708,N_4641,N_4627);
or U4709 (N_4709,N_4609,N_4648);
and U4710 (N_4710,N_4640,N_4650);
nand U4711 (N_4711,N_4603,N_4677);
and U4712 (N_4712,N_4656,N_4643);
xor U4713 (N_4713,N_4671,N_4634);
xor U4714 (N_4714,N_4697,N_4661);
and U4715 (N_4715,N_4644,N_4611);
and U4716 (N_4716,N_4689,N_4600);
nor U4717 (N_4717,N_4631,N_4675);
nor U4718 (N_4718,N_4651,N_4608);
xnor U4719 (N_4719,N_4637,N_4676);
and U4720 (N_4720,N_4610,N_4678);
nand U4721 (N_4721,N_4618,N_4687);
nand U4722 (N_4722,N_4602,N_4669);
nand U4723 (N_4723,N_4621,N_4659);
nor U4724 (N_4724,N_4636,N_4607);
and U4725 (N_4725,N_4664,N_4623);
nand U4726 (N_4726,N_4690,N_4657);
nand U4727 (N_4727,N_4673,N_4624);
nand U4728 (N_4728,N_4681,N_4684);
nor U4729 (N_4729,N_4688,N_4696);
xor U4730 (N_4730,N_4616,N_4653);
nand U4731 (N_4731,N_4612,N_4667);
nand U4732 (N_4732,N_4628,N_4683);
or U4733 (N_4733,N_4699,N_4626);
nand U4734 (N_4734,N_4655,N_4658);
and U4735 (N_4735,N_4692,N_4682);
and U4736 (N_4736,N_4617,N_4601);
nand U4737 (N_4737,N_4642,N_4694);
or U4738 (N_4738,N_4606,N_4663);
or U4739 (N_4739,N_4647,N_4672);
or U4740 (N_4740,N_4649,N_4662);
nand U4741 (N_4741,N_4605,N_4674);
xor U4742 (N_4742,N_4635,N_4691);
nand U4743 (N_4743,N_4633,N_4668);
xnor U4744 (N_4744,N_4693,N_4614);
xor U4745 (N_4745,N_4639,N_4646);
nor U4746 (N_4746,N_4620,N_4629);
or U4747 (N_4747,N_4670,N_4619);
and U4748 (N_4748,N_4630,N_4679);
or U4749 (N_4749,N_4660,N_4613);
or U4750 (N_4750,N_4606,N_4612);
nor U4751 (N_4751,N_4681,N_4626);
or U4752 (N_4752,N_4614,N_4695);
nand U4753 (N_4753,N_4623,N_4629);
xor U4754 (N_4754,N_4606,N_4642);
and U4755 (N_4755,N_4621,N_4606);
nor U4756 (N_4756,N_4692,N_4659);
nand U4757 (N_4757,N_4637,N_4688);
and U4758 (N_4758,N_4628,N_4671);
and U4759 (N_4759,N_4639,N_4653);
and U4760 (N_4760,N_4699,N_4682);
nand U4761 (N_4761,N_4699,N_4603);
or U4762 (N_4762,N_4658,N_4605);
nor U4763 (N_4763,N_4673,N_4653);
or U4764 (N_4764,N_4618,N_4640);
or U4765 (N_4765,N_4678,N_4688);
or U4766 (N_4766,N_4682,N_4647);
xor U4767 (N_4767,N_4682,N_4636);
nand U4768 (N_4768,N_4633,N_4603);
xor U4769 (N_4769,N_4683,N_4641);
nand U4770 (N_4770,N_4662,N_4619);
nand U4771 (N_4771,N_4629,N_4699);
and U4772 (N_4772,N_4665,N_4697);
xnor U4773 (N_4773,N_4696,N_4609);
or U4774 (N_4774,N_4613,N_4625);
nor U4775 (N_4775,N_4651,N_4616);
and U4776 (N_4776,N_4682,N_4657);
nor U4777 (N_4777,N_4662,N_4669);
or U4778 (N_4778,N_4657,N_4626);
and U4779 (N_4779,N_4634,N_4674);
xnor U4780 (N_4780,N_4651,N_4680);
xnor U4781 (N_4781,N_4683,N_4658);
nor U4782 (N_4782,N_4628,N_4602);
nand U4783 (N_4783,N_4643,N_4684);
xnor U4784 (N_4784,N_4681,N_4658);
or U4785 (N_4785,N_4639,N_4674);
and U4786 (N_4786,N_4616,N_4637);
nor U4787 (N_4787,N_4687,N_4633);
nand U4788 (N_4788,N_4630,N_4671);
nor U4789 (N_4789,N_4609,N_4695);
and U4790 (N_4790,N_4631,N_4656);
and U4791 (N_4791,N_4670,N_4666);
xnor U4792 (N_4792,N_4641,N_4666);
nand U4793 (N_4793,N_4678,N_4605);
nor U4794 (N_4794,N_4681,N_4662);
or U4795 (N_4795,N_4685,N_4644);
xnor U4796 (N_4796,N_4674,N_4632);
nand U4797 (N_4797,N_4697,N_4655);
and U4798 (N_4798,N_4697,N_4614);
nor U4799 (N_4799,N_4683,N_4649);
nand U4800 (N_4800,N_4760,N_4797);
and U4801 (N_4801,N_4742,N_4749);
nor U4802 (N_4802,N_4743,N_4788);
nand U4803 (N_4803,N_4753,N_4783);
nor U4804 (N_4804,N_4734,N_4771);
nor U4805 (N_4805,N_4764,N_4772);
xor U4806 (N_4806,N_4735,N_4766);
xnor U4807 (N_4807,N_4785,N_4718);
xor U4808 (N_4808,N_4730,N_4754);
and U4809 (N_4809,N_4723,N_4793);
nand U4810 (N_4810,N_4712,N_4711);
xnor U4811 (N_4811,N_4729,N_4722);
nor U4812 (N_4812,N_4781,N_4702);
and U4813 (N_4813,N_4791,N_4717);
nor U4814 (N_4814,N_4778,N_4709);
nand U4815 (N_4815,N_4782,N_4755);
nand U4816 (N_4816,N_4768,N_4794);
nor U4817 (N_4817,N_4728,N_4724);
nor U4818 (N_4818,N_4741,N_4798);
nand U4819 (N_4819,N_4715,N_4732);
xor U4820 (N_4820,N_4727,N_4770);
and U4821 (N_4821,N_4745,N_4796);
nand U4822 (N_4822,N_4719,N_4787);
or U4823 (N_4823,N_4747,N_4744);
and U4824 (N_4824,N_4759,N_4750);
nand U4825 (N_4825,N_4773,N_4765);
and U4826 (N_4826,N_4762,N_4733);
or U4827 (N_4827,N_4795,N_4777);
or U4828 (N_4828,N_4720,N_4799);
xor U4829 (N_4829,N_4751,N_4700);
nor U4830 (N_4830,N_4701,N_4761);
nand U4831 (N_4831,N_4779,N_4721);
or U4832 (N_4832,N_4763,N_4737);
nor U4833 (N_4833,N_4708,N_4710);
xor U4834 (N_4834,N_4767,N_4706);
xnor U4835 (N_4835,N_4774,N_4769);
nor U4836 (N_4836,N_4736,N_4705);
nor U4837 (N_4837,N_4775,N_4756);
nand U4838 (N_4838,N_4740,N_4784);
or U4839 (N_4839,N_4725,N_4758);
nor U4840 (N_4840,N_4739,N_4789);
nor U4841 (N_4841,N_4790,N_4748);
or U4842 (N_4842,N_4776,N_4780);
xnor U4843 (N_4843,N_4713,N_4786);
nand U4844 (N_4844,N_4752,N_4738);
and U4845 (N_4845,N_4703,N_4757);
nand U4846 (N_4846,N_4716,N_4714);
xnor U4847 (N_4847,N_4746,N_4726);
or U4848 (N_4848,N_4792,N_4707);
or U4849 (N_4849,N_4704,N_4731);
and U4850 (N_4850,N_4703,N_4750);
nand U4851 (N_4851,N_4745,N_4789);
nand U4852 (N_4852,N_4740,N_4767);
nand U4853 (N_4853,N_4770,N_4776);
nand U4854 (N_4854,N_4721,N_4702);
and U4855 (N_4855,N_4796,N_4765);
xor U4856 (N_4856,N_4751,N_4765);
and U4857 (N_4857,N_4768,N_4775);
nor U4858 (N_4858,N_4713,N_4711);
nor U4859 (N_4859,N_4761,N_4792);
and U4860 (N_4860,N_4799,N_4736);
or U4861 (N_4861,N_4789,N_4729);
or U4862 (N_4862,N_4758,N_4784);
xnor U4863 (N_4863,N_4706,N_4775);
or U4864 (N_4864,N_4756,N_4786);
or U4865 (N_4865,N_4797,N_4736);
nand U4866 (N_4866,N_4722,N_4736);
and U4867 (N_4867,N_4772,N_4721);
nor U4868 (N_4868,N_4741,N_4711);
and U4869 (N_4869,N_4707,N_4757);
and U4870 (N_4870,N_4715,N_4734);
or U4871 (N_4871,N_4717,N_4790);
nand U4872 (N_4872,N_4786,N_4782);
nand U4873 (N_4873,N_4702,N_4754);
xnor U4874 (N_4874,N_4738,N_4773);
and U4875 (N_4875,N_4734,N_4764);
nor U4876 (N_4876,N_4714,N_4726);
and U4877 (N_4877,N_4796,N_4748);
xor U4878 (N_4878,N_4796,N_4702);
nor U4879 (N_4879,N_4752,N_4748);
xor U4880 (N_4880,N_4771,N_4797);
or U4881 (N_4881,N_4723,N_4719);
nor U4882 (N_4882,N_4708,N_4795);
and U4883 (N_4883,N_4752,N_4774);
or U4884 (N_4884,N_4710,N_4792);
xor U4885 (N_4885,N_4769,N_4781);
nand U4886 (N_4886,N_4793,N_4722);
nand U4887 (N_4887,N_4747,N_4771);
nor U4888 (N_4888,N_4751,N_4740);
xor U4889 (N_4889,N_4721,N_4791);
nor U4890 (N_4890,N_4702,N_4711);
nor U4891 (N_4891,N_4722,N_4796);
or U4892 (N_4892,N_4761,N_4785);
and U4893 (N_4893,N_4713,N_4710);
nor U4894 (N_4894,N_4792,N_4725);
nor U4895 (N_4895,N_4721,N_4747);
and U4896 (N_4896,N_4764,N_4703);
or U4897 (N_4897,N_4730,N_4776);
nand U4898 (N_4898,N_4743,N_4725);
xnor U4899 (N_4899,N_4707,N_4763);
nand U4900 (N_4900,N_4834,N_4892);
xor U4901 (N_4901,N_4870,N_4809);
and U4902 (N_4902,N_4841,N_4865);
nand U4903 (N_4903,N_4803,N_4884);
and U4904 (N_4904,N_4857,N_4853);
nor U4905 (N_4905,N_4813,N_4807);
xor U4906 (N_4906,N_4808,N_4833);
nor U4907 (N_4907,N_4872,N_4888);
and U4908 (N_4908,N_4844,N_4826);
and U4909 (N_4909,N_4804,N_4859);
xnor U4910 (N_4910,N_4867,N_4835);
nor U4911 (N_4911,N_4810,N_4825);
nor U4912 (N_4912,N_4818,N_4881);
xor U4913 (N_4913,N_4893,N_4838);
nor U4914 (N_4914,N_4815,N_4828);
nand U4915 (N_4915,N_4819,N_4851);
and U4916 (N_4916,N_4877,N_4847);
nand U4917 (N_4917,N_4891,N_4899);
nand U4918 (N_4918,N_4822,N_4855);
nand U4919 (N_4919,N_4862,N_4875);
nand U4920 (N_4920,N_4842,N_4852);
nand U4921 (N_4921,N_4801,N_4845);
nand U4922 (N_4922,N_4800,N_4883);
nor U4923 (N_4923,N_4821,N_4868);
nor U4924 (N_4924,N_4864,N_4816);
and U4925 (N_4925,N_4806,N_4837);
and U4926 (N_4926,N_4839,N_4887);
and U4927 (N_4927,N_4858,N_4850);
and U4928 (N_4928,N_4805,N_4848);
and U4929 (N_4929,N_4878,N_4811);
or U4930 (N_4930,N_4880,N_4879);
xor U4931 (N_4931,N_4843,N_4886);
nand U4932 (N_4932,N_4894,N_4863);
nand U4933 (N_4933,N_4824,N_4876);
xnor U4934 (N_4934,N_4895,N_4871);
nor U4935 (N_4935,N_4885,N_4854);
nor U4936 (N_4936,N_4874,N_4889);
xnor U4937 (N_4937,N_4861,N_4897);
nand U4938 (N_4938,N_4814,N_4823);
or U4939 (N_4939,N_4830,N_4869);
or U4940 (N_4940,N_4827,N_4890);
nor U4941 (N_4941,N_4831,N_4856);
and U4942 (N_4942,N_4817,N_4873);
or U4943 (N_4943,N_4896,N_4866);
nand U4944 (N_4944,N_4829,N_4898);
nor U4945 (N_4945,N_4836,N_4840);
or U4946 (N_4946,N_4882,N_4812);
or U4947 (N_4947,N_4832,N_4802);
and U4948 (N_4948,N_4860,N_4846);
xnor U4949 (N_4949,N_4820,N_4849);
or U4950 (N_4950,N_4829,N_4849);
xnor U4951 (N_4951,N_4826,N_4836);
or U4952 (N_4952,N_4855,N_4870);
and U4953 (N_4953,N_4837,N_4894);
or U4954 (N_4954,N_4893,N_4862);
nor U4955 (N_4955,N_4856,N_4819);
xor U4956 (N_4956,N_4827,N_4849);
nor U4957 (N_4957,N_4824,N_4831);
and U4958 (N_4958,N_4830,N_4871);
or U4959 (N_4959,N_4847,N_4817);
xnor U4960 (N_4960,N_4822,N_4863);
or U4961 (N_4961,N_4861,N_4841);
nand U4962 (N_4962,N_4850,N_4804);
xnor U4963 (N_4963,N_4878,N_4884);
and U4964 (N_4964,N_4877,N_4859);
nor U4965 (N_4965,N_4857,N_4811);
nand U4966 (N_4966,N_4898,N_4828);
xnor U4967 (N_4967,N_4866,N_4833);
nand U4968 (N_4968,N_4886,N_4890);
xnor U4969 (N_4969,N_4870,N_4858);
xor U4970 (N_4970,N_4807,N_4873);
or U4971 (N_4971,N_4811,N_4894);
or U4972 (N_4972,N_4866,N_4843);
and U4973 (N_4973,N_4860,N_4897);
nand U4974 (N_4974,N_4850,N_4843);
xnor U4975 (N_4975,N_4801,N_4853);
nand U4976 (N_4976,N_4883,N_4835);
and U4977 (N_4977,N_4819,N_4869);
nand U4978 (N_4978,N_4863,N_4889);
xor U4979 (N_4979,N_4882,N_4814);
or U4980 (N_4980,N_4864,N_4822);
xor U4981 (N_4981,N_4865,N_4878);
nand U4982 (N_4982,N_4829,N_4806);
nand U4983 (N_4983,N_4843,N_4807);
and U4984 (N_4984,N_4808,N_4840);
nand U4985 (N_4985,N_4885,N_4883);
and U4986 (N_4986,N_4816,N_4833);
or U4987 (N_4987,N_4867,N_4825);
xor U4988 (N_4988,N_4808,N_4823);
and U4989 (N_4989,N_4828,N_4800);
nor U4990 (N_4990,N_4857,N_4833);
and U4991 (N_4991,N_4804,N_4825);
nand U4992 (N_4992,N_4870,N_4816);
or U4993 (N_4993,N_4878,N_4857);
nand U4994 (N_4994,N_4872,N_4804);
xnor U4995 (N_4995,N_4877,N_4899);
or U4996 (N_4996,N_4843,N_4884);
and U4997 (N_4997,N_4846,N_4826);
nor U4998 (N_4998,N_4852,N_4807);
xor U4999 (N_4999,N_4875,N_4828);
nand UO_0 (O_0,N_4986,N_4906);
nor UO_1 (O_1,N_4917,N_4946);
nand UO_2 (O_2,N_4964,N_4947);
nand UO_3 (O_3,N_4968,N_4904);
or UO_4 (O_4,N_4919,N_4921);
and UO_5 (O_5,N_4950,N_4927);
nand UO_6 (O_6,N_4928,N_4996);
or UO_7 (O_7,N_4990,N_4952);
xor UO_8 (O_8,N_4912,N_4987);
nor UO_9 (O_9,N_4918,N_4959);
nand UO_10 (O_10,N_4966,N_4960);
nor UO_11 (O_11,N_4981,N_4970);
or UO_12 (O_12,N_4967,N_4943);
nand UO_13 (O_13,N_4998,N_4988);
xor UO_14 (O_14,N_4931,N_4938);
xnor UO_15 (O_15,N_4973,N_4936);
nand UO_16 (O_16,N_4991,N_4969);
nor UO_17 (O_17,N_4903,N_4940);
and UO_18 (O_18,N_4908,N_4965);
and UO_19 (O_19,N_4954,N_4978);
or UO_20 (O_20,N_4929,N_4980);
nand UO_21 (O_21,N_4920,N_4900);
nor UO_22 (O_22,N_4974,N_4923);
and UO_23 (O_23,N_4922,N_4924);
and UO_24 (O_24,N_4957,N_4956);
and UO_25 (O_25,N_4901,N_4933);
xor UO_26 (O_26,N_4913,N_4911);
and UO_27 (O_27,N_4984,N_4909);
nor UO_28 (O_28,N_4902,N_4910);
or UO_29 (O_29,N_4945,N_4948);
nand UO_30 (O_30,N_4993,N_4992);
and UO_31 (O_31,N_4999,N_4949);
nand UO_32 (O_32,N_4982,N_4997);
nand UO_33 (O_33,N_4995,N_4905);
and UO_34 (O_34,N_4983,N_4951);
or UO_35 (O_35,N_4975,N_4937);
and UO_36 (O_36,N_4979,N_4915);
nand UO_37 (O_37,N_4914,N_4916);
xnor UO_38 (O_38,N_4926,N_4962);
and UO_39 (O_39,N_4932,N_4976);
nor UO_40 (O_40,N_4944,N_4958);
or UO_41 (O_41,N_4942,N_4989);
nor UO_42 (O_42,N_4972,N_4925);
or UO_43 (O_43,N_4934,N_4953);
nor UO_44 (O_44,N_4930,N_4963);
xnor UO_45 (O_45,N_4955,N_4941);
or UO_46 (O_46,N_4977,N_4971);
xnor UO_47 (O_47,N_4994,N_4935);
or UO_48 (O_48,N_4961,N_4907);
and UO_49 (O_49,N_4985,N_4939);
nor UO_50 (O_50,N_4995,N_4919);
xnor UO_51 (O_51,N_4928,N_4978);
and UO_52 (O_52,N_4942,N_4995);
nand UO_53 (O_53,N_4920,N_4948);
xor UO_54 (O_54,N_4988,N_4921);
or UO_55 (O_55,N_4938,N_4959);
and UO_56 (O_56,N_4954,N_4988);
and UO_57 (O_57,N_4975,N_4945);
or UO_58 (O_58,N_4926,N_4999);
or UO_59 (O_59,N_4922,N_4906);
nor UO_60 (O_60,N_4912,N_4911);
nor UO_61 (O_61,N_4956,N_4960);
nor UO_62 (O_62,N_4980,N_4924);
nand UO_63 (O_63,N_4945,N_4936);
and UO_64 (O_64,N_4902,N_4946);
and UO_65 (O_65,N_4909,N_4963);
xnor UO_66 (O_66,N_4947,N_4924);
nand UO_67 (O_67,N_4972,N_4953);
and UO_68 (O_68,N_4901,N_4920);
xnor UO_69 (O_69,N_4932,N_4916);
nand UO_70 (O_70,N_4988,N_4967);
nor UO_71 (O_71,N_4964,N_4910);
xor UO_72 (O_72,N_4981,N_4968);
and UO_73 (O_73,N_4989,N_4931);
xnor UO_74 (O_74,N_4939,N_4981);
and UO_75 (O_75,N_4954,N_4906);
and UO_76 (O_76,N_4906,N_4983);
nor UO_77 (O_77,N_4927,N_4991);
nor UO_78 (O_78,N_4960,N_4953);
nor UO_79 (O_79,N_4962,N_4906);
xnor UO_80 (O_80,N_4921,N_4952);
xnor UO_81 (O_81,N_4971,N_4965);
nand UO_82 (O_82,N_4994,N_4997);
or UO_83 (O_83,N_4955,N_4958);
xor UO_84 (O_84,N_4908,N_4901);
xnor UO_85 (O_85,N_4958,N_4900);
xor UO_86 (O_86,N_4917,N_4988);
nor UO_87 (O_87,N_4983,N_4989);
and UO_88 (O_88,N_4935,N_4974);
nand UO_89 (O_89,N_4987,N_4962);
nor UO_90 (O_90,N_4997,N_4951);
or UO_91 (O_91,N_4902,N_4934);
or UO_92 (O_92,N_4934,N_4928);
nand UO_93 (O_93,N_4995,N_4959);
or UO_94 (O_94,N_4966,N_4927);
or UO_95 (O_95,N_4930,N_4912);
nor UO_96 (O_96,N_4923,N_4947);
nor UO_97 (O_97,N_4975,N_4962);
nor UO_98 (O_98,N_4914,N_4932);
or UO_99 (O_99,N_4961,N_4981);
nand UO_100 (O_100,N_4914,N_4958);
nor UO_101 (O_101,N_4938,N_4905);
nor UO_102 (O_102,N_4938,N_4974);
xnor UO_103 (O_103,N_4926,N_4910);
or UO_104 (O_104,N_4959,N_4976);
xor UO_105 (O_105,N_4961,N_4920);
or UO_106 (O_106,N_4949,N_4938);
and UO_107 (O_107,N_4938,N_4978);
and UO_108 (O_108,N_4968,N_4944);
nand UO_109 (O_109,N_4963,N_4905);
xnor UO_110 (O_110,N_4962,N_4999);
and UO_111 (O_111,N_4922,N_4978);
or UO_112 (O_112,N_4912,N_4998);
or UO_113 (O_113,N_4922,N_4975);
or UO_114 (O_114,N_4973,N_4946);
nand UO_115 (O_115,N_4983,N_4939);
or UO_116 (O_116,N_4900,N_4912);
nand UO_117 (O_117,N_4971,N_4958);
nor UO_118 (O_118,N_4985,N_4981);
and UO_119 (O_119,N_4946,N_4976);
or UO_120 (O_120,N_4930,N_4984);
nand UO_121 (O_121,N_4955,N_4908);
xor UO_122 (O_122,N_4999,N_4934);
nor UO_123 (O_123,N_4993,N_4952);
xnor UO_124 (O_124,N_4988,N_4973);
nor UO_125 (O_125,N_4926,N_4908);
nor UO_126 (O_126,N_4978,N_4951);
nand UO_127 (O_127,N_4995,N_4963);
nor UO_128 (O_128,N_4990,N_4971);
nor UO_129 (O_129,N_4904,N_4924);
and UO_130 (O_130,N_4904,N_4942);
and UO_131 (O_131,N_4962,N_4941);
nand UO_132 (O_132,N_4958,N_4964);
or UO_133 (O_133,N_4992,N_4949);
nand UO_134 (O_134,N_4929,N_4958);
and UO_135 (O_135,N_4904,N_4962);
nand UO_136 (O_136,N_4970,N_4960);
nor UO_137 (O_137,N_4927,N_4931);
and UO_138 (O_138,N_4965,N_4921);
nor UO_139 (O_139,N_4936,N_4978);
nor UO_140 (O_140,N_4987,N_4963);
nand UO_141 (O_141,N_4918,N_4901);
xor UO_142 (O_142,N_4921,N_4986);
and UO_143 (O_143,N_4995,N_4962);
or UO_144 (O_144,N_4998,N_4920);
and UO_145 (O_145,N_4922,N_4919);
nor UO_146 (O_146,N_4957,N_4993);
or UO_147 (O_147,N_4975,N_4920);
nor UO_148 (O_148,N_4926,N_4951);
or UO_149 (O_149,N_4934,N_4903);
and UO_150 (O_150,N_4987,N_4990);
nand UO_151 (O_151,N_4948,N_4982);
and UO_152 (O_152,N_4936,N_4982);
nand UO_153 (O_153,N_4973,N_4938);
or UO_154 (O_154,N_4958,N_4923);
and UO_155 (O_155,N_4914,N_4923);
and UO_156 (O_156,N_4928,N_4972);
xnor UO_157 (O_157,N_4943,N_4901);
xor UO_158 (O_158,N_4945,N_4957);
or UO_159 (O_159,N_4928,N_4968);
and UO_160 (O_160,N_4933,N_4957);
nor UO_161 (O_161,N_4997,N_4946);
or UO_162 (O_162,N_4966,N_4950);
or UO_163 (O_163,N_4903,N_4955);
or UO_164 (O_164,N_4996,N_4995);
or UO_165 (O_165,N_4991,N_4923);
nor UO_166 (O_166,N_4982,N_4905);
xor UO_167 (O_167,N_4920,N_4947);
or UO_168 (O_168,N_4912,N_4924);
nor UO_169 (O_169,N_4995,N_4900);
nor UO_170 (O_170,N_4990,N_4928);
xor UO_171 (O_171,N_4922,N_4910);
nor UO_172 (O_172,N_4952,N_4908);
nor UO_173 (O_173,N_4996,N_4905);
nor UO_174 (O_174,N_4905,N_4927);
nand UO_175 (O_175,N_4916,N_4960);
or UO_176 (O_176,N_4921,N_4951);
nor UO_177 (O_177,N_4913,N_4996);
nand UO_178 (O_178,N_4917,N_4977);
nor UO_179 (O_179,N_4930,N_4970);
and UO_180 (O_180,N_4941,N_4934);
xor UO_181 (O_181,N_4971,N_4981);
xnor UO_182 (O_182,N_4908,N_4960);
or UO_183 (O_183,N_4904,N_4995);
and UO_184 (O_184,N_4902,N_4987);
xnor UO_185 (O_185,N_4997,N_4947);
xnor UO_186 (O_186,N_4912,N_4965);
nor UO_187 (O_187,N_4949,N_4927);
nor UO_188 (O_188,N_4962,N_4940);
or UO_189 (O_189,N_4941,N_4968);
nand UO_190 (O_190,N_4977,N_4900);
and UO_191 (O_191,N_4920,N_4911);
nand UO_192 (O_192,N_4945,N_4953);
or UO_193 (O_193,N_4950,N_4911);
xnor UO_194 (O_194,N_4970,N_4992);
and UO_195 (O_195,N_4917,N_4994);
nand UO_196 (O_196,N_4913,N_4904);
and UO_197 (O_197,N_4983,N_4949);
and UO_198 (O_198,N_4937,N_4995);
xnor UO_199 (O_199,N_4902,N_4952);
and UO_200 (O_200,N_4901,N_4989);
nor UO_201 (O_201,N_4902,N_4992);
nand UO_202 (O_202,N_4959,N_4999);
and UO_203 (O_203,N_4957,N_4969);
nand UO_204 (O_204,N_4925,N_4983);
nor UO_205 (O_205,N_4910,N_4906);
nor UO_206 (O_206,N_4967,N_4958);
or UO_207 (O_207,N_4907,N_4967);
nand UO_208 (O_208,N_4998,N_4936);
or UO_209 (O_209,N_4935,N_4919);
or UO_210 (O_210,N_4969,N_4906);
and UO_211 (O_211,N_4956,N_4918);
nor UO_212 (O_212,N_4948,N_4987);
nand UO_213 (O_213,N_4951,N_4966);
and UO_214 (O_214,N_4936,N_4990);
and UO_215 (O_215,N_4931,N_4984);
nor UO_216 (O_216,N_4909,N_4919);
or UO_217 (O_217,N_4987,N_4991);
xnor UO_218 (O_218,N_4985,N_4957);
nor UO_219 (O_219,N_4942,N_4940);
and UO_220 (O_220,N_4975,N_4980);
nand UO_221 (O_221,N_4933,N_4909);
nor UO_222 (O_222,N_4987,N_4969);
xor UO_223 (O_223,N_4961,N_4985);
nand UO_224 (O_224,N_4921,N_4944);
nor UO_225 (O_225,N_4973,N_4998);
nor UO_226 (O_226,N_4997,N_4955);
nand UO_227 (O_227,N_4931,N_4998);
nand UO_228 (O_228,N_4928,N_4967);
xor UO_229 (O_229,N_4986,N_4900);
nor UO_230 (O_230,N_4949,N_4916);
or UO_231 (O_231,N_4967,N_4965);
or UO_232 (O_232,N_4909,N_4974);
xor UO_233 (O_233,N_4994,N_4974);
xor UO_234 (O_234,N_4954,N_4992);
and UO_235 (O_235,N_4910,N_4996);
nor UO_236 (O_236,N_4944,N_4989);
and UO_237 (O_237,N_4940,N_4964);
nor UO_238 (O_238,N_4941,N_4982);
or UO_239 (O_239,N_4993,N_4949);
xor UO_240 (O_240,N_4954,N_4907);
nor UO_241 (O_241,N_4989,N_4952);
and UO_242 (O_242,N_4963,N_4931);
and UO_243 (O_243,N_4932,N_4997);
nand UO_244 (O_244,N_4940,N_4935);
or UO_245 (O_245,N_4956,N_4963);
xor UO_246 (O_246,N_4947,N_4996);
xor UO_247 (O_247,N_4960,N_4937);
and UO_248 (O_248,N_4993,N_4939);
or UO_249 (O_249,N_4916,N_4908);
xor UO_250 (O_250,N_4985,N_4945);
nand UO_251 (O_251,N_4941,N_4926);
xor UO_252 (O_252,N_4964,N_4924);
xnor UO_253 (O_253,N_4944,N_4992);
or UO_254 (O_254,N_4943,N_4948);
and UO_255 (O_255,N_4948,N_4957);
and UO_256 (O_256,N_4930,N_4975);
nor UO_257 (O_257,N_4936,N_4972);
nor UO_258 (O_258,N_4932,N_4992);
nor UO_259 (O_259,N_4979,N_4900);
or UO_260 (O_260,N_4913,N_4905);
nor UO_261 (O_261,N_4918,N_4961);
and UO_262 (O_262,N_4915,N_4947);
or UO_263 (O_263,N_4943,N_4913);
and UO_264 (O_264,N_4916,N_4944);
nand UO_265 (O_265,N_4961,N_4958);
nand UO_266 (O_266,N_4923,N_4927);
or UO_267 (O_267,N_4900,N_4993);
nor UO_268 (O_268,N_4966,N_4991);
or UO_269 (O_269,N_4945,N_4962);
or UO_270 (O_270,N_4952,N_4957);
and UO_271 (O_271,N_4918,N_4958);
and UO_272 (O_272,N_4982,N_4949);
nor UO_273 (O_273,N_4983,N_4940);
nand UO_274 (O_274,N_4911,N_4993);
and UO_275 (O_275,N_4969,N_4994);
nor UO_276 (O_276,N_4937,N_4941);
nand UO_277 (O_277,N_4951,N_4945);
xor UO_278 (O_278,N_4948,N_4965);
and UO_279 (O_279,N_4999,N_4946);
xor UO_280 (O_280,N_4972,N_4974);
or UO_281 (O_281,N_4961,N_4925);
xnor UO_282 (O_282,N_4981,N_4974);
nor UO_283 (O_283,N_4962,N_4946);
or UO_284 (O_284,N_4957,N_4907);
or UO_285 (O_285,N_4915,N_4986);
nor UO_286 (O_286,N_4931,N_4924);
nor UO_287 (O_287,N_4907,N_4965);
or UO_288 (O_288,N_4986,N_4952);
xor UO_289 (O_289,N_4933,N_4972);
nand UO_290 (O_290,N_4910,N_4962);
nor UO_291 (O_291,N_4947,N_4934);
xnor UO_292 (O_292,N_4914,N_4985);
nand UO_293 (O_293,N_4971,N_4989);
nor UO_294 (O_294,N_4911,N_4963);
xnor UO_295 (O_295,N_4986,N_4973);
nor UO_296 (O_296,N_4966,N_4935);
xnor UO_297 (O_297,N_4910,N_4942);
or UO_298 (O_298,N_4984,N_4925);
nor UO_299 (O_299,N_4915,N_4963);
nor UO_300 (O_300,N_4952,N_4956);
and UO_301 (O_301,N_4919,N_4977);
or UO_302 (O_302,N_4909,N_4968);
or UO_303 (O_303,N_4949,N_4950);
and UO_304 (O_304,N_4995,N_4941);
or UO_305 (O_305,N_4959,N_4947);
xnor UO_306 (O_306,N_4910,N_4965);
nor UO_307 (O_307,N_4996,N_4967);
xor UO_308 (O_308,N_4929,N_4924);
nand UO_309 (O_309,N_4940,N_4921);
and UO_310 (O_310,N_4937,N_4913);
and UO_311 (O_311,N_4964,N_4928);
xor UO_312 (O_312,N_4994,N_4936);
and UO_313 (O_313,N_4958,N_4939);
or UO_314 (O_314,N_4972,N_4979);
or UO_315 (O_315,N_4930,N_4948);
xnor UO_316 (O_316,N_4948,N_4961);
or UO_317 (O_317,N_4906,N_4991);
xor UO_318 (O_318,N_4946,N_4964);
nand UO_319 (O_319,N_4956,N_4904);
nand UO_320 (O_320,N_4950,N_4999);
nor UO_321 (O_321,N_4923,N_4975);
xor UO_322 (O_322,N_4938,N_4958);
xor UO_323 (O_323,N_4989,N_4990);
nand UO_324 (O_324,N_4947,N_4953);
xnor UO_325 (O_325,N_4936,N_4985);
or UO_326 (O_326,N_4931,N_4951);
and UO_327 (O_327,N_4934,N_4944);
xor UO_328 (O_328,N_4933,N_4956);
nor UO_329 (O_329,N_4990,N_4991);
and UO_330 (O_330,N_4984,N_4960);
xor UO_331 (O_331,N_4984,N_4994);
or UO_332 (O_332,N_4950,N_4961);
nor UO_333 (O_333,N_4958,N_4992);
or UO_334 (O_334,N_4916,N_4955);
and UO_335 (O_335,N_4920,N_4949);
or UO_336 (O_336,N_4986,N_4997);
nor UO_337 (O_337,N_4918,N_4941);
and UO_338 (O_338,N_4972,N_4902);
or UO_339 (O_339,N_4996,N_4909);
nor UO_340 (O_340,N_4946,N_4956);
nor UO_341 (O_341,N_4942,N_4900);
and UO_342 (O_342,N_4956,N_4922);
xnor UO_343 (O_343,N_4977,N_4913);
nand UO_344 (O_344,N_4916,N_4936);
or UO_345 (O_345,N_4946,N_4985);
xnor UO_346 (O_346,N_4964,N_4997);
or UO_347 (O_347,N_4998,N_4929);
nand UO_348 (O_348,N_4946,N_4948);
nand UO_349 (O_349,N_4910,N_4933);
nand UO_350 (O_350,N_4912,N_4953);
or UO_351 (O_351,N_4983,N_4982);
nor UO_352 (O_352,N_4933,N_4923);
or UO_353 (O_353,N_4980,N_4957);
and UO_354 (O_354,N_4916,N_4930);
nor UO_355 (O_355,N_4951,N_4908);
xor UO_356 (O_356,N_4977,N_4916);
nand UO_357 (O_357,N_4943,N_4906);
and UO_358 (O_358,N_4971,N_4914);
and UO_359 (O_359,N_4999,N_4924);
and UO_360 (O_360,N_4987,N_4997);
nand UO_361 (O_361,N_4961,N_4954);
nor UO_362 (O_362,N_4950,N_4941);
xor UO_363 (O_363,N_4968,N_4995);
xnor UO_364 (O_364,N_4955,N_4944);
nor UO_365 (O_365,N_4991,N_4988);
and UO_366 (O_366,N_4915,N_4966);
or UO_367 (O_367,N_4910,N_4905);
or UO_368 (O_368,N_4926,N_4996);
xor UO_369 (O_369,N_4990,N_4970);
and UO_370 (O_370,N_4910,N_4967);
xnor UO_371 (O_371,N_4998,N_4904);
and UO_372 (O_372,N_4906,N_4953);
and UO_373 (O_373,N_4985,N_4975);
xor UO_374 (O_374,N_4914,N_4988);
nor UO_375 (O_375,N_4923,N_4980);
or UO_376 (O_376,N_4981,N_4902);
or UO_377 (O_377,N_4978,N_4943);
xor UO_378 (O_378,N_4938,N_4937);
xor UO_379 (O_379,N_4949,N_4958);
nand UO_380 (O_380,N_4953,N_4983);
or UO_381 (O_381,N_4985,N_4976);
xnor UO_382 (O_382,N_4954,N_4959);
and UO_383 (O_383,N_4965,N_4906);
or UO_384 (O_384,N_4974,N_4920);
and UO_385 (O_385,N_4949,N_4918);
nor UO_386 (O_386,N_4929,N_4941);
nand UO_387 (O_387,N_4949,N_4942);
xor UO_388 (O_388,N_4972,N_4946);
xnor UO_389 (O_389,N_4930,N_4934);
nand UO_390 (O_390,N_4974,N_4946);
xor UO_391 (O_391,N_4903,N_4987);
nor UO_392 (O_392,N_4973,N_4923);
nand UO_393 (O_393,N_4901,N_4983);
or UO_394 (O_394,N_4981,N_4945);
xnor UO_395 (O_395,N_4985,N_4916);
xnor UO_396 (O_396,N_4918,N_4952);
and UO_397 (O_397,N_4970,N_4947);
xor UO_398 (O_398,N_4956,N_4924);
and UO_399 (O_399,N_4960,N_4938);
nand UO_400 (O_400,N_4905,N_4976);
nor UO_401 (O_401,N_4934,N_4969);
or UO_402 (O_402,N_4908,N_4984);
xor UO_403 (O_403,N_4918,N_4919);
and UO_404 (O_404,N_4961,N_4909);
and UO_405 (O_405,N_4976,N_4917);
xor UO_406 (O_406,N_4969,N_4950);
or UO_407 (O_407,N_4978,N_4911);
nor UO_408 (O_408,N_4917,N_4964);
xor UO_409 (O_409,N_4996,N_4929);
nor UO_410 (O_410,N_4977,N_4997);
or UO_411 (O_411,N_4981,N_4944);
and UO_412 (O_412,N_4934,N_4913);
nor UO_413 (O_413,N_4991,N_4938);
xor UO_414 (O_414,N_4985,N_4974);
nand UO_415 (O_415,N_4994,N_4991);
and UO_416 (O_416,N_4970,N_4920);
nor UO_417 (O_417,N_4935,N_4913);
or UO_418 (O_418,N_4905,N_4906);
or UO_419 (O_419,N_4957,N_4914);
or UO_420 (O_420,N_4939,N_4933);
xnor UO_421 (O_421,N_4926,N_4950);
nor UO_422 (O_422,N_4950,N_4932);
and UO_423 (O_423,N_4936,N_4950);
or UO_424 (O_424,N_4920,N_4950);
nand UO_425 (O_425,N_4940,N_4955);
nand UO_426 (O_426,N_4939,N_4982);
xnor UO_427 (O_427,N_4992,N_4935);
nor UO_428 (O_428,N_4944,N_4978);
or UO_429 (O_429,N_4957,N_4994);
and UO_430 (O_430,N_4992,N_4989);
xor UO_431 (O_431,N_4934,N_4948);
nor UO_432 (O_432,N_4974,N_4963);
xor UO_433 (O_433,N_4942,N_4905);
xor UO_434 (O_434,N_4997,N_4930);
xnor UO_435 (O_435,N_4965,N_4983);
or UO_436 (O_436,N_4996,N_4935);
and UO_437 (O_437,N_4914,N_4921);
nor UO_438 (O_438,N_4986,N_4953);
and UO_439 (O_439,N_4998,N_4933);
xor UO_440 (O_440,N_4900,N_4939);
and UO_441 (O_441,N_4925,N_4934);
or UO_442 (O_442,N_4955,N_4945);
or UO_443 (O_443,N_4974,N_4919);
nor UO_444 (O_444,N_4976,N_4962);
nor UO_445 (O_445,N_4998,N_4902);
or UO_446 (O_446,N_4905,N_4948);
or UO_447 (O_447,N_4911,N_4971);
nor UO_448 (O_448,N_4960,N_4905);
xnor UO_449 (O_449,N_4996,N_4978);
xor UO_450 (O_450,N_4947,N_4948);
nand UO_451 (O_451,N_4963,N_4946);
xnor UO_452 (O_452,N_4973,N_4953);
nand UO_453 (O_453,N_4927,N_4967);
nor UO_454 (O_454,N_4993,N_4921);
and UO_455 (O_455,N_4907,N_4924);
nand UO_456 (O_456,N_4921,N_4931);
and UO_457 (O_457,N_4935,N_4941);
or UO_458 (O_458,N_4907,N_4966);
xor UO_459 (O_459,N_4914,N_4982);
or UO_460 (O_460,N_4926,N_4905);
and UO_461 (O_461,N_4951,N_4985);
xnor UO_462 (O_462,N_4979,N_4909);
and UO_463 (O_463,N_4985,N_4964);
nand UO_464 (O_464,N_4941,N_4957);
or UO_465 (O_465,N_4977,N_4935);
nand UO_466 (O_466,N_4984,N_4935);
nor UO_467 (O_467,N_4908,N_4963);
xor UO_468 (O_468,N_4906,N_4927);
xor UO_469 (O_469,N_4914,N_4937);
or UO_470 (O_470,N_4993,N_4959);
and UO_471 (O_471,N_4999,N_4958);
xnor UO_472 (O_472,N_4914,N_4909);
or UO_473 (O_473,N_4912,N_4996);
nor UO_474 (O_474,N_4923,N_4998);
xor UO_475 (O_475,N_4968,N_4980);
nor UO_476 (O_476,N_4902,N_4923);
or UO_477 (O_477,N_4997,N_4972);
xnor UO_478 (O_478,N_4903,N_4923);
nor UO_479 (O_479,N_4913,N_4951);
nor UO_480 (O_480,N_4995,N_4997);
nand UO_481 (O_481,N_4950,N_4971);
nand UO_482 (O_482,N_4943,N_4987);
or UO_483 (O_483,N_4966,N_4937);
xnor UO_484 (O_484,N_4921,N_4912);
nand UO_485 (O_485,N_4982,N_4992);
and UO_486 (O_486,N_4968,N_4920);
nand UO_487 (O_487,N_4945,N_4997);
nand UO_488 (O_488,N_4920,N_4918);
and UO_489 (O_489,N_4948,N_4972);
nand UO_490 (O_490,N_4921,N_4977);
xor UO_491 (O_491,N_4994,N_4932);
xnor UO_492 (O_492,N_4959,N_4984);
or UO_493 (O_493,N_4911,N_4926);
nor UO_494 (O_494,N_4901,N_4966);
xnor UO_495 (O_495,N_4942,N_4955);
nand UO_496 (O_496,N_4996,N_4959);
and UO_497 (O_497,N_4945,N_4970);
and UO_498 (O_498,N_4921,N_4927);
nand UO_499 (O_499,N_4924,N_4923);
or UO_500 (O_500,N_4915,N_4904);
and UO_501 (O_501,N_4913,N_4923);
xnor UO_502 (O_502,N_4976,N_4914);
and UO_503 (O_503,N_4964,N_4988);
or UO_504 (O_504,N_4970,N_4902);
nand UO_505 (O_505,N_4913,N_4950);
or UO_506 (O_506,N_4917,N_4918);
and UO_507 (O_507,N_4952,N_4916);
nand UO_508 (O_508,N_4972,N_4917);
xor UO_509 (O_509,N_4985,N_4923);
or UO_510 (O_510,N_4951,N_4911);
or UO_511 (O_511,N_4912,N_4964);
nand UO_512 (O_512,N_4961,N_4903);
nand UO_513 (O_513,N_4960,N_4971);
or UO_514 (O_514,N_4974,N_4988);
nor UO_515 (O_515,N_4906,N_4945);
and UO_516 (O_516,N_4908,N_4907);
nand UO_517 (O_517,N_4949,N_4966);
xor UO_518 (O_518,N_4940,N_4924);
xnor UO_519 (O_519,N_4960,N_4929);
nand UO_520 (O_520,N_4900,N_4926);
nand UO_521 (O_521,N_4955,N_4987);
nor UO_522 (O_522,N_4968,N_4994);
xor UO_523 (O_523,N_4980,N_4941);
nor UO_524 (O_524,N_4904,N_4932);
or UO_525 (O_525,N_4959,N_4934);
and UO_526 (O_526,N_4937,N_4998);
xor UO_527 (O_527,N_4958,N_4972);
or UO_528 (O_528,N_4917,N_4958);
or UO_529 (O_529,N_4971,N_4949);
nand UO_530 (O_530,N_4906,N_4941);
nand UO_531 (O_531,N_4957,N_4981);
and UO_532 (O_532,N_4900,N_4911);
nor UO_533 (O_533,N_4977,N_4958);
and UO_534 (O_534,N_4960,N_4967);
or UO_535 (O_535,N_4907,N_4927);
or UO_536 (O_536,N_4964,N_4948);
and UO_537 (O_537,N_4906,N_4940);
and UO_538 (O_538,N_4903,N_4957);
nand UO_539 (O_539,N_4933,N_4913);
nor UO_540 (O_540,N_4966,N_4923);
nor UO_541 (O_541,N_4984,N_4913);
and UO_542 (O_542,N_4985,N_4910);
or UO_543 (O_543,N_4915,N_4958);
or UO_544 (O_544,N_4912,N_4933);
or UO_545 (O_545,N_4962,N_4933);
xnor UO_546 (O_546,N_4910,N_4908);
nand UO_547 (O_547,N_4944,N_4974);
nand UO_548 (O_548,N_4964,N_4976);
nor UO_549 (O_549,N_4960,N_4991);
or UO_550 (O_550,N_4990,N_4988);
nor UO_551 (O_551,N_4927,N_4933);
and UO_552 (O_552,N_4918,N_4936);
xnor UO_553 (O_553,N_4937,N_4959);
xnor UO_554 (O_554,N_4985,N_4921);
xnor UO_555 (O_555,N_4963,N_4910);
or UO_556 (O_556,N_4901,N_4938);
and UO_557 (O_557,N_4927,N_4953);
xor UO_558 (O_558,N_4988,N_4922);
or UO_559 (O_559,N_4941,N_4993);
or UO_560 (O_560,N_4921,N_4923);
nand UO_561 (O_561,N_4941,N_4989);
nand UO_562 (O_562,N_4934,N_4997);
xor UO_563 (O_563,N_4974,N_4936);
xor UO_564 (O_564,N_4906,N_4974);
nor UO_565 (O_565,N_4947,N_4940);
nor UO_566 (O_566,N_4924,N_4937);
or UO_567 (O_567,N_4910,N_4921);
nor UO_568 (O_568,N_4995,N_4934);
xnor UO_569 (O_569,N_4942,N_4933);
xnor UO_570 (O_570,N_4945,N_4978);
and UO_571 (O_571,N_4911,N_4937);
nor UO_572 (O_572,N_4975,N_4902);
nand UO_573 (O_573,N_4986,N_4927);
nand UO_574 (O_574,N_4984,N_4900);
and UO_575 (O_575,N_4949,N_4991);
nor UO_576 (O_576,N_4981,N_4900);
xnor UO_577 (O_577,N_4977,N_4915);
or UO_578 (O_578,N_4903,N_4911);
nor UO_579 (O_579,N_4990,N_4920);
or UO_580 (O_580,N_4934,N_4968);
and UO_581 (O_581,N_4959,N_4992);
xor UO_582 (O_582,N_4981,N_4977);
xor UO_583 (O_583,N_4979,N_4980);
nor UO_584 (O_584,N_4946,N_4931);
nor UO_585 (O_585,N_4966,N_4988);
nor UO_586 (O_586,N_4901,N_4960);
nor UO_587 (O_587,N_4985,N_4980);
and UO_588 (O_588,N_4932,N_4947);
xnor UO_589 (O_589,N_4983,N_4909);
or UO_590 (O_590,N_4922,N_4983);
nand UO_591 (O_591,N_4920,N_4999);
nand UO_592 (O_592,N_4981,N_4925);
and UO_593 (O_593,N_4961,N_4994);
nor UO_594 (O_594,N_4922,N_4918);
nor UO_595 (O_595,N_4955,N_4965);
nor UO_596 (O_596,N_4941,N_4958);
nor UO_597 (O_597,N_4903,N_4988);
and UO_598 (O_598,N_4945,N_4933);
or UO_599 (O_599,N_4904,N_4914);
nor UO_600 (O_600,N_4977,N_4911);
and UO_601 (O_601,N_4991,N_4986);
nor UO_602 (O_602,N_4910,N_4975);
nor UO_603 (O_603,N_4925,N_4997);
and UO_604 (O_604,N_4994,N_4921);
xor UO_605 (O_605,N_4994,N_4941);
xnor UO_606 (O_606,N_4944,N_4922);
nand UO_607 (O_607,N_4948,N_4998);
and UO_608 (O_608,N_4914,N_4952);
xnor UO_609 (O_609,N_4925,N_4965);
xnor UO_610 (O_610,N_4997,N_4900);
nand UO_611 (O_611,N_4995,N_4927);
nand UO_612 (O_612,N_4992,N_4957);
xor UO_613 (O_613,N_4968,N_4987);
nand UO_614 (O_614,N_4936,N_4991);
nor UO_615 (O_615,N_4918,N_4923);
nand UO_616 (O_616,N_4952,N_4961);
or UO_617 (O_617,N_4910,N_4955);
and UO_618 (O_618,N_4914,N_4959);
nor UO_619 (O_619,N_4959,N_4985);
nor UO_620 (O_620,N_4946,N_4945);
or UO_621 (O_621,N_4924,N_4981);
nand UO_622 (O_622,N_4911,N_4916);
nand UO_623 (O_623,N_4976,N_4906);
xnor UO_624 (O_624,N_4942,N_4957);
xor UO_625 (O_625,N_4975,N_4907);
xor UO_626 (O_626,N_4984,N_4907);
nand UO_627 (O_627,N_4960,N_4959);
or UO_628 (O_628,N_4957,N_4967);
xor UO_629 (O_629,N_4973,N_4927);
or UO_630 (O_630,N_4996,N_4904);
nand UO_631 (O_631,N_4970,N_4979);
or UO_632 (O_632,N_4935,N_4948);
or UO_633 (O_633,N_4989,N_4940);
xor UO_634 (O_634,N_4988,N_4969);
xnor UO_635 (O_635,N_4956,N_4907);
nor UO_636 (O_636,N_4933,N_4926);
xnor UO_637 (O_637,N_4994,N_4937);
nor UO_638 (O_638,N_4999,N_4947);
and UO_639 (O_639,N_4995,N_4994);
nor UO_640 (O_640,N_4951,N_4965);
and UO_641 (O_641,N_4919,N_4978);
or UO_642 (O_642,N_4997,N_4992);
xnor UO_643 (O_643,N_4980,N_4906);
nor UO_644 (O_644,N_4967,N_4993);
xor UO_645 (O_645,N_4950,N_4963);
nor UO_646 (O_646,N_4987,N_4901);
nand UO_647 (O_647,N_4934,N_4938);
nor UO_648 (O_648,N_4978,N_4903);
nand UO_649 (O_649,N_4968,N_4913);
xnor UO_650 (O_650,N_4983,N_4979);
xnor UO_651 (O_651,N_4944,N_4987);
nor UO_652 (O_652,N_4991,N_4924);
nand UO_653 (O_653,N_4977,N_4969);
nor UO_654 (O_654,N_4986,N_4917);
or UO_655 (O_655,N_4974,N_4964);
or UO_656 (O_656,N_4910,N_4928);
xor UO_657 (O_657,N_4940,N_4998);
and UO_658 (O_658,N_4975,N_4961);
nor UO_659 (O_659,N_4947,N_4901);
and UO_660 (O_660,N_4947,N_4976);
nand UO_661 (O_661,N_4991,N_4941);
nand UO_662 (O_662,N_4967,N_4933);
and UO_663 (O_663,N_4900,N_4937);
nor UO_664 (O_664,N_4995,N_4991);
nand UO_665 (O_665,N_4967,N_4966);
nand UO_666 (O_666,N_4976,N_4902);
nand UO_667 (O_667,N_4950,N_4931);
or UO_668 (O_668,N_4914,N_4990);
nor UO_669 (O_669,N_4962,N_4938);
nand UO_670 (O_670,N_4931,N_4941);
or UO_671 (O_671,N_4998,N_4987);
or UO_672 (O_672,N_4939,N_4912);
xnor UO_673 (O_673,N_4932,N_4946);
xor UO_674 (O_674,N_4989,N_4953);
nor UO_675 (O_675,N_4913,N_4995);
and UO_676 (O_676,N_4900,N_4972);
or UO_677 (O_677,N_4944,N_4919);
xnor UO_678 (O_678,N_4999,N_4943);
or UO_679 (O_679,N_4921,N_4909);
xnor UO_680 (O_680,N_4984,N_4922);
and UO_681 (O_681,N_4912,N_4997);
or UO_682 (O_682,N_4997,N_4960);
or UO_683 (O_683,N_4957,N_4900);
nor UO_684 (O_684,N_4907,N_4968);
nand UO_685 (O_685,N_4908,N_4969);
xor UO_686 (O_686,N_4990,N_4973);
nand UO_687 (O_687,N_4951,N_4998);
nand UO_688 (O_688,N_4933,N_4929);
nor UO_689 (O_689,N_4938,N_4980);
or UO_690 (O_690,N_4974,N_4952);
or UO_691 (O_691,N_4936,N_4913);
nand UO_692 (O_692,N_4915,N_4988);
nor UO_693 (O_693,N_4951,N_4964);
xor UO_694 (O_694,N_4985,N_4996);
nand UO_695 (O_695,N_4998,N_4975);
nor UO_696 (O_696,N_4952,N_4970);
xor UO_697 (O_697,N_4985,N_4931);
nand UO_698 (O_698,N_4949,N_4963);
xor UO_699 (O_699,N_4991,N_4993);
or UO_700 (O_700,N_4952,N_4940);
nand UO_701 (O_701,N_4919,N_4917);
or UO_702 (O_702,N_4946,N_4918);
or UO_703 (O_703,N_4978,N_4940);
xor UO_704 (O_704,N_4938,N_4971);
nand UO_705 (O_705,N_4951,N_4946);
and UO_706 (O_706,N_4924,N_4906);
nor UO_707 (O_707,N_4975,N_4993);
nor UO_708 (O_708,N_4966,N_4977);
nor UO_709 (O_709,N_4920,N_4969);
xor UO_710 (O_710,N_4946,N_4983);
nor UO_711 (O_711,N_4974,N_4970);
xor UO_712 (O_712,N_4915,N_4935);
xor UO_713 (O_713,N_4906,N_4904);
xnor UO_714 (O_714,N_4942,N_4966);
xnor UO_715 (O_715,N_4921,N_4991);
nand UO_716 (O_716,N_4957,N_4998);
nand UO_717 (O_717,N_4991,N_4915);
nand UO_718 (O_718,N_4922,N_4907);
nor UO_719 (O_719,N_4983,N_4931);
nor UO_720 (O_720,N_4968,N_4960);
xnor UO_721 (O_721,N_4929,N_4985);
and UO_722 (O_722,N_4987,N_4910);
nand UO_723 (O_723,N_4985,N_4962);
nor UO_724 (O_724,N_4921,N_4970);
nand UO_725 (O_725,N_4970,N_4922);
and UO_726 (O_726,N_4998,N_4980);
nor UO_727 (O_727,N_4908,N_4964);
nand UO_728 (O_728,N_4961,N_4957);
nand UO_729 (O_729,N_4914,N_4991);
nand UO_730 (O_730,N_4912,N_4975);
nand UO_731 (O_731,N_4952,N_4965);
xor UO_732 (O_732,N_4951,N_4944);
nand UO_733 (O_733,N_4900,N_4904);
or UO_734 (O_734,N_4960,N_4935);
nand UO_735 (O_735,N_4934,N_4963);
and UO_736 (O_736,N_4982,N_4970);
and UO_737 (O_737,N_4917,N_4953);
or UO_738 (O_738,N_4981,N_4928);
nand UO_739 (O_739,N_4948,N_4949);
or UO_740 (O_740,N_4950,N_4942);
nand UO_741 (O_741,N_4928,N_4955);
xnor UO_742 (O_742,N_4948,N_4926);
xor UO_743 (O_743,N_4991,N_4905);
xor UO_744 (O_744,N_4957,N_4928);
nand UO_745 (O_745,N_4977,N_4944);
nor UO_746 (O_746,N_4987,N_4993);
or UO_747 (O_747,N_4992,N_4924);
and UO_748 (O_748,N_4938,N_4951);
nor UO_749 (O_749,N_4996,N_4914);
nand UO_750 (O_750,N_4936,N_4986);
nand UO_751 (O_751,N_4969,N_4965);
nand UO_752 (O_752,N_4942,N_4911);
and UO_753 (O_753,N_4919,N_4986);
nor UO_754 (O_754,N_4924,N_4967);
or UO_755 (O_755,N_4990,N_4942);
nand UO_756 (O_756,N_4975,N_4927);
or UO_757 (O_757,N_4913,N_4938);
nand UO_758 (O_758,N_4971,N_4919);
nor UO_759 (O_759,N_4960,N_4954);
nor UO_760 (O_760,N_4921,N_4996);
and UO_761 (O_761,N_4991,N_4989);
nand UO_762 (O_762,N_4974,N_4977);
nor UO_763 (O_763,N_4998,N_4909);
nand UO_764 (O_764,N_4997,N_4919);
xor UO_765 (O_765,N_4943,N_4907);
and UO_766 (O_766,N_4901,N_4911);
and UO_767 (O_767,N_4939,N_4969);
nor UO_768 (O_768,N_4961,N_4917);
nand UO_769 (O_769,N_4993,N_4917);
nor UO_770 (O_770,N_4920,N_4914);
and UO_771 (O_771,N_4904,N_4991);
nor UO_772 (O_772,N_4952,N_4909);
nor UO_773 (O_773,N_4963,N_4990);
xnor UO_774 (O_774,N_4989,N_4922);
nor UO_775 (O_775,N_4930,N_4966);
xor UO_776 (O_776,N_4933,N_4973);
and UO_777 (O_777,N_4947,N_4946);
nand UO_778 (O_778,N_4982,N_4938);
nor UO_779 (O_779,N_4979,N_4981);
and UO_780 (O_780,N_4967,N_4977);
xnor UO_781 (O_781,N_4947,N_4902);
xnor UO_782 (O_782,N_4955,N_4951);
nand UO_783 (O_783,N_4958,N_4989);
nor UO_784 (O_784,N_4961,N_4916);
and UO_785 (O_785,N_4938,N_4910);
nand UO_786 (O_786,N_4928,N_4915);
and UO_787 (O_787,N_4992,N_4921);
nor UO_788 (O_788,N_4998,N_4921);
nand UO_789 (O_789,N_4923,N_4963);
xnor UO_790 (O_790,N_4957,N_4931);
nor UO_791 (O_791,N_4964,N_4916);
nor UO_792 (O_792,N_4978,N_4948);
and UO_793 (O_793,N_4961,N_4911);
nor UO_794 (O_794,N_4957,N_4950);
xor UO_795 (O_795,N_4993,N_4969);
xor UO_796 (O_796,N_4971,N_4927);
and UO_797 (O_797,N_4920,N_4913);
and UO_798 (O_798,N_4961,N_4913);
or UO_799 (O_799,N_4920,N_4907);
and UO_800 (O_800,N_4944,N_4963);
or UO_801 (O_801,N_4984,N_4903);
and UO_802 (O_802,N_4992,N_4977);
xor UO_803 (O_803,N_4926,N_4972);
and UO_804 (O_804,N_4919,N_4943);
xnor UO_805 (O_805,N_4977,N_4996);
and UO_806 (O_806,N_4994,N_4981);
xnor UO_807 (O_807,N_4949,N_4939);
nor UO_808 (O_808,N_4947,N_4900);
xor UO_809 (O_809,N_4940,N_4963);
nor UO_810 (O_810,N_4904,N_4981);
and UO_811 (O_811,N_4945,N_4912);
xor UO_812 (O_812,N_4915,N_4921);
or UO_813 (O_813,N_4972,N_4991);
or UO_814 (O_814,N_4985,N_4967);
nor UO_815 (O_815,N_4920,N_4973);
nor UO_816 (O_816,N_4949,N_4946);
and UO_817 (O_817,N_4958,N_4959);
and UO_818 (O_818,N_4925,N_4956);
xor UO_819 (O_819,N_4915,N_4974);
and UO_820 (O_820,N_4989,N_4936);
nor UO_821 (O_821,N_4951,N_4949);
and UO_822 (O_822,N_4937,N_4908);
nor UO_823 (O_823,N_4965,N_4961);
xor UO_824 (O_824,N_4906,N_4929);
and UO_825 (O_825,N_4960,N_4939);
nor UO_826 (O_826,N_4921,N_4961);
nand UO_827 (O_827,N_4912,N_4940);
and UO_828 (O_828,N_4904,N_4922);
and UO_829 (O_829,N_4983,N_4959);
and UO_830 (O_830,N_4940,N_4957);
and UO_831 (O_831,N_4956,N_4936);
nor UO_832 (O_832,N_4998,N_4981);
xor UO_833 (O_833,N_4939,N_4946);
nor UO_834 (O_834,N_4977,N_4912);
nor UO_835 (O_835,N_4910,N_4956);
nor UO_836 (O_836,N_4923,N_4946);
nand UO_837 (O_837,N_4915,N_4975);
nor UO_838 (O_838,N_4958,N_4942);
and UO_839 (O_839,N_4970,N_4924);
or UO_840 (O_840,N_4907,N_4923);
or UO_841 (O_841,N_4942,N_4956);
nor UO_842 (O_842,N_4963,N_4920);
and UO_843 (O_843,N_4932,N_4905);
and UO_844 (O_844,N_4972,N_4995);
or UO_845 (O_845,N_4918,N_4910);
xor UO_846 (O_846,N_4958,N_4957);
or UO_847 (O_847,N_4974,N_4991);
and UO_848 (O_848,N_4982,N_4972);
or UO_849 (O_849,N_4957,N_4968);
or UO_850 (O_850,N_4999,N_4925);
or UO_851 (O_851,N_4979,N_4901);
or UO_852 (O_852,N_4983,N_4935);
nand UO_853 (O_853,N_4929,N_4907);
or UO_854 (O_854,N_4974,N_4914);
xor UO_855 (O_855,N_4900,N_4962);
nor UO_856 (O_856,N_4954,N_4990);
or UO_857 (O_857,N_4968,N_4901);
or UO_858 (O_858,N_4932,N_4961);
nand UO_859 (O_859,N_4994,N_4938);
nand UO_860 (O_860,N_4950,N_4928);
nor UO_861 (O_861,N_4924,N_4915);
xor UO_862 (O_862,N_4956,N_4917);
xor UO_863 (O_863,N_4960,N_4917);
nor UO_864 (O_864,N_4981,N_4927);
nand UO_865 (O_865,N_4949,N_4933);
nand UO_866 (O_866,N_4954,N_4905);
xor UO_867 (O_867,N_4943,N_4960);
or UO_868 (O_868,N_4911,N_4986);
or UO_869 (O_869,N_4939,N_4924);
nor UO_870 (O_870,N_4941,N_4953);
and UO_871 (O_871,N_4924,N_4984);
nand UO_872 (O_872,N_4951,N_4979);
xor UO_873 (O_873,N_4915,N_4936);
and UO_874 (O_874,N_4943,N_4990);
nand UO_875 (O_875,N_4974,N_4913);
nor UO_876 (O_876,N_4914,N_4930);
xor UO_877 (O_877,N_4903,N_4935);
xnor UO_878 (O_878,N_4916,N_4902);
or UO_879 (O_879,N_4979,N_4945);
and UO_880 (O_880,N_4916,N_4965);
nand UO_881 (O_881,N_4956,N_4969);
or UO_882 (O_882,N_4955,N_4980);
or UO_883 (O_883,N_4932,N_4990);
and UO_884 (O_884,N_4994,N_4978);
nand UO_885 (O_885,N_4958,N_4908);
and UO_886 (O_886,N_4926,N_4967);
or UO_887 (O_887,N_4974,N_4951);
or UO_888 (O_888,N_4909,N_4924);
xor UO_889 (O_889,N_4985,N_4934);
and UO_890 (O_890,N_4947,N_4936);
and UO_891 (O_891,N_4978,N_4990);
nand UO_892 (O_892,N_4985,N_4937);
nor UO_893 (O_893,N_4922,N_4914);
and UO_894 (O_894,N_4900,N_4903);
nor UO_895 (O_895,N_4956,N_4927);
nor UO_896 (O_896,N_4971,N_4996);
nand UO_897 (O_897,N_4991,N_4902);
and UO_898 (O_898,N_4905,N_4907);
nor UO_899 (O_899,N_4949,N_4987);
xor UO_900 (O_900,N_4948,N_4913);
and UO_901 (O_901,N_4958,N_4998);
nand UO_902 (O_902,N_4982,N_4907);
nand UO_903 (O_903,N_4920,N_4903);
nor UO_904 (O_904,N_4974,N_4933);
nand UO_905 (O_905,N_4996,N_4920);
nor UO_906 (O_906,N_4991,N_4959);
and UO_907 (O_907,N_4912,N_4958);
xnor UO_908 (O_908,N_4988,N_4970);
nor UO_909 (O_909,N_4911,N_4955);
xnor UO_910 (O_910,N_4957,N_4984);
nand UO_911 (O_911,N_4988,N_4927);
or UO_912 (O_912,N_4966,N_4973);
and UO_913 (O_913,N_4965,N_4994);
nand UO_914 (O_914,N_4911,N_4946);
and UO_915 (O_915,N_4949,N_4922);
or UO_916 (O_916,N_4982,N_4937);
and UO_917 (O_917,N_4923,N_4953);
or UO_918 (O_918,N_4921,N_4995);
xnor UO_919 (O_919,N_4993,N_4962);
and UO_920 (O_920,N_4929,N_4919);
nor UO_921 (O_921,N_4924,N_4910);
nor UO_922 (O_922,N_4901,N_4982);
and UO_923 (O_923,N_4907,N_4983);
or UO_924 (O_924,N_4985,N_4984);
xnor UO_925 (O_925,N_4993,N_4902);
nor UO_926 (O_926,N_4935,N_4973);
xnor UO_927 (O_927,N_4940,N_4919);
xor UO_928 (O_928,N_4958,N_4974);
nor UO_929 (O_929,N_4966,N_4992);
nand UO_930 (O_930,N_4939,N_4910);
nand UO_931 (O_931,N_4954,N_4935);
xor UO_932 (O_932,N_4960,N_4909);
nand UO_933 (O_933,N_4997,N_4969);
nor UO_934 (O_934,N_4980,N_4946);
nand UO_935 (O_935,N_4920,N_4941);
xor UO_936 (O_936,N_4957,N_4904);
xor UO_937 (O_937,N_4951,N_4994);
and UO_938 (O_938,N_4947,N_4903);
nand UO_939 (O_939,N_4940,N_4960);
xnor UO_940 (O_940,N_4926,N_4960);
or UO_941 (O_941,N_4973,N_4987);
xor UO_942 (O_942,N_4929,N_4947);
or UO_943 (O_943,N_4954,N_4914);
xor UO_944 (O_944,N_4912,N_4908);
nand UO_945 (O_945,N_4915,N_4946);
nand UO_946 (O_946,N_4968,N_4955);
xor UO_947 (O_947,N_4975,N_4957);
or UO_948 (O_948,N_4979,N_4995);
or UO_949 (O_949,N_4930,N_4951);
nor UO_950 (O_950,N_4981,N_4955);
or UO_951 (O_951,N_4907,N_4911);
and UO_952 (O_952,N_4993,N_4980);
nand UO_953 (O_953,N_4974,N_4912);
xnor UO_954 (O_954,N_4928,N_4959);
nor UO_955 (O_955,N_4956,N_4929);
and UO_956 (O_956,N_4921,N_4934);
nor UO_957 (O_957,N_4987,N_4942);
or UO_958 (O_958,N_4986,N_4947);
nand UO_959 (O_959,N_4902,N_4982);
xnor UO_960 (O_960,N_4989,N_4907);
nor UO_961 (O_961,N_4905,N_4980);
nor UO_962 (O_962,N_4915,N_4933);
xnor UO_963 (O_963,N_4958,N_4901);
nor UO_964 (O_964,N_4913,N_4964);
or UO_965 (O_965,N_4989,N_4951);
xnor UO_966 (O_966,N_4990,N_4933);
and UO_967 (O_967,N_4948,N_4906);
and UO_968 (O_968,N_4941,N_4996);
nor UO_969 (O_969,N_4931,N_4906);
nor UO_970 (O_970,N_4925,N_4915);
xnor UO_971 (O_971,N_4977,N_4928);
nand UO_972 (O_972,N_4937,N_4965);
nand UO_973 (O_973,N_4992,N_4936);
and UO_974 (O_974,N_4987,N_4917);
xnor UO_975 (O_975,N_4963,N_4961);
or UO_976 (O_976,N_4959,N_4906);
or UO_977 (O_977,N_4962,N_4971);
and UO_978 (O_978,N_4952,N_4904);
and UO_979 (O_979,N_4936,N_4911);
nand UO_980 (O_980,N_4929,N_4961);
and UO_981 (O_981,N_4979,N_4924);
xor UO_982 (O_982,N_4921,N_4908);
and UO_983 (O_983,N_4928,N_4953);
nand UO_984 (O_984,N_4944,N_4966);
nor UO_985 (O_985,N_4930,N_4940);
xnor UO_986 (O_986,N_4970,N_4993);
xor UO_987 (O_987,N_4907,N_4919);
or UO_988 (O_988,N_4955,N_4989);
nor UO_989 (O_989,N_4935,N_4979);
or UO_990 (O_990,N_4959,N_4957);
nor UO_991 (O_991,N_4903,N_4971);
nor UO_992 (O_992,N_4902,N_4985);
and UO_993 (O_993,N_4970,N_4904);
nand UO_994 (O_994,N_4907,N_4906);
and UO_995 (O_995,N_4926,N_4971);
nand UO_996 (O_996,N_4933,N_4940);
nor UO_997 (O_997,N_4963,N_4999);
nor UO_998 (O_998,N_4980,N_4932);
and UO_999 (O_999,N_4957,N_4972);
endmodule