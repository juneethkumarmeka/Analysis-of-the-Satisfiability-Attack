module basic_500_3000_500_3_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_81,In_56);
xnor U1 (N_1,In_398,In_440);
nand U2 (N_2,In_225,In_18);
nor U3 (N_3,In_90,In_7);
nor U4 (N_4,In_142,In_251);
and U5 (N_5,In_60,In_252);
nor U6 (N_6,In_190,In_394);
and U7 (N_7,In_278,In_391);
and U8 (N_8,In_285,In_408);
xor U9 (N_9,In_293,In_307);
nor U10 (N_10,In_448,In_26);
or U11 (N_11,In_355,In_465);
nor U12 (N_12,In_462,In_491);
xnor U13 (N_13,In_42,In_434);
nand U14 (N_14,In_55,In_373);
or U15 (N_15,In_486,In_33);
nor U16 (N_16,In_400,In_148);
nor U17 (N_17,In_354,In_405);
xnor U18 (N_18,In_195,In_356);
or U19 (N_19,In_302,In_29);
nand U20 (N_20,In_139,In_374);
or U21 (N_21,In_265,In_165);
nor U22 (N_22,In_143,In_468);
and U23 (N_23,In_368,In_85);
xnor U24 (N_24,In_79,In_464);
and U25 (N_25,In_97,In_48);
nor U26 (N_26,In_212,In_270);
xor U27 (N_27,In_4,In_403);
and U28 (N_28,In_235,In_104);
and U29 (N_29,In_3,In_473);
nor U30 (N_30,In_396,In_58);
nor U31 (N_31,In_99,In_122);
nand U32 (N_32,In_5,In_358);
and U33 (N_33,In_210,In_247);
and U34 (N_34,In_301,In_484);
xor U35 (N_35,In_427,In_232);
or U36 (N_36,In_53,In_315);
xor U37 (N_37,In_207,In_277);
xnor U38 (N_38,In_414,In_321);
xor U39 (N_39,In_96,In_250);
xor U40 (N_40,In_429,In_112);
xnor U41 (N_41,In_279,In_311);
nor U42 (N_42,In_337,In_351);
xor U43 (N_43,In_272,In_375);
and U44 (N_44,In_98,In_146);
nand U45 (N_45,In_13,In_449);
nand U46 (N_46,In_173,In_40);
xnor U47 (N_47,In_490,In_357);
and U48 (N_48,In_64,In_494);
nor U49 (N_49,In_213,In_0);
or U50 (N_50,In_482,In_336);
nand U51 (N_51,In_128,In_231);
nand U52 (N_52,In_20,In_6);
xor U53 (N_53,In_199,In_228);
nand U54 (N_54,In_348,In_492);
or U55 (N_55,In_230,In_281);
nor U56 (N_56,In_350,In_498);
nand U57 (N_57,In_153,In_262);
nand U58 (N_58,In_380,In_92);
or U59 (N_59,In_94,In_211);
nor U60 (N_60,In_91,In_168);
nor U61 (N_61,In_383,In_273);
and U62 (N_62,In_149,In_203);
xnor U63 (N_63,In_319,In_297);
or U64 (N_64,In_450,In_162);
or U65 (N_65,In_157,In_197);
or U66 (N_66,In_282,In_268);
nor U67 (N_67,In_187,In_331);
or U68 (N_68,In_127,In_38);
nor U69 (N_69,In_349,In_2);
xor U70 (N_70,In_344,In_343);
and U71 (N_71,In_107,In_339);
and U72 (N_72,In_335,In_25);
or U73 (N_73,In_275,In_223);
nor U74 (N_74,In_249,In_150);
and U75 (N_75,In_36,In_101);
nor U76 (N_76,In_341,In_177);
and U77 (N_77,In_392,In_50);
and U78 (N_78,In_410,In_239);
nor U79 (N_79,In_152,In_244);
xor U80 (N_80,In_109,In_167);
nand U81 (N_81,In_118,In_180);
and U82 (N_82,In_322,In_292);
or U83 (N_83,In_418,In_216);
and U84 (N_84,In_453,In_433);
nand U85 (N_85,In_372,In_46);
and U86 (N_86,In_169,In_1);
nand U87 (N_87,In_266,In_489);
and U88 (N_88,In_182,In_54);
and U89 (N_89,In_314,In_474);
and U90 (N_90,In_328,In_442);
nand U91 (N_91,In_352,In_136);
nand U92 (N_92,In_393,In_14);
or U93 (N_93,In_488,In_218);
or U94 (N_94,In_236,In_8);
or U95 (N_95,In_111,In_439);
and U96 (N_96,In_382,In_243);
and U97 (N_97,In_52,In_451);
and U98 (N_98,In_57,In_445);
nand U99 (N_99,In_255,In_360);
or U100 (N_100,In_455,In_27);
xnor U101 (N_101,In_367,In_176);
or U102 (N_102,In_209,In_318);
xnor U103 (N_103,In_110,In_78);
xnor U104 (N_104,In_459,In_191);
or U105 (N_105,In_181,In_446);
xor U106 (N_106,In_495,In_134);
nor U107 (N_107,In_271,In_144);
and U108 (N_108,In_208,In_407);
nand U109 (N_109,In_158,In_82);
nand U110 (N_110,In_346,In_59);
nand U111 (N_111,In_179,In_483);
xnor U112 (N_112,In_145,In_30);
xor U113 (N_113,In_411,In_276);
nand U114 (N_114,In_196,In_304);
and U115 (N_115,In_163,In_332);
or U116 (N_116,In_133,In_409);
nand U117 (N_117,In_456,In_204);
and U118 (N_118,In_245,In_119);
or U119 (N_119,In_184,In_366);
or U120 (N_120,In_469,In_34);
xnor U121 (N_121,In_37,In_384);
nor U122 (N_122,In_61,In_246);
nor U123 (N_123,In_39,In_379);
nor U124 (N_124,In_466,In_83);
or U125 (N_125,In_198,In_386);
or U126 (N_126,In_103,In_487);
and U127 (N_127,In_481,In_329);
nor U128 (N_128,In_364,In_217);
nand U129 (N_129,In_269,In_214);
nor U130 (N_130,In_71,In_288);
nand U131 (N_131,In_219,In_88);
xnor U132 (N_132,In_74,In_330);
xnor U133 (N_133,In_299,In_77);
nand U134 (N_134,In_406,In_256);
and U135 (N_135,In_140,In_447);
nor U136 (N_136,In_416,In_41);
xnor U137 (N_137,In_241,In_261);
or U138 (N_138,In_114,In_159);
nand U139 (N_139,In_108,In_189);
or U140 (N_140,In_397,In_477);
xor U141 (N_141,In_258,In_294);
xor U142 (N_142,In_417,In_170);
nor U143 (N_143,In_234,In_338);
and U144 (N_144,In_345,In_404);
xnor U145 (N_145,In_395,In_415);
nor U146 (N_146,In_308,In_160);
nand U147 (N_147,In_84,In_117);
and U148 (N_148,In_436,In_254);
nand U149 (N_149,In_151,In_296);
nand U150 (N_150,In_93,In_22);
xor U151 (N_151,In_444,In_267);
xnor U152 (N_152,In_385,In_432);
xnor U153 (N_153,In_284,In_206);
nand U154 (N_154,In_295,In_95);
nor U155 (N_155,In_132,In_124);
or U156 (N_156,In_12,In_125);
or U157 (N_157,In_342,In_120);
nand U158 (N_158,In_363,In_326);
nor U159 (N_159,In_376,In_479);
and U160 (N_160,In_70,In_28);
and U161 (N_161,In_340,In_161);
and U162 (N_162,In_290,In_80);
nor U163 (N_163,In_166,In_200);
or U164 (N_164,In_260,In_237);
and U165 (N_165,In_31,In_298);
and U166 (N_166,In_420,In_381);
or U167 (N_167,In_437,In_316);
or U168 (N_168,In_389,In_471);
nor U169 (N_169,In_129,In_300);
or U170 (N_170,In_113,In_23);
nand U171 (N_171,In_257,In_226);
nor U172 (N_172,In_478,In_493);
nor U173 (N_173,In_135,In_248);
and U174 (N_174,In_47,In_362);
xnor U175 (N_175,In_106,In_467);
nor U176 (N_176,In_460,In_105);
nand U177 (N_177,In_194,In_229);
and U178 (N_178,In_202,In_480);
or U179 (N_179,In_361,In_221);
or U180 (N_180,In_185,In_240);
xnor U181 (N_181,In_353,In_115);
or U182 (N_182,In_175,In_421);
and U183 (N_183,In_401,In_21);
nand U184 (N_184,In_438,In_121);
nand U185 (N_185,In_126,In_192);
or U186 (N_186,In_72,In_16);
nand U187 (N_187,In_238,In_320);
or U188 (N_188,In_422,In_323);
and U189 (N_189,In_388,In_306);
nand U190 (N_190,In_51,In_224);
xor U191 (N_191,In_164,In_220);
nand U192 (N_192,In_334,In_15);
and U193 (N_193,In_499,In_174);
nor U194 (N_194,In_123,In_274);
and U195 (N_195,In_371,In_86);
xnor U196 (N_196,In_201,In_222);
nor U197 (N_197,In_419,In_280);
nand U198 (N_198,In_309,In_283);
and U199 (N_199,In_67,In_65);
nand U200 (N_200,In_470,In_89);
and U201 (N_201,In_141,In_264);
nand U202 (N_202,In_413,In_378);
nand U203 (N_203,In_312,In_412);
nand U204 (N_204,In_443,In_155);
xnor U205 (N_205,In_172,In_327);
or U206 (N_206,In_313,In_171);
nor U207 (N_207,In_156,In_333);
or U208 (N_208,In_215,In_259);
nor U209 (N_209,In_325,In_11);
xnor U210 (N_210,In_497,In_423);
and U211 (N_211,In_66,In_45);
nor U212 (N_212,In_178,In_63);
xnor U213 (N_213,In_454,In_205);
nand U214 (N_214,In_377,In_359);
nor U215 (N_215,In_475,In_43);
xnor U216 (N_216,In_476,In_435);
nand U217 (N_217,In_472,In_147);
xnor U218 (N_218,In_87,In_365);
and U219 (N_219,In_263,In_289);
xor U220 (N_220,In_305,In_227);
and U221 (N_221,In_138,In_102);
and U222 (N_222,In_369,In_116);
and U223 (N_223,In_100,In_324);
nand U224 (N_224,In_463,In_183);
xnor U225 (N_225,In_452,In_390);
and U226 (N_226,In_253,In_287);
and U227 (N_227,In_242,In_399);
xnor U228 (N_228,In_10,In_17);
or U229 (N_229,In_458,In_49);
xor U230 (N_230,In_430,In_426);
nand U231 (N_231,In_69,In_24);
nand U232 (N_232,In_76,In_19);
xor U233 (N_233,In_233,In_154);
and U234 (N_234,In_370,In_424);
nand U235 (N_235,In_387,In_496);
nand U236 (N_236,In_286,In_186);
nand U237 (N_237,In_425,In_317);
and U238 (N_238,In_62,In_32);
nor U239 (N_239,In_441,In_68);
nand U240 (N_240,In_291,In_485);
or U241 (N_241,In_431,In_73);
or U242 (N_242,In_35,In_457);
and U243 (N_243,In_303,In_9);
nor U244 (N_244,In_131,In_130);
and U245 (N_245,In_402,In_137);
nand U246 (N_246,In_193,In_310);
nor U247 (N_247,In_347,In_75);
or U248 (N_248,In_44,In_428);
xnor U249 (N_249,In_188,In_461);
xor U250 (N_250,In_223,In_474);
or U251 (N_251,In_368,In_9);
and U252 (N_252,In_453,In_302);
or U253 (N_253,In_277,In_366);
and U254 (N_254,In_337,In_144);
xnor U255 (N_255,In_248,In_151);
nand U256 (N_256,In_428,In_142);
nand U257 (N_257,In_111,In_6);
xor U258 (N_258,In_426,In_258);
or U259 (N_259,In_287,In_202);
and U260 (N_260,In_287,In_151);
and U261 (N_261,In_216,In_299);
or U262 (N_262,In_101,In_486);
nor U263 (N_263,In_77,In_84);
xnor U264 (N_264,In_423,In_195);
nor U265 (N_265,In_490,In_459);
nor U266 (N_266,In_304,In_37);
xnor U267 (N_267,In_410,In_302);
or U268 (N_268,In_328,In_3);
nor U269 (N_269,In_307,In_74);
xor U270 (N_270,In_24,In_339);
nand U271 (N_271,In_52,In_388);
or U272 (N_272,In_205,In_35);
nand U273 (N_273,In_13,In_84);
nand U274 (N_274,In_226,In_261);
xor U275 (N_275,In_462,In_399);
nor U276 (N_276,In_142,In_471);
nor U277 (N_277,In_76,In_169);
nand U278 (N_278,In_29,In_173);
and U279 (N_279,In_179,In_77);
and U280 (N_280,In_63,In_317);
xnor U281 (N_281,In_365,In_106);
or U282 (N_282,In_31,In_93);
and U283 (N_283,In_495,In_298);
nand U284 (N_284,In_115,In_202);
and U285 (N_285,In_301,In_211);
nand U286 (N_286,In_43,In_448);
nand U287 (N_287,In_69,In_266);
xor U288 (N_288,In_97,In_429);
nand U289 (N_289,In_131,In_454);
xor U290 (N_290,In_432,In_47);
nor U291 (N_291,In_29,In_132);
or U292 (N_292,In_220,In_459);
or U293 (N_293,In_297,In_321);
xor U294 (N_294,In_487,In_287);
or U295 (N_295,In_366,In_143);
and U296 (N_296,In_124,In_329);
and U297 (N_297,In_392,In_482);
xor U298 (N_298,In_19,In_12);
nand U299 (N_299,In_428,In_380);
or U300 (N_300,In_393,In_194);
nand U301 (N_301,In_211,In_285);
and U302 (N_302,In_150,In_390);
nor U303 (N_303,In_449,In_450);
nor U304 (N_304,In_218,In_285);
and U305 (N_305,In_269,In_56);
xor U306 (N_306,In_268,In_239);
nor U307 (N_307,In_431,In_164);
and U308 (N_308,In_118,In_177);
or U309 (N_309,In_100,In_187);
nand U310 (N_310,In_447,In_309);
nor U311 (N_311,In_264,In_122);
nand U312 (N_312,In_420,In_48);
nand U313 (N_313,In_295,In_331);
nor U314 (N_314,In_352,In_184);
or U315 (N_315,In_467,In_237);
or U316 (N_316,In_331,In_365);
xor U317 (N_317,In_39,In_347);
and U318 (N_318,In_89,In_116);
and U319 (N_319,In_354,In_448);
nand U320 (N_320,In_494,In_449);
and U321 (N_321,In_428,In_208);
and U322 (N_322,In_153,In_2);
nand U323 (N_323,In_174,In_39);
or U324 (N_324,In_23,In_398);
or U325 (N_325,In_47,In_148);
or U326 (N_326,In_55,In_263);
nor U327 (N_327,In_121,In_204);
and U328 (N_328,In_135,In_6);
nand U329 (N_329,In_380,In_178);
xnor U330 (N_330,In_211,In_0);
xnor U331 (N_331,In_276,In_402);
nor U332 (N_332,In_105,In_389);
and U333 (N_333,In_267,In_493);
xnor U334 (N_334,In_221,In_113);
and U335 (N_335,In_231,In_300);
or U336 (N_336,In_342,In_232);
and U337 (N_337,In_275,In_347);
nor U338 (N_338,In_367,In_37);
xor U339 (N_339,In_350,In_488);
nand U340 (N_340,In_471,In_122);
xor U341 (N_341,In_279,In_173);
and U342 (N_342,In_219,In_296);
xnor U343 (N_343,In_316,In_346);
or U344 (N_344,In_339,In_95);
nor U345 (N_345,In_176,In_315);
nand U346 (N_346,In_391,In_129);
nor U347 (N_347,In_202,In_332);
nor U348 (N_348,In_279,In_410);
and U349 (N_349,In_411,In_264);
nor U350 (N_350,In_155,In_230);
and U351 (N_351,In_381,In_243);
or U352 (N_352,In_120,In_150);
or U353 (N_353,In_301,In_403);
xor U354 (N_354,In_152,In_7);
nor U355 (N_355,In_85,In_78);
nand U356 (N_356,In_367,In_83);
or U357 (N_357,In_209,In_414);
nor U358 (N_358,In_212,In_46);
and U359 (N_359,In_106,In_286);
or U360 (N_360,In_0,In_67);
and U361 (N_361,In_202,In_351);
and U362 (N_362,In_88,In_54);
nand U363 (N_363,In_339,In_280);
xnor U364 (N_364,In_456,In_153);
or U365 (N_365,In_302,In_467);
nor U366 (N_366,In_58,In_7);
xor U367 (N_367,In_75,In_325);
nor U368 (N_368,In_203,In_355);
nor U369 (N_369,In_56,In_12);
xor U370 (N_370,In_323,In_145);
nand U371 (N_371,In_354,In_350);
nor U372 (N_372,In_49,In_270);
xor U373 (N_373,In_66,In_357);
nand U374 (N_374,In_216,In_9);
xnor U375 (N_375,In_291,In_113);
xor U376 (N_376,In_175,In_246);
xor U377 (N_377,In_258,In_199);
or U378 (N_378,In_185,In_147);
nand U379 (N_379,In_469,In_19);
and U380 (N_380,In_143,In_354);
nor U381 (N_381,In_246,In_318);
xor U382 (N_382,In_177,In_185);
and U383 (N_383,In_309,In_17);
nor U384 (N_384,In_300,In_183);
xor U385 (N_385,In_175,In_406);
and U386 (N_386,In_182,In_27);
nor U387 (N_387,In_43,In_144);
or U388 (N_388,In_300,In_444);
nand U389 (N_389,In_386,In_202);
nor U390 (N_390,In_7,In_190);
nand U391 (N_391,In_99,In_220);
nor U392 (N_392,In_464,In_357);
and U393 (N_393,In_354,In_266);
xor U394 (N_394,In_302,In_359);
xnor U395 (N_395,In_353,In_306);
and U396 (N_396,In_364,In_106);
nand U397 (N_397,In_420,In_331);
and U398 (N_398,In_322,In_122);
and U399 (N_399,In_449,In_140);
nor U400 (N_400,In_86,In_208);
nand U401 (N_401,In_19,In_47);
xnor U402 (N_402,In_293,In_394);
or U403 (N_403,In_330,In_474);
and U404 (N_404,In_314,In_51);
nor U405 (N_405,In_307,In_179);
nand U406 (N_406,In_7,In_73);
nor U407 (N_407,In_241,In_221);
or U408 (N_408,In_157,In_133);
and U409 (N_409,In_398,In_24);
nand U410 (N_410,In_354,In_292);
or U411 (N_411,In_465,In_471);
and U412 (N_412,In_93,In_141);
nor U413 (N_413,In_341,In_258);
nor U414 (N_414,In_240,In_172);
xor U415 (N_415,In_106,In_339);
xor U416 (N_416,In_265,In_211);
or U417 (N_417,In_18,In_497);
or U418 (N_418,In_203,In_154);
nand U419 (N_419,In_49,In_229);
nand U420 (N_420,In_401,In_367);
and U421 (N_421,In_326,In_306);
nor U422 (N_422,In_259,In_491);
or U423 (N_423,In_237,In_198);
or U424 (N_424,In_60,In_393);
nand U425 (N_425,In_126,In_356);
nor U426 (N_426,In_297,In_231);
and U427 (N_427,In_445,In_260);
xor U428 (N_428,In_447,In_284);
or U429 (N_429,In_477,In_391);
and U430 (N_430,In_204,In_168);
nand U431 (N_431,In_15,In_137);
nor U432 (N_432,In_134,In_91);
nor U433 (N_433,In_159,In_50);
nand U434 (N_434,In_169,In_168);
nand U435 (N_435,In_176,In_422);
and U436 (N_436,In_250,In_483);
or U437 (N_437,In_391,In_393);
nor U438 (N_438,In_26,In_315);
nand U439 (N_439,In_103,In_435);
xnor U440 (N_440,In_162,In_329);
nor U441 (N_441,In_249,In_381);
or U442 (N_442,In_398,In_457);
and U443 (N_443,In_423,In_116);
and U444 (N_444,In_82,In_238);
and U445 (N_445,In_96,In_236);
xnor U446 (N_446,In_465,In_166);
nor U447 (N_447,In_403,In_333);
or U448 (N_448,In_53,In_6);
nor U449 (N_449,In_381,In_205);
and U450 (N_450,In_70,In_468);
or U451 (N_451,In_370,In_87);
nand U452 (N_452,In_221,In_118);
nand U453 (N_453,In_351,In_84);
and U454 (N_454,In_464,In_479);
nor U455 (N_455,In_201,In_233);
and U456 (N_456,In_295,In_164);
or U457 (N_457,In_117,In_357);
nor U458 (N_458,In_405,In_319);
and U459 (N_459,In_139,In_372);
xnor U460 (N_460,In_167,In_146);
nand U461 (N_461,In_371,In_419);
xnor U462 (N_462,In_350,In_327);
nor U463 (N_463,In_56,In_336);
and U464 (N_464,In_472,In_360);
and U465 (N_465,In_178,In_475);
nor U466 (N_466,In_365,In_191);
nor U467 (N_467,In_326,In_435);
nand U468 (N_468,In_304,In_30);
and U469 (N_469,In_76,In_364);
nand U470 (N_470,In_9,In_22);
xnor U471 (N_471,In_446,In_328);
xnor U472 (N_472,In_309,In_360);
and U473 (N_473,In_113,In_294);
and U474 (N_474,In_408,In_1);
xnor U475 (N_475,In_157,In_478);
xor U476 (N_476,In_46,In_165);
and U477 (N_477,In_258,In_288);
nor U478 (N_478,In_77,In_457);
nand U479 (N_479,In_276,In_90);
nand U480 (N_480,In_361,In_202);
and U481 (N_481,In_124,In_296);
and U482 (N_482,In_481,In_99);
or U483 (N_483,In_308,In_205);
nand U484 (N_484,In_296,In_125);
or U485 (N_485,In_355,In_23);
and U486 (N_486,In_358,In_82);
xor U487 (N_487,In_358,In_219);
or U488 (N_488,In_300,In_60);
or U489 (N_489,In_103,In_65);
xor U490 (N_490,In_41,In_117);
or U491 (N_491,In_478,In_292);
and U492 (N_492,In_261,In_486);
xnor U493 (N_493,In_320,In_101);
nand U494 (N_494,In_157,In_240);
xnor U495 (N_495,In_263,In_494);
xor U496 (N_496,In_198,In_453);
nand U497 (N_497,In_114,In_260);
nor U498 (N_498,In_277,In_402);
nor U499 (N_499,In_364,In_188);
nor U500 (N_500,In_202,In_148);
nor U501 (N_501,In_374,In_396);
nand U502 (N_502,In_318,In_121);
or U503 (N_503,In_470,In_384);
xnor U504 (N_504,In_80,In_269);
nor U505 (N_505,In_112,In_348);
xnor U506 (N_506,In_378,In_270);
or U507 (N_507,In_493,In_354);
or U508 (N_508,In_132,In_100);
xnor U509 (N_509,In_384,In_41);
and U510 (N_510,In_98,In_442);
or U511 (N_511,In_5,In_45);
nand U512 (N_512,In_247,In_303);
nor U513 (N_513,In_351,In_454);
or U514 (N_514,In_200,In_141);
xor U515 (N_515,In_352,In_162);
and U516 (N_516,In_89,In_171);
nand U517 (N_517,In_302,In_80);
xor U518 (N_518,In_115,In_472);
nor U519 (N_519,In_37,In_85);
and U520 (N_520,In_395,In_365);
nor U521 (N_521,In_112,In_21);
and U522 (N_522,In_244,In_350);
and U523 (N_523,In_217,In_331);
xor U524 (N_524,In_146,In_497);
or U525 (N_525,In_206,In_447);
nor U526 (N_526,In_39,In_1);
xnor U527 (N_527,In_228,In_241);
nand U528 (N_528,In_102,In_180);
xnor U529 (N_529,In_310,In_257);
nand U530 (N_530,In_474,In_379);
nand U531 (N_531,In_358,In_435);
xor U532 (N_532,In_25,In_331);
nand U533 (N_533,In_273,In_238);
or U534 (N_534,In_455,In_36);
or U535 (N_535,In_405,In_362);
nor U536 (N_536,In_294,In_307);
and U537 (N_537,In_489,In_145);
nand U538 (N_538,In_5,In_403);
and U539 (N_539,In_118,In_466);
or U540 (N_540,In_386,In_271);
or U541 (N_541,In_209,In_372);
xnor U542 (N_542,In_471,In_348);
or U543 (N_543,In_106,In_300);
and U544 (N_544,In_302,In_456);
nand U545 (N_545,In_490,In_317);
xor U546 (N_546,In_244,In_298);
and U547 (N_547,In_284,In_462);
and U548 (N_548,In_64,In_467);
nand U549 (N_549,In_105,In_321);
and U550 (N_550,In_417,In_357);
nor U551 (N_551,In_265,In_77);
or U552 (N_552,In_205,In_184);
nand U553 (N_553,In_245,In_454);
and U554 (N_554,In_105,In_490);
nor U555 (N_555,In_125,In_298);
nand U556 (N_556,In_38,In_249);
nor U557 (N_557,In_495,In_267);
and U558 (N_558,In_93,In_235);
xor U559 (N_559,In_394,In_176);
xor U560 (N_560,In_219,In_120);
and U561 (N_561,In_262,In_79);
nand U562 (N_562,In_269,In_18);
and U563 (N_563,In_465,In_291);
or U564 (N_564,In_329,In_420);
or U565 (N_565,In_333,In_458);
xnor U566 (N_566,In_407,In_147);
and U567 (N_567,In_11,In_62);
or U568 (N_568,In_267,In_134);
and U569 (N_569,In_39,In_385);
or U570 (N_570,In_52,In_85);
nand U571 (N_571,In_442,In_23);
nand U572 (N_572,In_23,In_297);
nor U573 (N_573,In_87,In_374);
nand U574 (N_574,In_29,In_338);
xor U575 (N_575,In_301,In_321);
or U576 (N_576,In_392,In_428);
nor U577 (N_577,In_488,In_11);
and U578 (N_578,In_248,In_380);
or U579 (N_579,In_107,In_121);
or U580 (N_580,In_34,In_496);
nor U581 (N_581,In_407,In_212);
xor U582 (N_582,In_50,In_81);
nand U583 (N_583,In_100,In_129);
and U584 (N_584,In_319,In_291);
nor U585 (N_585,In_40,In_238);
or U586 (N_586,In_177,In_46);
xnor U587 (N_587,In_62,In_60);
xor U588 (N_588,In_213,In_267);
or U589 (N_589,In_139,In_213);
and U590 (N_590,In_450,In_292);
or U591 (N_591,In_148,In_73);
nand U592 (N_592,In_354,In_123);
nor U593 (N_593,In_351,In_261);
and U594 (N_594,In_430,In_347);
and U595 (N_595,In_467,In_271);
xor U596 (N_596,In_347,In_481);
xnor U597 (N_597,In_9,In_424);
nor U598 (N_598,In_185,In_199);
nand U599 (N_599,In_398,In_162);
nor U600 (N_600,In_253,In_237);
and U601 (N_601,In_131,In_135);
xnor U602 (N_602,In_3,In_341);
nor U603 (N_603,In_358,In_151);
or U604 (N_604,In_265,In_354);
xnor U605 (N_605,In_185,In_277);
or U606 (N_606,In_109,In_300);
nor U607 (N_607,In_223,In_59);
nor U608 (N_608,In_238,In_482);
and U609 (N_609,In_290,In_348);
or U610 (N_610,In_320,In_316);
nand U611 (N_611,In_449,In_467);
xnor U612 (N_612,In_460,In_319);
nand U613 (N_613,In_449,In_369);
xor U614 (N_614,In_285,In_231);
or U615 (N_615,In_425,In_287);
or U616 (N_616,In_215,In_407);
nand U617 (N_617,In_173,In_167);
nor U618 (N_618,In_439,In_221);
nand U619 (N_619,In_29,In_270);
nand U620 (N_620,In_395,In_280);
nand U621 (N_621,In_462,In_402);
xnor U622 (N_622,In_175,In_498);
nand U623 (N_623,In_319,In_56);
nor U624 (N_624,In_356,In_77);
or U625 (N_625,In_459,In_322);
or U626 (N_626,In_489,In_235);
nor U627 (N_627,In_180,In_478);
nand U628 (N_628,In_353,In_297);
or U629 (N_629,In_143,In_128);
xor U630 (N_630,In_225,In_323);
or U631 (N_631,In_64,In_262);
xor U632 (N_632,In_32,In_276);
and U633 (N_633,In_93,In_243);
or U634 (N_634,In_48,In_276);
and U635 (N_635,In_188,In_127);
nand U636 (N_636,In_349,In_262);
nand U637 (N_637,In_78,In_108);
xnor U638 (N_638,In_53,In_360);
nand U639 (N_639,In_74,In_263);
nand U640 (N_640,In_17,In_407);
nand U641 (N_641,In_399,In_286);
or U642 (N_642,In_103,In_109);
or U643 (N_643,In_498,In_89);
and U644 (N_644,In_217,In_263);
xor U645 (N_645,In_1,In_103);
or U646 (N_646,In_40,In_206);
and U647 (N_647,In_265,In_177);
nand U648 (N_648,In_144,In_483);
nand U649 (N_649,In_128,In_214);
or U650 (N_650,In_0,In_140);
and U651 (N_651,In_7,In_236);
and U652 (N_652,In_311,In_360);
nand U653 (N_653,In_347,In_336);
and U654 (N_654,In_415,In_341);
or U655 (N_655,In_38,In_331);
and U656 (N_656,In_351,In_438);
nand U657 (N_657,In_230,In_414);
xor U658 (N_658,In_50,In_465);
nor U659 (N_659,In_172,In_443);
or U660 (N_660,In_199,In_311);
nand U661 (N_661,In_283,In_421);
xor U662 (N_662,In_161,In_261);
or U663 (N_663,In_476,In_191);
and U664 (N_664,In_432,In_54);
nand U665 (N_665,In_43,In_400);
nand U666 (N_666,In_436,In_413);
or U667 (N_667,In_483,In_491);
nand U668 (N_668,In_252,In_85);
or U669 (N_669,In_234,In_26);
nand U670 (N_670,In_38,In_372);
nand U671 (N_671,In_275,In_317);
xnor U672 (N_672,In_25,In_391);
nor U673 (N_673,In_448,In_437);
or U674 (N_674,In_363,In_385);
and U675 (N_675,In_6,In_305);
or U676 (N_676,In_431,In_65);
xor U677 (N_677,In_149,In_414);
nand U678 (N_678,In_76,In_109);
xor U679 (N_679,In_308,In_456);
or U680 (N_680,In_486,In_129);
xnor U681 (N_681,In_360,In_73);
xor U682 (N_682,In_60,In_109);
nand U683 (N_683,In_62,In_285);
nor U684 (N_684,In_425,In_331);
nor U685 (N_685,In_31,In_265);
nand U686 (N_686,In_352,In_145);
nand U687 (N_687,In_459,In_111);
and U688 (N_688,In_301,In_455);
nand U689 (N_689,In_61,In_496);
nand U690 (N_690,In_386,In_168);
or U691 (N_691,In_98,In_161);
and U692 (N_692,In_393,In_181);
nor U693 (N_693,In_185,In_342);
nand U694 (N_694,In_69,In_57);
xor U695 (N_695,In_435,In_229);
xnor U696 (N_696,In_106,In_337);
nand U697 (N_697,In_44,In_423);
nand U698 (N_698,In_70,In_64);
nor U699 (N_699,In_108,In_274);
nor U700 (N_700,In_491,In_52);
xor U701 (N_701,In_154,In_63);
xnor U702 (N_702,In_50,In_355);
and U703 (N_703,In_402,In_412);
xnor U704 (N_704,In_59,In_342);
xor U705 (N_705,In_202,In_424);
and U706 (N_706,In_323,In_397);
and U707 (N_707,In_196,In_166);
xor U708 (N_708,In_226,In_154);
xnor U709 (N_709,In_81,In_152);
and U710 (N_710,In_391,In_315);
xnor U711 (N_711,In_327,In_469);
or U712 (N_712,In_20,In_247);
or U713 (N_713,In_30,In_73);
xor U714 (N_714,In_346,In_488);
and U715 (N_715,In_249,In_15);
xor U716 (N_716,In_33,In_85);
and U717 (N_717,In_342,In_83);
or U718 (N_718,In_317,In_469);
or U719 (N_719,In_38,In_288);
or U720 (N_720,In_360,In_257);
xnor U721 (N_721,In_427,In_74);
nor U722 (N_722,In_134,In_211);
and U723 (N_723,In_48,In_79);
or U724 (N_724,In_467,In_338);
nand U725 (N_725,In_406,In_18);
xor U726 (N_726,In_289,In_484);
or U727 (N_727,In_417,In_281);
xor U728 (N_728,In_223,In_413);
or U729 (N_729,In_210,In_316);
xor U730 (N_730,In_62,In_292);
and U731 (N_731,In_280,In_13);
or U732 (N_732,In_192,In_266);
xnor U733 (N_733,In_277,In_376);
and U734 (N_734,In_221,In_286);
nor U735 (N_735,In_30,In_440);
nand U736 (N_736,In_157,In_369);
nand U737 (N_737,In_5,In_352);
xnor U738 (N_738,In_160,In_36);
and U739 (N_739,In_367,In_70);
and U740 (N_740,In_367,In_212);
and U741 (N_741,In_488,In_194);
nand U742 (N_742,In_439,In_249);
nand U743 (N_743,In_328,In_20);
or U744 (N_744,In_198,In_329);
xor U745 (N_745,In_282,In_12);
xor U746 (N_746,In_103,In_499);
and U747 (N_747,In_356,In_266);
and U748 (N_748,In_152,In_22);
nand U749 (N_749,In_330,In_407);
nor U750 (N_750,In_108,In_112);
or U751 (N_751,In_467,In_136);
or U752 (N_752,In_462,In_92);
and U753 (N_753,In_29,In_437);
xnor U754 (N_754,In_400,In_287);
or U755 (N_755,In_62,In_112);
or U756 (N_756,In_140,In_165);
nor U757 (N_757,In_24,In_28);
nor U758 (N_758,In_312,In_76);
xor U759 (N_759,In_393,In_229);
and U760 (N_760,In_111,In_97);
xnor U761 (N_761,In_164,In_94);
nand U762 (N_762,In_458,In_147);
xor U763 (N_763,In_206,In_470);
or U764 (N_764,In_469,In_121);
nor U765 (N_765,In_368,In_7);
and U766 (N_766,In_175,In_83);
xor U767 (N_767,In_236,In_430);
and U768 (N_768,In_170,In_325);
or U769 (N_769,In_420,In_408);
and U770 (N_770,In_302,In_203);
or U771 (N_771,In_19,In_335);
or U772 (N_772,In_208,In_228);
xor U773 (N_773,In_13,In_399);
xnor U774 (N_774,In_420,In_56);
nor U775 (N_775,In_442,In_452);
xnor U776 (N_776,In_134,In_227);
xnor U777 (N_777,In_74,In_72);
nor U778 (N_778,In_109,In_148);
nor U779 (N_779,In_302,In_161);
and U780 (N_780,In_362,In_305);
xnor U781 (N_781,In_354,In_196);
or U782 (N_782,In_82,In_371);
and U783 (N_783,In_378,In_131);
nand U784 (N_784,In_32,In_367);
nor U785 (N_785,In_172,In_405);
nor U786 (N_786,In_431,In_194);
or U787 (N_787,In_314,In_293);
nand U788 (N_788,In_58,In_195);
nor U789 (N_789,In_62,In_58);
or U790 (N_790,In_401,In_257);
or U791 (N_791,In_298,In_345);
and U792 (N_792,In_228,In_25);
xor U793 (N_793,In_40,In_112);
nor U794 (N_794,In_183,In_351);
nor U795 (N_795,In_175,In_329);
or U796 (N_796,In_400,In_371);
and U797 (N_797,In_39,In_170);
or U798 (N_798,In_108,In_136);
nand U799 (N_799,In_259,In_495);
and U800 (N_800,In_404,In_265);
nor U801 (N_801,In_392,In_380);
xnor U802 (N_802,In_142,In_406);
nor U803 (N_803,In_124,In_300);
and U804 (N_804,In_380,In_294);
nor U805 (N_805,In_126,In_94);
xnor U806 (N_806,In_292,In_78);
and U807 (N_807,In_264,In_140);
xnor U808 (N_808,In_59,In_153);
xnor U809 (N_809,In_414,In_236);
xor U810 (N_810,In_2,In_407);
or U811 (N_811,In_401,In_190);
nor U812 (N_812,In_400,In_257);
nand U813 (N_813,In_190,In_224);
or U814 (N_814,In_43,In_488);
nor U815 (N_815,In_241,In_216);
and U816 (N_816,In_237,In_148);
nand U817 (N_817,In_329,In_185);
xor U818 (N_818,In_208,In_0);
nand U819 (N_819,In_79,In_438);
xnor U820 (N_820,In_496,In_485);
nand U821 (N_821,In_362,In_212);
nand U822 (N_822,In_25,In_183);
xor U823 (N_823,In_41,In_140);
nor U824 (N_824,In_68,In_158);
and U825 (N_825,In_486,In_344);
or U826 (N_826,In_432,In_153);
or U827 (N_827,In_463,In_250);
nand U828 (N_828,In_248,In_29);
or U829 (N_829,In_190,In_230);
or U830 (N_830,In_289,In_215);
nor U831 (N_831,In_46,In_209);
and U832 (N_832,In_142,In_336);
or U833 (N_833,In_323,In_166);
nand U834 (N_834,In_143,In_444);
nand U835 (N_835,In_436,In_356);
or U836 (N_836,In_454,In_133);
or U837 (N_837,In_119,In_243);
nand U838 (N_838,In_168,In_422);
xor U839 (N_839,In_355,In_338);
nor U840 (N_840,In_190,In_360);
or U841 (N_841,In_274,In_97);
or U842 (N_842,In_164,In_152);
xor U843 (N_843,In_335,In_229);
nand U844 (N_844,In_481,In_226);
nand U845 (N_845,In_441,In_89);
nand U846 (N_846,In_347,In_116);
or U847 (N_847,In_409,In_419);
xor U848 (N_848,In_373,In_312);
xnor U849 (N_849,In_177,In_17);
nor U850 (N_850,In_5,In_51);
xor U851 (N_851,In_184,In_477);
nand U852 (N_852,In_169,In_266);
nor U853 (N_853,In_171,In_275);
nor U854 (N_854,In_372,In_159);
nor U855 (N_855,In_490,In_495);
nor U856 (N_856,In_364,In_101);
nand U857 (N_857,In_153,In_351);
nor U858 (N_858,In_278,In_454);
xor U859 (N_859,In_86,In_327);
nand U860 (N_860,In_233,In_275);
nand U861 (N_861,In_309,In_57);
and U862 (N_862,In_164,In_268);
and U863 (N_863,In_325,In_430);
nand U864 (N_864,In_62,In_427);
and U865 (N_865,In_204,In_220);
and U866 (N_866,In_92,In_327);
xnor U867 (N_867,In_306,In_423);
xor U868 (N_868,In_433,In_398);
nor U869 (N_869,In_361,In_51);
and U870 (N_870,In_323,In_341);
or U871 (N_871,In_76,In_220);
nor U872 (N_872,In_292,In_420);
or U873 (N_873,In_293,In_58);
nor U874 (N_874,In_455,In_351);
nand U875 (N_875,In_447,In_464);
nor U876 (N_876,In_59,In_407);
and U877 (N_877,In_113,In_404);
xnor U878 (N_878,In_46,In_205);
nor U879 (N_879,In_79,In_237);
xnor U880 (N_880,In_42,In_189);
or U881 (N_881,In_250,In_328);
nand U882 (N_882,In_5,In_3);
or U883 (N_883,In_286,In_41);
xnor U884 (N_884,In_468,In_344);
nand U885 (N_885,In_321,In_403);
xor U886 (N_886,In_173,In_240);
nand U887 (N_887,In_241,In_159);
and U888 (N_888,In_218,In_336);
nand U889 (N_889,In_65,In_147);
nand U890 (N_890,In_216,In_149);
nand U891 (N_891,In_411,In_349);
or U892 (N_892,In_378,In_394);
and U893 (N_893,In_106,In_11);
nor U894 (N_894,In_423,In_11);
or U895 (N_895,In_379,In_42);
nor U896 (N_896,In_340,In_318);
and U897 (N_897,In_427,In_356);
xnor U898 (N_898,In_133,In_399);
xnor U899 (N_899,In_361,In_473);
nand U900 (N_900,In_128,In_274);
nor U901 (N_901,In_131,In_201);
nor U902 (N_902,In_309,In_383);
and U903 (N_903,In_307,In_14);
nor U904 (N_904,In_305,In_492);
xor U905 (N_905,In_226,In_479);
nor U906 (N_906,In_345,In_45);
and U907 (N_907,In_253,In_395);
and U908 (N_908,In_304,In_215);
nor U909 (N_909,In_183,In_315);
xnor U910 (N_910,In_441,In_317);
nand U911 (N_911,In_371,In_223);
nand U912 (N_912,In_234,In_416);
nor U913 (N_913,In_119,In_277);
nand U914 (N_914,In_459,In_420);
and U915 (N_915,In_235,In_245);
or U916 (N_916,In_497,In_449);
and U917 (N_917,In_289,In_28);
and U918 (N_918,In_258,In_397);
xnor U919 (N_919,In_447,In_340);
or U920 (N_920,In_444,In_72);
nor U921 (N_921,In_74,In_140);
nor U922 (N_922,In_322,In_294);
or U923 (N_923,In_341,In_372);
and U924 (N_924,In_269,In_47);
nand U925 (N_925,In_346,In_256);
and U926 (N_926,In_319,In_94);
nor U927 (N_927,In_249,In_250);
or U928 (N_928,In_353,In_396);
xor U929 (N_929,In_111,In_409);
nor U930 (N_930,In_18,In_322);
and U931 (N_931,In_105,In_207);
and U932 (N_932,In_205,In_96);
nor U933 (N_933,In_114,In_14);
or U934 (N_934,In_480,In_297);
or U935 (N_935,In_222,In_227);
and U936 (N_936,In_480,In_111);
and U937 (N_937,In_136,In_368);
nand U938 (N_938,In_126,In_165);
nor U939 (N_939,In_428,In_388);
and U940 (N_940,In_417,In_388);
nor U941 (N_941,In_55,In_382);
or U942 (N_942,In_386,In_183);
and U943 (N_943,In_3,In_359);
nand U944 (N_944,In_3,In_240);
xnor U945 (N_945,In_63,In_171);
xnor U946 (N_946,In_65,In_195);
nand U947 (N_947,In_450,In_93);
or U948 (N_948,In_432,In_18);
nor U949 (N_949,In_184,In_319);
and U950 (N_950,In_2,In_209);
nor U951 (N_951,In_35,In_464);
nor U952 (N_952,In_375,In_114);
nand U953 (N_953,In_184,In_103);
nor U954 (N_954,In_220,In_26);
and U955 (N_955,In_496,In_255);
xor U956 (N_956,In_7,In_40);
nor U957 (N_957,In_183,In_337);
or U958 (N_958,In_426,In_410);
nor U959 (N_959,In_86,In_201);
nand U960 (N_960,In_365,In_8);
and U961 (N_961,In_317,In_141);
nand U962 (N_962,In_224,In_302);
or U963 (N_963,In_39,In_461);
xnor U964 (N_964,In_454,In_126);
or U965 (N_965,In_259,In_125);
and U966 (N_966,In_205,In_141);
and U967 (N_967,In_8,In_377);
xnor U968 (N_968,In_265,In_104);
and U969 (N_969,In_17,In_65);
and U970 (N_970,In_139,In_30);
and U971 (N_971,In_431,In_64);
or U972 (N_972,In_264,In_253);
or U973 (N_973,In_50,In_35);
or U974 (N_974,In_72,In_389);
xor U975 (N_975,In_251,In_400);
nor U976 (N_976,In_31,In_330);
nor U977 (N_977,In_352,In_445);
xnor U978 (N_978,In_195,In_312);
and U979 (N_979,In_434,In_291);
nand U980 (N_980,In_477,In_423);
and U981 (N_981,In_60,In_451);
and U982 (N_982,In_176,In_321);
or U983 (N_983,In_402,In_186);
nor U984 (N_984,In_207,In_75);
or U985 (N_985,In_324,In_164);
nand U986 (N_986,In_340,In_301);
xnor U987 (N_987,In_383,In_487);
nand U988 (N_988,In_252,In_392);
nand U989 (N_989,In_215,In_439);
and U990 (N_990,In_437,In_352);
or U991 (N_991,In_402,In_54);
nand U992 (N_992,In_480,In_8);
or U993 (N_993,In_92,In_455);
or U994 (N_994,In_49,In_118);
nand U995 (N_995,In_335,In_148);
nand U996 (N_996,In_76,In_337);
xnor U997 (N_997,In_112,In_472);
and U998 (N_998,In_97,In_244);
nor U999 (N_999,In_458,In_295);
nand U1000 (N_1000,N_945,N_307);
nor U1001 (N_1001,N_28,N_296);
nand U1002 (N_1002,N_348,N_255);
nand U1003 (N_1003,N_525,N_57);
xor U1004 (N_1004,N_672,N_333);
xnor U1005 (N_1005,N_218,N_682);
or U1006 (N_1006,N_852,N_631);
nand U1007 (N_1007,N_85,N_858);
or U1008 (N_1008,N_980,N_961);
xnor U1009 (N_1009,N_718,N_179);
xor U1010 (N_1010,N_287,N_897);
nor U1011 (N_1011,N_605,N_160);
nor U1012 (N_1012,N_840,N_647);
or U1013 (N_1013,N_502,N_624);
xor U1014 (N_1014,N_51,N_925);
and U1015 (N_1015,N_668,N_708);
and U1016 (N_1016,N_377,N_974);
nor U1017 (N_1017,N_664,N_954);
nor U1018 (N_1018,N_913,N_893);
xor U1019 (N_1019,N_448,N_723);
xor U1020 (N_1020,N_544,N_40);
nand U1021 (N_1021,N_338,N_120);
nand U1022 (N_1022,N_522,N_595);
nor U1023 (N_1023,N_275,N_78);
or U1024 (N_1024,N_152,N_282);
xnor U1025 (N_1025,N_562,N_217);
nand U1026 (N_1026,N_311,N_417);
and U1027 (N_1027,N_48,N_155);
nand U1028 (N_1028,N_13,N_79);
or U1029 (N_1029,N_905,N_839);
xnor U1030 (N_1030,N_995,N_910);
nand U1031 (N_1031,N_540,N_446);
xor U1032 (N_1032,N_583,N_104);
nand U1033 (N_1033,N_399,N_439);
and U1034 (N_1034,N_342,N_259);
or U1035 (N_1035,N_742,N_687);
nor U1036 (N_1036,N_126,N_843);
nor U1037 (N_1037,N_942,N_329);
or U1038 (N_1038,N_151,N_731);
nand U1039 (N_1039,N_716,N_875);
xnor U1040 (N_1040,N_855,N_239);
or U1041 (N_1041,N_350,N_321);
nor U1042 (N_1042,N_557,N_187);
or U1043 (N_1043,N_89,N_570);
or U1044 (N_1044,N_582,N_988);
or U1045 (N_1045,N_52,N_827);
xor U1046 (N_1046,N_382,N_242);
xor U1047 (N_1047,N_671,N_116);
nand U1048 (N_1048,N_632,N_435);
or U1049 (N_1049,N_128,N_186);
and U1050 (N_1050,N_495,N_757);
xor U1051 (N_1051,N_626,N_467);
or U1052 (N_1052,N_358,N_931);
xnor U1053 (N_1053,N_712,N_533);
nand U1054 (N_1054,N_824,N_394);
nand U1055 (N_1055,N_33,N_704);
or U1056 (N_1056,N_740,N_414);
and U1057 (N_1057,N_825,N_418);
or U1058 (N_1058,N_387,N_136);
nor U1059 (N_1059,N_654,N_482);
or U1060 (N_1060,N_21,N_328);
xor U1061 (N_1061,N_987,N_706);
nor U1062 (N_1062,N_971,N_106);
nor U1063 (N_1063,N_376,N_617);
nand U1064 (N_1064,N_650,N_593);
nand U1065 (N_1065,N_304,N_235);
or U1066 (N_1066,N_696,N_741);
or U1067 (N_1067,N_277,N_792);
and U1068 (N_1068,N_949,N_31);
nor U1069 (N_1069,N_972,N_2);
or U1070 (N_1070,N_395,N_123);
and U1071 (N_1071,N_319,N_604);
or U1072 (N_1072,N_880,N_280);
xor U1073 (N_1073,N_519,N_503);
nor U1074 (N_1074,N_977,N_653);
or U1075 (N_1075,N_762,N_561);
nand U1076 (N_1076,N_144,N_734);
or U1077 (N_1077,N_895,N_676);
xor U1078 (N_1078,N_845,N_941);
and U1079 (N_1079,N_80,N_20);
or U1080 (N_1080,N_699,N_178);
nor U1081 (N_1081,N_442,N_543);
xnor U1082 (N_1082,N_669,N_229);
nand U1083 (N_1083,N_787,N_226);
and U1084 (N_1084,N_766,N_252);
nor U1085 (N_1085,N_428,N_231);
and U1086 (N_1086,N_0,N_15);
xnor U1087 (N_1087,N_985,N_420);
and U1088 (N_1088,N_526,N_142);
nand U1089 (N_1089,N_565,N_691);
xnor U1090 (N_1090,N_459,N_819);
xnor U1091 (N_1091,N_665,N_63);
and U1092 (N_1092,N_135,N_683);
xnor U1093 (N_1093,N_585,N_460);
or U1094 (N_1094,N_685,N_550);
or U1095 (N_1095,N_59,N_68);
or U1096 (N_1096,N_962,N_641);
or U1097 (N_1097,N_602,N_894);
or U1098 (N_1098,N_814,N_363);
xor U1099 (N_1099,N_554,N_84);
or U1100 (N_1100,N_464,N_714);
nand U1101 (N_1101,N_125,N_938);
and U1102 (N_1102,N_891,N_421);
and U1103 (N_1103,N_37,N_438);
nand U1104 (N_1104,N_310,N_536);
xnor U1105 (N_1105,N_161,N_574);
nand U1106 (N_1106,N_474,N_838);
and U1107 (N_1107,N_518,N_705);
xor U1108 (N_1108,N_462,N_23);
xnor U1109 (N_1109,N_403,N_480);
xor U1110 (N_1110,N_269,N_968);
xor U1111 (N_1111,N_429,N_586);
nand U1112 (N_1112,N_223,N_378);
nand U1113 (N_1113,N_517,N_274);
nand U1114 (N_1114,N_456,N_608);
xnor U1115 (N_1115,N_288,N_956);
xor U1116 (N_1116,N_778,N_272);
or U1117 (N_1117,N_302,N_933);
nor U1118 (N_1118,N_204,N_717);
nor U1119 (N_1119,N_208,N_849);
xor U1120 (N_1120,N_681,N_733);
xor U1121 (N_1121,N_896,N_802);
and U1122 (N_1122,N_69,N_334);
and U1123 (N_1123,N_870,N_422);
nor U1124 (N_1124,N_86,N_915);
nand U1125 (N_1125,N_391,N_828);
and U1126 (N_1126,N_514,N_473);
xor U1127 (N_1127,N_332,N_424);
and U1128 (N_1128,N_447,N_864);
and U1129 (N_1129,N_297,N_984);
xnor U1130 (N_1130,N_633,N_240);
nor U1131 (N_1131,N_575,N_39);
xnor U1132 (N_1132,N_983,N_188);
and U1133 (N_1133,N_901,N_598);
and U1134 (N_1134,N_657,N_236);
xor U1135 (N_1135,N_746,N_344);
or U1136 (N_1136,N_597,N_196);
xnor U1137 (N_1137,N_744,N_49);
or U1138 (N_1138,N_96,N_710);
and U1139 (N_1139,N_673,N_207);
xnor U1140 (N_1140,N_258,N_851);
or U1141 (N_1141,N_817,N_871);
and U1142 (N_1142,N_92,N_472);
and U1143 (N_1143,N_400,N_779);
nor U1144 (N_1144,N_552,N_553);
and U1145 (N_1145,N_628,N_791);
nand U1146 (N_1146,N_56,N_754);
or U1147 (N_1147,N_539,N_782);
and U1148 (N_1148,N_73,N_939);
or U1149 (N_1149,N_684,N_469);
and U1150 (N_1150,N_584,N_764);
xor U1151 (N_1151,N_100,N_692);
or U1152 (N_1152,N_773,N_789);
xnor U1153 (N_1153,N_923,N_173);
nand U1154 (N_1154,N_351,N_959);
nor U1155 (N_1155,N_786,N_580);
or U1156 (N_1156,N_103,N_195);
xor U1157 (N_1157,N_232,N_709);
nand U1158 (N_1158,N_529,N_268);
nor U1159 (N_1159,N_308,N_730);
nor U1160 (N_1160,N_753,N_879);
xnor U1161 (N_1161,N_569,N_406);
nand U1162 (N_1162,N_166,N_499);
xnor U1163 (N_1163,N_261,N_674);
nor U1164 (N_1164,N_803,N_504);
nor U1165 (N_1165,N_955,N_212);
xor U1166 (N_1166,N_171,N_892);
and U1167 (N_1167,N_200,N_981);
or U1168 (N_1168,N_32,N_774);
nor U1169 (N_1169,N_121,N_369);
or U1170 (N_1170,N_283,N_105);
and U1171 (N_1171,N_132,N_156);
xor U1172 (N_1172,N_112,N_12);
nor U1173 (N_1173,N_868,N_450);
or U1174 (N_1174,N_246,N_784);
or U1175 (N_1175,N_620,N_325);
nand U1176 (N_1176,N_413,N_867);
nor U1177 (N_1177,N_800,N_603);
and U1178 (N_1178,N_22,N_410);
xor U1179 (N_1179,N_976,N_199);
nor U1180 (N_1180,N_114,N_113);
nor U1181 (N_1181,N_262,N_943);
nor U1182 (N_1182,N_181,N_159);
nand U1183 (N_1183,N_630,N_430);
nor U1184 (N_1184,N_541,N_70);
xor U1185 (N_1185,N_621,N_122);
xor U1186 (N_1186,N_281,N_381);
nand U1187 (N_1187,N_238,N_524);
xnor U1188 (N_1188,N_759,N_36);
xnor U1189 (N_1189,N_45,N_154);
and U1190 (N_1190,N_549,N_614);
and U1191 (N_1191,N_625,N_370);
or U1192 (N_1192,N_990,N_91);
nor U1193 (N_1193,N_737,N_916);
nor U1194 (N_1194,N_129,N_433);
nor U1195 (N_1195,N_373,N_935);
nor U1196 (N_1196,N_865,N_443);
nor U1197 (N_1197,N_809,N_776);
and U1198 (N_1198,N_876,N_578);
or U1199 (N_1199,N_516,N_861);
xnor U1200 (N_1200,N_563,N_266);
nor U1201 (N_1201,N_306,N_224);
or U1202 (N_1202,N_965,N_627);
or U1203 (N_1203,N_646,N_873);
xnor U1204 (N_1204,N_798,N_975);
and U1205 (N_1205,N_911,N_639);
nand U1206 (N_1206,N_997,N_374);
nor U1207 (N_1207,N_610,N_793);
xnor U1208 (N_1208,N_835,N_451);
nor U1209 (N_1209,N_313,N_457);
and U1210 (N_1210,N_643,N_54);
or U1211 (N_1211,N_425,N_361);
xnor U1212 (N_1212,N_375,N_137);
or U1213 (N_1213,N_176,N_427);
xnor U1214 (N_1214,N_476,N_149);
nand U1215 (N_1215,N_559,N_906);
nor U1216 (N_1216,N_366,N_886);
and U1217 (N_1217,N_512,N_41);
nor U1218 (N_1218,N_315,N_645);
nor U1219 (N_1219,N_950,N_483);
nor U1220 (N_1220,N_359,N_728);
nand U1221 (N_1221,N_201,N_286);
nand U1222 (N_1222,N_108,N_326);
nor U1223 (N_1223,N_478,N_209);
xor U1224 (N_1224,N_379,N_276);
or U1225 (N_1225,N_158,N_253);
nand U1226 (N_1226,N_888,N_978);
nand U1227 (N_1227,N_532,N_528);
and U1228 (N_1228,N_926,N_648);
nand U1229 (N_1229,N_183,N_772);
or U1230 (N_1230,N_924,N_211);
nor U1231 (N_1231,N_993,N_656);
nor U1232 (N_1232,N_497,N_545);
and U1233 (N_1233,N_747,N_316);
and U1234 (N_1234,N_944,N_619);
xor U1235 (N_1235,N_175,N_330);
nor U1236 (N_1236,N_47,N_383);
xor U1237 (N_1237,N_95,N_177);
nand U1238 (N_1238,N_479,N_862);
xnor U1239 (N_1239,N_635,N_899);
or U1240 (N_1240,N_752,N_119);
or U1241 (N_1241,N_659,N_58);
xor U1242 (N_1242,N_715,N_243);
nor U1243 (N_1243,N_572,N_324);
nor U1244 (N_1244,N_440,N_700);
nand U1245 (N_1245,N_638,N_842);
xnor U1246 (N_1246,N_146,N_542);
nor U1247 (N_1247,N_402,N_419);
nand U1248 (N_1248,N_994,N_408);
or U1249 (N_1249,N_165,N_898);
nand U1250 (N_1250,N_719,N_436);
and U1251 (N_1251,N_341,N_761);
or U1252 (N_1252,N_206,N_343);
xor U1253 (N_1253,N_571,N_535);
or U1254 (N_1254,N_885,N_616);
nor U1255 (N_1255,N_477,N_735);
or U1256 (N_1256,N_750,N_481);
and U1257 (N_1257,N_856,N_127);
and U1258 (N_1258,N_301,N_854);
xor U1259 (N_1259,N_725,N_812);
and U1260 (N_1260,N_180,N_568);
nor U1261 (N_1261,N_748,N_292);
nand U1262 (N_1262,N_853,N_857);
nand U1263 (N_1263,N_458,N_928);
nor U1264 (N_1264,N_29,N_927);
xor U1265 (N_1265,N_680,N_966);
xor U1266 (N_1266,N_210,N_601);
and U1267 (N_1267,N_948,N_808);
nor U1268 (N_1268,N_312,N_290);
nor U1269 (N_1269,N_19,N_556);
nand U1270 (N_1270,N_694,N_111);
nand U1271 (N_1271,N_203,N_256);
nor U1272 (N_1272,N_567,N_743);
and U1273 (N_1273,N_498,N_887);
nand U1274 (N_1274,N_958,N_577);
nor U1275 (N_1275,N_153,N_139);
or U1276 (N_1276,N_768,N_751);
nand U1277 (N_1277,N_71,N_546);
nor U1278 (N_1278,N_174,N_437);
or U1279 (N_1279,N_279,N_141);
xor U1280 (N_1280,N_763,N_506);
and U1281 (N_1281,N_547,N_555);
xnor U1282 (N_1282,N_10,N_415);
nand U1283 (N_1283,N_220,N_331);
and U1284 (N_1284,N_140,N_703);
xor U1285 (N_1285,N_385,N_147);
and U1286 (N_1286,N_38,N_726);
nor U1287 (N_1287,N_689,N_225);
nor U1288 (N_1288,N_515,N_340);
nor U1289 (N_1289,N_531,N_769);
nor U1290 (N_1290,N_805,N_693);
xor U1291 (N_1291,N_431,N_110);
xor U1292 (N_1292,N_986,N_783);
nor U1293 (N_1293,N_736,N_432);
nor U1294 (N_1294,N_903,N_520);
xor U1295 (N_1295,N_788,N_833);
nand U1296 (N_1296,N_914,N_991);
nor U1297 (N_1297,N_722,N_882);
xor U1298 (N_1298,N_576,N_816);
and U1299 (N_1299,N_521,N_309);
and U1300 (N_1300,N_27,N_507);
nor U1301 (N_1301,N_335,N_530);
nor U1302 (N_1302,N_488,N_866);
and U1303 (N_1303,N_198,N_831);
nand U1304 (N_1304,N_953,N_219);
or U1305 (N_1305,N_613,N_505);
and U1306 (N_1306,N_162,N_690);
nor U1307 (N_1307,N_401,N_946);
nand U1308 (N_1308,N_493,N_794);
and U1309 (N_1309,N_72,N_591);
or U1310 (N_1310,N_169,N_285);
nor U1311 (N_1311,N_454,N_444);
xnor U1312 (N_1312,N_213,N_337);
nand U1313 (N_1313,N_182,N_202);
and U1314 (N_1314,N_347,N_471);
xnor U1315 (N_1315,N_53,N_234);
nor U1316 (N_1316,N_947,N_797);
nand U1317 (N_1317,N_724,N_799);
or U1318 (N_1318,N_560,N_1);
or U1319 (N_1319,N_729,N_8);
nor U1320 (N_1320,N_491,N_339);
or U1321 (N_1321,N_216,N_964);
and U1322 (N_1322,N_907,N_660);
nor U1323 (N_1323,N_960,N_42);
or U1324 (N_1324,N_83,N_581);
nand U1325 (N_1325,N_936,N_695);
nor U1326 (N_1326,N_661,N_929);
nor U1327 (N_1327,N_996,N_228);
nand U1328 (N_1328,N_484,N_951);
or U1329 (N_1329,N_273,N_969);
xnor U1330 (N_1330,N_396,N_257);
or U1331 (N_1331,N_859,N_801);
or U1332 (N_1332,N_131,N_409);
xnor U1333 (N_1333,N_623,N_404);
and U1334 (N_1334,N_35,N_249);
or U1335 (N_1335,N_434,N_461);
and U1336 (N_1336,N_465,N_815);
and U1337 (N_1337,N_323,N_636);
xnor U1338 (N_1338,N_999,N_470);
and U1339 (N_1339,N_368,N_150);
and U1340 (N_1340,N_922,N_489);
and U1341 (N_1341,N_662,N_806);
or U1342 (N_1342,N_713,N_599);
nand U1343 (N_1343,N_6,N_205);
xnor U1344 (N_1344,N_98,N_398);
nand U1345 (N_1345,N_711,N_566);
xnor U1346 (N_1346,N_18,N_117);
xnor U1347 (N_1347,N_970,N_115);
or U1348 (N_1348,N_293,N_829);
nand U1349 (N_1349,N_14,N_168);
and U1350 (N_1350,N_185,N_362);
nor U1351 (N_1351,N_93,N_670);
nand U1352 (N_1352,N_237,N_284);
or U1353 (N_1353,N_908,N_492);
xnor U1354 (N_1354,N_508,N_322);
or U1355 (N_1355,N_775,N_538);
nor U1356 (N_1356,N_392,N_919);
xor U1357 (N_1357,N_634,N_832);
nor U1358 (N_1358,N_148,N_157);
nor U1359 (N_1359,N_822,N_130);
nand U1360 (N_1360,N_644,N_836);
and U1361 (N_1361,N_590,N_606);
xnor U1362 (N_1362,N_371,N_609);
xor U1363 (N_1363,N_967,N_221);
xnor U1364 (N_1364,N_732,N_318);
nand U1365 (N_1365,N_874,N_412);
or U1366 (N_1366,N_386,N_755);
and U1367 (N_1367,N_918,N_989);
or U1368 (N_1368,N_17,N_558);
or U1369 (N_1369,N_940,N_527);
and U1370 (N_1370,N_998,N_739);
and U1371 (N_1371,N_46,N_878);
xnor U1372 (N_1372,N_87,N_118);
xor U1373 (N_1373,N_837,N_449);
nand U1374 (N_1374,N_16,N_55);
nand U1375 (N_1375,N_600,N_615);
and U1376 (N_1376,N_767,N_76);
xor U1377 (N_1377,N_61,N_75);
nand U1378 (N_1378,N_134,N_50);
and U1379 (N_1379,N_170,N_364);
nand U1380 (N_1380,N_263,N_26);
or U1381 (N_1381,N_510,N_222);
xnor U1382 (N_1382,N_124,N_534);
xor U1383 (N_1383,N_830,N_548);
and U1384 (N_1384,N_889,N_345);
or U1385 (N_1385,N_780,N_902);
xnor U1386 (N_1386,N_320,N_230);
or U1387 (N_1387,N_64,N_702);
and U1388 (N_1388,N_405,N_81);
nand U1389 (N_1389,N_640,N_883);
xor U1390 (N_1390,N_270,N_327);
and U1391 (N_1391,N_138,N_189);
and U1392 (N_1392,N_679,N_245);
xnor U1393 (N_1393,N_807,N_172);
nor U1394 (N_1394,N_790,N_133);
xor U1395 (N_1395,N_357,N_785);
nand U1396 (N_1396,N_197,N_74);
xnor U1397 (N_1397,N_88,N_869);
xor U1398 (N_1398,N_770,N_513);
nand U1399 (N_1399,N_537,N_190);
or U1400 (N_1400,N_367,N_511);
and U1401 (N_1401,N_771,N_912);
xnor U1402 (N_1402,N_611,N_300);
nand U1403 (N_1403,N_612,N_777);
or U1404 (N_1404,N_551,N_760);
xor U1405 (N_1405,N_490,N_265);
nand U1406 (N_1406,N_241,N_658);
and U1407 (N_1407,N_982,N_847);
nand U1408 (N_1408,N_445,N_486);
or U1409 (N_1409,N_360,N_194);
xnor U1410 (N_1410,N_67,N_500);
or U1411 (N_1411,N_846,N_592);
xor U1412 (N_1412,N_917,N_60);
xnor U1413 (N_1413,N_564,N_291);
nand U1414 (N_1414,N_192,N_463);
nand U1415 (N_1415,N_365,N_678);
or U1416 (N_1416,N_952,N_475);
nand U1417 (N_1417,N_30,N_305);
nand U1418 (N_1418,N_423,N_353);
nor U1419 (N_1419,N_109,N_251);
nand U1420 (N_1420,N_810,N_884);
and U1421 (N_1421,N_494,N_573);
and U1422 (N_1422,N_248,N_11);
nor U1423 (N_1423,N_94,N_663);
nor U1424 (N_1424,N_594,N_43);
or U1425 (N_1425,N_820,N_452);
nand U1426 (N_1426,N_3,N_841);
nor U1427 (N_1427,N_143,N_9);
xnor U1428 (N_1428,N_407,N_466);
and U1429 (N_1429,N_727,N_82);
and U1430 (N_1430,N_688,N_749);
xor U1431 (N_1431,N_649,N_745);
and U1432 (N_1432,N_992,N_215);
or U1433 (N_1433,N_468,N_487);
xor U1434 (N_1434,N_356,N_411);
and U1435 (N_1435,N_655,N_588);
xnor U1436 (N_1436,N_298,N_637);
and U1437 (N_1437,N_804,N_314);
and U1438 (N_1438,N_101,N_813);
or U1439 (N_1439,N_107,N_686);
nor U1440 (N_1440,N_349,N_397);
xnor U1441 (N_1441,N_227,N_920);
and U1442 (N_1442,N_65,N_4);
and U1443 (N_1443,N_675,N_7);
nor U1444 (N_1444,N_163,N_393);
nand U1445 (N_1445,N_247,N_622);
or U1446 (N_1446,N_34,N_289);
xor U1447 (N_1447,N_795,N_677);
xnor U1448 (N_1448,N_589,N_271);
and U1449 (N_1449,N_388,N_441);
xor U1450 (N_1450,N_264,N_295);
and U1451 (N_1451,N_317,N_877);
and U1452 (N_1452,N_167,N_250);
nand U1453 (N_1453,N_25,N_629);
and U1454 (N_1454,N_453,N_701);
nor U1455 (N_1455,N_666,N_848);
or U1456 (N_1456,N_587,N_24);
xnor U1457 (N_1457,N_909,N_90);
nor U1458 (N_1458,N_697,N_720);
nand U1459 (N_1459,N_233,N_834);
and U1460 (N_1460,N_900,N_579);
nor U1461 (N_1461,N_826,N_721);
and U1462 (N_1462,N_652,N_485);
nand U1463 (N_1463,N_145,N_979);
or U1464 (N_1464,N_352,N_818);
and U1465 (N_1465,N_642,N_509);
or U1466 (N_1466,N_850,N_765);
xnor U1467 (N_1467,N_607,N_164);
nand U1468 (N_1468,N_355,N_934);
nor U1469 (N_1469,N_667,N_380);
xor U1470 (N_1470,N_890,N_930);
and U1471 (N_1471,N_390,N_973);
nor U1472 (N_1472,N_426,N_99);
xor U1473 (N_1473,N_758,N_596);
nand U1474 (N_1474,N_294,N_863);
or U1475 (N_1475,N_254,N_354);
and U1476 (N_1476,N_5,N_389);
or U1477 (N_1477,N_738,N_821);
or U1478 (N_1478,N_872,N_336);
xnor U1479 (N_1479,N_904,N_651);
nand U1480 (N_1480,N_618,N_191);
or U1481 (N_1481,N_193,N_963);
and U1482 (N_1482,N_102,N_844);
nor U1483 (N_1483,N_455,N_932);
or U1484 (N_1484,N_781,N_303);
nor U1485 (N_1485,N_44,N_707);
nor U1486 (N_1486,N_260,N_957);
xnor U1487 (N_1487,N_756,N_823);
and U1488 (N_1488,N_523,N_937);
nand U1489 (N_1489,N_77,N_184);
nand U1490 (N_1490,N_921,N_811);
nor U1491 (N_1491,N_416,N_97);
and U1492 (N_1492,N_299,N_384);
nand U1493 (N_1493,N_796,N_501);
nor U1494 (N_1494,N_881,N_66);
or U1495 (N_1495,N_214,N_346);
nor U1496 (N_1496,N_267,N_698);
nor U1497 (N_1497,N_496,N_860);
or U1498 (N_1498,N_372,N_278);
nand U1499 (N_1499,N_244,N_62);
nand U1500 (N_1500,N_876,N_574);
or U1501 (N_1501,N_129,N_793);
nand U1502 (N_1502,N_18,N_58);
or U1503 (N_1503,N_919,N_875);
and U1504 (N_1504,N_913,N_543);
nor U1505 (N_1505,N_553,N_707);
xnor U1506 (N_1506,N_908,N_751);
or U1507 (N_1507,N_158,N_583);
or U1508 (N_1508,N_982,N_493);
nor U1509 (N_1509,N_110,N_427);
or U1510 (N_1510,N_304,N_232);
or U1511 (N_1511,N_106,N_176);
nand U1512 (N_1512,N_260,N_87);
nor U1513 (N_1513,N_637,N_279);
or U1514 (N_1514,N_448,N_411);
and U1515 (N_1515,N_277,N_660);
nand U1516 (N_1516,N_659,N_344);
and U1517 (N_1517,N_430,N_979);
xor U1518 (N_1518,N_643,N_321);
or U1519 (N_1519,N_917,N_200);
nor U1520 (N_1520,N_405,N_807);
nand U1521 (N_1521,N_424,N_706);
nor U1522 (N_1522,N_225,N_832);
nand U1523 (N_1523,N_731,N_297);
nor U1524 (N_1524,N_398,N_415);
or U1525 (N_1525,N_858,N_544);
or U1526 (N_1526,N_604,N_614);
xnor U1527 (N_1527,N_702,N_495);
or U1528 (N_1528,N_26,N_455);
and U1529 (N_1529,N_166,N_611);
nor U1530 (N_1530,N_733,N_192);
xnor U1531 (N_1531,N_554,N_324);
or U1532 (N_1532,N_99,N_289);
nor U1533 (N_1533,N_28,N_902);
or U1534 (N_1534,N_521,N_86);
xnor U1535 (N_1535,N_613,N_160);
and U1536 (N_1536,N_94,N_487);
or U1537 (N_1537,N_634,N_585);
nand U1538 (N_1538,N_377,N_547);
or U1539 (N_1539,N_878,N_785);
or U1540 (N_1540,N_164,N_33);
xor U1541 (N_1541,N_676,N_667);
or U1542 (N_1542,N_705,N_212);
nor U1543 (N_1543,N_934,N_107);
xor U1544 (N_1544,N_580,N_301);
or U1545 (N_1545,N_73,N_186);
and U1546 (N_1546,N_822,N_819);
or U1547 (N_1547,N_223,N_887);
nor U1548 (N_1548,N_666,N_163);
nand U1549 (N_1549,N_169,N_905);
nor U1550 (N_1550,N_309,N_218);
xor U1551 (N_1551,N_918,N_607);
nor U1552 (N_1552,N_48,N_296);
xnor U1553 (N_1553,N_207,N_321);
nor U1554 (N_1554,N_161,N_200);
and U1555 (N_1555,N_67,N_245);
and U1556 (N_1556,N_424,N_810);
and U1557 (N_1557,N_296,N_9);
nor U1558 (N_1558,N_586,N_478);
nor U1559 (N_1559,N_681,N_334);
and U1560 (N_1560,N_28,N_914);
xor U1561 (N_1561,N_70,N_54);
xor U1562 (N_1562,N_317,N_327);
xnor U1563 (N_1563,N_652,N_158);
and U1564 (N_1564,N_32,N_472);
or U1565 (N_1565,N_378,N_46);
or U1566 (N_1566,N_980,N_351);
nand U1567 (N_1567,N_895,N_816);
nand U1568 (N_1568,N_105,N_888);
nor U1569 (N_1569,N_877,N_464);
xor U1570 (N_1570,N_132,N_557);
or U1571 (N_1571,N_875,N_663);
and U1572 (N_1572,N_269,N_781);
nand U1573 (N_1573,N_234,N_15);
xnor U1574 (N_1574,N_417,N_957);
nor U1575 (N_1575,N_62,N_341);
and U1576 (N_1576,N_324,N_75);
nand U1577 (N_1577,N_112,N_217);
and U1578 (N_1578,N_149,N_671);
and U1579 (N_1579,N_579,N_991);
xnor U1580 (N_1580,N_632,N_284);
nand U1581 (N_1581,N_145,N_941);
or U1582 (N_1582,N_81,N_482);
nand U1583 (N_1583,N_388,N_513);
and U1584 (N_1584,N_819,N_20);
xor U1585 (N_1585,N_940,N_916);
nor U1586 (N_1586,N_712,N_524);
nand U1587 (N_1587,N_276,N_95);
or U1588 (N_1588,N_375,N_955);
xor U1589 (N_1589,N_726,N_990);
xnor U1590 (N_1590,N_620,N_254);
nand U1591 (N_1591,N_173,N_94);
and U1592 (N_1592,N_156,N_727);
or U1593 (N_1593,N_121,N_698);
or U1594 (N_1594,N_548,N_167);
or U1595 (N_1595,N_446,N_104);
nand U1596 (N_1596,N_786,N_808);
nand U1597 (N_1597,N_845,N_719);
xnor U1598 (N_1598,N_707,N_645);
and U1599 (N_1599,N_389,N_654);
nor U1600 (N_1600,N_142,N_753);
and U1601 (N_1601,N_74,N_417);
or U1602 (N_1602,N_839,N_402);
and U1603 (N_1603,N_914,N_241);
xnor U1604 (N_1604,N_633,N_107);
and U1605 (N_1605,N_625,N_423);
nand U1606 (N_1606,N_692,N_376);
xor U1607 (N_1607,N_788,N_166);
nor U1608 (N_1608,N_341,N_319);
xor U1609 (N_1609,N_873,N_973);
xnor U1610 (N_1610,N_646,N_925);
nor U1611 (N_1611,N_546,N_144);
or U1612 (N_1612,N_305,N_619);
xnor U1613 (N_1613,N_943,N_996);
xnor U1614 (N_1614,N_373,N_943);
and U1615 (N_1615,N_19,N_264);
and U1616 (N_1616,N_287,N_378);
nand U1617 (N_1617,N_484,N_588);
or U1618 (N_1618,N_51,N_503);
and U1619 (N_1619,N_262,N_936);
and U1620 (N_1620,N_424,N_159);
nand U1621 (N_1621,N_584,N_629);
and U1622 (N_1622,N_175,N_917);
or U1623 (N_1623,N_571,N_638);
and U1624 (N_1624,N_274,N_939);
and U1625 (N_1625,N_408,N_698);
or U1626 (N_1626,N_510,N_290);
or U1627 (N_1627,N_357,N_460);
nor U1628 (N_1628,N_833,N_341);
xnor U1629 (N_1629,N_535,N_440);
or U1630 (N_1630,N_463,N_541);
xnor U1631 (N_1631,N_759,N_938);
and U1632 (N_1632,N_697,N_375);
nand U1633 (N_1633,N_863,N_465);
nor U1634 (N_1634,N_134,N_290);
nor U1635 (N_1635,N_481,N_792);
xor U1636 (N_1636,N_873,N_663);
or U1637 (N_1637,N_787,N_336);
nand U1638 (N_1638,N_545,N_232);
xnor U1639 (N_1639,N_375,N_925);
or U1640 (N_1640,N_32,N_81);
and U1641 (N_1641,N_896,N_278);
or U1642 (N_1642,N_320,N_180);
nor U1643 (N_1643,N_938,N_62);
and U1644 (N_1644,N_662,N_884);
and U1645 (N_1645,N_415,N_399);
or U1646 (N_1646,N_399,N_133);
or U1647 (N_1647,N_631,N_412);
and U1648 (N_1648,N_906,N_771);
xnor U1649 (N_1649,N_978,N_541);
and U1650 (N_1650,N_461,N_169);
xor U1651 (N_1651,N_151,N_164);
nor U1652 (N_1652,N_225,N_142);
or U1653 (N_1653,N_902,N_661);
nor U1654 (N_1654,N_595,N_448);
xor U1655 (N_1655,N_726,N_307);
and U1656 (N_1656,N_999,N_116);
or U1657 (N_1657,N_517,N_799);
nor U1658 (N_1658,N_39,N_474);
nor U1659 (N_1659,N_234,N_968);
nor U1660 (N_1660,N_227,N_343);
nand U1661 (N_1661,N_992,N_564);
or U1662 (N_1662,N_380,N_958);
and U1663 (N_1663,N_745,N_683);
and U1664 (N_1664,N_691,N_857);
and U1665 (N_1665,N_531,N_723);
or U1666 (N_1666,N_838,N_920);
and U1667 (N_1667,N_862,N_562);
xnor U1668 (N_1668,N_411,N_49);
nor U1669 (N_1669,N_787,N_619);
nand U1670 (N_1670,N_763,N_7);
and U1671 (N_1671,N_32,N_916);
and U1672 (N_1672,N_926,N_361);
or U1673 (N_1673,N_248,N_117);
nor U1674 (N_1674,N_661,N_589);
xnor U1675 (N_1675,N_121,N_641);
or U1676 (N_1676,N_295,N_791);
and U1677 (N_1677,N_625,N_768);
nor U1678 (N_1678,N_812,N_67);
or U1679 (N_1679,N_953,N_801);
xor U1680 (N_1680,N_314,N_800);
and U1681 (N_1681,N_679,N_826);
or U1682 (N_1682,N_496,N_268);
nor U1683 (N_1683,N_503,N_516);
nor U1684 (N_1684,N_479,N_625);
and U1685 (N_1685,N_874,N_398);
and U1686 (N_1686,N_177,N_222);
nand U1687 (N_1687,N_62,N_694);
nor U1688 (N_1688,N_634,N_776);
or U1689 (N_1689,N_889,N_46);
or U1690 (N_1690,N_279,N_452);
or U1691 (N_1691,N_440,N_508);
or U1692 (N_1692,N_807,N_45);
and U1693 (N_1693,N_673,N_62);
or U1694 (N_1694,N_22,N_611);
nand U1695 (N_1695,N_224,N_522);
nor U1696 (N_1696,N_555,N_734);
or U1697 (N_1697,N_984,N_290);
and U1698 (N_1698,N_929,N_61);
nand U1699 (N_1699,N_145,N_385);
nor U1700 (N_1700,N_861,N_591);
nand U1701 (N_1701,N_888,N_452);
xor U1702 (N_1702,N_74,N_977);
or U1703 (N_1703,N_143,N_149);
and U1704 (N_1704,N_657,N_431);
or U1705 (N_1705,N_738,N_152);
nor U1706 (N_1706,N_487,N_589);
and U1707 (N_1707,N_324,N_26);
and U1708 (N_1708,N_78,N_207);
nor U1709 (N_1709,N_137,N_912);
nand U1710 (N_1710,N_402,N_838);
xnor U1711 (N_1711,N_620,N_561);
nor U1712 (N_1712,N_312,N_982);
nand U1713 (N_1713,N_140,N_41);
xor U1714 (N_1714,N_96,N_817);
nor U1715 (N_1715,N_630,N_853);
nand U1716 (N_1716,N_882,N_723);
nand U1717 (N_1717,N_171,N_262);
nor U1718 (N_1718,N_342,N_12);
xor U1719 (N_1719,N_134,N_958);
or U1720 (N_1720,N_306,N_402);
and U1721 (N_1721,N_592,N_316);
and U1722 (N_1722,N_841,N_357);
nor U1723 (N_1723,N_922,N_297);
nand U1724 (N_1724,N_243,N_537);
nand U1725 (N_1725,N_403,N_598);
and U1726 (N_1726,N_864,N_590);
nor U1727 (N_1727,N_868,N_975);
nand U1728 (N_1728,N_706,N_840);
and U1729 (N_1729,N_335,N_206);
nor U1730 (N_1730,N_284,N_898);
nor U1731 (N_1731,N_88,N_445);
xor U1732 (N_1732,N_968,N_603);
xor U1733 (N_1733,N_577,N_937);
xnor U1734 (N_1734,N_871,N_181);
or U1735 (N_1735,N_571,N_492);
xor U1736 (N_1736,N_788,N_39);
nand U1737 (N_1737,N_673,N_578);
xnor U1738 (N_1738,N_624,N_910);
nor U1739 (N_1739,N_910,N_246);
nor U1740 (N_1740,N_498,N_150);
nor U1741 (N_1741,N_689,N_244);
and U1742 (N_1742,N_339,N_724);
xnor U1743 (N_1743,N_443,N_976);
nand U1744 (N_1744,N_313,N_24);
and U1745 (N_1745,N_205,N_827);
xnor U1746 (N_1746,N_825,N_341);
or U1747 (N_1747,N_207,N_636);
xor U1748 (N_1748,N_63,N_922);
nand U1749 (N_1749,N_879,N_663);
nor U1750 (N_1750,N_354,N_973);
xnor U1751 (N_1751,N_262,N_420);
xor U1752 (N_1752,N_179,N_294);
xor U1753 (N_1753,N_352,N_0);
xor U1754 (N_1754,N_460,N_935);
xor U1755 (N_1755,N_498,N_969);
xnor U1756 (N_1756,N_16,N_190);
and U1757 (N_1757,N_174,N_392);
nand U1758 (N_1758,N_841,N_737);
and U1759 (N_1759,N_495,N_750);
or U1760 (N_1760,N_624,N_441);
xnor U1761 (N_1761,N_594,N_408);
or U1762 (N_1762,N_910,N_847);
nor U1763 (N_1763,N_653,N_830);
nand U1764 (N_1764,N_745,N_180);
xor U1765 (N_1765,N_972,N_337);
and U1766 (N_1766,N_639,N_637);
nand U1767 (N_1767,N_723,N_10);
and U1768 (N_1768,N_637,N_253);
or U1769 (N_1769,N_27,N_394);
xnor U1770 (N_1770,N_535,N_570);
or U1771 (N_1771,N_222,N_202);
nor U1772 (N_1772,N_636,N_796);
xor U1773 (N_1773,N_696,N_532);
and U1774 (N_1774,N_657,N_798);
nor U1775 (N_1775,N_76,N_494);
or U1776 (N_1776,N_108,N_15);
and U1777 (N_1777,N_399,N_808);
nand U1778 (N_1778,N_246,N_40);
and U1779 (N_1779,N_324,N_230);
nand U1780 (N_1780,N_996,N_406);
and U1781 (N_1781,N_22,N_980);
xor U1782 (N_1782,N_604,N_444);
or U1783 (N_1783,N_370,N_558);
and U1784 (N_1784,N_84,N_163);
xor U1785 (N_1785,N_514,N_994);
nor U1786 (N_1786,N_728,N_342);
and U1787 (N_1787,N_477,N_659);
and U1788 (N_1788,N_836,N_739);
xnor U1789 (N_1789,N_208,N_415);
and U1790 (N_1790,N_394,N_204);
and U1791 (N_1791,N_908,N_725);
nand U1792 (N_1792,N_953,N_163);
nand U1793 (N_1793,N_66,N_91);
nand U1794 (N_1794,N_865,N_792);
nor U1795 (N_1795,N_943,N_117);
and U1796 (N_1796,N_862,N_455);
or U1797 (N_1797,N_549,N_765);
nand U1798 (N_1798,N_0,N_178);
and U1799 (N_1799,N_248,N_201);
or U1800 (N_1800,N_541,N_387);
or U1801 (N_1801,N_183,N_241);
and U1802 (N_1802,N_360,N_47);
or U1803 (N_1803,N_822,N_277);
nor U1804 (N_1804,N_669,N_903);
and U1805 (N_1805,N_300,N_270);
xnor U1806 (N_1806,N_509,N_845);
nand U1807 (N_1807,N_642,N_377);
nor U1808 (N_1808,N_665,N_202);
nor U1809 (N_1809,N_745,N_23);
nand U1810 (N_1810,N_525,N_755);
nor U1811 (N_1811,N_589,N_455);
nand U1812 (N_1812,N_984,N_511);
nor U1813 (N_1813,N_36,N_614);
xor U1814 (N_1814,N_798,N_494);
or U1815 (N_1815,N_159,N_513);
and U1816 (N_1816,N_402,N_659);
or U1817 (N_1817,N_51,N_691);
or U1818 (N_1818,N_930,N_342);
nor U1819 (N_1819,N_526,N_735);
nand U1820 (N_1820,N_928,N_561);
and U1821 (N_1821,N_173,N_870);
and U1822 (N_1822,N_744,N_2);
and U1823 (N_1823,N_875,N_28);
xnor U1824 (N_1824,N_270,N_825);
and U1825 (N_1825,N_914,N_183);
or U1826 (N_1826,N_31,N_85);
nand U1827 (N_1827,N_514,N_289);
nand U1828 (N_1828,N_766,N_954);
or U1829 (N_1829,N_510,N_492);
nor U1830 (N_1830,N_727,N_835);
nor U1831 (N_1831,N_255,N_121);
nor U1832 (N_1832,N_815,N_691);
or U1833 (N_1833,N_60,N_617);
nor U1834 (N_1834,N_482,N_194);
nor U1835 (N_1835,N_405,N_729);
nor U1836 (N_1836,N_536,N_427);
or U1837 (N_1837,N_453,N_824);
xnor U1838 (N_1838,N_8,N_517);
and U1839 (N_1839,N_318,N_11);
nand U1840 (N_1840,N_86,N_948);
xnor U1841 (N_1841,N_86,N_222);
xnor U1842 (N_1842,N_247,N_836);
and U1843 (N_1843,N_180,N_378);
xnor U1844 (N_1844,N_467,N_903);
xor U1845 (N_1845,N_425,N_59);
and U1846 (N_1846,N_857,N_531);
xor U1847 (N_1847,N_301,N_636);
xor U1848 (N_1848,N_588,N_478);
nand U1849 (N_1849,N_831,N_369);
and U1850 (N_1850,N_69,N_687);
nand U1851 (N_1851,N_43,N_530);
nand U1852 (N_1852,N_559,N_144);
xnor U1853 (N_1853,N_981,N_818);
nor U1854 (N_1854,N_507,N_886);
and U1855 (N_1855,N_865,N_894);
or U1856 (N_1856,N_312,N_21);
nand U1857 (N_1857,N_871,N_895);
nor U1858 (N_1858,N_829,N_747);
and U1859 (N_1859,N_279,N_834);
nor U1860 (N_1860,N_892,N_208);
nand U1861 (N_1861,N_319,N_574);
xor U1862 (N_1862,N_161,N_682);
xnor U1863 (N_1863,N_616,N_767);
or U1864 (N_1864,N_679,N_228);
and U1865 (N_1865,N_698,N_894);
xor U1866 (N_1866,N_728,N_788);
xor U1867 (N_1867,N_690,N_472);
xor U1868 (N_1868,N_812,N_557);
xor U1869 (N_1869,N_682,N_834);
or U1870 (N_1870,N_301,N_136);
xor U1871 (N_1871,N_150,N_454);
nor U1872 (N_1872,N_825,N_230);
or U1873 (N_1873,N_661,N_766);
nor U1874 (N_1874,N_905,N_217);
nand U1875 (N_1875,N_124,N_911);
or U1876 (N_1876,N_583,N_253);
xor U1877 (N_1877,N_880,N_973);
xnor U1878 (N_1878,N_121,N_466);
nor U1879 (N_1879,N_482,N_563);
and U1880 (N_1880,N_242,N_90);
or U1881 (N_1881,N_902,N_920);
and U1882 (N_1882,N_494,N_159);
nand U1883 (N_1883,N_807,N_949);
and U1884 (N_1884,N_607,N_173);
or U1885 (N_1885,N_792,N_127);
nand U1886 (N_1886,N_430,N_4);
or U1887 (N_1887,N_275,N_247);
nand U1888 (N_1888,N_536,N_919);
or U1889 (N_1889,N_30,N_907);
and U1890 (N_1890,N_527,N_503);
or U1891 (N_1891,N_561,N_659);
nand U1892 (N_1892,N_553,N_445);
or U1893 (N_1893,N_88,N_276);
nand U1894 (N_1894,N_139,N_889);
and U1895 (N_1895,N_702,N_468);
and U1896 (N_1896,N_27,N_79);
and U1897 (N_1897,N_660,N_408);
xnor U1898 (N_1898,N_824,N_787);
and U1899 (N_1899,N_849,N_734);
nor U1900 (N_1900,N_153,N_388);
and U1901 (N_1901,N_893,N_826);
xor U1902 (N_1902,N_236,N_783);
nor U1903 (N_1903,N_817,N_324);
nand U1904 (N_1904,N_399,N_494);
nor U1905 (N_1905,N_313,N_298);
or U1906 (N_1906,N_223,N_51);
xnor U1907 (N_1907,N_847,N_94);
nand U1908 (N_1908,N_210,N_291);
nor U1909 (N_1909,N_492,N_848);
or U1910 (N_1910,N_595,N_409);
or U1911 (N_1911,N_180,N_821);
xnor U1912 (N_1912,N_72,N_607);
nor U1913 (N_1913,N_331,N_614);
or U1914 (N_1914,N_287,N_635);
nor U1915 (N_1915,N_982,N_820);
or U1916 (N_1916,N_316,N_790);
xor U1917 (N_1917,N_908,N_568);
and U1918 (N_1918,N_29,N_805);
or U1919 (N_1919,N_584,N_683);
nand U1920 (N_1920,N_15,N_404);
xor U1921 (N_1921,N_762,N_63);
nand U1922 (N_1922,N_764,N_556);
and U1923 (N_1923,N_654,N_714);
nand U1924 (N_1924,N_665,N_698);
xor U1925 (N_1925,N_743,N_944);
xor U1926 (N_1926,N_548,N_627);
and U1927 (N_1927,N_266,N_979);
xnor U1928 (N_1928,N_26,N_896);
and U1929 (N_1929,N_336,N_626);
or U1930 (N_1930,N_178,N_327);
or U1931 (N_1931,N_424,N_323);
nand U1932 (N_1932,N_518,N_837);
xor U1933 (N_1933,N_521,N_458);
nand U1934 (N_1934,N_966,N_352);
nand U1935 (N_1935,N_940,N_507);
xnor U1936 (N_1936,N_502,N_616);
and U1937 (N_1937,N_238,N_10);
or U1938 (N_1938,N_583,N_377);
nand U1939 (N_1939,N_46,N_128);
and U1940 (N_1940,N_108,N_451);
and U1941 (N_1941,N_447,N_610);
nand U1942 (N_1942,N_187,N_859);
or U1943 (N_1943,N_830,N_61);
xor U1944 (N_1944,N_619,N_291);
nand U1945 (N_1945,N_215,N_183);
and U1946 (N_1946,N_668,N_489);
or U1947 (N_1947,N_651,N_655);
xor U1948 (N_1948,N_712,N_159);
xor U1949 (N_1949,N_34,N_954);
nor U1950 (N_1950,N_87,N_93);
and U1951 (N_1951,N_617,N_220);
or U1952 (N_1952,N_62,N_735);
nor U1953 (N_1953,N_660,N_359);
and U1954 (N_1954,N_671,N_284);
xnor U1955 (N_1955,N_891,N_99);
nor U1956 (N_1956,N_36,N_40);
nand U1957 (N_1957,N_568,N_107);
nand U1958 (N_1958,N_27,N_425);
nor U1959 (N_1959,N_930,N_524);
nor U1960 (N_1960,N_501,N_639);
nand U1961 (N_1961,N_726,N_866);
and U1962 (N_1962,N_516,N_702);
nor U1963 (N_1963,N_178,N_258);
nand U1964 (N_1964,N_517,N_231);
or U1965 (N_1965,N_898,N_470);
and U1966 (N_1966,N_8,N_871);
or U1967 (N_1967,N_96,N_57);
xnor U1968 (N_1968,N_865,N_202);
nor U1969 (N_1969,N_509,N_936);
nand U1970 (N_1970,N_594,N_823);
and U1971 (N_1971,N_464,N_87);
and U1972 (N_1972,N_355,N_806);
xnor U1973 (N_1973,N_804,N_413);
xnor U1974 (N_1974,N_611,N_456);
or U1975 (N_1975,N_947,N_432);
nand U1976 (N_1976,N_651,N_329);
xor U1977 (N_1977,N_850,N_307);
and U1978 (N_1978,N_126,N_55);
nand U1979 (N_1979,N_837,N_705);
nor U1980 (N_1980,N_699,N_674);
and U1981 (N_1981,N_762,N_354);
xnor U1982 (N_1982,N_439,N_307);
nand U1983 (N_1983,N_964,N_649);
nor U1984 (N_1984,N_928,N_367);
nand U1985 (N_1985,N_235,N_8);
nand U1986 (N_1986,N_745,N_178);
nand U1987 (N_1987,N_991,N_120);
nand U1988 (N_1988,N_297,N_348);
nor U1989 (N_1989,N_800,N_230);
xnor U1990 (N_1990,N_157,N_96);
nor U1991 (N_1991,N_465,N_746);
and U1992 (N_1992,N_418,N_38);
or U1993 (N_1993,N_428,N_494);
xor U1994 (N_1994,N_448,N_591);
or U1995 (N_1995,N_537,N_693);
nand U1996 (N_1996,N_222,N_584);
nor U1997 (N_1997,N_613,N_932);
and U1998 (N_1998,N_291,N_237);
nand U1999 (N_1999,N_203,N_29);
nor U2000 (N_2000,N_1726,N_1448);
nor U2001 (N_2001,N_1586,N_1662);
nand U2002 (N_2002,N_1568,N_1090);
nand U2003 (N_2003,N_1794,N_1139);
nand U2004 (N_2004,N_1634,N_1954);
nand U2005 (N_2005,N_1089,N_1515);
nor U2006 (N_2006,N_1289,N_1135);
and U2007 (N_2007,N_1440,N_1364);
xnor U2008 (N_2008,N_1035,N_1078);
nand U2009 (N_2009,N_1298,N_1658);
and U2010 (N_2010,N_1183,N_1282);
xor U2011 (N_2011,N_1710,N_1732);
xor U2012 (N_2012,N_1761,N_1245);
nor U2013 (N_2013,N_1885,N_1288);
or U2014 (N_2014,N_1018,N_1454);
xor U2015 (N_2015,N_1682,N_1964);
nor U2016 (N_2016,N_1113,N_1124);
and U2017 (N_2017,N_1354,N_1397);
nor U2018 (N_2018,N_1565,N_1343);
nand U2019 (N_2019,N_1914,N_1898);
nor U2020 (N_2020,N_1540,N_1164);
nand U2021 (N_2021,N_1916,N_1866);
and U2022 (N_2022,N_1766,N_1203);
nor U2023 (N_2023,N_1153,N_1152);
and U2024 (N_2024,N_1535,N_1082);
nand U2025 (N_2025,N_1337,N_1383);
xnor U2026 (N_2026,N_1935,N_1671);
xnor U2027 (N_2027,N_1297,N_1229);
and U2028 (N_2028,N_1753,N_1497);
nor U2029 (N_2029,N_1776,N_1132);
xnor U2030 (N_2030,N_1640,N_1429);
nand U2031 (N_2031,N_1011,N_1999);
nor U2032 (N_2032,N_1594,N_1121);
nand U2033 (N_2033,N_1752,N_1254);
nor U2034 (N_2034,N_1698,N_1032);
nand U2035 (N_2035,N_1517,N_1412);
nor U2036 (N_2036,N_1686,N_1111);
or U2037 (N_2037,N_1697,N_1617);
nand U2038 (N_2038,N_1899,N_1555);
or U2039 (N_2039,N_1562,N_1770);
nor U2040 (N_2040,N_1079,N_1377);
or U2041 (N_2041,N_1232,N_1211);
or U2042 (N_2042,N_1248,N_1253);
nor U2043 (N_2043,N_1906,N_1739);
or U2044 (N_2044,N_1528,N_1342);
xor U2045 (N_2045,N_1822,N_1845);
and U2046 (N_2046,N_1039,N_1496);
xor U2047 (N_2047,N_1600,N_1743);
and U2048 (N_2048,N_1595,N_1989);
nand U2049 (N_2049,N_1106,N_1873);
nand U2050 (N_2050,N_1509,N_1174);
and U2051 (N_2051,N_1792,N_1054);
xnor U2052 (N_2052,N_1775,N_1416);
nand U2053 (N_2053,N_1001,N_1042);
and U2054 (N_2054,N_1307,N_1733);
xor U2055 (N_2055,N_1053,N_1745);
xor U2056 (N_2056,N_1579,N_1228);
xnor U2057 (N_2057,N_1591,N_1273);
nand U2058 (N_2058,N_1738,N_1214);
nand U2059 (N_2059,N_1327,N_1684);
and U2060 (N_2060,N_1049,N_1172);
and U2061 (N_2061,N_1966,N_1843);
nand U2062 (N_2062,N_1829,N_1905);
nor U2063 (N_2063,N_1016,N_1353);
and U2064 (N_2064,N_1073,N_1541);
xor U2065 (N_2065,N_1126,N_1865);
and U2066 (N_2066,N_1584,N_1551);
nor U2067 (N_2067,N_1453,N_1668);
nand U2068 (N_2068,N_1476,N_1376);
nor U2069 (N_2069,N_1015,N_1570);
nand U2070 (N_2070,N_1473,N_1860);
xor U2071 (N_2071,N_1886,N_1799);
or U2072 (N_2072,N_1646,N_1270);
xor U2073 (N_2073,N_1455,N_1945);
or U2074 (N_2074,N_1031,N_1261);
or U2075 (N_2075,N_1560,N_1785);
and U2076 (N_2076,N_1236,N_1810);
and U2077 (N_2077,N_1177,N_1355);
nor U2078 (N_2078,N_1787,N_1240);
nor U2079 (N_2079,N_1890,N_1471);
and U2080 (N_2080,N_1045,N_1501);
and U2081 (N_2081,N_1825,N_1449);
nand U2082 (N_2082,N_1303,N_1877);
nand U2083 (N_2083,N_1086,N_1013);
nor U2084 (N_2084,N_1813,N_1610);
xor U2085 (N_2085,N_1424,N_1107);
and U2086 (N_2086,N_1009,N_1176);
nand U2087 (N_2087,N_1285,N_1181);
nand U2088 (N_2088,N_1818,N_1936);
nand U2089 (N_2089,N_1173,N_1774);
nand U2090 (N_2090,N_1201,N_1474);
or U2091 (N_2091,N_1022,N_1536);
nor U2092 (N_2092,N_1834,N_1573);
xor U2093 (N_2093,N_1499,N_1044);
nand U2094 (N_2094,N_1324,N_1731);
nor U2095 (N_2095,N_1724,N_1614);
or U2096 (N_2096,N_1826,N_1838);
nand U2097 (N_2097,N_1928,N_1812);
and U2098 (N_2098,N_1048,N_1421);
or U2099 (N_2099,N_1159,N_1213);
nand U2100 (N_2100,N_1538,N_1025);
nand U2101 (N_2101,N_1309,N_1790);
nor U2102 (N_2102,N_1814,N_1876);
or U2103 (N_2103,N_1242,N_1204);
or U2104 (N_2104,N_1464,N_1589);
nor U2105 (N_2105,N_1329,N_1328);
nor U2106 (N_2106,N_1479,N_1407);
nand U2107 (N_2107,N_1360,N_1757);
or U2108 (N_2108,N_1123,N_1807);
xnor U2109 (N_2109,N_1007,N_1508);
or U2110 (N_2110,N_1179,N_1104);
and U2111 (N_2111,N_1017,N_1868);
nand U2112 (N_2112,N_1892,N_1112);
nand U2113 (N_2113,N_1149,N_1639);
or U2114 (N_2114,N_1701,N_1771);
nor U2115 (N_2115,N_1058,N_1260);
and U2116 (N_2116,N_1144,N_1991);
nor U2117 (N_2117,N_1861,N_1587);
and U2118 (N_2118,N_1224,N_1549);
nor U2119 (N_2119,N_1628,N_1756);
nor U2120 (N_2120,N_1712,N_1849);
and U2121 (N_2121,N_1626,N_1599);
nor U2122 (N_2122,N_1005,N_1506);
nand U2123 (N_2123,N_1206,N_1024);
nor U2124 (N_2124,N_1396,N_1041);
and U2125 (N_2125,N_1488,N_1323);
nor U2126 (N_2126,N_1801,N_1809);
nor U2127 (N_2127,N_1403,N_1931);
nor U2128 (N_2128,N_1118,N_1981);
xnor U2129 (N_2129,N_1484,N_1797);
and U2130 (N_2130,N_1744,N_1333);
nand U2131 (N_2131,N_1675,N_1166);
or U2132 (N_2132,N_1727,N_1398);
and U2133 (N_2133,N_1767,N_1184);
xnor U2134 (N_2134,N_1883,N_1678);
xor U2135 (N_2135,N_1023,N_1037);
nor U2136 (N_2136,N_1315,N_1490);
nor U2137 (N_2137,N_1585,N_1577);
and U2138 (N_2138,N_1957,N_1059);
xor U2139 (N_2139,N_1714,N_1102);
xor U2140 (N_2140,N_1027,N_1197);
or U2141 (N_2141,N_1299,N_1817);
or U2142 (N_2142,N_1857,N_1721);
xnor U2143 (N_2143,N_1320,N_1163);
nor U2144 (N_2144,N_1859,N_1393);
or U2145 (N_2145,N_1477,N_1363);
or U2146 (N_2146,N_1511,N_1483);
and U2147 (N_2147,N_1489,N_1846);
nor U2148 (N_2148,N_1938,N_1103);
or U2149 (N_2149,N_1359,N_1379);
nor U2150 (N_2150,N_1125,N_1075);
xnor U2151 (N_2151,N_1130,N_1613);
nand U2152 (N_2152,N_1217,N_1661);
and U2153 (N_2153,N_1556,N_1858);
xnor U2154 (N_2154,N_1704,N_1108);
or U2155 (N_2155,N_1604,N_1066);
or U2156 (N_2156,N_1388,N_1872);
nor U2157 (N_2157,N_1820,N_1271);
nor U2158 (N_2158,N_1976,N_1644);
and U2159 (N_2159,N_1955,N_1993);
and U2160 (N_2160,N_1510,N_1447);
or U2161 (N_2161,N_1904,N_1940);
xnor U2162 (N_2162,N_1070,N_1390);
xor U2163 (N_2163,N_1332,N_1485);
and U2164 (N_2164,N_1021,N_1142);
nand U2165 (N_2165,N_1093,N_1347);
nor U2166 (N_2166,N_1322,N_1863);
and U2167 (N_2167,N_1420,N_1705);
or U2168 (N_2168,N_1947,N_1458);
nand U2169 (N_2169,N_1654,N_1350);
and U2170 (N_2170,N_1052,N_1576);
nor U2171 (N_2171,N_1395,N_1029);
nand U2172 (N_2172,N_1085,N_1856);
nor U2173 (N_2173,N_1074,N_1580);
nor U2174 (N_2174,N_1830,N_1855);
nand U2175 (N_2175,N_1523,N_1765);
or U2176 (N_2176,N_1735,N_1308);
nor U2177 (N_2177,N_1956,N_1729);
nand U2178 (N_2178,N_1965,N_1806);
and U2179 (N_2179,N_1609,N_1902);
or U2180 (N_2180,N_1268,N_1175);
nand U2181 (N_2181,N_1625,N_1716);
or U2182 (N_2182,N_1472,N_1050);
nor U2183 (N_2183,N_1795,N_1864);
xnor U2184 (N_2184,N_1321,N_1800);
nor U2185 (N_2185,N_1356,N_1294);
nand U2186 (N_2186,N_1046,N_1338);
and U2187 (N_2187,N_1318,N_1612);
and U2188 (N_2188,N_1798,N_1432);
xnor U2189 (N_2189,N_1690,N_1117);
nor U2190 (N_2190,N_1504,N_1038);
xor U2191 (N_2191,N_1419,N_1227);
xor U2192 (N_2192,N_1962,N_1193);
nor U2193 (N_2193,N_1894,N_1569);
and U2194 (N_2194,N_1871,N_1664);
xor U2195 (N_2195,N_1451,N_1572);
or U2196 (N_2196,N_1210,N_1707);
nand U2197 (N_2197,N_1428,N_1061);
nand U2198 (N_2198,N_1437,N_1832);
and U2199 (N_2199,N_1653,N_1546);
xor U2200 (N_2200,N_1629,N_1366);
nand U2201 (N_2201,N_1975,N_1215);
nor U2202 (N_2202,N_1647,N_1408);
and U2203 (N_2203,N_1747,N_1438);
nand U2204 (N_2204,N_1824,N_1505);
nor U2205 (N_2205,N_1719,N_1346);
xor U2206 (N_2206,N_1919,N_1486);
nor U2207 (N_2207,N_1689,N_1374);
xor U2208 (N_2208,N_1137,N_1205);
nor U2209 (N_2209,N_1150,N_1764);
nand U2210 (N_2210,N_1833,N_1115);
xor U2211 (N_2211,N_1951,N_1693);
xnor U2212 (N_2212,N_1839,N_1641);
nor U2213 (N_2213,N_1695,N_1122);
xor U2214 (N_2214,N_1889,N_1119);
xnor U2215 (N_2215,N_1095,N_1722);
xnor U2216 (N_2216,N_1401,N_1060);
or U2217 (N_2217,N_1971,N_1441);
nor U2218 (N_2218,N_1340,N_1406);
or U2219 (N_2219,N_1136,N_1385);
nor U2220 (N_2220,N_1683,N_1921);
nand U2221 (N_2221,N_1469,N_1944);
and U2222 (N_2222,N_1618,N_1493);
nor U2223 (N_2223,N_1051,N_1357);
xnor U2224 (N_2224,N_1207,N_1043);
nand U2225 (N_2225,N_1548,N_1526);
or U2226 (N_2226,N_1537,N_1450);
nand U2227 (N_2227,N_1847,N_1788);
nor U2228 (N_2228,N_1417,N_1141);
nor U2229 (N_2229,N_1762,N_1623);
nor U2230 (N_2230,N_1881,N_1632);
or U2231 (N_2231,N_1769,N_1445);
or U2232 (N_2232,N_1578,N_1430);
and U2233 (N_2233,N_1367,N_1442);
and U2234 (N_2234,N_1272,N_1274);
and U2235 (N_2235,N_1554,N_1837);
xnor U2236 (N_2236,N_1468,N_1287);
and U2237 (N_2237,N_1423,N_1778);
or U2238 (N_2238,N_1257,N_1312);
xor U2239 (N_2239,N_1998,N_1942);
nand U2240 (N_2240,N_1265,N_1186);
or U2241 (N_2241,N_1922,N_1602);
or U2242 (N_2242,N_1140,N_1913);
xnor U2243 (N_2243,N_1960,N_1606);
xor U2244 (N_2244,N_1087,N_1633);
xnor U2245 (N_2245,N_1495,N_1984);
nand U2246 (N_2246,N_1802,N_1997);
nor U2247 (N_2247,N_1558,N_1221);
or U2248 (N_2248,N_1256,N_1590);
or U2249 (N_2249,N_1763,N_1821);
nand U2250 (N_2250,N_1258,N_1751);
nor U2251 (N_2251,N_1734,N_1083);
xor U2252 (N_2252,N_1384,N_1741);
nor U2253 (N_2253,N_1462,N_1370);
nor U2254 (N_2254,N_1185,N_1827);
and U2255 (N_2255,N_1657,N_1676);
and U2256 (N_2256,N_1219,N_1963);
nand U2257 (N_2257,N_1055,N_1399);
or U2258 (N_2258,N_1598,N_1518);
or U2259 (N_2259,N_1316,N_1637);
or U2260 (N_2260,N_1311,N_1171);
nand U2261 (N_2261,N_1708,N_1004);
and U2262 (N_2262,N_1995,N_1842);
and U2263 (N_2263,N_1241,N_1068);
or U2264 (N_2264,N_1387,N_1725);
nor U2265 (N_2265,N_1869,N_1992);
nor U2266 (N_2266,N_1685,N_1878);
or U2267 (N_2267,N_1665,N_1758);
xnor U2268 (N_2268,N_1198,N_1335);
nor U2269 (N_2269,N_1696,N_1952);
xnor U2270 (N_2270,N_1677,N_1169);
nand U2271 (N_2271,N_1267,N_1557);
and U2272 (N_2272,N_1187,N_1252);
nand U2273 (N_2273,N_1290,N_1230);
or U2274 (N_2274,N_1099,N_1514);
xor U2275 (N_2275,N_1953,N_1231);
or U2276 (N_2276,N_1915,N_1434);
nand U2277 (N_2277,N_1702,N_1681);
and U2278 (N_2278,N_1389,N_1543);
and U2279 (N_2279,N_1645,N_1351);
or U2280 (N_2280,N_1939,N_1870);
xnor U2281 (N_2281,N_1791,N_1460);
xor U2282 (N_2282,N_1244,N_1912);
xor U2283 (N_2283,N_1978,N_1619);
nand U2284 (N_2284,N_1190,N_1310);
and U2285 (N_2285,N_1828,N_1012);
xor U2286 (N_2286,N_1715,N_1165);
or U2287 (N_2287,N_1196,N_1854);
and U2288 (N_2288,N_1679,N_1131);
xor U2289 (N_2289,N_1974,N_1611);
nand U2290 (N_2290,N_1969,N_1239);
nor U2291 (N_2291,N_1850,N_1603);
xor U2292 (N_2292,N_1909,N_1893);
nor U2293 (N_2293,N_1092,N_1411);
or U2294 (N_2294,N_1313,N_1552);
xor U2295 (N_2295,N_1918,N_1404);
and U2296 (N_2296,N_1276,N_1669);
or U2297 (N_2297,N_1154,N_1133);
or U2298 (N_2298,N_1280,N_1266);
nor U2299 (N_2299,N_1607,N_1680);
nor U2300 (N_2300,N_1970,N_1180);
and U2301 (N_2301,N_1925,N_1780);
nand U2302 (N_2302,N_1415,N_1063);
or U2303 (N_2303,N_1391,N_1740);
xnor U2304 (N_2304,N_1002,N_1286);
nor U2305 (N_2305,N_1973,N_1760);
xor U2306 (N_2306,N_1443,N_1178);
nand U2307 (N_2307,N_1781,N_1815);
or U2308 (N_2308,N_1982,N_1901);
or U2309 (N_2309,N_1655,N_1128);
nand U2310 (N_2310,N_1672,N_1065);
or U2311 (N_2311,N_1492,N_1375);
nand U2312 (N_2312,N_1717,N_1067);
or U2313 (N_2313,N_1161,N_1779);
nor U2314 (N_2314,N_1694,N_1097);
xor U2315 (N_2315,N_1003,N_1987);
xnor U2316 (N_2316,N_1786,N_1251);
and U2317 (N_2317,N_1803,N_1519);
nand U2318 (N_2318,N_1129,N_1804);
or U2319 (N_2319,N_1369,N_1218);
or U2320 (N_2320,N_1888,N_1848);
nor U2321 (N_2321,N_1006,N_1223);
and U2322 (N_2322,N_1782,N_1648);
nor U2323 (N_2323,N_1972,N_1927);
and U2324 (N_2324,N_1138,N_1371);
nor U2325 (N_2325,N_1279,N_1673);
nor U2326 (N_2326,N_1608,N_1147);
xor U2327 (N_2327,N_1295,N_1530);
nand U2328 (N_2328,N_1575,N_1937);
nand U2329 (N_2329,N_1642,N_1621);
nand U2330 (N_2330,N_1402,N_1891);
nor U2331 (N_2331,N_1202,N_1088);
nor U2332 (N_2332,N_1636,N_1533);
xnor U2333 (N_2333,N_1348,N_1284);
nor U2334 (N_2334,N_1302,N_1336);
xnor U2335 (N_2335,N_1674,N_1326);
nand U2336 (N_2336,N_1875,N_1895);
nand U2337 (N_2337,N_1596,N_1026);
nand U2338 (N_2338,N_1200,N_1170);
xor U2339 (N_2339,N_1713,N_1365);
xor U2340 (N_2340,N_1582,N_1344);
nand U2341 (N_2341,N_1525,N_1539);
xnor U2342 (N_2342,N_1475,N_1564);
nand U2343 (N_2343,N_1110,N_1819);
xnor U2344 (N_2344,N_1304,N_1498);
xor U2345 (N_2345,N_1941,N_1158);
and U2346 (N_2346,N_1456,N_1567);
nand U2347 (N_2347,N_1522,N_1884);
or U2348 (N_2348,N_1482,N_1480);
xor U2349 (N_2349,N_1494,N_1091);
or U2350 (N_2350,N_1247,N_1189);
and U2351 (N_2351,N_1487,N_1789);
xor U2352 (N_2352,N_1728,N_1840);
nor U2353 (N_2353,N_1768,N_1571);
nor U2354 (N_2354,N_1793,N_1467);
and U2355 (N_2355,N_1077,N_1699);
nor U2356 (N_2356,N_1461,N_1278);
nor U2357 (N_2357,N_1317,N_1422);
nand U2358 (N_2358,N_1334,N_1911);
and U2359 (N_2359,N_1652,N_1831);
and U2360 (N_2360,N_1746,N_1853);
nor U2361 (N_2361,N_1100,N_1930);
nor U2362 (N_2362,N_1275,N_1980);
or U2363 (N_2363,N_1306,N_1362);
xor U2364 (N_2364,N_1358,N_1742);
nand U2365 (N_2365,N_1056,N_1431);
xor U2366 (N_2366,N_1028,N_1507);
xor U2367 (N_2367,N_1926,N_1116);
xor U2368 (N_2368,N_1638,N_1862);
nand U2369 (N_2369,N_1841,N_1529);
nor U2370 (N_2370,N_1188,N_1319);
and U2371 (N_2371,N_1723,N_1920);
nor U2372 (N_2372,N_1923,N_1392);
nor U2373 (N_2373,N_1996,N_1605);
xnor U2374 (N_2374,N_1851,N_1934);
and U2375 (N_2375,N_1929,N_1019);
or U2376 (N_2376,N_1896,N_1410);
xor U2377 (N_2377,N_1381,N_1465);
xor U2378 (N_2378,N_1933,N_1151);
or U2379 (N_2379,N_1650,N_1405);
nor U2380 (N_2380,N_1062,N_1544);
nor U2381 (N_2381,N_1156,N_1882);
or U2382 (N_2382,N_1076,N_1627);
or U2383 (N_2383,N_1811,N_1314);
nand U2384 (N_2384,N_1084,N_1264);
and U2385 (N_2385,N_1532,N_1143);
or U2386 (N_2386,N_1805,N_1667);
nand U2387 (N_2387,N_1720,N_1553);
xnor U2388 (N_2388,N_1292,N_1755);
nand U2389 (N_2389,N_1737,N_1209);
or U2390 (N_2390,N_1730,N_1439);
or U2391 (N_2391,N_1120,N_1014);
and U2392 (N_2392,N_1703,N_1101);
or U2393 (N_2393,N_1146,N_1624);
nor U2394 (N_2394,N_1670,N_1736);
nand U2395 (N_2395,N_1000,N_1783);
nor U2396 (N_2396,N_1109,N_1466);
and U2397 (N_2397,N_1622,N_1220);
and U2398 (N_2398,N_1691,N_1759);
nor U2399 (N_2399,N_1545,N_1643);
xor U2400 (N_2400,N_1503,N_1008);
nor U2401 (N_2401,N_1225,N_1547);
or U2402 (N_2402,N_1243,N_1649);
nor U2403 (N_2403,N_1836,N_1666);
or U2404 (N_2404,N_1057,N_1773);
nand U2405 (N_2405,N_1948,N_1500);
or U2406 (N_2406,N_1887,N_1990);
xnor U2407 (N_2407,N_1520,N_1823);
nor U2408 (N_2408,N_1979,N_1226);
or U2409 (N_2409,N_1081,N_1418);
or U2410 (N_2410,N_1784,N_1296);
nand U2411 (N_2411,N_1444,N_1134);
nor U2412 (N_2412,N_1542,N_1330);
xnor U2413 (N_2413,N_1033,N_1433);
and U2414 (N_2414,N_1581,N_1816);
or U2415 (N_2415,N_1047,N_1331);
nand U2416 (N_2416,N_1709,N_1985);
or U2417 (N_2417,N_1959,N_1446);
nand U2418 (N_2418,N_1660,N_1096);
and U2419 (N_2419,N_1597,N_1182);
xor U2420 (N_2420,N_1457,N_1349);
nand U2421 (N_2421,N_1234,N_1212);
xor U2422 (N_2422,N_1932,N_1656);
nand U2423 (N_2423,N_1277,N_1692);
nor U2424 (N_2424,N_1852,N_1534);
xnor U2425 (N_2425,N_1237,N_1373);
and U2426 (N_2426,N_1249,N_1098);
or U2427 (N_2427,N_1233,N_1907);
xor U2428 (N_2428,N_1835,N_1195);
or U2429 (N_2429,N_1345,N_1293);
and U2430 (N_2430,N_1867,N_1512);
or U2431 (N_2431,N_1259,N_1601);
nor U2432 (N_2432,N_1339,N_1879);
xor U2433 (N_2433,N_1036,N_1986);
xnor U2434 (N_2434,N_1114,N_1238);
xnor U2435 (N_2435,N_1436,N_1967);
nor U2436 (N_2436,N_1064,N_1157);
xor U2437 (N_2437,N_1382,N_1903);
and U2438 (N_2438,N_1325,N_1235);
nand U2439 (N_2439,N_1105,N_1291);
nor U2440 (N_2440,N_1531,N_1949);
and U2441 (N_2441,N_1900,N_1513);
xor U2442 (N_2442,N_1559,N_1145);
nand U2443 (N_2443,N_1192,N_1502);
xnor U2444 (N_2444,N_1844,N_1414);
or U2445 (N_2445,N_1961,N_1635);
xnor U2446 (N_2446,N_1413,N_1977);
nand U2447 (N_2447,N_1615,N_1958);
nand U2448 (N_2448,N_1750,N_1478);
nand U2449 (N_2449,N_1435,N_1563);
xor U2450 (N_2450,N_1168,N_1030);
xnor U2451 (N_2451,N_1368,N_1663);
nand U2452 (N_2452,N_1593,N_1283);
nor U2453 (N_2453,N_1409,N_1777);
and U2454 (N_2454,N_1687,N_1988);
xnor U2455 (N_2455,N_1550,N_1160);
xor U2456 (N_2456,N_1167,N_1094);
and U2457 (N_2457,N_1080,N_1255);
or U2458 (N_2458,N_1688,N_1194);
and U2459 (N_2459,N_1208,N_1749);
or U2460 (N_2460,N_1352,N_1946);
and U2461 (N_2461,N_1216,N_1246);
and U2462 (N_2462,N_1341,N_1968);
xor U2463 (N_2463,N_1620,N_1394);
or U2464 (N_2464,N_1191,N_1706);
or U2465 (N_2465,N_1994,N_1583);
nor U2466 (N_2466,N_1281,N_1772);
nor U2467 (N_2467,N_1400,N_1425);
xor U2468 (N_2468,N_1711,N_1561);
nand U2469 (N_2469,N_1263,N_1269);
and U2470 (N_2470,N_1659,N_1162);
and U2471 (N_2471,N_1426,N_1199);
nand U2472 (N_2472,N_1521,N_1072);
or U2473 (N_2473,N_1943,N_1491);
and U2474 (N_2474,N_1592,N_1380);
xor U2475 (N_2475,N_1300,N_1524);
nand U2476 (N_2476,N_1020,N_1718);
and U2477 (N_2477,N_1301,N_1262);
xnor U2478 (N_2478,N_1010,N_1880);
nor U2479 (N_2479,N_1459,N_1897);
and U2480 (N_2480,N_1566,N_1481);
and U2481 (N_2481,N_1910,N_1917);
xnor U2482 (N_2482,N_1155,N_1574);
nor U2483 (N_2483,N_1372,N_1908);
or U2484 (N_2484,N_1470,N_1631);
nor U2485 (N_2485,N_1924,N_1071);
and U2486 (N_2486,N_1630,N_1305);
nor U2487 (N_2487,N_1452,N_1034);
nand U2488 (N_2488,N_1427,N_1386);
nor U2489 (N_2489,N_1796,N_1616);
and U2490 (N_2490,N_1127,N_1808);
or U2491 (N_2491,N_1148,N_1950);
and U2492 (N_2492,N_1748,N_1516);
and U2493 (N_2493,N_1754,N_1983);
xor U2494 (N_2494,N_1700,N_1463);
and U2495 (N_2495,N_1378,N_1250);
xnor U2496 (N_2496,N_1361,N_1588);
nand U2497 (N_2497,N_1527,N_1069);
xor U2498 (N_2498,N_1874,N_1222);
nand U2499 (N_2499,N_1040,N_1651);
and U2500 (N_2500,N_1713,N_1910);
xor U2501 (N_2501,N_1050,N_1611);
nand U2502 (N_2502,N_1387,N_1835);
xor U2503 (N_2503,N_1254,N_1835);
nand U2504 (N_2504,N_1423,N_1539);
nor U2505 (N_2505,N_1904,N_1985);
or U2506 (N_2506,N_1775,N_1073);
nor U2507 (N_2507,N_1719,N_1751);
nand U2508 (N_2508,N_1559,N_1280);
xnor U2509 (N_2509,N_1577,N_1660);
nand U2510 (N_2510,N_1884,N_1333);
nand U2511 (N_2511,N_1025,N_1553);
xor U2512 (N_2512,N_1939,N_1453);
and U2513 (N_2513,N_1526,N_1448);
xor U2514 (N_2514,N_1324,N_1511);
xnor U2515 (N_2515,N_1701,N_1351);
nand U2516 (N_2516,N_1116,N_1583);
nand U2517 (N_2517,N_1927,N_1130);
or U2518 (N_2518,N_1149,N_1461);
nand U2519 (N_2519,N_1742,N_1020);
or U2520 (N_2520,N_1556,N_1378);
nand U2521 (N_2521,N_1958,N_1549);
nor U2522 (N_2522,N_1538,N_1912);
or U2523 (N_2523,N_1731,N_1839);
nand U2524 (N_2524,N_1917,N_1288);
xor U2525 (N_2525,N_1380,N_1792);
xor U2526 (N_2526,N_1817,N_1131);
xor U2527 (N_2527,N_1243,N_1527);
nand U2528 (N_2528,N_1670,N_1556);
xor U2529 (N_2529,N_1522,N_1834);
or U2530 (N_2530,N_1595,N_1341);
xnor U2531 (N_2531,N_1239,N_1798);
and U2532 (N_2532,N_1736,N_1790);
xnor U2533 (N_2533,N_1533,N_1491);
and U2534 (N_2534,N_1364,N_1526);
nand U2535 (N_2535,N_1836,N_1039);
nor U2536 (N_2536,N_1396,N_1631);
xor U2537 (N_2537,N_1823,N_1595);
and U2538 (N_2538,N_1366,N_1191);
nor U2539 (N_2539,N_1036,N_1013);
and U2540 (N_2540,N_1927,N_1773);
nand U2541 (N_2541,N_1447,N_1068);
and U2542 (N_2542,N_1410,N_1435);
xor U2543 (N_2543,N_1064,N_1367);
and U2544 (N_2544,N_1268,N_1634);
xnor U2545 (N_2545,N_1063,N_1773);
nand U2546 (N_2546,N_1500,N_1952);
or U2547 (N_2547,N_1065,N_1064);
nor U2548 (N_2548,N_1054,N_1738);
and U2549 (N_2549,N_1985,N_1054);
xnor U2550 (N_2550,N_1912,N_1471);
nor U2551 (N_2551,N_1170,N_1087);
nand U2552 (N_2552,N_1664,N_1448);
nand U2553 (N_2553,N_1629,N_1887);
xnor U2554 (N_2554,N_1267,N_1355);
nor U2555 (N_2555,N_1726,N_1731);
nor U2556 (N_2556,N_1265,N_1903);
and U2557 (N_2557,N_1705,N_1170);
or U2558 (N_2558,N_1891,N_1306);
xor U2559 (N_2559,N_1056,N_1818);
and U2560 (N_2560,N_1521,N_1151);
nor U2561 (N_2561,N_1428,N_1168);
nand U2562 (N_2562,N_1232,N_1877);
and U2563 (N_2563,N_1411,N_1397);
and U2564 (N_2564,N_1042,N_1064);
nor U2565 (N_2565,N_1075,N_1773);
and U2566 (N_2566,N_1352,N_1471);
or U2567 (N_2567,N_1766,N_1813);
nor U2568 (N_2568,N_1049,N_1010);
xnor U2569 (N_2569,N_1969,N_1907);
or U2570 (N_2570,N_1425,N_1282);
nor U2571 (N_2571,N_1493,N_1875);
or U2572 (N_2572,N_1774,N_1130);
nand U2573 (N_2573,N_1691,N_1251);
and U2574 (N_2574,N_1938,N_1228);
nor U2575 (N_2575,N_1536,N_1449);
or U2576 (N_2576,N_1383,N_1865);
nand U2577 (N_2577,N_1300,N_1678);
and U2578 (N_2578,N_1993,N_1748);
and U2579 (N_2579,N_1145,N_1299);
and U2580 (N_2580,N_1174,N_1130);
and U2581 (N_2581,N_1318,N_1420);
and U2582 (N_2582,N_1672,N_1087);
or U2583 (N_2583,N_1568,N_1081);
and U2584 (N_2584,N_1779,N_1364);
nand U2585 (N_2585,N_1723,N_1813);
and U2586 (N_2586,N_1933,N_1378);
nand U2587 (N_2587,N_1828,N_1857);
xor U2588 (N_2588,N_1944,N_1437);
or U2589 (N_2589,N_1200,N_1880);
nand U2590 (N_2590,N_1390,N_1117);
nor U2591 (N_2591,N_1622,N_1422);
nor U2592 (N_2592,N_1118,N_1338);
and U2593 (N_2593,N_1385,N_1273);
nand U2594 (N_2594,N_1607,N_1925);
or U2595 (N_2595,N_1479,N_1758);
nor U2596 (N_2596,N_1581,N_1704);
or U2597 (N_2597,N_1684,N_1559);
nand U2598 (N_2598,N_1904,N_1041);
nor U2599 (N_2599,N_1984,N_1336);
nor U2600 (N_2600,N_1031,N_1689);
and U2601 (N_2601,N_1436,N_1860);
nor U2602 (N_2602,N_1027,N_1549);
nand U2603 (N_2603,N_1848,N_1025);
nand U2604 (N_2604,N_1137,N_1787);
nor U2605 (N_2605,N_1617,N_1347);
or U2606 (N_2606,N_1998,N_1751);
nand U2607 (N_2607,N_1351,N_1407);
and U2608 (N_2608,N_1953,N_1964);
and U2609 (N_2609,N_1835,N_1381);
xor U2610 (N_2610,N_1597,N_1405);
nand U2611 (N_2611,N_1040,N_1616);
and U2612 (N_2612,N_1121,N_1099);
xor U2613 (N_2613,N_1939,N_1792);
or U2614 (N_2614,N_1533,N_1078);
or U2615 (N_2615,N_1590,N_1351);
and U2616 (N_2616,N_1373,N_1747);
and U2617 (N_2617,N_1801,N_1295);
or U2618 (N_2618,N_1373,N_1026);
nand U2619 (N_2619,N_1379,N_1265);
and U2620 (N_2620,N_1805,N_1185);
nand U2621 (N_2621,N_1530,N_1072);
and U2622 (N_2622,N_1265,N_1476);
nor U2623 (N_2623,N_1827,N_1132);
nor U2624 (N_2624,N_1275,N_1752);
and U2625 (N_2625,N_1012,N_1657);
nor U2626 (N_2626,N_1060,N_1041);
nor U2627 (N_2627,N_1263,N_1576);
or U2628 (N_2628,N_1897,N_1770);
nor U2629 (N_2629,N_1373,N_1319);
nor U2630 (N_2630,N_1068,N_1500);
nand U2631 (N_2631,N_1033,N_1875);
nand U2632 (N_2632,N_1593,N_1279);
nor U2633 (N_2633,N_1902,N_1803);
nand U2634 (N_2634,N_1952,N_1094);
nor U2635 (N_2635,N_1549,N_1597);
xnor U2636 (N_2636,N_1807,N_1691);
and U2637 (N_2637,N_1176,N_1181);
nor U2638 (N_2638,N_1665,N_1313);
nand U2639 (N_2639,N_1511,N_1595);
or U2640 (N_2640,N_1344,N_1937);
nor U2641 (N_2641,N_1142,N_1863);
xnor U2642 (N_2642,N_1440,N_1613);
xnor U2643 (N_2643,N_1102,N_1019);
or U2644 (N_2644,N_1156,N_1525);
xor U2645 (N_2645,N_1574,N_1530);
and U2646 (N_2646,N_1522,N_1699);
and U2647 (N_2647,N_1124,N_1372);
nand U2648 (N_2648,N_1078,N_1994);
and U2649 (N_2649,N_1667,N_1884);
or U2650 (N_2650,N_1983,N_1323);
nand U2651 (N_2651,N_1176,N_1539);
nor U2652 (N_2652,N_1955,N_1028);
and U2653 (N_2653,N_1395,N_1544);
nand U2654 (N_2654,N_1534,N_1862);
nand U2655 (N_2655,N_1602,N_1191);
or U2656 (N_2656,N_1662,N_1212);
and U2657 (N_2657,N_1106,N_1691);
nor U2658 (N_2658,N_1247,N_1132);
nand U2659 (N_2659,N_1739,N_1434);
and U2660 (N_2660,N_1372,N_1911);
xor U2661 (N_2661,N_1263,N_1003);
nor U2662 (N_2662,N_1302,N_1734);
nor U2663 (N_2663,N_1904,N_1926);
nand U2664 (N_2664,N_1817,N_1892);
nand U2665 (N_2665,N_1859,N_1643);
or U2666 (N_2666,N_1664,N_1621);
xor U2667 (N_2667,N_1155,N_1876);
nor U2668 (N_2668,N_1331,N_1737);
xnor U2669 (N_2669,N_1974,N_1939);
nand U2670 (N_2670,N_1095,N_1474);
and U2671 (N_2671,N_1217,N_1054);
nor U2672 (N_2672,N_1681,N_1698);
or U2673 (N_2673,N_1826,N_1854);
xor U2674 (N_2674,N_1462,N_1510);
xnor U2675 (N_2675,N_1552,N_1231);
xor U2676 (N_2676,N_1934,N_1396);
and U2677 (N_2677,N_1252,N_1782);
nor U2678 (N_2678,N_1545,N_1488);
xor U2679 (N_2679,N_1936,N_1006);
nand U2680 (N_2680,N_1229,N_1233);
and U2681 (N_2681,N_1072,N_1397);
and U2682 (N_2682,N_1805,N_1616);
and U2683 (N_2683,N_1719,N_1611);
nor U2684 (N_2684,N_1863,N_1589);
nor U2685 (N_2685,N_1183,N_1121);
and U2686 (N_2686,N_1607,N_1173);
or U2687 (N_2687,N_1043,N_1237);
or U2688 (N_2688,N_1241,N_1179);
and U2689 (N_2689,N_1164,N_1282);
nand U2690 (N_2690,N_1954,N_1807);
nor U2691 (N_2691,N_1426,N_1216);
xor U2692 (N_2692,N_1098,N_1992);
or U2693 (N_2693,N_1195,N_1606);
xnor U2694 (N_2694,N_1656,N_1596);
or U2695 (N_2695,N_1336,N_1182);
nor U2696 (N_2696,N_1661,N_1479);
nand U2697 (N_2697,N_1627,N_1211);
xnor U2698 (N_2698,N_1859,N_1073);
or U2699 (N_2699,N_1933,N_1665);
and U2700 (N_2700,N_1081,N_1987);
and U2701 (N_2701,N_1933,N_1507);
or U2702 (N_2702,N_1961,N_1496);
and U2703 (N_2703,N_1695,N_1379);
nor U2704 (N_2704,N_1989,N_1137);
xor U2705 (N_2705,N_1888,N_1901);
nand U2706 (N_2706,N_1468,N_1505);
nor U2707 (N_2707,N_1784,N_1802);
nor U2708 (N_2708,N_1169,N_1194);
xor U2709 (N_2709,N_1577,N_1044);
nor U2710 (N_2710,N_1944,N_1164);
nand U2711 (N_2711,N_1934,N_1253);
xnor U2712 (N_2712,N_1576,N_1211);
or U2713 (N_2713,N_1179,N_1186);
nand U2714 (N_2714,N_1404,N_1202);
and U2715 (N_2715,N_1501,N_1759);
and U2716 (N_2716,N_1115,N_1349);
and U2717 (N_2717,N_1452,N_1759);
nand U2718 (N_2718,N_1982,N_1312);
xnor U2719 (N_2719,N_1537,N_1140);
nand U2720 (N_2720,N_1616,N_1608);
xor U2721 (N_2721,N_1296,N_1898);
and U2722 (N_2722,N_1070,N_1977);
nand U2723 (N_2723,N_1594,N_1197);
or U2724 (N_2724,N_1483,N_1207);
or U2725 (N_2725,N_1536,N_1531);
xor U2726 (N_2726,N_1428,N_1078);
and U2727 (N_2727,N_1651,N_1456);
or U2728 (N_2728,N_1093,N_1570);
nand U2729 (N_2729,N_1132,N_1067);
nor U2730 (N_2730,N_1706,N_1905);
nor U2731 (N_2731,N_1234,N_1650);
xor U2732 (N_2732,N_1865,N_1041);
xor U2733 (N_2733,N_1808,N_1920);
nor U2734 (N_2734,N_1149,N_1612);
nand U2735 (N_2735,N_1932,N_1750);
or U2736 (N_2736,N_1331,N_1955);
or U2737 (N_2737,N_1995,N_1864);
and U2738 (N_2738,N_1005,N_1753);
xnor U2739 (N_2739,N_1373,N_1889);
nor U2740 (N_2740,N_1631,N_1163);
nor U2741 (N_2741,N_1479,N_1512);
nand U2742 (N_2742,N_1459,N_1191);
xor U2743 (N_2743,N_1323,N_1585);
xor U2744 (N_2744,N_1225,N_1887);
or U2745 (N_2745,N_1352,N_1823);
or U2746 (N_2746,N_1742,N_1763);
and U2747 (N_2747,N_1192,N_1341);
xor U2748 (N_2748,N_1042,N_1626);
xor U2749 (N_2749,N_1928,N_1083);
xor U2750 (N_2750,N_1378,N_1619);
nand U2751 (N_2751,N_1519,N_1763);
and U2752 (N_2752,N_1942,N_1923);
and U2753 (N_2753,N_1833,N_1056);
or U2754 (N_2754,N_1683,N_1413);
and U2755 (N_2755,N_1261,N_1588);
xor U2756 (N_2756,N_1747,N_1192);
and U2757 (N_2757,N_1456,N_1857);
nand U2758 (N_2758,N_1602,N_1376);
and U2759 (N_2759,N_1860,N_1391);
nand U2760 (N_2760,N_1811,N_1694);
nor U2761 (N_2761,N_1939,N_1208);
and U2762 (N_2762,N_1095,N_1771);
xnor U2763 (N_2763,N_1212,N_1274);
nor U2764 (N_2764,N_1147,N_1703);
or U2765 (N_2765,N_1453,N_1514);
xnor U2766 (N_2766,N_1696,N_1259);
xnor U2767 (N_2767,N_1223,N_1816);
xnor U2768 (N_2768,N_1704,N_1960);
and U2769 (N_2769,N_1562,N_1687);
or U2770 (N_2770,N_1385,N_1388);
nand U2771 (N_2771,N_1904,N_1237);
xnor U2772 (N_2772,N_1947,N_1118);
or U2773 (N_2773,N_1234,N_1495);
nor U2774 (N_2774,N_1985,N_1119);
and U2775 (N_2775,N_1616,N_1113);
and U2776 (N_2776,N_1158,N_1362);
nor U2777 (N_2777,N_1094,N_1596);
xnor U2778 (N_2778,N_1407,N_1766);
nand U2779 (N_2779,N_1657,N_1534);
and U2780 (N_2780,N_1562,N_1933);
and U2781 (N_2781,N_1719,N_1829);
xnor U2782 (N_2782,N_1637,N_1420);
nor U2783 (N_2783,N_1329,N_1819);
xor U2784 (N_2784,N_1092,N_1456);
nor U2785 (N_2785,N_1052,N_1541);
xor U2786 (N_2786,N_1843,N_1731);
and U2787 (N_2787,N_1944,N_1473);
xnor U2788 (N_2788,N_1039,N_1952);
nand U2789 (N_2789,N_1788,N_1503);
or U2790 (N_2790,N_1662,N_1631);
or U2791 (N_2791,N_1316,N_1771);
nor U2792 (N_2792,N_1653,N_1683);
and U2793 (N_2793,N_1637,N_1535);
and U2794 (N_2794,N_1480,N_1392);
xnor U2795 (N_2795,N_1136,N_1972);
and U2796 (N_2796,N_1354,N_1365);
nand U2797 (N_2797,N_1653,N_1656);
xor U2798 (N_2798,N_1302,N_1882);
nand U2799 (N_2799,N_1956,N_1811);
nor U2800 (N_2800,N_1948,N_1947);
and U2801 (N_2801,N_1248,N_1359);
nor U2802 (N_2802,N_1453,N_1918);
and U2803 (N_2803,N_1476,N_1411);
and U2804 (N_2804,N_1321,N_1971);
and U2805 (N_2805,N_1030,N_1392);
or U2806 (N_2806,N_1514,N_1973);
nor U2807 (N_2807,N_1720,N_1497);
or U2808 (N_2808,N_1593,N_1663);
or U2809 (N_2809,N_1730,N_1321);
nand U2810 (N_2810,N_1284,N_1083);
or U2811 (N_2811,N_1011,N_1700);
xor U2812 (N_2812,N_1929,N_1910);
nand U2813 (N_2813,N_1036,N_1731);
xnor U2814 (N_2814,N_1329,N_1285);
nand U2815 (N_2815,N_1994,N_1062);
nor U2816 (N_2816,N_1468,N_1996);
nand U2817 (N_2817,N_1051,N_1323);
and U2818 (N_2818,N_1020,N_1180);
nand U2819 (N_2819,N_1250,N_1347);
nand U2820 (N_2820,N_1506,N_1749);
nand U2821 (N_2821,N_1661,N_1208);
nor U2822 (N_2822,N_1177,N_1834);
or U2823 (N_2823,N_1830,N_1765);
or U2824 (N_2824,N_1339,N_1046);
and U2825 (N_2825,N_1432,N_1862);
or U2826 (N_2826,N_1382,N_1038);
or U2827 (N_2827,N_1431,N_1473);
and U2828 (N_2828,N_1426,N_1463);
or U2829 (N_2829,N_1441,N_1184);
xor U2830 (N_2830,N_1152,N_1116);
nor U2831 (N_2831,N_1978,N_1647);
or U2832 (N_2832,N_1886,N_1065);
xnor U2833 (N_2833,N_1254,N_1855);
nand U2834 (N_2834,N_1666,N_1854);
nor U2835 (N_2835,N_1394,N_1784);
and U2836 (N_2836,N_1956,N_1360);
xor U2837 (N_2837,N_1560,N_1619);
xor U2838 (N_2838,N_1770,N_1685);
and U2839 (N_2839,N_1510,N_1852);
and U2840 (N_2840,N_1585,N_1795);
nand U2841 (N_2841,N_1314,N_1537);
and U2842 (N_2842,N_1850,N_1507);
nor U2843 (N_2843,N_1304,N_1497);
xnor U2844 (N_2844,N_1369,N_1720);
nor U2845 (N_2845,N_1578,N_1545);
xnor U2846 (N_2846,N_1351,N_1144);
and U2847 (N_2847,N_1515,N_1874);
nand U2848 (N_2848,N_1722,N_1098);
and U2849 (N_2849,N_1853,N_1407);
nand U2850 (N_2850,N_1551,N_1450);
nor U2851 (N_2851,N_1564,N_1788);
xnor U2852 (N_2852,N_1094,N_1400);
nand U2853 (N_2853,N_1759,N_1192);
xnor U2854 (N_2854,N_1668,N_1645);
and U2855 (N_2855,N_1296,N_1087);
nor U2856 (N_2856,N_1873,N_1956);
xor U2857 (N_2857,N_1249,N_1365);
and U2858 (N_2858,N_1022,N_1993);
nor U2859 (N_2859,N_1590,N_1440);
xor U2860 (N_2860,N_1471,N_1022);
nor U2861 (N_2861,N_1497,N_1646);
or U2862 (N_2862,N_1266,N_1187);
and U2863 (N_2863,N_1997,N_1376);
xor U2864 (N_2864,N_1360,N_1749);
xor U2865 (N_2865,N_1372,N_1982);
nor U2866 (N_2866,N_1122,N_1144);
and U2867 (N_2867,N_1480,N_1539);
nand U2868 (N_2868,N_1905,N_1913);
or U2869 (N_2869,N_1706,N_1552);
and U2870 (N_2870,N_1098,N_1906);
xnor U2871 (N_2871,N_1924,N_1392);
nor U2872 (N_2872,N_1880,N_1136);
or U2873 (N_2873,N_1879,N_1856);
xnor U2874 (N_2874,N_1931,N_1511);
nand U2875 (N_2875,N_1114,N_1974);
nor U2876 (N_2876,N_1549,N_1360);
nand U2877 (N_2877,N_1682,N_1083);
nor U2878 (N_2878,N_1407,N_1496);
xor U2879 (N_2879,N_1409,N_1788);
or U2880 (N_2880,N_1387,N_1195);
nor U2881 (N_2881,N_1375,N_1920);
nor U2882 (N_2882,N_1489,N_1322);
xor U2883 (N_2883,N_1986,N_1657);
nor U2884 (N_2884,N_1399,N_1340);
and U2885 (N_2885,N_1150,N_1798);
xor U2886 (N_2886,N_1691,N_1784);
xnor U2887 (N_2887,N_1491,N_1989);
nand U2888 (N_2888,N_1553,N_1295);
nand U2889 (N_2889,N_1291,N_1157);
and U2890 (N_2890,N_1946,N_1417);
and U2891 (N_2891,N_1301,N_1426);
xnor U2892 (N_2892,N_1912,N_1923);
xor U2893 (N_2893,N_1129,N_1565);
and U2894 (N_2894,N_1069,N_1386);
xor U2895 (N_2895,N_1410,N_1951);
or U2896 (N_2896,N_1233,N_1798);
and U2897 (N_2897,N_1030,N_1613);
or U2898 (N_2898,N_1301,N_1827);
and U2899 (N_2899,N_1921,N_1140);
or U2900 (N_2900,N_1455,N_1667);
or U2901 (N_2901,N_1921,N_1803);
and U2902 (N_2902,N_1490,N_1129);
or U2903 (N_2903,N_1845,N_1645);
and U2904 (N_2904,N_1577,N_1330);
and U2905 (N_2905,N_1558,N_1313);
or U2906 (N_2906,N_1981,N_1377);
and U2907 (N_2907,N_1841,N_1405);
or U2908 (N_2908,N_1478,N_1867);
nor U2909 (N_2909,N_1429,N_1187);
nor U2910 (N_2910,N_1018,N_1200);
nor U2911 (N_2911,N_1695,N_1312);
or U2912 (N_2912,N_1459,N_1487);
or U2913 (N_2913,N_1185,N_1633);
xor U2914 (N_2914,N_1143,N_1290);
nand U2915 (N_2915,N_1632,N_1715);
and U2916 (N_2916,N_1110,N_1822);
xor U2917 (N_2917,N_1337,N_1952);
xnor U2918 (N_2918,N_1930,N_1533);
xor U2919 (N_2919,N_1620,N_1095);
or U2920 (N_2920,N_1132,N_1539);
and U2921 (N_2921,N_1876,N_1087);
nor U2922 (N_2922,N_1908,N_1635);
nand U2923 (N_2923,N_1711,N_1459);
or U2924 (N_2924,N_1496,N_1045);
or U2925 (N_2925,N_1036,N_1257);
or U2926 (N_2926,N_1208,N_1775);
nor U2927 (N_2927,N_1403,N_1392);
or U2928 (N_2928,N_1470,N_1100);
xnor U2929 (N_2929,N_1097,N_1505);
xor U2930 (N_2930,N_1596,N_1542);
xnor U2931 (N_2931,N_1443,N_1119);
and U2932 (N_2932,N_1097,N_1905);
and U2933 (N_2933,N_1931,N_1988);
or U2934 (N_2934,N_1639,N_1234);
and U2935 (N_2935,N_1348,N_1279);
or U2936 (N_2936,N_1903,N_1858);
nor U2937 (N_2937,N_1329,N_1353);
nor U2938 (N_2938,N_1591,N_1512);
nor U2939 (N_2939,N_1916,N_1266);
and U2940 (N_2940,N_1416,N_1978);
and U2941 (N_2941,N_1467,N_1136);
and U2942 (N_2942,N_1486,N_1233);
nand U2943 (N_2943,N_1377,N_1059);
xor U2944 (N_2944,N_1891,N_1112);
nor U2945 (N_2945,N_1248,N_1845);
nand U2946 (N_2946,N_1278,N_1857);
xor U2947 (N_2947,N_1980,N_1514);
nor U2948 (N_2948,N_1417,N_1471);
and U2949 (N_2949,N_1056,N_1052);
xor U2950 (N_2950,N_1945,N_1884);
nor U2951 (N_2951,N_1482,N_1304);
and U2952 (N_2952,N_1153,N_1810);
xor U2953 (N_2953,N_1703,N_1095);
and U2954 (N_2954,N_1130,N_1960);
nor U2955 (N_2955,N_1354,N_1065);
nand U2956 (N_2956,N_1477,N_1846);
xnor U2957 (N_2957,N_1271,N_1140);
nand U2958 (N_2958,N_1277,N_1921);
nand U2959 (N_2959,N_1819,N_1918);
xor U2960 (N_2960,N_1128,N_1893);
nand U2961 (N_2961,N_1953,N_1662);
and U2962 (N_2962,N_1263,N_1603);
nor U2963 (N_2963,N_1315,N_1392);
nor U2964 (N_2964,N_1250,N_1474);
xnor U2965 (N_2965,N_1102,N_1537);
and U2966 (N_2966,N_1205,N_1363);
nand U2967 (N_2967,N_1433,N_1588);
nor U2968 (N_2968,N_1147,N_1692);
or U2969 (N_2969,N_1268,N_1410);
or U2970 (N_2970,N_1755,N_1632);
nand U2971 (N_2971,N_1070,N_1034);
and U2972 (N_2972,N_1125,N_1454);
or U2973 (N_2973,N_1192,N_1497);
nor U2974 (N_2974,N_1737,N_1090);
nor U2975 (N_2975,N_1413,N_1267);
nor U2976 (N_2976,N_1872,N_1392);
and U2977 (N_2977,N_1613,N_1719);
nand U2978 (N_2978,N_1252,N_1761);
xnor U2979 (N_2979,N_1235,N_1259);
and U2980 (N_2980,N_1228,N_1156);
and U2981 (N_2981,N_1108,N_1997);
nor U2982 (N_2982,N_1358,N_1238);
and U2983 (N_2983,N_1756,N_1549);
and U2984 (N_2984,N_1003,N_1800);
or U2985 (N_2985,N_1189,N_1894);
nor U2986 (N_2986,N_1940,N_1986);
xnor U2987 (N_2987,N_1579,N_1463);
nand U2988 (N_2988,N_1817,N_1230);
xor U2989 (N_2989,N_1168,N_1080);
nand U2990 (N_2990,N_1274,N_1316);
nand U2991 (N_2991,N_1341,N_1477);
and U2992 (N_2992,N_1824,N_1208);
or U2993 (N_2993,N_1235,N_1650);
nand U2994 (N_2994,N_1703,N_1079);
and U2995 (N_2995,N_1817,N_1655);
nand U2996 (N_2996,N_1036,N_1949);
nand U2997 (N_2997,N_1198,N_1919);
nand U2998 (N_2998,N_1942,N_1191);
or U2999 (N_2999,N_1755,N_1094);
nor UO_0 (O_0,N_2784,N_2421);
nor UO_1 (O_1,N_2074,N_2707);
or UO_2 (O_2,N_2390,N_2085);
nor UO_3 (O_3,N_2907,N_2975);
or UO_4 (O_4,N_2989,N_2949);
xnor UO_5 (O_5,N_2146,N_2035);
nand UO_6 (O_6,N_2003,N_2827);
nand UO_7 (O_7,N_2313,N_2518);
nand UO_8 (O_8,N_2498,N_2622);
nor UO_9 (O_9,N_2167,N_2550);
nand UO_10 (O_10,N_2316,N_2459);
and UO_11 (O_11,N_2774,N_2884);
nor UO_12 (O_12,N_2253,N_2575);
nor UO_13 (O_13,N_2903,N_2254);
nand UO_14 (O_14,N_2926,N_2299);
or UO_15 (O_15,N_2011,N_2291);
nand UO_16 (O_16,N_2327,N_2204);
nand UO_17 (O_17,N_2106,N_2581);
nand UO_18 (O_18,N_2611,N_2967);
or UO_19 (O_19,N_2377,N_2862);
or UO_20 (O_20,N_2047,N_2066);
nor UO_21 (O_21,N_2534,N_2198);
or UO_22 (O_22,N_2898,N_2173);
and UO_23 (O_23,N_2337,N_2803);
nor UO_24 (O_24,N_2347,N_2213);
or UO_25 (O_25,N_2778,N_2294);
xor UO_26 (O_26,N_2163,N_2469);
and UO_27 (O_27,N_2932,N_2295);
or UO_28 (O_28,N_2144,N_2482);
and UO_29 (O_29,N_2983,N_2491);
nor UO_30 (O_30,N_2570,N_2814);
xnor UO_31 (O_31,N_2566,N_2312);
nand UO_32 (O_32,N_2441,N_2950);
and UO_33 (O_33,N_2417,N_2571);
or UO_34 (O_34,N_2092,N_2252);
or UO_35 (O_35,N_2118,N_2639);
nand UO_36 (O_36,N_2798,N_2278);
nor UO_37 (O_37,N_2166,N_2634);
nand UO_38 (O_38,N_2062,N_2083);
or UO_39 (O_39,N_2483,N_2363);
or UO_40 (O_40,N_2378,N_2471);
nor UO_41 (O_41,N_2560,N_2045);
nor UO_42 (O_42,N_2015,N_2947);
and UO_43 (O_43,N_2265,N_2524);
nor UO_44 (O_44,N_2485,N_2138);
or UO_45 (O_45,N_2957,N_2473);
and UO_46 (O_46,N_2683,N_2755);
and UO_47 (O_47,N_2564,N_2461);
xor UO_48 (O_48,N_2296,N_2335);
nand UO_49 (O_49,N_2854,N_2197);
and UO_50 (O_50,N_2667,N_2355);
or UO_51 (O_51,N_2746,N_2897);
and UO_52 (O_52,N_2002,N_2311);
nor UO_53 (O_53,N_2585,N_2141);
nand UO_54 (O_54,N_2972,N_2952);
and UO_55 (O_55,N_2137,N_2054);
nand UO_56 (O_56,N_2855,N_2394);
nor UO_57 (O_57,N_2958,N_2598);
and UO_58 (O_58,N_2732,N_2470);
or UO_59 (O_59,N_2542,N_2124);
nor UO_60 (O_60,N_2492,N_2569);
or UO_61 (O_61,N_2314,N_2782);
nand UO_62 (O_62,N_2224,N_2336);
xor UO_63 (O_63,N_2259,N_2438);
nor UO_64 (O_64,N_2371,N_2572);
nor UO_65 (O_65,N_2848,N_2966);
and UO_66 (O_66,N_2396,N_2332);
nand UO_67 (O_67,N_2097,N_2077);
or UO_68 (O_68,N_2935,N_2899);
and UO_69 (O_69,N_2747,N_2728);
nor UO_70 (O_70,N_2619,N_2623);
nor UO_71 (O_71,N_2756,N_2554);
nand UO_72 (O_72,N_2496,N_2889);
nand UO_73 (O_73,N_2751,N_2970);
nor UO_74 (O_74,N_2817,N_2001);
nand UO_75 (O_75,N_2271,N_2123);
xor UO_76 (O_76,N_2754,N_2519);
nand UO_77 (O_77,N_2229,N_2646);
nand UO_78 (O_78,N_2494,N_2551);
or UO_79 (O_79,N_2759,N_2275);
and UO_80 (O_80,N_2321,N_2087);
or UO_81 (O_81,N_2068,N_2109);
nor UO_82 (O_82,N_2257,N_2379);
xnor UO_83 (O_83,N_2160,N_2238);
xnor UO_84 (O_84,N_2822,N_2537);
xnor UO_85 (O_85,N_2320,N_2049);
nand UO_86 (O_86,N_2654,N_2940);
nand UO_87 (O_87,N_2480,N_2221);
nand UO_88 (O_88,N_2834,N_2162);
xor UO_89 (O_89,N_2497,N_2158);
or UO_90 (O_90,N_2752,N_2093);
and UO_91 (O_91,N_2693,N_2182);
nor UO_92 (O_92,N_2446,N_2681);
nand UO_93 (O_93,N_2445,N_2710);
xor UO_94 (O_94,N_2112,N_2069);
and UO_95 (O_95,N_2214,N_2104);
nor UO_96 (O_96,N_2770,N_2578);
nor UO_97 (O_97,N_2994,N_2190);
nor UO_98 (O_98,N_2308,N_2328);
xor UO_99 (O_99,N_2895,N_2736);
and UO_100 (O_100,N_2535,N_2247);
nand UO_101 (O_101,N_2196,N_2200);
and UO_102 (O_102,N_2960,N_2946);
xor UO_103 (O_103,N_2334,N_2339);
and UO_104 (O_104,N_2107,N_2908);
or UO_105 (O_105,N_2301,N_2342);
or UO_106 (O_106,N_2050,N_2912);
xnor UO_107 (O_107,N_2995,N_2303);
xnor UO_108 (O_108,N_2630,N_2323);
nand UO_109 (O_109,N_2694,N_2892);
xor UO_110 (O_110,N_2675,N_2169);
nand UO_111 (O_111,N_2715,N_2526);
nand UO_112 (O_112,N_2738,N_2719);
xor UO_113 (O_113,N_2217,N_2875);
nor UO_114 (O_114,N_2815,N_2464);
nand UO_115 (O_115,N_2955,N_2711);
or UO_116 (O_116,N_2629,N_2541);
and UO_117 (O_117,N_2743,N_2375);
nor UO_118 (O_118,N_2772,N_2090);
or UO_119 (O_119,N_2165,N_2527);
and UO_120 (O_120,N_2962,N_2409);
xnor UO_121 (O_121,N_2650,N_2555);
or UO_122 (O_122,N_2448,N_2606);
or UO_123 (O_123,N_2603,N_2757);
xor UO_124 (O_124,N_2724,N_2310);
or UO_125 (O_125,N_2956,N_2830);
or UO_126 (O_126,N_2988,N_2913);
and UO_127 (O_127,N_2319,N_2270);
and UO_128 (O_128,N_2763,N_2382);
and UO_129 (O_129,N_2626,N_2997);
xnor UO_130 (O_130,N_2023,N_2134);
or UO_131 (O_131,N_2348,N_2804);
nor UO_132 (O_132,N_2258,N_2920);
nand UO_133 (O_133,N_2722,N_2070);
xnor UO_134 (O_134,N_2510,N_2644);
nand UO_135 (O_135,N_2432,N_2261);
nor UO_136 (O_136,N_2289,N_2837);
nand UO_137 (O_137,N_2628,N_2168);
or UO_138 (O_138,N_2234,N_2431);
xnor UO_139 (O_139,N_2358,N_2742);
xnor UO_140 (O_140,N_2621,N_2596);
nor UO_141 (O_141,N_2099,N_2574);
or UO_142 (O_142,N_2018,N_2937);
or UO_143 (O_143,N_2553,N_2027);
nor UO_144 (O_144,N_2672,N_2691);
nor UO_145 (O_145,N_2102,N_2178);
or UO_146 (O_146,N_2914,N_2515);
xor UO_147 (O_147,N_2051,N_2543);
and UO_148 (O_148,N_2364,N_2076);
nand UO_149 (O_149,N_2046,N_2256);
nand UO_150 (O_150,N_2523,N_2468);
nand UO_151 (O_151,N_2304,N_2863);
nand UO_152 (O_152,N_2305,N_2108);
xnor UO_153 (O_153,N_2893,N_2272);
and UO_154 (O_154,N_2489,N_2887);
xor UO_155 (O_155,N_2591,N_2548);
or UO_156 (O_156,N_2031,N_2058);
xnor UO_157 (O_157,N_2655,N_2164);
xor UO_158 (O_158,N_2996,N_2269);
nand UO_159 (O_159,N_2451,N_2645);
nand UO_160 (O_160,N_2762,N_2367);
nand UO_161 (O_161,N_2096,N_2404);
nand UO_162 (O_162,N_2232,N_2333);
nor UO_163 (O_163,N_2401,N_2831);
xnor UO_164 (O_164,N_2065,N_2936);
nor UO_165 (O_165,N_2450,N_2007);
and UO_166 (O_166,N_2943,N_2882);
xor UO_167 (O_167,N_2153,N_2495);
nor UO_168 (O_168,N_2505,N_2544);
or UO_169 (O_169,N_2813,N_2753);
xor UO_170 (O_170,N_2359,N_2260);
and UO_171 (O_171,N_2536,N_2079);
and UO_172 (O_172,N_2465,N_2857);
nor UO_173 (O_173,N_2040,N_2666);
or UO_174 (O_174,N_2717,N_2398);
and UO_175 (O_175,N_2520,N_2663);
nand UO_176 (O_176,N_2389,N_2900);
and UO_177 (O_177,N_2845,N_2749);
or UO_178 (O_178,N_2171,N_2352);
nand UO_179 (O_179,N_2905,N_2048);
and UO_180 (O_180,N_2677,N_2640);
and UO_181 (O_181,N_2826,N_2791);
xor UO_182 (O_182,N_2664,N_2730);
nor UO_183 (O_183,N_2142,N_2540);
or UO_184 (O_184,N_2608,N_2202);
or UO_185 (O_185,N_2959,N_2727);
nor UO_186 (O_186,N_2739,N_2503);
nor UO_187 (O_187,N_2825,N_2678);
and UO_188 (O_188,N_2865,N_2514);
and UO_189 (O_189,N_2979,N_2929);
xnor UO_190 (O_190,N_2277,N_2248);
or UO_191 (O_191,N_2411,N_2105);
nand UO_192 (O_192,N_2840,N_2467);
and UO_193 (O_193,N_2869,N_2181);
and UO_194 (O_194,N_2705,N_2546);
nand UO_195 (O_195,N_2241,N_2531);
nor UO_196 (O_196,N_2635,N_2405);
xnor UO_197 (O_197,N_2227,N_2853);
or UO_198 (O_198,N_2129,N_2004);
xnor UO_199 (O_199,N_2590,N_2504);
and UO_200 (O_200,N_2251,N_2901);
or UO_201 (O_201,N_2407,N_2356);
and UO_202 (O_202,N_2330,N_2156);
and UO_203 (O_203,N_2750,N_2010);
nor UO_204 (O_204,N_2442,N_2285);
xor UO_205 (O_205,N_2891,N_2595);
nand UO_206 (O_206,N_2264,N_2673);
and UO_207 (O_207,N_2557,N_2340);
nor UO_208 (O_208,N_2771,N_2916);
nor UO_209 (O_209,N_2435,N_2648);
xor UO_210 (O_210,N_2075,N_2582);
nor UO_211 (O_211,N_2951,N_2013);
or UO_212 (O_212,N_2506,N_2682);
nor UO_213 (O_213,N_2766,N_2306);
xor UO_214 (O_214,N_2043,N_2059);
nor UO_215 (O_215,N_2974,N_2419);
or UO_216 (O_216,N_2687,N_2381);
nand UO_217 (O_217,N_2369,N_2858);
nor UO_218 (O_218,N_2529,N_2346);
and UO_219 (O_219,N_2242,N_2315);
nand UO_220 (O_220,N_2343,N_2511);
xor UO_221 (O_221,N_2872,N_2636);
nand UO_222 (O_222,N_2244,N_2216);
nand UO_223 (O_223,N_2767,N_2425);
or UO_224 (O_224,N_2126,N_2685);
xor UO_225 (O_225,N_2835,N_2925);
or UO_226 (O_226,N_2478,N_2326);
xnor UO_227 (O_227,N_2282,N_2273);
or UO_228 (O_228,N_2225,N_2917);
and UO_229 (O_229,N_2063,N_2741);
nor UO_230 (O_230,N_2362,N_2758);
xnor UO_231 (O_231,N_2292,N_2584);
nor UO_232 (O_232,N_2185,N_2233);
and UO_233 (O_233,N_2987,N_2056);
nand UO_234 (O_234,N_2808,N_2860);
or UO_235 (O_235,N_2821,N_2931);
nand UO_236 (O_236,N_2424,N_2796);
and UO_237 (O_237,N_2942,N_2006);
nand UO_238 (O_238,N_2880,N_2787);
nor UO_239 (O_239,N_2964,N_2961);
nand UO_240 (O_240,N_2816,N_2706);
nor UO_241 (O_241,N_2368,N_2061);
nor UO_242 (O_242,N_2392,N_2802);
nor UO_243 (O_243,N_2288,N_2680);
xnor UO_244 (O_244,N_2921,N_2737);
and UO_245 (O_245,N_2973,N_2426);
nor UO_246 (O_246,N_2610,N_2674);
or UO_247 (O_247,N_2600,N_2721);
and UO_248 (O_248,N_2302,N_2226);
xor UO_249 (O_249,N_2422,N_2761);
and UO_250 (O_250,N_2945,N_2360);
nand UO_251 (O_251,N_2692,N_2089);
or UO_252 (O_252,N_2053,N_2953);
nor UO_253 (O_253,N_2274,N_2859);
nand UO_254 (O_254,N_2558,N_2184);
and UO_255 (O_255,N_2602,N_2904);
nor UO_256 (O_256,N_2538,N_2911);
xnor UO_257 (O_257,N_2243,N_2532);
nand UO_258 (O_258,N_2206,N_2397);
nand UO_259 (O_259,N_2509,N_2688);
xnor UO_260 (O_260,N_2818,N_2843);
nand UO_261 (O_261,N_2179,N_2652);
nor UO_262 (O_262,N_2170,N_2266);
or UO_263 (O_263,N_2748,N_2086);
and UO_264 (O_264,N_2765,N_2522);
and UO_265 (O_265,N_2466,N_2698);
nand UO_266 (O_266,N_2573,N_2344);
nor UO_267 (O_267,N_2117,N_2428);
and UO_268 (O_268,N_2856,N_2395);
or UO_269 (O_269,N_2740,N_2189);
and UO_270 (O_270,N_2712,N_2811);
nor UO_271 (O_271,N_2601,N_2030);
xor UO_272 (O_272,N_2130,N_2172);
or UO_273 (O_273,N_2684,N_2769);
or UO_274 (O_274,N_2161,N_2850);
or UO_275 (O_275,N_2472,N_2177);
nor UO_276 (O_276,N_2071,N_2923);
nand UO_277 (O_277,N_2453,N_2976);
nor UO_278 (O_278,N_2607,N_2038);
and UO_279 (O_279,N_2157,N_2841);
nor UO_280 (O_280,N_2508,N_2576);
nand UO_281 (O_281,N_2174,N_2094);
or UO_282 (O_282,N_2187,N_2708);
xor UO_283 (O_283,N_2113,N_2036);
nor UO_284 (O_284,N_2776,N_2999);
or UO_285 (O_285,N_2888,N_2110);
and UO_286 (O_286,N_2434,N_2080);
nor UO_287 (O_287,N_2222,N_2462);
nand UO_288 (O_288,N_2703,N_2833);
or UO_289 (O_289,N_2014,N_2021);
or UO_290 (O_290,N_2842,N_2350);
nand UO_291 (O_291,N_2883,N_2902);
nand UO_292 (O_292,N_2832,N_2781);
or UO_293 (O_293,N_2298,N_2205);
nor UO_294 (O_294,N_2279,N_2500);
nor UO_295 (O_295,N_2072,N_2060);
or UO_296 (O_296,N_2809,N_2208);
nand UO_297 (O_297,N_2345,N_2481);
nand UO_298 (O_298,N_2443,N_2121);
and UO_299 (O_299,N_2354,N_2414);
or UO_300 (O_300,N_2250,N_2718);
or UO_301 (O_301,N_2868,N_2433);
or UO_302 (O_302,N_2111,N_2410);
nor UO_303 (O_303,N_2331,N_2662);
and UO_304 (O_304,N_2773,N_2486);
and UO_305 (O_305,N_2507,N_2985);
nand UO_306 (O_306,N_2700,N_2649);
nor UO_307 (O_307,N_2246,N_2633);
nand UO_308 (O_308,N_2016,N_2638);
xor UO_309 (O_309,N_2659,N_2183);
xnor UO_310 (O_310,N_2729,N_2287);
xnor UO_311 (O_311,N_2436,N_2372);
or UO_312 (O_312,N_2262,N_2982);
or UO_313 (O_313,N_2230,N_2317);
nand UO_314 (O_314,N_2695,N_2801);
and UO_315 (O_315,N_2552,N_2697);
nand UO_316 (O_316,N_2679,N_2454);
nor UO_317 (O_317,N_2968,N_2119);
nand UO_318 (O_318,N_2012,N_2657);
and UO_319 (O_319,N_2406,N_2792);
or UO_320 (O_320,N_2563,N_2642);
xnor UO_321 (O_321,N_2670,N_2586);
or UO_322 (O_322,N_2874,N_2627);
and UO_323 (O_323,N_2567,N_2122);
and UO_324 (O_324,N_2026,N_2267);
and UO_325 (O_325,N_2487,N_2440);
nand UO_326 (O_326,N_2151,N_2095);
nor UO_327 (O_327,N_2993,N_2041);
xor UO_328 (O_328,N_2699,N_2651);
nand UO_329 (O_329,N_2374,N_2823);
and UO_330 (O_330,N_2385,N_2039);
or UO_331 (O_331,N_2415,N_2188);
xor UO_332 (O_332,N_2399,N_2307);
and UO_333 (O_333,N_2203,N_2604);
xor UO_334 (O_334,N_2449,N_2133);
nand UO_335 (O_335,N_2668,N_2788);
and UO_336 (O_336,N_2579,N_2702);
and UO_337 (O_337,N_2933,N_2701);
nor UO_338 (O_338,N_2484,N_2290);
nor UO_339 (O_339,N_2139,N_2790);
or UO_340 (O_340,N_2365,N_2609);
nand UO_341 (O_341,N_2829,N_2067);
xor UO_342 (O_342,N_2851,N_2806);
and UO_343 (O_343,N_2844,N_2616);
nor UO_344 (O_344,N_2615,N_2896);
xor UO_345 (O_345,N_2427,N_2159);
nor UO_346 (O_346,N_2044,N_2280);
and UO_347 (O_347,N_2998,N_2236);
nand UO_348 (O_348,N_2284,N_2879);
nor UO_349 (O_349,N_2091,N_2735);
xor UO_350 (O_350,N_2559,N_2000);
and UO_351 (O_351,N_2025,N_2073);
nor UO_352 (O_352,N_2034,N_2132);
nand UO_353 (O_353,N_2231,N_2114);
or UO_354 (O_354,N_2775,N_2941);
nor UO_355 (O_355,N_2383,N_2218);
nand UO_356 (O_356,N_2605,N_2812);
and UO_357 (O_357,N_2599,N_2587);
nor UO_358 (O_358,N_2211,N_2733);
xor UO_359 (O_359,N_2881,N_2475);
nand UO_360 (O_360,N_2393,N_2447);
or UO_361 (O_361,N_2556,N_2631);
and UO_362 (O_362,N_2704,N_2847);
and UO_363 (O_363,N_2136,N_2992);
or UO_364 (O_364,N_2660,N_2521);
xor UO_365 (O_365,N_2493,N_2934);
or UO_366 (O_366,N_2361,N_2918);
and UO_367 (O_367,N_2191,N_2836);
nand UO_368 (O_368,N_2785,N_2539);
nor UO_369 (O_369,N_2223,N_2263);
and UO_370 (O_370,N_2871,N_2488);
nor UO_371 (O_371,N_2661,N_2696);
xor UO_372 (O_372,N_2780,N_2318);
xnor UO_373 (O_373,N_2745,N_2686);
nand UO_374 (O_374,N_2910,N_2437);
nand UO_375 (O_375,N_2986,N_2131);
or UO_376 (O_376,N_2807,N_2512);
and UO_377 (O_377,N_2789,N_2873);
and UO_378 (O_378,N_2005,N_2212);
xor UO_379 (O_379,N_2653,N_2456);
and UO_380 (O_380,N_2810,N_2423);
nor UO_381 (O_381,N_2846,N_2154);
nand UO_382 (O_382,N_2176,N_2516);
and UO_383 (O_383,N_2199,N_2209);
or UO_384 (O_384,N_2547,N_2180);
or UO_385 (O_385,N_2017,N_2255);
xor UO_386 (O_386,N_2101,N_2408);
xnor UO_387 (O_387,N_2530,N_2786);
and UO_388 (O_388,N_2418,N_2624);
nor UO_389 (O_389,N_2870,N_2944);
and UO_390 (O_390,N_2613,N_2924);
nor UO_391 (O_391,N_2145,N_2477);
nand UO_392 (O_392,N_2939,N_2819);
and UO_393 (O_393,N_2890,N_2460);
xnor UO_394 (O_394,N_2400,N_2720);
nand UO_395 (O_395,N_2797,N_2768);
xnor UO_396 (O_396,N_2948,N_2391);
or UO_397 (O_397,N_2990,N_2353);
nor UO_398 (O_398,N_2828,N_2024);
and UO_399 (O_399,N_2341,N_2052);
xor UO_400 (O_400,N_2127,N_2637);
xnor UO_401 (O_401,N_2577,N_2386);
nand UO_402 (O_402,N_2594,N_2713);
nand UO_403 (O_403,N_2963,N_2245);
and UO_404 (O_404,N_2632,N_2193);
or UO_405 (O_405,N_2689,N_2019);
and UO_406 (O_406,N_2115,N_2351);
nor UO_407 (O_407,N_2954,N_2877);
or UO_408 (O_408,N_2726,N_2370);
and UO_409 (O_409,N_2593,N_2658);
xnor UO_410 (O_410,N_2501,N_2457);
xnor UO_411 (O_411,N_2149,N_2349);
nand UO_412 (O_412,N_2420,N_2731);
or UO_413 (O_413,N_2612,N_2201);
nor UO_414 (O_414,N_2867,N_2777);
and UO_415 (O_415,N_2444,N_2479);
nor UO_416 (O_416,N_2592,N_2366);
or UO_417 (O_417,N_2978,N_2597);
and UO_418 (O_418,N_2965,N_2324);
nand UO_419 (O_419,N_2140,N_2517);
and UO_420 (O_420,N_2714,N_2671);
nand UO_421 (O_421,N_2103,N_2981);
xnor UO_422 (O_422,N_2276,N_2458);
xnor UO_423 (O_423,N_2565,N_2502);
and UO_424 (O_424,N_2549,N_2866);
nand UO_425 (O_425,N_2152,N_2969);
or UO_426 (O_426,N_2793,N_2143);
nand UO_427 (O_427,N_2885,N_2894);
or UO_428 (O_428,N_2413,N_2135);
xor UO_429 (O_429,N_2033,N_2525);
xnor UO_430 (O_430,N_2322,N_2228);
and UO_431 (O_431,N_2128,N_2744);
and UO_432 (O_432,N_2064,N_2081);
or UO_433 (O_433,N_2150,N_2915);
xnor UO_434 (O_434,N_2991,N_2838);
nor UO_435 (O_435,N_2240,N_2120);
and UO_436 (O_436,N_2971,N_2620);
or UO_437 (O_437,N_2373,N_2416);
and UO_438 (O_438,N_2009,N_2309);
and UO_439 (O_439,N_2820,N_2561);
and UO_440 (O_440,N_2864,N_2568);
xnor UO_441 (O_441,N_2676,N_2919);
nand UO_442 (O_442,N_2799,N_2100);
xor UO_443 (O_443,N_2452,N_2618);
and UO_444 (O_444,N_2562,N_2429);
nor UO_445 (O_445,N_2037,N_2906);
xor UO_446 (O_446,N_2283,N_2928);
xor UO_447 (O_447,N_2078,N_2116);
nor UO_448 (O_448,N_2499,N_2725);
nor UO_449 (O_449,N_2249,N_2032);
or UO_450 (O_450,N_2617,N_2125);
nand UO_451 (O_451,N_2474,N_2175);
xnor UO_452 (O_452,N_2220,N_2210);
or UO_453 (O_453,N_2656,N_2380);
nand UO_454 (O_454,N_2088,N_2297);
nand UO_455 (O_455,N_2357,N_2082);
nand UO_456 (O_456,N_2665,N_2455);
and UO_457 (O_457,N_2148,N_2824);
nand UO_458 (O_458,N_2300,N_2528);
xor UO_459 (O_459,N_2186,N_2977);
and UO_460 (O_460,N_2057,N_2690);
nor UO_461 (O_461,N_2403,N_2876);
or UO_462 (O_462,N_2641,N_2476);
nor UO_463 (O_463,N_2839,N_2192);
nor UO_464 (O_464,N_2022,N_2764);
or UO_465 (O_465,N_2194,N_2338);
nor UO_466 (O_466,N_2878,N_2388);
or UO_467 (O_467,N_2195,N_2028);
nand UO_468 (O_468,N_2439,N_2580);
or UO_469 (O_469,N_2589,N_2029);
nor UO_470 (O_470,N_2042,N_2215);
or UO_471 (O_471,N_2909,N_2155);
nand UO_472 (O_472,N_2643,N_2545);
nor UO_473 (O_473,N_2625,N_2760);
nor UO_474 (O_474,N_2861,N_2239);
nor UO_475 (O_475,N_2513,N_2779);
xnor UO_476 (O_476,N_2723,N_2583);
nand UO_477 (O_477,N_2533,N_2852);
xnor UO_478 (O_478,N_2376,N_2235);
nor UO_479 (O_479,N_2055,N_2805);
nand UO_480 (O_480,N_2794,N_2147);
nand UO_481 (O_481,N_2980,N_2084);
xnor UO_482 (O_482,N_2849,N_2927);
nor UO_483 (O_483,N_2647,N_2886);
xor UO_484 (O_484,N_2938,N_2384);
nor UO_485 (O_485,N_2329,N_2281);
nand UO_486 (O_486,N_2207,N_2098);
and UO_487 (O_487,N_2387,N_2219);
nand UO_488 (O_488,N_2268,N_2463);
or UO_489 (O_489,N_2402,N_2286);
or UO_490 (O_490,N_2734,N_2716);
nand UO_491 (O_491,N_2293,N_2795);
or UO_492 (O_492,N_2412,N_2800);
or UO_493 (O_493,N_2430,N_2930);
xnor UO_494 (O_494,N_2237,N_2008);
or UO_495 (O_495,N_2922,N_2669);
and UO_496 (O_496,N_2588,N_2325);
nand UO_497 (O_497,N_2709,N_2984);
or UO_498 (O_498,N_2783,N_2020);
and UO_499 (O_499,N_2490,N_2614);
endmodule