module basic_2000_20000_2500_80_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_416,In_1752);
nor U1 (N_1,In_437,In_155);
nand U2 (N_2,In_674,In_1546);
and U3 (N_3,In_1204,In_275);
or U4 (N_4,In_915,In_803);
nor U5 (N_5,In_1938,In_693);
and U6 (N_6,In_448,In_1469);
and U7 (N_7,In_341,In_1838);
xor U8 (N_8,In_852,In_1506);
and U9 (N_9,In_862,In_1231);
nor U10 (N_10,In_549,In_1848);
xnor U11 (N_11,In_1061,In_1819);
nor U12 (N_12,In_978,In_1889);
and U13 (N_13,In_1324,In_1842);
or U14 (N_14,In_991,In_1120);
nor U15 (N_15,In_547,In_1106);
nand U16 (N_16,In_53,In_347);
or U17 (N_17,In_1937,In_1530);
and U18 (N_18,In_1568,In_114);
nand U19 (N_19,In_624,In_376);
and U20 (N_20,In_1222,In_1843);
or U21 (N_21,In_491,In_112);
or U22 (N_22,In_1456,In_946);
xor U23 (N_23,In_1095,In_1719);
or U24 (N_24,In_717,In_1683);
nand U25 (N_25,In_378,In_1959);
nand U26 (N_26,In_1646,In_144);
nor U27 (N_27,In_1053,In_696);
and U28 (N_28,In_1138,In_1229);
nand U29 (N_29,In_1513,In_1969);
nand U30 (N_30,In_1825,In_1031);
and U31 (N_31,In_392,In_983);
xnor U32 (N_32,In_1894,In_1987);
nor U33 (N_33,In_1455,In_1201);
nand U34 (N_34,In_1339,In_75);
nand U35 (N_35,In_6,In_922);
nand U36 (N_36,In_1474,In_1774);
nor U37 (N_37,In_1385,In_499);
xor U38 (N_38,In_1706,In_359);
xor U39 (N_39,In_50,In_286);
and U40 (N_40,In_1746,In_641);
nand U41 (N_41,In_1160,In_1432);
nand U42 (N_42,In_1383,In_526);
nor U43 (N_43,In_1214,In_365);
or U44 (N_44,In_1321,In_633);
nor U45 (N_45,In_1915,In_190);
and U46 (N_46,In_408,In_889);
nor U47 (N_47,In_330,In_1495);
xor U48 (N_48,In_737,In_686);
nor U49 (N_49,In_1558,In_1669);
nor U50 (N_50,In_412,In_1805);
or U51 (N_51,In_615,In_593);
nand U52 (N_52,In_403,In_968);
nor U53 (N_53,In_800,In_1493);
or U54 (N_54,In_1491,In_896);
and U55 (N_55,In_1677,In_524);
or U56 (N_56,In_1426,In_82);
and U57 (N_57,In_1407,In_644);
and U58 (N_58,In_570,In_996);
nor U59 (N_59,In_442,In_296);
xnor U60 (N_60,In_1598,In_1145);
and U61 (N_61,In_473,In_1640);
and U62 (N_62,In_785,In_1500);
nor U63 (N_63,In_1166,In_1748);
xnor U64 (N_64,In_1662,In_1689);
nor U65 (N_65,In_1760,In_701);
nor U66 (N_66,In_332,In_1566);
or U67 (N_67,In_668,In_1139);
or U68 (N_68,In_346,In_804);
nor U69 (N_69,In_35,In_1823);
nand U70 (N_70,In_410,In_1860);
and U71 (N_71,In_1758,In_367);
nand U72 (N_72,In_481,In_160);
nor U73 (N_73,In_444,In_979);
xnor U74 (N_74,In_1944,In_1520);
and U75 (N_75,In_154,In_1236);
nor U76 (N_76,In_1319,In_1745);
nor U77 (N_77,In_81,In_1991);
or U78 (N_78,In_1129,In_1384);
or U79 (N_79,In_368,In_1526);
and U80 (N_80,In_370,In_828);
or U81 (N_81,In_1173,In_1066);
and U82 (N_82,In_727,In_1377);
xnor U83 (N_83,In_1498,In_1639);
nand U84 (N_84,In_363,In_1503);
and U85 (N_85,In_987,In_925);
or U86 (N_86,In_892,In_1133);
and U87 (N_87,In_322,In_1092);
nor U88 (N_88,In_298,In_1686);
nor U89 (N_89,In_579,In_1291);
nand U90 (N_90,In_1835,In_1128);
or U91 (N_91,In_2,In_169);
and U92 (N_92,In_1325,In_1056);
or U93 (N_93,In_1542,In_588);
or U94 (N_94,In_1370,In_167);
xnor U95 (N_95,In_951,In_245);
or U96 (N_96,In_1365,In_117);
and U97 (N_97,In_916,In_1684);
and U98 (N_98,In_517,In_1673);
or U99 (N_99,In_1518,In_261);
and U100 (N_100,In_1397,In_1100);
or U101 (N_101,In_1089,In_1911);
xnor U102 (N_102,In_890,In_699);
or U103 (N_103,In_501,In_1146);
xnor U104 (N_104,In_830,In_116);
and U105 (N_105,In_119,In_1647);
or U106 (N_106,In_527,In_1317);
nand U107 (N_107,In_113,In_23);
and U108 (N_108,In_1876,In_1747);
or U109 (N_109,In_1586,In_465);
xnor U110 (N_110,In_1979,In_533);
nor U111 (N_111,In_125,In_789);
nor U112 (N_112,In_1466,In_1151);
xor U113 (N_113,In_1625,In_1094);
and U114 (N_114,In_1282,In_352);
nor U115 (N_115,In_1452,In_54);
nor U116 (N_116,In_1135,In_515);
nand U117 (N_117,In_761,In_1014);
nor U118 (N_118,In_1028,In_536);
nand U119 (N_119,In_1414,In_1970);
and U120 (N_120,In_1112,In_1699);
xnor U121 (N_121,In_1104,In_1641);
nor U122 (N_122,In_1223,In_430);
or U123 (N_123,In_1696,In_1334);
xor U124 (N_124,In_159,In_120);
xnor U125 (N_125,In_1422,In_1951);
nand U126 (N_126,In_1117,In_815);
nand U127 (N_127,In_1124,In_999);
and U128 (N_128,In_10,In_939);
and U129 (N_129,In_1517,In_1965);
or U130 (N_130,In_1603,In_426);
and U131 (N_131,In_1863,In_1582);
xnor U132 (N_132,In_1181,In_288);
or U133 (N_133,In_1149,In_1921);
nand U134 (N_134,In_49,In_602);
nand U135 (N_135,In_1333,In_314);
xnor U136 (N_136,In_324,In_1490);
and U137 (N_137,In_1896,In_19);
nor U138 (N_138,In_1875,In_1999);
nand U139 (N_139,In_351,In_630);
nor U140 (N_140,In_1026,In_1754);
or U141 (N_141,In_395,In_1849);
xnor U142 (N_142,In_1962,In_257);
nand U143 (N_143,In_512,In_886);
or U144 (N_144,In_301,In_1034);
nand U145 (N_145,In_1961,In_1424);
nor U146 (N_146,In_1230,In_59);
nand U147 (N_147,In_1008,In_210);
xor U148 (N_148,In_1556,In_614);
nand U149 (N_149,In_580,In_379);
nor U150 (N_150,In_1733,In_72);
and U151 (N_151,In_755,In_763);
nand U152 (N_152,In_1868,In_46);
or U153 (N_153,In_640,In_1926);
nand U154 (N_154,In_265,In_1039);
nand U155 (N_155,In_1716,In_438);
or U156 (N_156,In_1033,In_254);
xnor U157 (N_157,In_1820,In_20);
or U158 (N_158,In_478,In_173);
or U159 (N_159,In_813,In_1903);
xor U160 (N_160,In_494,In_213);
xor U161 (N_161,In_855,In_903);
nor U162 (N_162,In_1459,In_1775);
xnor U163 (N_163,In_1076,In_511);
nor U164 (N_164,In_217,In_94);
xnor U165 (N_165,In_793,In_425);
nor U166 (N_166,In_1182,In_260);
nor U167 (N_167,In_1416,In_711);
nor U168 (N_168,In_1001,In_1580);
and U169 (N_169,In_394,In_1990);
nand U170 (N_170,In_1192,In_1943);
xor U171 (N_171,In_1612,In_543);
and U172 (N_172,In_887,In_777);
or U173 (N_173,In_1679,In_1275);
xnor U174 (N_174,In_456,In_1931);
nor U175 (N_175,In_1750,In_1137);
or U176 (N_176,In_17,In_436);
xnor U177 (N_177,In_269,In_719);
nand U178 (N_178,In_1090,In_1767);
nand U179 (N_179,In_566,In_441);
nand U180 (N_180,In_1537,In_486);
nand U181 (N_181,In_816,In_1572);
xnor U182 (N_182,In_534,In_1188);
or U183 (N_183,In_710,In_1815);
nand U184 (N_184,In_608,In_1308);
nor U185 (N_185,In_1501,In_1457);
nand U186 (N_186,In_1349,In_728);
nand U187 (N_187,In_1912,In_37);
nor U188 (N_188,In_594,In_483);
nor U189 (N_189,In_328,In_1358);
xnor U190 (N_190,In_241,In_1771);
nor U191 (N_191,In_1839,In_1300);
or U192 (N_192,In_1854,In_1132);
or U193 (N_193,In_1707,In_1957);
xor U194 (N_194,In_956,In_1796);
xnor U195 (N_195,In_1030,In_986);
xor U196 (N_196,In_949,In_846);
or U197 (N_197,In_1035,In_1613);
xnor U198 (N_198,In_636,In_222);
nor U199 (N_199,In_786,In_1272);
xor U200 (N_200,In_598,In_1451);
and U201 (N_201,In_1899,In_869);
nor U202 (N_202,In_1263,In_135);
nand U203 (N_203,In_1447,In_329);
and U204 (N_204,In_1007,In_805);
xnor U205 (N_205,In_387,In_1461);
nand U206 (N_206,In_1338,In_545);
nor U207 (N_207,In_750,In_1917);
nor U208 (N_208,In_758,In_958);
or U209 (N_209,In_305,In_888);
xnor U210 (N_210,In_860,In_858);
nor U211 (N_211,In_504,In_854);
or U212 (N_212,In_694,In_548);
or U213 (N_213,In_802,In_1477);
xnor U214 (N_214,In_205,In_1265);
xor U215 (N_215,In_1108,In_791);
or U216 (N_216,In_1623,In_386);
nor U217 (N_217,In_518,In_964);
xnor U218 (N_218,In_492,In_1994);
nor U219 (N_219,In_1665,In_33);
nand U220 (N_220,In_1786,In_1968);
and U221 (N_221,In_661,In_1430);
nand U222 (N_222,In_965,In_1855);
and U223 (N_223,In_1354,In_1885);
xor U224 (N_224,In_189,In_1788);
nand U225 (N_225,In_1023,In_806);
xnor U226 (N_226,In_311,In_4);
nand U227 (N_227,In_1102,In_262);
nand U228 (N_228,In_204,In_43);
xor U229 (N_229,In_271,In_1293);
and U230 (N_230,In_377,In_1794);
nand U231 (N_231,In_884,In_1276);
and U232 (N_232,In_1438,In_402);
or U233 (N_233,In_1434,In_629);
nor U234 (N_234,In_1605,In_1047);
or U235 (N_235,In_1922,In_1828);
or U236 (N_236,In_894,In_954);
nand U237 (N_237,In_603,In_1059);
or U238 (N_238,In_1392,In_1867);
nand U239 (N_239,In_1267,In_775);
and U240 (N_240,In_1727,In_776);
nand U241 (N_241,In_52,In_1080);
and U242 (N_242,In_1806,In_199);
or U243 (N_243,In_1783,In_1992);
xnor U244 (N_244,In_509,In_1525);
and U245 (N_245,In_864,In_132);
nor U246 (N_246,In_1978,In_667);
and U247 (N_247,In_1675,In_1790);
and U248 (N_248,In_475,In_826);
or U249 (N_249,In_1661,In_1870);
xnor U250 (N_250,N_92,In_1123);
xor U251 (N_251,In_631,In_682);
nand U252 (N_252,In_91,In_867);
or U253 (N_253,In_539,In_1589);
and U254 (N_254,In_1178,In_1423);
nor U255 (N_255,In_1939,In_1751);
xor U256 (N_256,In_39,In_875);
xor U257 (N_257,In_673,In_568);
or U258 (N_258,In_357,In_1258);
and U259 (N_259,In_303,In_798);
nand U260 (N_260,In_57,In_1200);
nand U261 (N_261,In_1509,In_1685);
or U262 (N_262,In_809,In_1928);
nor U263 (N_263,N_173,In_1184);
xnor U264 (N_264,In_1793,N_158);
or U265 (N_265,In_807,In_449);
or U266 (N_266,In_1194,In_948);
nor U267 (N_267,In_1410,In_1906);
or U268 (N_268,In_871,In_1453);
or U269 (N_269,In_1655,In_842);
and U270 (N_270,In_385,N_231);
nand U271 (N_271,In_1924,In_103);
nand U272 (N_272,In_784,In_748);
nand U273 (N_273,In_971,In_1141);
nor U274 (N_274,In_353,In_1721);
xor U275 (N_275,N_76,N_90);
xor U276 (N_276,In_302,In_947);
nor U277 (N_277,In_1219,In_609);
nor U278 (N_278,N_2,In_1499);
and U279 (N_279,In_1134,In_1011);
nand U280 (N_280,In_264,In_812);
and U281 (N_281,In_1652,In_1162);
and U282 (N_282,In_1887,In_764);
or U283 (N_283,In_520,In_1578);
or U284 (N_284,In_1749,In_464);
or U285 (N_285,N_219,In_969);
nor U286 (N_286,In_1882,In_531);
or U287 (N_287,In_1631,In_1645);
nand U288 (N_288,In_234,In_1824);
xor U289 (N_289,In_762,In_1676);
xor U290 (N_290,In_1826,In_100);
and U291 (N_291,In_1487,N_225);
nor U292 (N_292,N_236,N_131);
nor U293 (N_293,In_839,In_1695);
nor U294 (N_294,In_924,In_1672);
and U295 (N_295,In_709,In_1404);
or U296 (N_296,In_835,In_532);
xnor U297 (N_297,In_1533,In_1394);
xnor U298 (N_298,In_734,In_1780);
nand U299 (N_299,In_1329,N_179);
nor U300 (N_300,In_142,In_1369);
and U301 (N_301,In_747,In_110);
nand U302 (N_302,In_1844,In_1981);
xor U303 (N_303,In_1073,In_577);
nand U304 (N_304,N_1,N_112);
nand U305 (N_305,In_1440,N_169);
and U306 (N_306,In_731,In_477);
or U307 (N_307,In_446,In_55);
xnor U308 (N_308,In_1901,In_977);
nand U309 (N_309,In_1055,In_1697);
nor U310 (N_310,In_195,In_398);
or U311 (N_311,In_1712,In_1409);
and U312 (N_312,In_1973,N_238);
nor U313 (N_313,In_1361,In_38);
xnor U314 (N_314,In_782,In_697);
xor U315 (N_315,In_1861,N_84);
and U316 (N_316,N_220,In_1168);
or U317 (N_317,In_233,In_604);
or U318 (N_318,In_44,In_1210);
nor U319 (N_319,In_470,N_130);
nand U320 (N_320,In_1193,In_730);
or U321 (N_321,N_23,In_930);
nor U322 (N_322,In_1602,In_244);
or U323 (N_323,In_1551,In_1761);
nor U324 (N_324,In_1021,In_771);
xnor U325 (N_325,N_99,In_1180);
and U326 (N_326,In_849,N_229);
and U327 (N_327,In_180,In_1765);
nand U328 (N_328,In_1437,In_1682);
or U329 (N_329,In_1831,In_1131);
nor U330 (N_330,In_256,In_601);
or U331 (N_331,In_12,In_1834);
xnor U332 (N_332,In_140,In_1036);
nor U333 (N_333,In_1743,In_1985);
or U334 (N_334,N_239,In_1975);
nand U335 (N_335,In_1933,In_1164);
nor U336 (N_336,In_1653,In_1054);
nand U337 (N_337,N_30,In_1615);
or U338 (N_338,N_249,In_1773);
nor U339 (N_339,In_156,In_1785);
or U340 (N_340,In_790,In_396);
and U341 (N_341,In_863,In_687);
xor U342 (N_342,In_7,In_121);
or U343 (N_343,In_1764,In_348);
nand U344 (N_344,In_3,In_489);
nor U345 (N_345,In_510,N_136);
or U346 (N_346,In_859,In_404);
nor U347 (N_347,In_970,In_381);
nor U348 (N_348,In_1348,In_1373);
or U349 (N_349,N_212,In_1351);
nand U350 (N_350,In_419,In_612);
or U351 (N_351,In_484,In_850);
nand U352 (N_352,In_1170,N_175);
xnor U353 (N_353,In_98,In_79);
nand U354 (N_354,In_228,In_759);
xnor U355 (N_355,In_767,In_1042);
or U356 (N_356,In_276,In_1420);
nand U357 (N_357,In_325,In_1051);
and U358 (N_358,In_1574,In_40);
nor U359 (N_359,In_1065,In_1101);
or U360 (N_360,N_151,In_289);
and U361 (N_361,In_60,In_1691);
nand U362 (N_362,N_58,In_1171);
or U363 (N_363,N_188,In_554);
nor U364 (N_364,N_177,In_421);
or U365 (N_365,In_1154,In_27);
nand U366 (N_366,In_108,In_290);
xor U367 (N_367,N_150,In_1538);
nand U368 (N_368,In_974,In_1216);
xnor U369 (N_369,N_217,In_1175);
xnor U370 (N_370,In_1739,In_866);
xnor U371 (N_371,In_1949,In_268);
nor U372 (N_372,In_203,In_364);
xor U373 (N_373,In_1475,N_63);
nand U374 (N_374,In_1412,In_952);
nand U375 (N_375,In_781,N_104);
and U376 (N_376,In_90,In_354);
and U377 (N_377,In_1442,In_498);
or U378 (N_378,In_794,In_133);
or U379 (N_379,In_1998,In_1472);
nand U380 (N_380,N_83,In_1983);
nand U381 (N_381,In_130,In_1596);
nand U382 (N_382,In_1594,In_1585);
xnor U383 (N_383,In_375,In_171);
xnor U384 (N_384,In_148,N_46);
xor U385 (N_385,N_247,In_193);
nand U386 (N_386,In_1371,In_1157);
and U387 (N_387,N_126,In_1081);
nand U388 (N_388,In_327,In_1428);
nand U389 (N_389,In_1980,In_1634);
nor U390 (N_390,In_1411,N_156);
xnor U391 (N_391,In_1576,In_623);
and U392 (N_392,In_753,In_997);
and U393 (N_393,In_834,In_172);
or U394 (N_394,N_78,In_811);
nand U395 (N_395,N_24,In_1237);
or U396 (N_396,N_128,In_136);
nand U397 (N_397,N_116,N_121);
and U398 (N_398,In_1232,N_118);
and U399 (N_399,In_1618,In_649);
or U400 (N_400,In_1711,In_1260);
and U401 (N_401,In_1262,In_1984);
nor U402 (N_402,In_1601,In_1344);
xnor U403 (N_403,In_1235,In_1881);
xor U404 (N_404,In_333,N_95);
xor U405 (N_405,In_122,In_1243);
nor U406 (N_406,In_1522,In_882);
nor U407 (N_407,In_1326,In_321);
xnor U408 (N_408,In_51,N_108);
nor U409 (N_409,In_1337,In_1865);
nor U410 (N_410,In_1731,In_1241);
xor U411 (N_411,In_1710,In_1777);
and U412 (N_412,In_1253,In_745);
nand U413 (N_413,In_787,N_66);
nor U414 (N_414,N_43,In_1709);
nor U415 (N_415,In_902,In_891);
nor U416 (N_416,In_1136,In_655);
xnor U417 (N_417,In_561,In_591);
xor U418 (N_418,In_1660,In_1779);
xnor U419 (N_419,In_792,In_878);
or U420 (N_420,In_610,In_343);
nor U421 (N_421,N_68,In_315);
xor U422 (N_422,In_41,In_1391);
xor U423 (N_423,In_1017,In_1559);
nand U424 (N_424,In_246,N_240);
xnor U425 (N_425,In_48,In_277);
nor U426 (N_426,In_856,In_1494);
nand U427 (N_427,In_868,In_1555);
and U428 (N_428,In_1019,In_1708);
nor U429 (N_429,In_932,In_841);
nand U430 (N_430,In_1798,In_11);
or U431 (N_431,N_230,In_1953);
xnor U432 (N_432,In_529,In_1830);
nand U433 (N_433,In_1087,In_13);
and U434 (N_434,N_227,In_1044);
xor U435 (N_435,In_166,In_1722);
nand U436 (N_436,In_188,In_736);
nand U437 (N_437,In_931,In_525);
or U438 (N_438,In_187,In_877);
and U439 (N_439,In_1629,In_617);
or U440 (N_440,In_1484,In_291);
nand U441 (N_441,In_69,In_1914);
nor U442 (N_442,In_1252,In_71);
and U443 (N_443,In_407,In_1945);
or U444 (N_444,In_349,In_162);
nor U445 (N_445,In_1841,In_1762);
nand U446 (N_446,In_1583,In_1006);
nand U447 (N_447,N_216,In_1822);
nor U448 (N_448,In_823,In_1085);
and U449 (N_449,In_393,In_1846);
and U450 (N_450,In_1504,In_1795);
and U451 (N_451,N_117,In_1197);
nor U452 (N_452,In_1360,In_1562);
and U453 (N_453,N_10,In_285);
nand U454 (N_454,In_587,In_752);
and U455 (N_455,N_67,In_1872);
or U456 (N_456,In_558,In_503);
nor U457 (N_457,In_1429,In_1567);
nand U458 (N_458,In_1818,In_1755);
nor U459 (N_459,In_1769,In_1890);
or U460 (N_460,In_420,In_982);
nor U461 (N_461,In_1209,In_307);
nand U462 (N_462,In_1255,N_138);
or U463 (N_463,In_350,In_1186);
xor U464 (N_464,N_146,N_75);
and U465 (N_465,In_985,In_83);
nor U466 (N_466,In_1187,In_1220);
nor U467 (N_467,In_1700,In_1315);
and U468 (N_468,N_49,In_1837);
or U469 (N_469,In_1930,In_1427);
and U470 (N_470,In_797,In_1814);
or U471 (N_471,In_1657,In_485);
and U472 (N_472,In_1462,In_1565);
xnor U473 (N_473,In_356,In_1936);
or U474 (N_474,In_1986,In_817);
and U475 (N_475,In_1038,In_880);
or U476 (N_476,In_1862,N_39);
nor U477 (N_477,In_1355,In_1570);
nand U478 (N_478,In_1488,In_1633);
xor U479 (N_479,In_873,In_1345);
nand U480 (N_480,In_218,In_1212);
or U481 (N_481,In_429,In_1359);
nor U482 (N_482,In_451,In_270);
nand U483 (N_483,In_961,In_917);
xor U484 (N_484,In_1995,In_88);
nor U485 (N_485,N_207,In_1833);
xnor U486 (N_486,In_1934,In_772);
nand U487 (N_487,In_123,In_1483);
and U488 (N_488,In_1376,N_139);
nor U489 (N_489,In_1877,N_40);
and U490 (N_490,In_1246,In_1925);
or U491 (N_491,In_1964,N_52);
nand U492 (N_492,In_1853,In_1630);
xnor U493 (N_493,In_1037,In_872);
nor U494 (N_494,In_77,In_102);
xor U495 (N_495,In_1622,In_1069);
and U496 (N_496,In_1155,In_1480);
and U497 (N_497,In_1142,In_336);
or U498 (N_498,In_1072,In_1163);
or U499 (N_499,In_220,In_1549);
or U500 (N_500,In_326,N_193);
and U501 (N_501,In_606,In_1481);
or U502 (N_502,In_833,In_1595);
nand U503 (N_503,In_1290,In_544);
nand U504 (N_504,In_61,N_241);
nor U505 (N_505,In_192,In_723);
and U506 (N_506,In_1667,N_142);
or U507 (N_507,In_1597,In_8);
or U508 (N_508,In_716,In_1264);
nand U509 (N_509,In_911,N_431);
nor U510 (N_510,In_1372,N_383);
nand U511 (N_511,N_18,In_1531);
nand U512 (N_512,In_936,In_207);
xnor U513 (N_513,In_109,In_1398);
or U514 (N_514,In_1801,In_824);
xnor U515 (N_515,N_465,In_1205);
nand U516 (N_516,N_201,In_905);
xnor U517 (N_517,In_185,In_235);
nor U518 (N_518,N_346,In_1283);
and U519 (N_519,In_1127,In_1356);
nor U520 (N_520,N_362,N_246);
or U521 (N_521,In_1118,In_1314);
nor U522 (N_522,In_1553,In_80);
nand U523 (N_523,In_161,In_25);
nand U524 (N_524,N_423,N_145);
xnor U525 (N_525,In_1024,N_427);
xor U526 (N_526,In_1508,In_1413);
nand U527 (N_527,In_1271,In_1408);
nor U528 (N_528,In_904,In_292);
or U529 (N_529,In_1148,In_1643);
xor U530 (N_530,In_1176,In_1800);
and U531 (N_531,N_245,In_1636);
or U532 (N_532,N_373,In_732);
nand U533 (N_533,In_1489,N_473);
nand U534 (N_534,In_1935,N_395);
xor U535 (N_535,N_244,In_31);
xor U536 (N_536,In_1628,In_1227);
or U537 (N_537,N_55,In_1374);
xnor U538 (N_538,In_908,In_1624);
nor U539 (N_539,In_1581,N_276);
nor U540 (N_540,In_30,In_1946);
xor U541 (N_541,In_462,In_1368);
nor U542 (N_542,N_407,N_182);
xor U543 (N_543,N_17,In_1305);
xor U544 (N_544,In_844,In_1294);
nand U545 (N_545,N_413,N_483);
and U546 (N_546,N_267,N_178);
nor U547 (N_547,In_56,In_689);
nand U548 (N_548,In_1010,In_65);
nand U549 (N_549,In_513,N_261);
and U550 (N_550,In_1736,In_150);
xor U551 (N_551,In_1419,In_141);
nand U552 (N_552,N_277,In_455);
nand U553 (N_553,In_676,In_695);
and U554 (N_554,In_1063,In_310);
xor U555 (N_555,In_1857,N_149);
and U556 (N_556,In_458,In_1421);
nand U557 (N_557,N_35,In_984);
nor U558 (N_558,N_496,In_196);
xor U559 (N_559,In_1381,In_308);
nand U560 (N_560,In_1514,In_496);
and U561 (N_561,In_502,N_88);
and U562 (N_562,N_318,N_489);
nor U563 (N_563,In_551,N_198);
nor U564 (N_564,N_471,In_1067);
nand U565 (N_565,In_1963,In_1606);
and U566 (N_566,In_778,In_1169);
or U567 (N_567,In_92,In_1571);
or U568 (N_568,In_214,N_255);
xor U569 (N_569,In_1213,N_401);
and U570 (N_570,In_1941,N_436);
nand U571 (N_571,In_106,In_990);
or U572 (N_572,In_783,N_301);
nand U573 (N_573,In_621,In_1803);
xor U574 (N_574,In_1250,In_648);
nand U575 (N_575,In_1738,In_32);
nand U576 (N_576,N_153,In_768);
or U577 (N_577,N_302,N_105);
xnor U578 (N_578,In_1816,In_26);
nand U579 (N_579,In_766,N_159);
nand U580 (N_580,In_1766,N_367);
nor U581 (N_581,In_250,In_1296);
nand U582 (N_582,In_1974,N_60);
and U583 (N_583,In_323,N_485);
nor U584 (N_584,In_366,In_433);
nor U585 (N_585,In_1560,In_1664);
and U586 (N_586,In_818,In_1119);
xor U587 (N_587,In_372,In_1809);
xnor U588 (N_588,In_770,In_232);
nor U589 (N_589,In_1892,N_414);
and U590 (N_590,N_36,In_913);
nand U591 (N_591,In_1729,In_1405);
and U592 (N_592,In_293,In_413);
and U593 (N_593,In_1544,In_934);
and U594 (N_594,In_206,In_440);
and U595 (N_595,In_746,In_463);
xnor U596 (N_596,N_248,N_332);
nand U597 (N_597,N_351,N_22);
xnor U598 (N_598,In_1718,In_1203);
xor U599 (N_599,In_1454,In_705);
and U600 (N_600,In_953,In_1958);
xor U601 (N_601,In_1366,N_80);
and U602 (N_602,In_28,N_298);
xnor U603 (N_603,In_1971,N_317);
or U604 (N_604,N_37,N_396);
xor U605 (N_605,In_1563,In_1111);
and U606 (N_606,N_163,In_1569);
and U607 (N_607,In_1357,In_1916);
nand U608 (N_608,In_1040,In_1808);
nor U609 (N_609,N_102,N_97);
xnor U610 (N_610,In_1086,N_228);
nor U611 (N_611,In_683,In_93);
nor U612 (N_612,N_450,In_313);
xnor U613 (N_613,In_202,In_626);
nor U614 (N_614,In_937,N_167);
xnor U615 (N_615,N_444,In_1879);
and U616 (N_616,In_679,In_1590);
nand U617 (N_617,In_1431,N_319);
or U618 (N_618,In_278,N_7);
nor U619 (N_619,N_443,In_774);
nand U620 (N_620,In_70,In_1579);
xnor U621 (N_621,In_620,In_1759);
xor U622 (N_622,In_1982,In_1768);
xnor U623 (N_623,In_382,In_935);
xnor U624 (N_624,In_1648,In_1448);
nor U625 (N_625,In_355,In_1720);
xnor U626 (N_626,In_1940,N_137);
nand U627 (N_627,In_788,In_1287);
xnor U628 (N_628,N_333,In_1847);
or U629 (N_629,In_1068,In_1389);
nand U630 (N_630,In_197,In_578);
and U631 (N_631,In_521,In_312);
nor U632 (N_632,In_1523,N_113);
nor U633 (N_633,In_796,N_34);
nor U634 (N_634,In_1864,In_1144);
xnor U635 (N_635,In_1658,In_1046);
nand U636 (N_636,N_202,In_453);
and U637 (N_637,In_596,N_428);
nand U638 (N_638,In_749,In_597);
xnor U639 (N_639,N_71,In_1107);
and U640 (N_640,N_425,In_1198);
and U641 (N_641,In_714,In_1744);
and U642 (N_642,N_381,In_1776);
nand U643 (N_643,In_567,In_0);
and U644 (N_644,N_252,In_452);
nor U645 (N_645,In_1379,In_105);
nand U646 (N_646,In_1238,In_988);
nor U647 (N_647,In_225,In_1435);
or U648 (N_648,In_901,N_256);
and U649 (N_649,N_307,In_600);
xnor U650 (N_650,In_1703,N_366);
and U651 (N_651,In_1730,In_550);
xor U652 (N_652,In_981,N_268);
and U653 (N_653,In_319,In_1919);
xnor U654 (N_654,N_143,N_161);
nor U655 (N_655,N_61,In_1740);
nand U656 (N_656,In_450,In_1143);
nand U657 (N_657,In_1390,In_757);
and U658 (N_658,In_1536,In_967);
nand U659 (N_659,In_1540,In_457);
xor U660 (N_660,N_440,In_1091);
nor U661 (N_661,In_1274,In_836);
xor U662 (N_662,In_1077,In_482);
nand U663 (N_663,N_115,In_1741);
nor U664 (N_664,N_269,In_182);
xor U665 (N_665,N_462,In_1070);
or U666 (N_666,In_21,N_274);
nand U667 (N_667,In_1280,In_447);
nand U668 (N_668,N_38,N_481);
and U669 (N_669,In_658,N_472);
nand U670 (N_670,In_1609,In_179);
nand U671 (N_671,In_459,In_1852);
and U672 (N_672,N_103,In_176);
xor U673 (N_673,N_144,In_1350);
xnor U674 (N_674,In_68,In_832);
and U675 (N_675,In_1202,In_1032);
xor U676 (N_676,In_435,In_825);
or U677 (N_677,In_1380,In_1723);
xor U678 (N_678,In_1909,In_1927);
nor U679 (N_679,In_1550,N_59);
or U680 (N_680,N_345,In_247);
and U681 (N_681,In_1449,N_387);
nor U682 (N_682,In_853,In_1693);
nor U683 (N_683,In_1199,In_1417);
or U684 (N_684,N_323,In_201);
nor U685 (N_685,In_1150,In_838);
xor U686 (N_686,In_1401,In_1015);
or U687 (N_687,N_226,N_403);
nor U688 (N_688,In_431,In_1817);
nand U689 (N_689,N_123,In_1320);
or U690 (N_690,In_1269,In_995);
nand U691 (N_691,In_1932,In_744);
xnor U692 (N_692,In_943,In_505);
or U693 (N_693,In_1948,In_1895);
nand U694 (N_694,In_259,In_848);
and U695 (N_695,In_124,In_662);
nand U696 (N_696,N_495,N_299);
and U697 (N_697,N_251,In_263);
or U698 (N_698,N_275,In_85);
xor U699 (N_699,In_1878,In_702);
nor U700 (N_700,In_1529,In_467);
or U701 (N_701,N_295,N_215);
xor U702 (N_702,In_1856,In_1116);
nand U703 (N_703,N_487,In_575);
xnor U704 (N_704,In_1097,In_497);
nor U705 (N_705,In_211,N_0);
xnor U706 (N_706,In_1545,N_498);
and U707 (N_707,In_1907,In_992);
nand U708 (N_708,In_742,In_1353);
xor U709 (N_709,In_468,In_1115);
nor U710 (N_710,N_265,N_221);
nand U711 (N_711,In_1336,In_1406);
nor U712 (N_712,N_402,N_451);
xnor U713 (N_713,In_1725,In_240);
nor U714 (N_714,In_1666,In_318);
and U715 (N_715,In_1463,In_474);
or U716 (N_716,In_87,N_466);
or U717 (N_717,N_296,In_309);
xnor U718 (N_718,In_1465,N_203);
and U719 (N_719,N_223,In_666);
nand U720 (N_720,In_553,In_1735);
or U721 (N_721,In_720,In_769);
or U722 (N_722,In_1496,In_1728);
xor U723 (N_723,In_1242,In_1929);
and U724 (N_724,In_1908,N_433);
xor U725 (N_725,In_1217,In_417);
and U726 (N_726,In_1505,In_227);
or U727 (N_727,In_1811,N_57);
nor U728 (N_728,In_829,In_1827);
nor U729 (N_729,N_214,N_87);
or U730 (N_730,In_678,In_1224);
or U731 (N_731,In_1060,In_1627);
nor U732 (N_732,In_63,N_426);
or U733 (N_733,N_349,N_488);
xnor U734 (N_734,In_1577,N_494);
xnor U735 (N_735,In_966,In_184);
xnor U736 (N_736,In_338,In_1724);
or U737 (N_737,In_369,In_1395);
nand U738 (N_738,N_288,In_507);
and U739 (N_739,In_651,N_461);
nor U740 (N_740,In_78,N_180);
nor U741 (N_741,N_310,N_455);
nand U742 (N_742,N_257,N_8);
nand U743 (N_743,In_76,In_1233);
nand U744 (N_744,In_780,In_881);
and U745 (N_745,In_1303,In_1637);
nand U746 (N_746,In_1874,In_1649);
or U747 (N_747,In_1954,In_933);
or U748 (N_748,In_151,In_170);
xor U749 (N_749,N_280,In_1020);
nand U750 (N_750,In_1897,In_99);
and U751 (N_751,In_585,N_120);
nand U752 (N_752,In_1486,In_906);
or U753 (N_753,N_541,N_19);
nand U754 (N_754,N_185,N_691);
xor U755 (N_755,In_306,In_1443);
nor U756 (N_756,In_1910,N_710);
nor U757 (N_757,In_73,In_1165);
and U758 (N_758,N_48,N_463);
or U759 (N_759,N_421,In_921);
nand U760 (N_760,N_673,In_1000);
and U761 (N_761,In_1393,In_1763);
nor U762 (N_762,In_950,In_691);
nor U763 (N_763,N_478,In_1704);
nor U764 (N_764,N_576,In_1352);
nand U765 (N_765,N_460,In_267);
xor U766 (N_766,In_304,N_243);
or U767 (N_767,In_64,In_861);
nand U768 (N_768,In_665,In_1084);
xnor U769 (N_769,In_287,In_706);
nor U770 (N_770,In_1626,In_1737);
or U771 (N_771,In_900,In_1122);
and U772 (N_772,In_1698,In_371);
nor U773 (N_773,N_132,In_1742);
or U774 (N_774,N_446,N_692);
and U775 (N_775,In_1614,In_1311);
xor U776 (N_776,N_622,N_166);
or U777 (N_777,N_232,N_570);
nand U778 (N_778,In_729,In_1458);
and U779 (N_779,N_721,N_676);
and U780 (N_780,N_467,N_618);
xor U781 (N_781,N_631,In_1920);
and U782 (N_782,N_386,In_751);
nand U783 (N_783,N_565,In_1898);
and U784 (N_784,In_1304,N_533);
nand U785 (N_785,In_1322,In_619);
and U786 (N_786,N_689,N_361);
nand U787 (N_787,N_655,N_680);
xnor U788 (N_788,N_342,In_1439);
nand U789 (N_789,In_145,N_675);
or U790 (N_790,In_1362,In_1778);
nor U791 (N_791,N_665,In_495);
xnor U792 (N_792,N_633,In_1273);
nand U793 (N_793,In_1191,N_662);
nand U794 (N_794,In_1851,In_1328);
or U795 (N_795,N_98,In_994);
nor U796 (N_796,N_100,N_632);
nor U797 (N_797,N_140,In_1158);
nor U798 (N_798,N_343,N_572);
nor U799 (N_799,In_388,In_1312);
nand U800 (N_800,In_555,In_1396);
xor U801 (N_801,N_643,In_684);
nand U802 (N_802,In_274,In_692);
nand U803 (N_803,In_516,In_380);
and U804 (N_804,In_384,In_1335);
nand U805 (N_805,In_115,N_612);
or U806 (N_806,N_677,N_331);
xnor U807 (N_807,N_597,N_94);
and U808 (N_808,In_605,In_592);
or U809 (N_809,In_1656,In_1893);
xnor U810 (N_810,In_1045,In_960);
and U811 (N_811,N_107,In_183);
nor U812 (N_812,N_152,In_1593);
nand U813 (N_813,In_847,N_282);
xnor U814 (N_814,N_611,In_1346);
xnor U815 (N_815,N_171,N_50);
nor U816 (N_816,In_941,In_837);
xnor U817 (N_817,In_1680,In_795);
xor U818 (N_818,N_649,In_36);
or U819 (N_819,In_1297,In_400);
or U820 (N_820,N_365,In_528);
nand U821 (N_821,N_51,N_419);
xnor U822 (N_822,In_741,N_567);
or U823 (N_823,In_126,N_638);
nand U824 (N_824,In_143,N_441);
nand U825 (N_825,N_81,N_263);
and U826 (N_826,In_1156,In_1298);
xor U827 (N_827,In_111,In_724);
nor U828 (N_828,In_560,N_626);
and U829 (N_829,In_712,In_1923);
xnor U830 (N_830,In_1659,In_718);
nand U831 (N_831,In_1668,N_16);
and U832 (N_832,N_89,In_657);
or U833 (N_833,N_605,N_25);
nand U834 (N_834,In_460,N_45);
and U835 (N_835,N_549,In_149);
and U836 (N_836,In_1650,In_584);
and U837 (N_837,In_208,N_147);
nor U838 (N_838,N_399,In_660);
nor U839 (N_839,In_1342,N_727);
xnor U840 (N_840,N_506,N_189);
or U841 (N_841,In_1770,In_998);
xnor U842 (N_842,In_1239,In_1418);
nand U843 (N_843,N_368,In_1470);
and U844 (N_844,N_187,N_685);
or U845 (N_845,N_540,In_476);
and U846 (N_846,N_196,In_1485);
and U847 (N_847,N_300,N_716);
xnor U848 (N_848,In_1049,In_1450);
or U849 (N_849,In_411,In_299);
nand U850 (N_850,N_378,N_438);
xnor U851 (N_851,In_643,In_1254);
or U852 (N_852,In_955,N_474);
or U853 (N_853,In_556,N_279);
and U854 (N_854,In_1378,N_543);
and U855 (N_855,N_573,In_1226);
xor U856 (N_856,In_1433,In_344);
nor U857 (N_857,In_703,In_1195);
nor U858 (N_858,In_573,In_1285);
and U859 (N_859,In_479,In_283);
xnor U860 (N_860,In_390,N_579);
or U861 (N_861,In_1510,In_1972);
xnor U862 (N_862,In_581,N_729);
or U863 (N_863,In_801,In_1988);
xor U864 (N_864,N_29,In_637);
or U865 (N_865,In_993,In_680);
or U866 (N_866,In_134,N_254);
nand U867 (N_867,N_602,N_449);
nor U868 (N_868,N_294,In_1547);
xnor U869 (N_869,N_379,N_133);
and U870 (N_870,N_273,In_740);
xor U871 (N_871,In_1511,N_635);
nand U872 (N_872,N_434,N_539);
xnor U873 (N_873,In_45,N_96);
nor U874 (N_874,N_520,In_383);
or U875 (N_875,In_557,In_923);
and U876 (N_876,N_656,N_728);
and U877 (N_877,N_730,In_607);
xnor U878 (N_878,In_1121,N_595);
and U879 (N_879,N_311,In_564);
and U880 (N_880,N_686,In_1554);
nor U881 (N_881,In_519,In_221);
nor U882 (N_882,N_258,In_480);
nand U883 (N_883,In_1172,N_424);
nor U884 (N_884,In_164,In_677);
or U885 (N_885,In_1588,In_1681);
nor U886 (N_886,N_259,In_226);
xor U887 (N_887,N_157,In_1886);
xnor U888 (N_888,In_434,In_1147);
and U889 (N_889,In_1792,In_1292);
nor U890 (N_890,N_518,In_1130);
xnor U891 (N_891,N_523,In_704);
or U892 (N_892,In_1114,N_697);
nand U893 (N_893,In_754,N_555);
nor U894 (N_894,In_530,N_500);
nand U895 (N_895,N_648,N_736);
nor U896 (N_896,N_437,N_501);
and U897 (N_897,N_375,In_1638);
and U898 (N_898,In_1813,In_1281);
xnor U899 (N_899,In_652,In_725);
and U900 (N_900,N_553,N_719);
and U901 (N_901,N_464,In_29);
nor U902 (N_902,N_698,N_693);
xnor U903 (N_903,In_628,In_883);
xnor U904 (N_904,In_1584,In_1905);
and U905 (N_905,N_505,In_1561);
and U906 (N_906,N_4,N_213);
nor U907 (N_907,N_370,In_104);
nand U908 (N_908,In_439,N_199);
nand U909 (N_909,In_1753,In_1050);
or U910 (N_910,In_1635,N_604);
nor U911 (N_911,In_845,N_512);
nor U912 (N_912,In_224,N_400);
xor U913 (N_913,In_1821,In_1996);
nand U914 (N_914,In_1075,N_234);
xor U915 (N_915,In_1009,In_1278);
xor U916 (N_916,N_344,N_508);
nor U917 (N_917,N_575,In_461);
nand U918 (N_918,N_645,N_526);
or U919 (N_919,N_706,N_694);
xor U920 (N_920,In_5,In_345);
or U921 (N_921,In_865,In_86);
or U922 (N_922,N_493,N_591);
nand U923 (N_923,In_362,N_314);
and U924 (N_924,In_1340,N_9);
or U925 (N_925,N_290,N_468);
or U926 (N_926,In_537,In_1110);
and U927 (N_927,In_1573,N_313);
xor U928 (N_928,In_107,In_1057);
or U929 (N_929,In_599,In_625);
nand U930 (N_930,N_713,In_1240);
nor U931 (N_931,N_625,N_408);
xor U932 (N_932,In_89,In_1464);
or U933 (N_933,N_718,In_443);
xor U934 (N_934,In_1621,In_779);
nor U935 (N_935,In_1083,N_636);
nor U936 (N_936,N_409,N_209);
nor U937 (N_937,In_820,In_137);
or U938 (N_938,N_134,In_893);
xnor U939 (N_939,N_456,N_210);
and U940 (N_940,N_590,N_669);
nand U941 (N_941,N_748,N_27);
xnor U942 (N_942,N_13,N_497);
and U943 (N_943,In_174,In_238);
or U944 (N_944,N_197,N_101);
or U945 (N_945,N_235,In_1900);
and U946 (N_946,In_360,N_388);
or U947 (N_947,In_563,In_945);
and U948 (N_948,In_1471,In_1367);
nor U949 (N_949,N_724,N_566);
nor U950 (N_950,In_1866,N_47);
or U951 (N_951,In_1259,In_918);
nand U952 (N_952,In_282,N_714);
nand U953 (N_953,In_1221,N_341);
and U954 (N_954,N_272,N_554);
and U955 (N_955,In_153,In_1064);
or U956 (N_956,N_587,In_1688);
and U957 (N_957,N_416,In_198);
nand U958 (N_958,In_611,N_172);
nand U959 (N_959,N_568,N_162);
xor U960 (N_960,In_1327,In_540);
xnor U961 (N_961,In_670,N_363);
nor U962 (N_962,In_1548,N_679);
xor U963 (N_963,In_663,In_669);
nand U964 (N_964,In_1153,In_919);
xor U965 (N_965,In_1502,N_492);
nand U966 (N_966,In_1479,N_322);
nand U967 (N_967,N_699,N_297);
nor U968 (N_968,N_544,N_336);
xnor U969 (N_969,N_482,N_746);
and U970 (N_970,In_972,In_535);
nand U971 (N_971,N_668,In_1873);
xor U972 (N_972,In_1692,In_1674);
nor U973 (N_973,In_1185,N_82);
nor U974 (N_974,N_316,N_194);
or U975 (N_975,N_260,N_703);
and U976 (N_976,In_1918,N_641);
nand U977 (N_977,N_513,In_1670);
and U978 (N_978,N_684,N_391);
and U979 (N_979,N_560,In_1714);
or U980 (N_980,In_571,N_382);
or U981 (N_981,In_1103,N_320);
nor U982 (N_982,In_1772,In_1247);
xnor U983 (N_983,N_722,N_535);
xnor U984 (N_984,N_119,In_739);
or U985 (N_985,In_1206,N_470);
nand U986 (N_986,In_415,In_959);
nor U987 (N_987,In_1891,In_1663);
nor U988 (N_988,N_530,N_702);
nand U989 (N_989,N_479,In_1415);
or U990 (N_990,In_414,In_423);
xor U991 (N_991,In_62,In_1074);
xor U992 (N_992,In_1295,N_737);
or U993 (N_993,N_583,N_733);
or U994 (N_994,In_84,In_743);
and U995 (N_995,N_135,In_237);
nor U996 (N_996,N_262,In_1791);
or U997 (N_997,In_574,N_54);
nand U998 (N_998,N_525,In_342);
or U999 (N_999,In_1524,N_192);
nand U1000 (N_1000,N_868,In_295);
or U1001 (N_1001,In_760,In_1782);
or U1002 (N_1002,N_867,N_56);
nor U1003 (N_1003,N_854,N_805);
and U1004 (N_1004,N_91,In_822);
xor U1005 (N_1005,In_1177,In_831);
and U1006 (N_1006,In_1330,N_977);
or U1007 (N_1007,In_1318,N_974);
and U1008 (N_1008,N_581,N_892);
nand U1009 (N_1009,In_589,In_1557);
and U1010 (N_1010,In_1388,In_1476);
and U1011 (N_1011,In_1654,N_26);
xor U1012 (N_1012,N_965,N_890);
or U1013 (N_1013,N_981,In_733);
nand U1014 (N_1014,N_211,In_821);
xnor U1015 (N_1015,In_1829,N_561);
nor U1016 (N_1016,In_1266,In_1781);
or U1017 (N_1017,N_983,N_393);
nor U1018 (N_1018,N_771,N_762);
xnor U1019 (N_1019,N_206,In_944);
nor U1020 (N_1020,In_1078,N_784);
and U1021 (N_1021,N_780,N_847);
nor U1022 (N_1022,In_405,In_1587);
xnor U1023 (N_1023,In_857,In_1787);
and U1024 (N_1024,In_1997,N_767);
nand U1025 (N_1025,In_1286,N_624);
nand U1026 (N_1026,N_174,N_283);
nand U1027 (N_1027,N_350,In_738);
and U1028 (N_1028,In_973,In_1313);
and U1029 (N_1029,N_903,N_871);
or U1030 (N_1030,N_12,In_216);
nor U1031 (N_1031,N_747,N_608);
xor U1032 (N_1032,N_667,N_990);
or U1033 (N_1033,In_1079,In_765);
nand U1034 (N_1034,N_340,N_825);
nand U1035 (N_1035,In_940,N_411);
nor U1036 (N_1036,N_930,N_709);
or U1037 (N_1037,N_164,In_1052);
xor U1038 (N_1038,In_672,N_933);
xnor U1039 (N_1039,In_1884,In_1705);
or U1040 (N_1040,N_637,N_963);
or U1041 (N_1041,In_1288,In_659);
nor U1042 (N_1042,In_688,In_1836);
xor U1043 (N_1043,In_1516,N_330);
and U1044 (N_1044,N_835,In_843);
and U1045 (N_1045,N_129,N_740);
and U1046 (N_1046,In_675,In_522);
or U1047 (N_1047,N_938,In_127);
nor U1048 (N_1048,N_502,N_601);
nor U1049 (N_1049,In_1004,In_139);
nor U1050 (N_1050,N_532,In_1218);
or U1051 (N_1051,In_212,N_690);
and U1052 (N_1052,N_958,In_1196);
and U1053 (N_1053,In_248,N_289);
and U1054 (N_1054,In_1190,In_707);
and U1055 (N_1055,In_1207,N_148);
and U1056 (N_1056,N_964,In_129);
and U1057 (N_1057,N_758,N_757);
xor U1058 (N_1058,N_731,N_86);
nand U1059 (N_1059,N_359,In_469);
xor U1060 (N_1060,N_281,N_584);
nor U1061 (N_1061,N_997,In_1002);
nor U1062 (N_1062,N_682,N_838);
or U1063 (N_1063,N_810,N_355);
nand U1064 (N_1064,In_1632,N_883);
nand U1065 (N_1065,In_424,In_454);
xor U1066 (N_1066,N_768,In_1211);
nand U1067 (N_1067,N_430,N_752);
and U1068 (N_1068,In_1152,N_577);
or U1069 (N_1069,N_21,In_409);
or U1070 (N_1070,N_646,In_401);
xor U1071 (N_1071,In_163,In_1859);
and U1072 (N_1072,In_690,N_992);
nor U1073 (N_1073,N_183,In_1167);
or U1074 (N_1074,In_1460,N_936);
and U1075 (N_1075,In_335,N_909);
or U1076 (N_1076,In_251,In_320);
xnor U1077 (N_1077,N_947,In_899);
xnor U1078 (N_1078,In_1093,In_243);
nand U1079 (N_1079,In_639,In_1617);
xor U1080 (N_1080,In_1599,N_551);
and U1081 (N_1081,N_695,N_987);
or U1082 (N_1082,In_422,N_808);
nand U1083 (N_1083,In_929,In_316);
and U1084 (N_1084,In_1257,N_873);
or U1085 (N_1085,N_809,N_264);
or U1086 (N_1086,In_632,N_406);
xor U1087 (N_1087,In_962,N_807);
xnor U1088 (N_1088,In_229,N_790);
or U1089 (N_1089,N_205,N_910);
nor U1090 (N_1090,In_647,In_874);
or U1091 (N_1091,In_957,N_452);
nand U1092 (N_1092,In_1543,In_523);
nor U1093 (N_1093,N_594,N_851);
xor U1094 (N_1094,In_427,In_1307);
xnor U1095 (N_1095,N_907,N_900);
xor U1096 (N_1096,N_415,N_315);
or U1097 (N_1097,N_486,N_242);
or U1098 (N_1098,N_723,In_67);
or U1099 (N_1099,N_534,N_208);
nor U1100 (N_1100,In_1012,In_273);
or U1101 (N_1101,In_1812,N_122);
nand U1102 (N_1102,N_3,In_1726);
xnor U1103 (N_1103,N_377,N_522);
and U1104 (N_1104,In_1403,In_280);
or U1105 (N_1105,N_916,N_204);
or U1106 (N_1106,N_453,N_364);
and U1107 (N_1107,N_352,N_726);
or U1108 (N_1108,In_1048,In_1041);
or U1109 (N_1109,N_176,In_177);
and U1110 (N_1110,In_1678,N_574);
nor U1111 (N_1111,In_1802,In_1734);
nor U1112 (N_1112,In_1610,N_537);
xnor U1113 (N_1113,In_1088,N_324);
or U1114 (N_1114,In_1492,In_642);
nand U1115 (N_1115,N_995,In_1512);
nand U1116 (N_1116,In_34,In_266);
xor U1117 (N_1117,N_681,N_634);
and U1118 (N_1118,N_811,N_291);
nor U1119 (N_1119,In_215,N_940);
and U1120 (N_1120,In_279,In_942);
xnor U1121 (N_1121,N_754,N_966);
and U1122 (N_1122,In_147,In_1332);
nand U1123 (N_1123,N_617,N_293);
xor U1124 (N_1124,N_770,N_376);
nand U1125 (N_1125,In_1446,N_795);
and U1126 (N_1126,N_32,N_720);
and U1127 (N_1127,N_503,In_508);
nand U1128 (N_1128,N_374,N_329);
nand U1129 (N_1129,In_870,N_812);
xor U1130 (N_1130,In_131,In_445);
or U1131 (N_1131,N_418,N_893);
or U1132 (N_1132,N_884,In_546);
nor U1133 (N_1133,In_1883,N_968);
nor U1134 (N_1134,In_1756,N_813);
xnor U1135 (N_1135,N_270,In_700);
nand U1136 (N_1136,In_538,In_1306);
nor U1137 (N_1137,In_1025,N_42);
nand U1138 (N_1138,N_967,In_255);
nor U1139 (N_1139,In_1159,In_1270);
and U1140 (N_1140,In_1215,In_1098);
nand U1141 (N_1141,N_125,In_876);
nand U1142 (N_1142,N_619,N_979);
nor U1143 (N_1143,In_219,N_949);
nor U1144 (N_1144,N_861,In_1279);
nand U1145 (N_1145,In_595,In_1310);
nand U1146 (N_1146,N_872,N_609);
nand U1147 (N_1147,N_562,In_297);
nand U1148 (N_1148,N_774,In_42);
nor U1149 (N_1149,N_755,N_943);
nand U1150 (N_1150,In_634,N_945);
or U1151 (N_1151,N_993,N_787);
or U1152 (N_1152,In_1534,N_712);
and U1153 (N_1153,N_93,In_1402);
and U1154 (N_1154,N_127,N_889);
nor U1155 (N_1155,N_863,N_715);
and U1156 (N_1156,In_1400,N_546);
or U1157 (N_1157,N_666,In_840);
or U1158 (N_1158,N_287,In_152);
nor U1159 (N_1159,N_877,In_239);
nor U1160 (N_1160,N_988,In_1234);
xnor U1161 (N_1161,In_490,N_823);
and U1162 (N_1162,N_671,In_1687);
nor U1163 (N_1163,In_975,N_321);
xor U1164 (N_1164,In_1018,N_705);
nand U1165 (N_1165,In_178,In_1528);
and U1166 (N_1166,N_725,N_696);
nand U1167 (N_1167,In_586,N_586);
or U1168 (N_1168,In_284,N_917);
or U1169 (N_1169,N_732,N_849);
nor U1170 (N_1170,In_912,N_800);
nand U1171 (N_1171,N_28,N_886);
nand U1172 (N_1172,N_874,In_1869);
and U1173 (N_1173,N_547,N_31);
and U1174 (N_1174,N_678,N_880);
nand U1175 (N_1175,N_337,In_1592);
nand U1176 (N_1176,In_1113,In_1507);
nor U1177 (N_1177,In_487,N_422);
and U1178 (N_1178,N_960,In_938);
or U1179 (N_1179,In_101,N_976);
nor U1180 (N_1180,N_653,N_490);
or U1181 (N_1181,N_394,In_1694);
or U1182 (N_1182,In_1519,N_802);
nor U1183 (N_1183,N_542,N_844);
xor U1184 (N_1184,N_840,N_360);
xnor U1185 (N_1185,In_1467,N_410);
or U1186 (N_1186,N_898,In_756);
and U1187 (N_1187,In_418,In_656);
or U1188 (N_1188,In_1642,In_721);
or U1189 (N_1189,In_650,In_1966);
xnor U1190 (N_1190,N_948,N_339);
and U1191 (N_1191,N_519,In_646);
or U1192 (N_1192,In_1515,N_571);
and U1193 (N_1193,In_361,In_1784);
nor U1194 (N_1194,N_233,N_582);
nor U1195 (N_1195,In_1179,N_895);
nor U1196 (N_1196,N_901,In_1375);
nor U1197 (N_1197,In_685,N_913);
nand U1198 (N_1198,N_841,N_155);
nor U1199 (N_1199,N_869,In_230);
and U1200 (N_1200,N_842,In_1845);
and U1201 (N_1201,N_989,N_833);
xnor U1202 (N_1202,N_457,In_814);
or U1203 (N_1203,In_1717,N_515);
nand U1204 (N_1204,N_110,N_596);
or U1205 (N_1205,N_801,N_420);
xor U1206 (N_1206,N_764,N_781);
nor U1207 (N_1207,In_1277,In_500);
and U1208 (N_1208,N_657,In_1302);
nor U1209 (N_1209,N_610,In_200);
and U1210 (N_1210,N_445,N_891);
xor U1211 (N_1211,N_704,N_334);
nand U1212 (N_1212,N_778,N_791);
and U1213 (N_1213,In_1244,N_588);
nand U1214 (N_1214,In_1183,In_242);
and U1215 (N_1215,N_510,In_1027);
nor U1216 (N_1216,N_935,N_607);
nor U1217 (N_1217,N_432,N_865);
xnor U1218 (N_1218,N_824,N_536);
and U1219 (N_1219,N_578,In_910);
and U1220 (N_1220,N_372,In_300);
xnor U1221 (N_1221,N_934,In_406);
nor U1222 (N_1222,N_937,In_399);
and U1223 (N_1223,In_493,N_701);
nor U1224 (N_1224,N_356,N_664);
and U1225 (N_1225,In_810,In_1989);
or U1226 (N_1226,N_688,In_1126);
nor U1227 (N_1227,In_1386,In_1620);
nor U1228 (N_1228,In_1299,N_660);
nand U1229 (N_1229,In_231,In_1535);
xor U1230 (N_1230,In_541,In_18);
xnor U1231 (N_1231,N_794,In_1289);
nor U1232 (N_1232,In_1607,In_14);
nor U1233 (N_1233,N_286,N_994);
nand U1234 (N_1234,In_194,N_308);
nand U1235 (N_1235,N_846,N_932);
or U1236 (N_1236,In_294,N_477);
or U1237 (N_1237,In_97,N_782);
xor U1238 (N_1238,N_569,In_1161);
nand U1239 (N_1239,In_358,In_613);
nor U1240 (N_1240,N_303,N_922);
xor U1241 (N_1241,N_832,N_798);
nor U1242 (N_1242,In_576,In_1245);
and U1243 (N_1243,In_726,In_58);
nor U1244 (N_1244,In_1977,N_603);
xor U1245 (N_1245,N_745,N_527);
and U1246 (N_1246,In_158,N_925);
xnor U1247 (N_1247,N_475,In_118);
nor U1248 (N_1248,In_1807,N_902);
xnor U1249 (N_1249,N_124,N_888);
and U1250 (N_1250,N_448,N_1217);
and U1251 (N_1251,In_1,N_191);
nand U1252 (N_1252,N_1029,N_1228);
or U1253 (N_1253,In_1343,N_848);
xnor U1254 (N_1254,N_1131,In_339);
or U1255 (N_1255,In_616,N_1185);
nor U1256 (N_1256,N_1012,N_106);
nor U1257 (N_1257,In_146,N_866);
xor U1258 (N_1258,In_1810,N_999);
xor U1259 (N_1259,N_190,N_1054);
nand U1260 (N_1260,N_1208,N_970);
or U1261 (N_1261,N_1221,In_1347);
and U1262 (N_1262,N_1220,N_1127);
nor U1263 (N_1263,N_834,In_1690);
nand U1264 (N_1264,N_783,N_919);
or U1265 (N_1265,N_1032,N_1085);
xnor U1266 (N_1266,N_405,In_681);
and U1267 (N_1267,N_954,N_271);
nand U1268 (N_1268,In_15,N_1162);
or U1269 (N_1269,N_613,N_1199);
nor U1270 (N_1270,N_821,In_1363);
or U1271 (N_1271,N_973,N_991);
or U1272 (N_1272,N_1030,In_1099);
nor U1273 (N_1273,N_616,N_1070);
nor U1274 (N_1274,N_598,N_1041);
xor U1275 (N_1275,N_1049,N_879);
and U1276 (N_1276,N_348,N_1215);
xor U1277 (N_1277,In_542,N_548);
xnor U1278 (N_1278,N_1202,N_1109);
and U1279 (N_1279,N_931,N_1059);
and U1280 (N_1280,N_1100,In_1251);
or U1281 (N_1281,N_1181,N_946);
nand U1282 (N_1282,N_1184,N_1018);
and U1283 (N_1283,N_1058,In_337);
nand U1284 (N_1284,N_168,In_1608);
or U1285 (N_1285,N_109,In_1616);
xnor U1286 (N_1286,In_1478,In_1003);
nand U1287 (N_1287,In_272,N_1246);
nand U1288 (N_1288,In_1619,N_628);
xnor U1289 (N_1289,N_385,In_128);
xnor U1290 (N_1290,N_1017,N_237);
nor U1291 (N_1291,In_1225,N_763);
xnor U1292 (N_1292,N_253,N_1237);
or U1293 (N_1293,In_373,N_70);
nand U1294 (N_1294,In_186,N_670);
or U1295 (N_1295,N_864,N_1105);
or U1296 (N_1296,N_882,N_614);
xnor U1297 (N_1297,N_620,N_514);
nor U1298 (N_1298,N_817,N_11);
nor U1299 (N_1299,In_1109,N_1243);
or U1300 (N_1300,N_1024,In_331);
nand U1301 (N_1301,In_1256,N_14);
or U1302 (N_1302,In_1880,N_1056);
nand U1303 (N_1303,N_663,In_1564);
nor U1304 (N_1304,N_1229,N_509);
and U1305 (N_1305,N_1027,N_1075);
or U1306 (N_1306,N_1089,In_488);
and U1307 (N_1307,N_1120,N_683);
and U1308 (N_1308,N_1174,In_1651);
nand U1309 (N_1309,N_1239,In_1713);
xnor U1310 (N_1310,N_1133,N_266);
and U1311 (N_1311,N_41,N_1212);
xnor U1312 (N_1312,N_803,N_1126);
or U1313 (N_1313,N_1216,In_562);
nand U1314 (N_1314,N_1214,N_1044);
nand U1315 (N_1315,N_956,N_1067);
and U1316 (N_1316,N_1065,In_95);
nor U1317 (N_1317,In_635,N_1233);
nand U1318 (N_1318,N_1159,N_165);
xor U1319 (N_1319,N_480,N_1128);
nor U1320 (N_1320,N_1028,N_831);
or U1321 (N_1321,N_1110,N_358);
nand U1322 (N_1322,N_971,In_506);
xnor U1323 (N_1323,N_1223,N_552);
xnor U1324 (N_1324,N_1234,N_600);
nand U1325 (N_1325,N_389,N_658);
and U1326 (N_1326,N_836,N_1203);
and U1327 (N_1327,N_1061,N_6);
or U1328 (N_1328,In_1942,N_839);
nor U1329 (N_1329,In_799,In_879);
xor U1330 (N_1330,N_529,In_582);
xnor U1331 (N_1331,N_654,N_850);
and U1332 (N_1332,N_64,In_47);
or U1333 (N_1333,In_209,In_157);
xor U1334 (N_1334,N_1153,N_380);
xnor U1335 (N_1335,N_1121,N_661);
and U1336 (N_1336,In_252,N_1198);
nor U1337 (N_1337,N_1062,N_743);
nand U1338 (N_1338,N_491,N_1063);
and U1339 (N_1339,N_384,N_1069);
and U1340 (N_1340,N_881,N_845);
nand U1341 (N_1341,N_1046,In_618);
xor U1342 (N_1342,In_1840,In_895);
and U1343 (N_1343,N_1037,N_1112);
or U1344 (N_1344,N_1057,N_1204);
nor U1345 (N_1345,N_820,In_773);
nor U1346 (N_1346,In_1952,N_1115);
xnor U1347 (N_1347,In_1436,N_511);
xor U1348 (N_1348,N_1164,In_583);
nor U1349 (N_1349,N_1172,In_1445);
xnor U1350 (N_1350,N_521,N_773);
or U1351 (N_1351,N_328,N_563);
or U1352 (N_1352,In_980,N_972);
and U1353 (N_1353,N_1145,In_1600);
xor U1354 (N_1354,N_796,In_664);
nand U1355 (N_1355,N_1156,N_1118);
xor U1356 (N_1356,N_929,N_826);
nand U1357 (N_1357,N_700,N_1014);
or U1358 (N_1358,In_1473,N_1242);
xnor U1359 (N_1359,N_181,N_1169);
xor U1360 (N_1360,N_822,N_1043);
nand U1361 (N_1361,N_1151,In_653);
nor U1362 (N_1362,N_312,N_1102);
or U1363 (N_1363,N_1008,N_1210);
nand U1364 (N_1364,N_996,N_738);
xor U1365 (N_1365,In_638,N_1178);
or U1366 (N_1366,In_1062,N_828);
xor U1367 (N_1367,N_550,N_1135);
nor U1368 (N_1368,In_1105,N_969);
nand U1369 (N_1369,N_761,N_186);
nand U1370 (N_1370,N_404,In_1956);
or U1371 (N_1371,N_1146,N_1015);
nand U1372 (N_1372,N_1188,N_1137);
nand U1373 (N_1373,N_799,N_659);
nand U1374 (N_1374,N_742,N_953);
xnor U1375 (N_1375,N_921,N_1073);
xor U1376 (N_1376,N_74,N_887);
nand U1377 (N_1377,In_317,N_284);
nor U1378 (N_1378,N_1175,N_357);
nor U1379 (N_1379,N_1147,N_73);
xor U1380 (N_1380,In_1904,N_652);
nand U1381 (N_1381,N_1114,In_66);
or U1382 (N_1382,In_1871,N_908);
or U1383 (N_1383,In_898,N_1087);
and U1384 (N_1384,N_1108,N_524);
nand U1385 (N_1385,N_304,N_1116);
or U1386 (N_1386,N_1084,N_1072);
or U1387 (N_1387,N_1196,In_1671);
or U1388 (N_1388,In_1043,N_33);
nand U1389 (N_1389,N_906,In_374);
nand U1390 (N_1390,N_184,N_912);
nor U1391 (N_1391,N_707,N_1230);
nor U1392 (N_1392,In_1950,In_654);
and U1393 (N_1393,In_927,In_1644);
xor U1394 (N_1394,N_1077,In_1701);
or U1395 (N_1395,N_1231,N_556);
nand U1396 (N_1396,N_816,In_926);
xnor U1397 (N_1397,N_1213,N_1094);
nor U1398 (N_1398,N_1139,N_327);
or U1399 (N_1399,N_114,N_751);
nand U1400 (N_1400,N_1152,N_1157);
nand U1401 (N_1401,N_914,N_1244);
nor U1402 (N_1402,N_1066,N_786);
nand U1403 (N_1403,N_856,N_775);
and U1404 (N_1404,N_1197,N_804);
nor U1405 (N_1405,In_907,N_390);
or U1406 (N_1406,N_772,N_793);
and U1407 (N_1407,In_1444,In_920);
xnor U1408 (N_1408,In_1468,N_1119);
nand U1409 (N_1409,N_623,N_354);
and U1410 (N_1410,N_819,N_250);
nor U1411 (N_1411,N_1019,N_717);
nor U1412 (N_1412,N_435,N_1107);
nor U1413 (N_1413,N_1142,In_1341);
nand U1414 (N_1414,N_1248,N_77);
or U1415 (N_1415,N_860,N_353);
xnor U1416 (N_1416,N_1141,N_44);
nand U1417 (N_1417,In_1797,N_1171);
and U1418 (N_1418,In_1591,N_1038);
nor U1419 (N_1419,In_432,N_1211);
or U1420 (N_1420,N_815,N_1103);
nor U1421 (N_1421,In_138,N_749);
nor U1422 (N_1422,N_1240,N_941);
nand U1423 (N_1423,N_218,N_885);
nor U1424 (N_1424,N_392,In_1993);
and U1425 (N_1425,N_69,N_639);
or U1426 (N_1426,N_986,N_797);
or U1427 (N_1427,N_753,N_952);
xnor U1428 (N_1428,N_1150,N_1106);
nand U1429 (N_1429,N_818,N_1039);
xnor U1430 (N_1430,N_674,N_20);
and U1431 (N_1431,In_1082,N_1098);
and U1432 (N_1432,N_1206,N_160);
xnor U1433 (N_1433,N_1140,N_170);
nand U1434 (N_1434,In_565,N_944);
xnor U1435 (N_1435,N_557,N_606);
and U1436 (N_1436,N_984,N_1193);
xor U1437 (N_1437,N_852,N_195);
and U1438 (N_1438,N_306,N_927);
nand U1439 (N_1439,N_1144,In_428);
and U1440 (N_1440,N_1083,N_1090);
xnor U1441 (N_1441,N_538,N_1051);
xnor U1442 (N_1442,N_439,N_499);
and U1443 (N_1443,In_1967,N_558);
or U1444 (N_1444,N_1060,N_1071);
or U1445 (N_1445,N_1022,N_1003);
xnor U1446 (N_1446,In_96,In_1125);
or U1447 (N_1447,In_559,N_875);
xor U1448 (N_1448,N_843,N_1096);
and U1449 (N_1449,N_429,N_15);
nor U1450 (N_1450,N_1124,N_1191);
and U1451 (N_1451,N_1088,N_292);
or U1452 (N_1452,N_894,N_779);
nand U1453 (N_1453,N_899,N_1036);
nand U1454 (N_1454,N_744,N_484);
and U1455 (N_1455,N_1183,In_391);
nor U1456 (N_1456,N_1200,In_622);
or U1457 (N_1457,In_851,N_756);
or U1458 (N_1458,N_923,In_168);
and U1459 (N_1459,N_1097,N_928);
or U1460 (N_1460,N_924,N_1117);
nand U1461 (N_1461,N_1190,N_1192);
nor U1462 (N_1462,N_1177,N_141);
nor U1463 (N_1463,N_285,N_1123);
nand U1464 (N_1464,N_65,N_1189);
nand U1465 (N_1465,N_1173,In_165);
xor U1466 (N_1466,N_644,N_1122);
or U1467 (N_1467,In_1947,In_249);
nor U1468 (N_1468,In_1497,N_1180);
nand U1469 (N_1469,N_580,N_1167);
xor U1470 (N_1470,N_1093,N_62);
nor U1471 (N_1471,N_325,N_858);
nor U1472 (N_1472,In_1323,In_236);
and U1473 (N_1473,In_1316,In_253);
nor U1474 (N_1474,In_1399,In_1482);
or U1475 (N_1475,N_1045,N_1021);
and U1476 (N_1476,In_827,In_1960);
nor U1477 (N_1477,N_951,N_766);
and U1478 (N_1478,In_340,In_808);
or U1479 (N_1479,N_1050,In_713);
nor U1480 (N_1480,In_627,N_1194);
or U1481 (N_1481,In_572,N_1130);
nor U1482 (N_1482,N_911,In_175);
nand U1483 (N_1483,N_629,N_870);
nor U1484 (N_1484,N_878,In_909);
xor U1485 (N_1485,N_1226,N_621);
nand U1486 (N_1486,In_181,N_777);
nand U1487 (N_1487,N_1149,N_1086);
nand U1488 (N_1488,N_224,N_647);
xor U1489 (N_1489,N_739,N_1179);
or U1490 (N_1490,N_672,In_1732);
and U1491 (N_1491,N_734,N_1138);
and U1492 (N_1492,N_458,N_1091);
nor U1493 (N_1493,N_1201,N_1195);
or U1494 (N_1494,N_857,In_1022);
xor U1495 (N_1495,N_1074,N_1010);
xnor U1496 (N_1496,N_759,In_1552);
xnor U1497 (N_1497,N_1236,N_920);
and U1498 (N_1498,N_559,N_1166);
xor U1499 (N_1499,N_454,N_1055);
and U1500 (N_1500,N_837,N_1489);
or U1501 (N_1501,N_1255,N_1272);
and U1502 (N_1502,In_722,N_545);
and U1503 (N_1503,N_814,N_412);
nor U1504 (N_1504,N_1047,N_1373);
nor U1505 (N_1505,N_1444,N_1431);
xor U1506 (N_1506,N_1472,In_1527);
or U1507 (N_1507,N_1443,In_1248);
nor U1508 (N_1508,In_1913,N_1414);
nor U1509 (N_1509,In_24,N_792);
nand U1510 (N_1510,N_1493,N_1318);
nand U1511 (N_1511,In_1521,N_1437);
and U1512 (N_1512,N_72,N_942);
and U1513 (N_1513,N_1005,In_1955);
nand U1514 (N_1514,N_1295,N_1366);
xnor U1515 (N_1515,N_1161,In_1850);
nor U1516 (N_1516,N_1483,N_1264);
nor U1517 (N_1517,N_1345,N_950);
nand U1518 (N_1518,N_1378,In_258);
xnor U1519 (N_1519,N_1446,N_1241);
nand U1520 (N_1520,N_827,N_1439);
xor U1521 (N_1521,In_1284,In_472);
nand U1522 (N_1522,N_516,N_1409);
nor U1523 (N_1523,N_1370,N_1297);
xor U1524 (N_1524,N_855,N_1315);
and U1525 (N_1525,N_1336,N_1485);
nand U1526 (N_1526,N_1249,N_1285);
xor U1527 (N_1527,N_1286,In_1757);
nand U1528 (N_1528,N_1325,N_1372);
nor U1529 (N_1529,N_1328,N_1284);
or U1530 (N_1530,N_338,N_1476);
and U1531 (N_1531,N_1379,N_1497);
and U1532 (N_1532,N_1434,N_1319);
nor U1533 (N_1533,N_978,N_599);
xnor U1534 (N_1534,In_514,N_1253);
xor U1535 (N_1535,N_1304,N_1256);
nor U1536 (N_1536,N_1321,N_1148);
nor U1537 (N_1537,N_1488,N_347);
xnor U1538 (N_1538,In_1140,In_74);
and U1539 (N_1539,N_1031,N_1491);
or U1540 (N_1540,N_1092,N_1270);
xnor U1541 (N_1541,N_853,N_1467);
nor U1542 (N_1542,N_1298,N_1251);
nor U1543 (N_1543,N_806,N_1362);
nand U1544 (N_1544,N_585,N_788);
or U1545 (N_1545,In_1016,N_397);
xnor U1546 (N_1546,In_1013,N_905);
or U1547 (N_1547,N_1368,N_1445);
and U1548 (N_1548,N_1397,N_85);
nor U1549 (N_1549,In_1804,N_1435);
nor U1550 (N_1550,In_1789,N_1388);
or U1551 (N_1551,N_1020,N_417);
nand U1552 (N_1552,In_708,N_642);
and U1553 (N_1553,N_1333,N_1398);
nor U1554 (N_1554,In_223,N_1099);
and U1555 (N_1555,N_1371,N_564);
and U1556 (N_1556,N_1068,N_1411);
or U1557 (N_1557,In_1309,N_1396);
nor U1558 (N_1558,In_1261,N_1104);
or U1559 (N_1559,N_1129,N_1430);
nor U1560 (N_1560,N_1267,N_1125);
xor U1561 (N_1561,In_1005,N_504);
and U1562 (N_1562,N_1222,N_528);
nor U1563 (N_1563,N_593,N_1487);
nand U1564 (N_1564,N_650,N_222);
nand U1565 (N_1565,N_1405,N_1323);
nand U1566 (N_1566,N_1335,In_1832);
nor U1567 (N_1567,N_1040,N_750);
nand U1568 (N_1568,N_1274,N_1235);
xor U1569 (N_1569,N_1425,N_1268);
nor U1570 (N_1570,N_1324,In_1715);
or U1571 (N_1571,N_531,N_1475);
or U1572 (N_1572,N_326,N_1498);
nand U1573 (N_1573,N_1064,N_1471);
nor U1574 (N_1574,N_962,N_1026);
xor U1575 (N_1575,In_1575,N_1095);
xnor U1576 (N_1576,N_1305,N_1224);
and U1577 (N_1577,N_1001,In_569);
xor U1578 (N_1578,N_1205,N_876);
nor U1579 (N_1579,In_466,In_1858);
or U1580 (N_1580,N_896,In_1539);
and U1581 (N_1581,In_590,N_1484);
or U1582 (N_1582,In_1888,N_1413);
or U1583 (N_1583,N_1299,N_1283);
and U1584 (N_1584,N_1386,N_1155);
and U1585 (N_1585,N_1355,N_1219);
nor U1586 (N_1586,N_1160,N_1410);
nor U1587 (N_1587,N_1207,N_1154);
nor U1588 (N_1588,N_1081,N_1495);
xor U1589 (N_1589,N_1348,In_645);
xnor U1590 (N_1590,N_640,N_1136);
nor U1591 (N_1591,In_928,N_1006);
xor U1592 (N_1592,N_1302,N_1269);
or U1593 (N_1593,N_1496,N_1265);
and U1594 (N_1594,N_1438,N_1310);
nor U1595 (N_1595,N_1399,N_1314);
and U1596 (N_1596,N_1352,N_1479);
or U1597 (N_1597,In_1301,N_1412);
nor U1598 (N_1598,N_1260,N_1327);
nor U1599 (N_1599,N_926,N_1347);
and U1600 (N_1600,N_1186,N_1307);
xor U1601 (N_1601,N_1406,N_1331);
nand U1602 (N_1602,N_615,In_1058);
nor U1603 (N_1603,N_1360,N_1428);
and U1604 (N_1604,N_1432,N_1048);
or U1605 (N_1605,In_1364,N_1025);
or U1606 (N_1606,N_1429,N_1261);
nand U1607 (N_1607,N_1400,In_671);
xnor U1608 (N_1608,N_1232,In_1249);
or U1609 (N_1609,N_1459,N_5);
nor U1610 (N_1610,N_1296,In_1189);
and U1611 (N_1611,In_715,N_1293);
or U1612 (N_1612,N_955,N_1004);
or U1613 (N_1613,N_200,In_1331);
nand U1614 (N_1614,N_278,N_79);
nand U1615 (N_1615,N_1344,N_630);
nor U1616 (N_1616,N_1341,N_1182);
xor U1617 (N_1617,N_1482,N_1433);
and U1618 (N_1618,N_1395,N_1292);
nor U1619 (N_1619,N_1225,In_1799);
nor U1620 (N_1620,N_1000,In_989);
or U1621 (N_1621,N_1374,N_1448);
nand U1622 (N_1622,N_1357,N_1458);
and U1623 (N_1623,N_1408,In_16);
and U1624 (N_1624,N_1455,N_507);
or U1625 (N_1625,N_1342,N_1440);
nor U1626 (N_1626,N_959,N_1453);
xnor U1627 (N_1627,N_1023,In_1425);
nand U1628 (N_1628,N_1394,N_651);
and U1629 (N_1629,N_1417,N_1474);
and U1630 (N_1630,In_1228,N_1277);
nand U1631 (N_1631,N_1490,N_1460);
and U1632 (N_1632,N_1011,N_589);
or U1633 (N_1633,N_1113,N_1282);
nor U1634 (N_1634,In_552,N_1415);
nor U1635 (N_1635,N_735,In_334);
xnor U1636 (N_1636,N_1381,N_1245);
or U1637 (N_1637,N_1387,N_517);
nor U1638 (N_1638,N_1257,N_1424);
or U1639 (N_1639,In_471,N_1078);
or U1640 (N_1640,In_1541,N_1404);
and U1641 (N_1641,N_708,In_1029);
nor U1642 (N_1642,N_1168,N_975);
or U1643 (N_1643,N_859,N_1421);
nand U1644 (N_1644,N_1499,N_1456);
nand U1645 (N_1645,N_1076,N_915);
or U1646 (N_1646,In_1268,N_1376);
or U1647 (N_1647,N_1053,N_1468);
nand U1648 (N_1648,In_397,N_1469);
nor U1649 (N_1649,N_53,In_698);
or U1650 (N_1650,N_1486,N_1457);
or U1651 (N_1651,In_735,In_1532);
or U1652 (N_1652,N_1402,N_1303);
nand U1653 (N_1653,N_1452,N_1393);
xnor U1654 (N_1654,N_1266,N_904);
or U1655 (N_1655,N_1392,N_1442);
xor U1656 (N_1656,N_627,N_1382);
and U1657 (N_1657,N_829,In_819);
and U1658 (N_1658,N_442,N_1111);
or U1659 (N_1659,N_459,N_1329);
or U1660 (N_1660,N_862,N_1466);
or U1661 (N_1661,N_1367,N_592);
or U1662 (N_1662,In_1208,N_1492);
or U1663 (N_1663,In_1611,N_1473);
or U1664 (N_1664,N_1470,N_1449);
nor U1665 (N_1665,N_1291,N_1290);
nor U1666 (N_1666,N_1422,In_897);
or U1667 (N_1667,N_1289,N_957);
nor U1668 (N_1668,N_687,N_1326);
nor U1669 (N_1669,N_1401,N_1300);
and U1670 (N_1670,N_469,In_1096);
or U1671 (N_1671,N_335,N_1481);
nor U1672 (N_1672,N_785,N_1377);
nand U1673 (N_1673,N_1306,N_1353);
xnor U1674 (N_1674,N_1238,N_1480);
nor U1675 (N_1675,N_305,N_1247);
or U1676 (N_1676,N_1317,N_1254);
or U1677 (N_1677,N_1407,N_1132);
and U1678 (N_1678,N_1101,N_1134);
xor U1679 (N_1679,N_1451,N_1350);
xor U1680 (N_1680,N_1450,N_1158);
xnor U1681 (N_1681,N_1013,N_765);
and U1682 (N_1682,In_885,N_1280);
nand U1683 (N_1683,N_1369,N_1187);
nand U1684 (N_1684,N_1351,N_1176);
xnor U1685 (N_1685,In_1976,N_1389);
nand U1686 (N_1686,N_1170,N_1494);
nand U1687 (N_1687,N_1227,N_309);
and U1688 (N_1688,N_1423,N_1454);
or U1689 (N_1689,N_1359,N_1034);
nand U1690 (N_1690,N_961,In_22);
and U1691 (N_1691,N_1294,N_711);
nor U1692 (N_1692,N_1312,N_1346);
nor U1693 (N_1693,N_1477,N_1320);
nor U1694 (N_1694,N_1384,N_1337);
or U1695 (N_1695,N_1079,N_1441);
and U1696 (N_1696,N_154,N_398);
and U1697 (N_1697,N_769,N_1276);
xor U1698 (N_1698,N_1271,N_1383);
or U1699 (N_1699,In_281,N_1316);
or U1700 (N_1700,N_1339,N_1082);
and U1701 (N_1701,N_985,N_1163);
and U1702 (N_1702,N_1349,N_1322);
or U1703 (N_1703,N_1016,N_1385);
nor U1704 (N_1704,N_1313,In_976);
nor U1705 (N_1705,N_1363,N_830);
and U1706 (N_1706,In_1702,N_1002);
and U1707 (N_1707,N_1165,In_389);
xor U1708 (N_1708,In_1604,In_1902);
and U1709 (N_1709,N_1009,In_1387);
nor U1710 (N_1710,N_1465,N_1143);
and U1711 (N_1711,N_447,N_1463);
xnor U1712 (N_1712,N_1426,N_1301);
and U1713 (N_1713,N_1042,N_1380);
and U1714 (N_1714,N_1287,N_1461);
and U1715 (N_1715,In_1382,In_1071);
nand U1716 (N_1716,N_1259,N_1262);
and U1717 (N_1717,N_982,In_191);
and U1718 (N_1718,N_1436,N_1288);
and U1719 (N_1719,N_1361,N_1334);
and U1720 (N_1720,N_1338,N_1464);
xor U1721 (N_1721,N_776,N_1364);
or U1722 (N_1722,N_1209,N_1250);
and U1723 (N_1723,N_1033,N_1447);
nand U1724 (N_1724,N_1332,N_1309);
and U1725 (N_1725,N_1007,In_914);
nor U1726 (N_1726,N_1308,N_897);
or U1727 (N_1727,In_963,N_1427);
and U1728 (N_1728,N_1218,N_1403);
or U1729 (N_1729,N_1281,N_1252);
nor U1730 (N_1730,N_789,N_1419);
nor U1731 (N_1731,N_111,N_939);
or U1732 (N_1732,N_1275,N_1420);
or U1733 (N_1733,N_1416,N_1340);
xor U1734 (N_1734,In_1441,N_1035);
or U1735 (N_1735,N_369,N_1052);
xor U1736 (N_1736,N_476,N_1258);
and U1737 (N_1737,N_1375,N_1358);
or U1738 (N_1738,N_1478,N_1080);
or U1739 (N_1739,N_1263,N_1418);
nor U1740 (N_1740,N_1330,N_998);
nand U1741 (N_1741,N_1273,N_1462);
xor U1742 (N_1742,N_1343,N_1279);
and U1743 (N_1743,N_760,N_1356);
nand U1744 (N_1744,N_1391,In_9);
xor U1745 (N_1745,N_1390,N_980);
and U1746 (N_1746,N_371,N_918);
and U1747 (N_1747,In_1174,N_1354);
nor U1748 (N_1748,N_1311,N_1278);
nand U1749 (N_1749,N_1365,N_741);
or U1750 (N_1750,N_1523,N_1589);
nor U1751 (N_1751,N_1609,N_1507);
nand U1752 (N_1752,N_1720,N_1729);
nand U1753 (N_1753,N_1695,N_1534);
or U1754 (N_1754,N_1651,N_1579);
xor U1755 (N_1755,N_1559,N_1600);
or U1756 (N_1756,N_1510,N_1558);
nand U1757 (N_1757,N_1658,N_1553);
nand U1758 (N_1758,N_1667,N_1554);
nor U1759 (N_1759,N_1563,N_1685);
xor U1760 (N_1760,N_1619,N_1670);
and U1761 (N_1761,N_1679,N_1546);
nand U1762 (N_1762,N_1728,N_1623);
or U1763 (N_1763,N_1578,N_1747);
and U1764 (N_1764,N_1624,N_1749);
and U1765 (N_1765,N_1731,N_1565);
xnor U1766 (N_1766,N_1644,N_1739);
xor U1767 (N_1767,N_1719,N_1687);
nand U1768 (N_1768,N_1590,N_1712);
nand U1769 (N_1769,N_1628,N_1723);
and U1770 (N_1770,N_1668,N_1528);
nand U1771 (N_1771,N_1652,N_1604);
nand U1772 (N_1772,N_1716,N_1606);
nor U1773 (N_1773,N_1694,N_1707);
nand U1774 (N_1774,N_1574,N_1616);
and U1775 (N_1775,N_1690,N_1625);
nor U1776 (N_1776,N_1557,N_1536);
nand U1777 (N_1777,N_1529,N_1708);
nand U1778 (N_1778,N_1602,N_1542);
and U1779 (N_1779,N_1673,N_1566);
and U1780 (N_1780,N_1521,N_1618);
or U1781 (N_1781,N_1552,N_1586);
and U1782 (N_1782,N_1741,N_1575);
xor U1783 (N_1783,N_1620,N_1517);
and U1784 (N_1784,N_1615,N_1656);
xor U1785 (N_1785,N_1700,N_1727);
or U1786 (N_1786,N_1539,N_1519);
xnor U1787 (N_1787,N_1568,N_1653);
xnor U1788 (N_1788,N_1648,N_1674);
or U1789 (N_1789,N_1631,N_1621);
nand U1790 (N_1790,N_1530,N_1540);
and U1791 (N_1791,N_1638,N_1664);
nand U1792 (N_1792,N_1655,N_1681);
xnor U1793 (N_1793,N_1743,N_1689);
nor U1794 (N_1794,N_1662,N_1630);
and U1795 (N_1795,N_1649,N_1748);
nor U1796 (N_1796,N_1520,N_1524);
or U1797 (N_1797,N_1587,N_1617);
nand U1798 (N_1798,N_1585,N_1646);
xor U1799 (N_1799,N_1550,N_1715);
nor U1800 (N_1800,N_1610,N_1663);
and U1801 (N_1801,N_1725,N_1561);
nor U1802 (N_1802,N_1556,N_1591);
nand U1803 (N_1803,N_1533,N_1698);
nand U1804 (N_1804,N_1746,N_1537);
nor U1805 (N_1805,N_1596,N_1511);
and U1806 (N_1806,N_1629,N_1726);
nand U1807 (N_1807,N_1669,N_1547);
and U1808 (N_1808,N_1732,N_1696);
nor U1809 (N_1809,N_1639,N_1583);
and U1810 (N_1810,N_1601,N_1595);
nor U1811 (N_1811,N_1582,N_1594);
or U1812 (N_1812,N_1612,N_1635);
nor U1813 (N_1813,N_1686,N_1714);
nand U1814 (N_1814,N_1541,N_1647);
nand U1815 (N_1815,N_1645,N_1675);
nor U1816 (N_1816,N_1730,N_1703);
nand U1817 (N_1817,N_1504,N_1665);
or U1818 (N_1818,N_1721,N_1622);
or U1819 (N_1819,N_1570,N_1581);
and U1820 (N_1820,N_1538,N_1508);
and U1821 (N_1821,N_1532,N_1598);
or U1822 (N_1822,N_1567,N_1682);
xor U1823 (N_1823,N_1643,N_1704);
xnor U1824 (N_1824,N_1505,N_1584);
and U1825 (N_1825,N_1642,N_1580);
nand U1826 (N_1826,N_1636,N_1509);
xor U1827 (N_1827,N_1683,N_1657);
nor U1828 (N_1828,N_1692,N_1611);
or U1829 (N_1829,N_1702,N_1503);
or U1830 (N_1830,N_1706,N_1734);
nand U1831 (N_1831,N_1603,N_1699);
nor U1832 (N_1832,N_1548,N_1733);
and U1833 (N_1833,N_1654,N_1684);
and U1834 (N_1834,N_1551,N_1576);
nand U1835 (N_1835,N_1697,N_1614);
xnor U1836 (N_1836,N_1597,N_1672);
nor U1837 (N_1837,N_1717,N_1560);
or U1838 (N_1838,N_1711,N_1626);
or U1839 (N_1839,N_1605,N_1713);
nor U1840 (N_1840,N_1738,N_1724);
or U1841 (N_1841,N_1593,N_1531);
nor U1842 (N_1842,N_1737,N_1709);
xor U1843 (N_1843,N_1502,N_1710);
nand U1844 (N_1844,N_1599,N_1627);
xnor U1845 (N_1845,N_1691,N_1588);
nand U1846 (N_1846,N_1513,N_1633);
and U1847 (N_1847,N_1564,N_1514);
nand U1848 (N_1848,N_1543,N_1634);
nand U1849 (N_1849,N_1677,N_1705);
xor U1850 (N_1850,N_1640,N_1592);
xnor U1851 (N_1851,N_1607,N_1659);
nand U1852 (N_1852,N_1577,N_1678);
nor U1853 (N_1853,N_1722,N_1506);
nor U1854 (N_1854,N_1525,N_1745);
and U1855 (N_1855,N_1718,N_1660);
xor U1856 (N_1856,N_1641,N_1744);
nand U1857 (N_1857,N_1736,N_1572);
nand U1858 (N_1858,N_1501,N_1637);
or U1859 (N_1859,N_1676,N_1512);
xor U1860 (N_1860,N_1545,N_1526);
xor U1861 (N_1861,N_1516,N_1742);
xor U1862 (N_1862,N_1544,N_1701);
or U1863 (N_1863,N_1518,N_1688);
nand U1864 (N_1864,N_1735,N_1680);
nand U1865 (N_1865,N_1515,N_1671);
nand U1866 (N_1866,N_1535,N_1522);
nor U1867 (N_1867,N_1573,N_1500);
nand U1868 (N_1868,N_1740,N_1569);
or U1869 (N_1869,N_1693,N_1608);
nand U1870 (N_1870,N_1555,N_1527);
and U1871 (N_1871,N_1650,N_1666);
xnor U1872 (N_1872,N_1562,N_1661);
nand U1873 (N_1873,N_1571,N_1549);
or U1874 (N_1874,N_1632,N_1613);
and U1875 (N_1875,N_1648,N_1657);
xor U1876 (N_1876,N_1720,N_1632);
and U1877 (N_1877,N_1693,N_1670);
or U1878 (N_1878,N_1615,N_1523);
or U1879 (N_1879,N_1588,N_1598);
or U1880 (N_1880,N_1742,N_1512);
nor U1881 (N_1881,N_1719,N_1713);
xnor U1882 (N_1882,N_1673,N_1589);
xor U1883 (N_1883,N_1515,N_1704);
and U1884 (N_1884,N_1561,N_1737);
nand U1885 (N_1885,N_1712,N_1701);
or U1886 (N_1886,N_1697,N_1601);
and U1887 (N_1887,N_1717,N_1680);
and U1888 (N_1888,N_1639,N_1570);
nand U1889 (N_1889,N_1748,N_1504);
xor U1890 (N_1890,N_1582,N_1565);
nor U1891 (N_1891,N_1724,N_1582);
xnor U1892 (N_1892,N_1568,N_1548);
and U1893 (N_1893,N_1627,N_1706);
xor U1894 (N_1894,N_1542,N_1721);
and U1895 (N_1895,N_1616,N_1556);
nand U1896 (N_1896,N_1649,N_1536);
or U1897 (N_1897,N_1511,N_1510);
or U1898 (N_1898,N_1635,N_1664);
and U1899 (N_1899,N_1581,N_1671);
xnor U1900 (N_1900,N_1611,N_1512);
nor U1901 (N_1901,N_1649,N_1702);
nand U1902 (N_1902,N_1622,N_1634);
nand U1903 (N_1903,N_1539,N_1647);
nor U1904 (N_1904,N_1672,N_1509);
xor U1905 (N_1905,N_1738,N_1549);
xnor U1906 (N_1906,N_1698,N_1563);
nand U1907 (N_1907,N_1653,N_1676);
or U1908 (N_1908,N_1629,N_1551);
or U1909 (N_1909,N_1684,N_1612);
or U1910 (N_1910,N_1530,N_1678);
nand U1911 (N_1911,N_1689,N_1520);
and U1912 (N_1912,N_1723,N_1587);
nor U1913 (N_1913,N_1622,N_1682);
nand U1914 (N_1914,N_1625,N_1684);
or U1915 (N_1915,N_1618,N_1732);
nor U1916 (N_1916,N_1634,N_1581);
xor U1917 (N_1917,N_1713,N_1746);
nor U1918 (N_1918,N_1741,N_1616);
nor U1919 (N_1919,N_1600,N_1649);
or U1920 (N_1920,N_1734,N_1717);
or U1921 (N_1921,N_1685,N_1730);
nand U1922 (N_1922,N_1634,N_1696);
and U1923 (N_1923,N_1570,N_1680);
xor U1924 (N_1924,N_1617,N_1719);
xor U1925 (N_1925,N_1578,N_1535);
nor U1926 (N_1926,N_1720,N_1556);
and U1927 (N_1927,N_1741,N_1577);
and U1928 (N_1928,N_1598,N_1559);
or U1929 (N_1929,N_1524,N_1570);
nand U1930 (N_1930,N_1510,N_1679);
xor U1931 (N_1931,N_1569,N_1586);
or U1932 (N_1932,N_1627,N_1519);
nand U1933 (N_1933,N_1508,N_1729);
and U1934 (N_1934,N_1588,N_1736);
and U1935 (N_1935,N_1651,N_1711);
and U1936 (N_1936,N_1672,N_1606);
nand U1937 (N_1937,N_1748,N_1608);
nor U1938 (N_1938,N_1615,N_1695);
xor U1939 (N_1939,N_1730,N_1668);
nor U1940 (N_1940,N_1594,N_1637);
xnor U1941 (N_1941,N_1559,N_1694);
or U1942 (N_1942,N_1658,N_1556);
xnor U1943 (N_1943,N_1744,N_1564);
and U1944 (N_1944,N_1735,N_1737);
and U1945 (N_1945,N_1551,N_1654);
xor U1946 (N_1946,N_1547,N_1665);
and U1947 (N_1947,N_1704,N_1529);
or U1948 (N_1948,N_1525,N_1513);
nor U1949 (N_1949,N_1642,N_1703);
or U1950 (N_1950,N_1504,N_1574);
xnor U1951 (N_1951,N_1692,N_1708);
and U1952 (N_1952,N_1649,N_1580);
nor U1953 (N_1953,N_1538,N_1676);
nand U1954 (N_1954,N_1544,N_1747);
or U1955 (N_1955,N_1618,N_1717);
or U1956 (N_1956,N_1665,N_1649);
xor U1957 (N_1957,N_1598,N_1547);
nand U1958 (N_1958,N_1531,N_1734);
xor U1959 (N_1959,N_1512,N_1715);
nor U1960 (N_1960,N_1643,N_1617);
and U1961 (N_1961,N_1745,N_1554);
nand U1962 (N_1962,N_1576,N_1675);
xor U1963 (N_1963,N_1631,N_1587);
nor U1964 (N_1964,N_1646,N_1679);
or U1965 (N_1965,N_1667,N_1726);
and U1966 (N_1966,N_1743,N_1716);
nand U1967 (N_1967,N_1646,N_1687);
nand U1968 (N_1968,N_1507,N_1697);
nand U1969 (N_1969,N_1725,N_1682);
and U1970 (N_1970,N_1747,N_1525);
nand U1971 (N_1971,N_1515,N_1591);
and U1972 (N_1972,N_1703,N_1561);
xor U1973 (N_1973,N_1610,N_1668);
and U1974 (N_1974,N_1636,N_1619);
nand U1975 (N_1975,N_1536,N_1734);
xnor U1976 (N_1976,N_1744,N_1548);
nor U1977 (N_1977,N_1595,N_1571);
nand U1978 (N_1978,N_1574,N_1698);
and U1979 (N_1979,N_1522,N_1605);
or U1980 (N_1980,N_1536,N_1743);
or U1981 (N_1981,N_1742,N_1565);
xnor U1982 (N_1982,N_1617,N_1545);
or U1983 (N_1983,N_1546,N_1733);
xnor U1984 (N_1984,N_1614,N_1744);
xor U1985 (N_1985,N_1700,N_1666);
nor U1986 (N_1986,N_1711,N_1740);
xnor U1987 (N_1987,N_1677,N_1525);
nor U1988 (N_1988,N_1592,N_1633);
xor U1989 (N_1989,N_1741,N_1615);
xnor U1990 (N_1990,N_1654,N_1527);
nand U1991 (N_1991,N_1562,N_1734);
nand U1992 (N_1992,N_1584,N_1659);
xor U1993 (N_1993,N_1710,N_1560);
nor U1994 (N_1994,N_1519,N_1684);
nand U1995 (N_1995,N_1733,N_1675);
xnor U1996 (N_1996,N_1642,N_1570);
nand U1997 (N_1997,N_1560,N_1700);
nand U1998 (N_1998,N_1536,N_1707);
and U1999 (N_1999,N_1685,N_1526);
xor U2000 (N_2000,N_1986,N_1762);
nor U2001 (N_2001,N_1993,N_1833);
or U2002 (N_2002,N_1752,N_1936);
xnor U2003 (N_2003,N_1763,N_1850);
and U2004 (N_2004,N_1807,N_1965);
or U2005 (N_2005,N_1854,N_1857);
and U2006 (N_2006,N_1921,N_1964);
nand U2007 (N_2007,N_1924,N_1975);
nor U2008 (N_2008,N_1751,N_1870);
and U2009 (N_2009,N_1816,N_1800);
or U2010 (N_2010,N_1979,N_1764);
xor U2011 (N_2011,N_1977,N_1983);
xor U2012 (N_2012,N_1848,N_1943);
or U2013 (N_2013,N_1847,N_1889);
and U2014 (N_2014,N_1892,N_1903);
or U2015 (N_2015,N_1830,N_1788);
xnor U2016 (N_2016,N_1840,N_1877);
and U2017 (N_2017,N_1786,N_1759);
or U2018 (N_2018,N_1799,N_1766);
xnor U2019 (N_2019,N_1996,N_1901);
nor U2020 (N_2020,N_1904,N_1770);
or U2021 (N_2021,N_1822,N_1789);
nor U2022 (N_2022,N_1970,N_1980);
nor U2023 (N_2023,N_1942,N_1930);
xnor U2024 (N_2024,N_1928,N_1905);
nand U2025 (N_2025,N_1793,N_1771);
nand U2026 (N_2026,N_1960,N_1939);
or U2027 (N_2027,N_1769,N_1869);
and U2028 (N_2028,N_1796,N_1785);
or U2029 (N_2029,N_1966,N_1932);
nor U2030 (N_2030,N_1864,N_1772);
nand U2031 (N_2031,N_1898,N_1909);
nand U2032 (N_2032,N_1838,N_1859);
or U2033 (N_2033,N_1837,N_1817);
and U2034 (N_2034,N_1866,N_1842);
and U2035 (N_2035,N_1795,N_1907);
or U2036 (N_2036,N_1856,N_1908);
xor U2037 (N_2037,N_1949,N_1841);
and U2038 (N_2038,N_1931,N_1805);
or U2039 (N_2039,N_1997,N_1897);
nor U2040 (N_2040,N_1821,N_1814);
nor U2041 (N_2041,N_1803,N_1792);
xnor U2042 (N_2042,N_1768,N_1999);
nor U2043 (N_2043,N_1899,N_1783);
or U2044 (N_2044,N_1961,N_1784);
nor U2045 (N_2045,N_1829,N_1948);
nand U2046 (N_2046,N_1982,N_1998);
and U2047 (N_2047,N_1990,N_1994);
and U2048 (N_2048,N_1851,N_1945);
and U2049 (N_2049,N_1860,N_1969);
xnor U2050 (N_2050,N_1956,N_1810);
nor U2051 (N_2051,N_1875,N_1826);
and U2052 (N_2052,N_1957,N_1801);
nand U2053 (N_2053,N_1972,N_1767);
and U2054 (N_2054,N_1765,N_1884);
nand U2055 (N_2055,N_1846,N_1887);
nand U2056 (N_2056,N_1828,N_1871);
nand U2057 (N_2057,N_1820,N_1872);
and U2058 (N_2058,N_1937,N_1926);
or U2059 (N_2059,N_1802,N_1813);
xnor U2060 (N_2060,N_1987,N_1849);
nand U2061 (N_2061,N_1776,N_1779);
xnor U2062 (N_2062,N_1865,N_1981);
nand U2063 (N_2063,N_1852,N_1912);
or U2064 (N_2064,N_1818,N_1873);
xnor U2065 (N_2065,N_1919,N_1750);
and U2066 (N_2066,N_1910,N_1955);
xnor U2067 (N_2067,N_1843,N_1882);
nand U2068 (N_2068,N_1973,N_1781);
and U2069 (N_2069,N_1774,N_1777);
and U2070 (N_2070,N_1918,N_1878);
xor U2071 (N_2071,N_1933,N_1985);
and U2072 (N_2072,N_1791,N_1946);
or U2073 (N_2073,N_1782,N_1974);
and U2074 (N_2074,N_1845,N_1809);
and U2075 (N_2075,N_1773,N_1855);
or U2076 (N_2076,N_1951,N_1927);
and U2077 (N_2077,N_1911,N_1940);
and U2078 (N_2078,N_1804,N_1893);
or U2079 (N_2079,N_1868,N_1885);
xor U2080 (N_2080,N_1760,N_1978);
and U2081 (N_2081,N_1950,N_1758);
or U2082 (N_2082,N_1929,N_1844);
xnor U2083 (N_2083,N_1883,N_1881);
or U2084 (N_2084,N_1958,N_1876);
nor U2085 (N_2085,N_1819,N_1995);
or U2086 (N_2086,N_1780,N_1963);
or U2087 (N_2087,N_1863,N_1823);
or U2088 (N_2088,N_1836,N_1879);
xor U2089 (N_2089,N_1935,N_1756);
nor U2090 (N_2090,N_1944,N_1811);
and U2091 (N_2091,N_1754,N_1874);
xor U2092 (N_2092,N_1976,N_1967);
nand U2093 (N_2093,N_1968,N_1984);
or U2094 (N_2094,N_1775,N_1920);
or U2095 (N_2095,N_1915,N_1954);
and U2096 (N_2096,N_1992,N_1839);
nand U2097 (N_2097,N_1886,N_1867);
or U2098 (N_2098,N_1971,N_1916);
nand U2099 (N_2099,N_1798,N_1894);
or U2100 (N_2100,N_1753,N_1806);
xor U2101 (N_2101,N_1991,N_1858);
or U2102 (N_2102,N_1896,N_1922);
and U2103 (N_2103,N_1962,N_1757);
or U2104 (N_2104,N_1988,N_1906);
xnor U2105 (N_2105,N_1890,N_1953);
nand U2106 (N_2106,N_1861,N_1835);
nor U2107 (N_2107,N_1941,N_1808);
nand U2108 (N_2108,N_1853,N_1934);
and U2109 (N_2109,N_1834,N_1880);
and U2110 (N_2110,N_1761,N_1815);
or U2111 (N_2111,N_1888,N_1900);
xnor U2112 (N_2112,N_1952,N_1925);
xnor U2113 (N_2113,N_1902,N_1959);
nand U2114 (N_2114,N_1923,N_1862);
or U2115 (N_2115,N_1790,N_1947);
or U2116 (N_2116,N_1825,N_1797);
xor U2117 (N_2117,N_1827,N_1778);
and U2118 (N_2118,N_1891,N_1914);
or U2119 (N_2119,N_1917,N_1824);
nand U2120 (N_2120,N_1812,N_1794);
nand U2121 (N_2121,N_1755,N_1938);
xnor U2122 (N_2122,N_1913,N_1831);
nand U2123 (N_2123,N_1989,N_1895);
nor U2124 (N_2124,N_1832,N_1787);
or U2125 (N_2125,N_1801,N_1895);
or U2126 (N_2126,N_1900,N_1916);
xnor U2127 (N_2127,N_1822,N_1811);
xnor U2128 (N_2128,N_1751,N_1774);
xnor U2129 (N_2129,N_1840,N_1889);
or U2130 (N_2130,N_1821,N_1806);
nor U2131 (N_2131,N_1817,N_1859);
nand U2132 (N_2132,N_1783,N_1939);
xnor U2133 (N_2133,N_1803,N_1800);
nand U2134 (N_2134,N_1825,N_1995);
xor U2135 (N_2135,N_1972,N_1915);
xor U2136 (N_2136,N_1947,N_1808);
nor U2137 (N_2137,N_1821,N_1824);
nand U2138 (N_2138,N_1905,N_1986);
and U2139 (N_2139,N_1903,N_1887);
nand U2140 (N_2140,N_1936,N_1814);
or U2141 (N_2141,N_1796,N_1849);
nor U2142 (N_2142,N_1772,N_1803);
nand U2143 (N_2143,N_1751,N_1780);
nor U2144 (N_2144,N_1979,N_1860);
or U2145 (N_2145,N_1818,N_1859);
or U2146 (N_2146,N_1804,N_1949);
nor U2147 (N_2147,N_1887,N_1895);
and U2148 (N_2148,N_1893,N_1967);
or U2149 (N_2149,N_1969,N_1888);
nand U2150 (N_2150,N_1915,N_1798);
xnor U2151 (N_2151,N_1956,N_1760);
or U2152 (N_2152,N_1833,N_1942);
or U2153 (N_2153,N_1821,N_1975);
nor U2154 (N_2154,N_1778,N_1799);
xor U2155 (N_2155,N_1886,N_1890);
nand U2156 (N_2156,N_1862,N_1891);
and U2157 (N_2157,N_1782,N_1928);
xnor U2158 (N_2158,N_1985,N_1823);
nor U2159 (N_2159,N_1956,N_1828);
or U2160 (N_2160,N_1778,N_1980);
xnor U2161 (N_2161,N_1845,N_1825);
nor U2162 (N_2162,N_1949,N_1954);
nor U2163 (N_2163,N_1963,N_1897);
or U2164 (N_2164,N_1941,N_1930);
or U2165 (N_2165,N_1963,N_1761);
and U2166 (N_2166,N_1869,N_1990);
xor U2167 (N_2167,N_1897,N_1931);
xor U2168 (N_2168,N_1997,N_1877);
xor U2169 (N_2169,N_1823,N_1798);
or U2170 (N_2170,N_1925,N_1934);
xor U2171 (N_2171,N_1872,N_1869);
nor U2172 (N_2172,N_1790,N_1768);
or U2173 (N_2173,N_1957,N_1848);
or U2174 (N_2174,N_1916,N_1771);
and U2175 (N_2175,N_1764,N_1925);
nand U2176 (N_2176,N_1923,N_1956);
nand U2177 (N_2177,N_1901,N_1962);
xor U2178 (N_2178,N_1811,N_1921);
xor U2179 (N_2179,N_1769,N_1806);
xnor U2180 (N_2180,N_1959,N_1858);
or U2181 (N_2181,N_1798,N_1877);
xnor U2182 (N_2182,N_1820,N_1857);
or U2183 (N_2183,N_1846,N_1978);
nand U2184 (N_2184,N_1750,N_1944);
or U2185 (N_2185,N_1965,N_1801);
xor U2186 (N_2186,N_1897,N_1763);
nand U2187 (N_2187,N_1759,N_1819);
nand U2188 (N_2188,N_1764,N_1863);
nand U2189 (N_2189,N_1925,N_1923);
nor U2190 (N_2190,N_1780,N_1944);
nor U2191 (N_2191,N_1905,N_1913);
nand U2192 (N_2192,N_1796,N_1952);
xnor U2193 (N_2193,N_1975,N_1921);
nand U2194 (N_2194,N_1910,N_1841);
xnor U2195 (N_2195,N_1913,N_1756);
or U2196 (N_2196,N_1756,N_1797);
and U2197 (N_2197,N_1912,N_1805);
nand U2198 (N_2198,N_1854,N_1856);
and U2199 (N_2199,N_1788,N_1808);
nor U2200 (N_2200,N_1938,N_1901);
or U2201 (N_2201,N_1964,N_1972);
nand U2202 (N_2202,N_1834,N_1890);
or U2203 (N_2203,N_1999,N_1818);
and U2204 (N_2204,N_1762,N_1897);
xor U2205 (N_2205,N_1960,N_1789);
nor U2206 (N_2206,N_1863,N_1957);
or U2207 (N_2207,N_1969,N_1965);
or U2208 (N_2208,N_1769,N_1800);
or U2209 (N_2209,N_1879,N_1983);
nor U2210 (N_2210,N_1968,N_1812);
xnor U2211 (N_2211,N_1980,N_1764);
and U2212 (N_2212,N_1895,N_1944);
and U2213 (N_2213,N_1905,N_1941);
nand U2214 (N_2214,N_1787,N_1960);
nand U2215 (N_2215,N_1971,N_1967);
and U2216 (N_2216,N_1975,N_1957);
nor U2217 (N_2217,N_1761,N_1854);
xor U2218 (N_2218,N_1774,N_1959);
or U2219 (N_2219,N_1972,N_1863);
and U2220 (N_2220,N_1989,N_1831);
or U2221 (N_2221,N_1866,N_1974);
nand U2222 (N_2222,N_1907,N_1992);
nor U2223 (N_2223,N_1876,N_1840);
xor U2224 (N_2224,N_1935,N_1885);
xnor U2225 (N_2225,N_1828,N_1902);
or U2226 (N_2226,N_1829,N_1862);
nand U2227 (N_2227,N_1987,N_1881);
nand U2228 (N_2228,N_1906,N_1763);
or U2229 (N_2229,N_1850,N_1844);
xnor U2230 (N_2230,N_1750,N_1902);
or U2231 (N_2231,N_1819,N_1912);
nand U2232 (N_2232,N_1932,N_1999);
and U2233 (N_2233,N_1773,N_1774);
xor U2234 (N_2234,N_1970,N_1988);
and U2235 (N_2235,N_1836,N_1822);
nand U2236 (N_2236,N_1832,N_1774);
nand U2237 (N_2237,N_1976,N_1754);
nand U2238 (N_2238,N_1892,N_1951);
xor U2239 (N_2239,N_1897,N_1872);
nor U2240 (N_2240,N_1891,N_1954);
or U2241 (N_2241,N_1972,N_1904);
xor U2242 (N_2242,N_1882,N_1946);
nand U2243 (N_2243,N_1849,N_1967);
or U2244 (N_2244,N_1899,N_1864);
or U2245 (N_2245,N_1793,N_1864);
nand U2246 (N_2246,N_1982,N_1972);
or U2247 (N_2247,N_1984,N_1787);
or U2248 (N_2248,N_1807,N_1978);
and U2249 (N_2249,N_1836,N_1943);
xor U2250 (N_2250,N_2151,N_2220);
xor U2251 (N_2251,N_2224,N_2006);
nor U2252 (N_2252,N_2127,N_2197);
and U2253 (N_2253,N_2155,N_2124);
or U2254 (N_2254,N_2175,N_2041);
xor U2255 (N_2255,N_2013,N_2085);
nor U2256 (N_2256,N_2071,N_2033);
xor U2257 (N_2257,N_2196,N_2183);
and U2258 (N_2258,N_2168,N_2156);
and U2259 (N_2259,N_2239,N_2027);
xnor U2260 (N_2260,N_2089,N_2055);
and U2261 (N_2261,N_2116,N_2083);
nand U2262 (N_2262,N_2024,N_2077);
xor U2263 (N_2263,N_2115,N_2218);
nor U2264 (N_2264,N_2081,N_2159);
and U2265 (N_2265,N_2130,N_2017);
or U2266 (N_2266,N_2063,N_2189);
nand U2267 (N_2267,N_2018,N_2091);
xnor U2268 (N_2268,N_2148,N_2019);
xnor U2269 (N_2269,N_2057,N_2074);
xor U2270 (N_2270,N_2061,N_2079);
or U2271 (N_2271,N_2160,N_2244);
nand U2272 (N_2272,N_2126,N_2051);
or U2273 (N_2273,N_2246,N_2180);
or U2274 (N_2274,N_2212,N_2075);
nand U2275 (N_2275,N_2119,N_2045);
and U2276 (N_2276,N_2170,N_2149);
nand U2277 (N_2277,N_2090,N_2078);
and U2278 (N_2278,N_2199,N_2167);
or U2279 (N_2279,N_2166,N_2191);
or U2280 (N_2280,N_2198,N_2144);
nor U2281 (N_2281,N_2137,N_2223);
and U2282 (N_2282,N_2094,N_2141);
xor U2283 (N_2283,N_2228,N_2248);
xnor U2284 (N_2284,N_2049,N_2125);
nor U2285 (N_2285,N_2139,N_2229);
nor U2286 (N_2286,N_2140,N_2046);
xnor U2287 (N_2287,N_2179,N_2206);
nor U2288 (N_2288,N_2120,N_2190);
or U2289 (N_2289,N_2186,N_2000);
nand U2290 (N_2290,N_2106,N_2087);
xor U2291 (N_2291,N_2009,N_2203);
nor U2292 (N_2292,N_2054,N_2242);
nor U2293 (N_2293,N_2042,N_2213);
nor U2294 (N_2294,N_2100,N_2164);
nor U2295 (N_2295,N_2038,N_2134);
nand U2296 (N_2296,N_2034,N_2172);
and U2297 (N_2297,N_2059,N_2030);
and U2298 (N_2298,N_2007,N_2010);
and U2299 (N_2299,N_2105,N_2211);
and U2300 (N_2300,N_2008,N_2112);
or U2301 (N_2301,N_2048,N_2145);
nor U2302 (N_2302,N_2240,N_2236);
xnor U2303 (N_2303,N_2247,N_2058);
nand U2304 (N_2304,N_2044,N_2073);
nor U2305 (N_2305,N_2020,N_2204);
or U2306 (N_2306,N_2084,N_2221);
and U2307 (N_2307,N_2110,N_2152);
nor U2308 (N_2308,N_2029,N_2052);
or U2309 (N_2309,N_2237,N_2205);
nand U2310 (N_2310,N_2118,N_2096);
nand U2311 (N_2311,N_2171,N_2249);
or U2312 (N_2312,N_2067,N_2104);
and U2313 (N_2313,N_2202,N_2114);
nor U2314 (N_2314,N_2080,N_2177);
nand U2315 (N_2315,N_2226,N_2210);
xor U2316 (N_2316,N_2113,N_2109);
and U2317 (N_2317,N_2178,N_2142);
and U2318 (N_2318,N_2003,N_2011);
nor U2319 (N_2319,N_2117,N_2016);
xor U2320 (N_2320,N_2238,N_2146);
and U2321 (N_2321,N_2157,N_2088);
nor U2322 (N_2322,N_2069,N_2014);
or U2323 (N_2323,N_2005,N_2022);
and U2324 (N_2324,N_2209,N_2219);
or U2325 (N_2325,N_2121,N_2215);
xor U2326 (N_2326,N_2173,N_2214);
and U2327 (N_2327,N_2193,N_2165);
and U2328 (N_2328,N_2241,N_2043);
nor U2329 (N_2329,N_2064,N_2195);
and U2330 (N_2330,N_2092,N_2101);
nand U2331 (N_2331,N_2185,N_2111);
nand U2332 (N_2332,N_2181,N_2047);
nand U2333 (N_2333,N_2216,N_2143);
xnor U2334 (N_2334,N_2086,N_2163);
xor U2335 (N_2335,N_2035,N_2093);
nor U2336 (N_2336,N_2053,N_2135);
nor U2337 (N_2337,N_2028,N_2200);
or U2338 (N_2338,N_2040,N_2245);
or U2339 (N_2339,N_2072,N_2023);
or U2340 (N_2340,N_2133,N_2026);
nor U2341 (N_2341,N_2129,N_2230);
xor U2342 (N_2342,N_2147,N_2066);
and U2343 (N_2343,N_2138,N_2076);
nand U2344 (N_2344,N_2187,N_2002);
nor U2345 (N_2345,N_2004,N_2231);
and U2346 (N_2346,N_2222,N_2182);
nor U2347 (N_2347,N_2184,N_2037);
nand U2348 (N_2348,N_2050,N_2031);
and U2349 (N_2349,N_2136,N_2001);
nand U2350 (N_2350,N_2161,N_2158);
xnor U2351 (N_2351,N_2103,N_2032);
and U2352 (N_2352,N_2056,N_2235);
and U2353 (N_2353,N_2068,N_2122);
xor U2354 (N_2354,N_2169,N_2107);
or U2355 (N_2355,N_2060,N_2123);
or U2356 (N_2356,N_2174,N_2097);
nor U2357 (N_2357,N_2025,N_2062);
xnor U2358 (N_2358,N_2012,N_2217);
and U2359 (N_2359,N_2201,N_2194);
nand U2360 (N_2360,N_2207,N_2225);
nand U2361 (N_2361,N_2015,N_2070);
xor U2362 (N_2362,N_2232,N_2102);
xnor U2363 (N_2363,N_2243,N_2036);
and U2364 (N_2364,N_2021,N_2098);
or U2365 (N_2365,N_2208,N_2162);
nor U2366 (N_2366,N_2082,N_2065);
nor U2367 (N_2367,N_2039,N_2234);
and U2368 (N_2368,N_2128,N_2095);
nand U2369 (N_2369,N_2099,N_2227);
xnor U2370 (N_2370,N_2153,N_2154);
nor U2371 (N_2371,N_2132,N_2108);
and U2372 (N_2372,N_2150,N_2176);
or U2373 (N_2373,N_2188,N_2233);
and U2374 (N_2374,N_2192,N_2131);
nand U2375 (N_2375,N_2055,N_2131);
and U2376 (N_2376,N_2178,N_2174);
nand U2377 (N_2377,N_2170,N_2083);
nor U2378 (N_2378,N_2064,N_2036);
and U2379 (N_2379,N_2235,N_2173);
nor U2380 (N_2380,N_2170,N_2017);
nand U2381 (N_2381,N_2121,N_2239);
or U2382 (N_2382,N_2104,N_2007);
xnor U2383 (N_2383,N_2171,N_2036);
or U2384 (N_2384,N_2234,N_2052);
and U2385 (N_2385,N_2219,N_2218);
nor U2386 (N_2386,N_2061,N_2060);
and U2387 (N_2387,N_2001,N_2162);
xnor U2388 (N_2388,N_2080,N_2182);
xor U2389 (N_2389,N_2130,N_2128);
nand U2390 (N_2390,N_2018,N_2236);
and U2391 (N_2391,N_2063,N_2158);
xor U2392 (N_2392,N_2214,N_2016);
xor U2393 (N_2393,N_2203,N_2099);
nor U2394 (N_2394,N_2011,N_2128);
nand U2395 (N_2395,N_2090,N_2214);
or U2396 (N_2396,N_2245,N_2239);
nor U2397 (N_2397,N_2058,N_2053);
or U2398 (N_2398,N_2015,N_2129);
nor U2399 (N_2399,N_2105,N_2157);
or U2400 (N_2400,N_2093,N_2063);
nor U2401 (N_2401,N_2209,N_2197);
and U2402 (N_2402,N_2175,N_2005);
nor U2403 (N_2403,N_2090,N_2216);
and U2404 (N_2404,N_2112,N_2142);
or U2405 (N_2405,N_2199,N_2194);
and U2406 (N_2406,N_2187,N_2082);
and U2407 (N_2407,N_2134,N_2069);
xor U2408 (N_2408,N_2177,N_2051);
or U2409 (N_2409,N_2067,N_2061);
nor U2410 (N_2410,N_2018,N_2036);
xnor U2411 (N_2411,N_2022,N_2042);
and U2412 (N_2412,N_2249,N_2077);
and U2413 (N_2413,N_2111,N_2093);
xor U2414 (N_2414,N_2071,N_2126);
nor U2415 (N_2415,N_2041,N_2238);
nor U2416 (N_2416,N_2041,N_2075);
nand U2417 (N_2417,N_2079,N_2170);
nand U2418 (N_2418,N_2188,N_2192);
or U2419 (N_2419,N_2018,N_2008);
or U2420 (N_2420,N_2148,N_2028);
nor U2421 (N_2421,N_2151,N_2143);
and U2422 (N_2422,N_2161,N_2051);
and U2423 (N_2423,N_2009,N_2145);
and U2424 (N_2424,N_2217,N_2138);
nor U2425 (N_2425,N_2109,N_2214);
and U2426 (N_2426,N_2161,N_2120);
nand U2427 (N_2427,N_2025,N_2090);
xor U2428 (N_2428,N_2027,N_2192);
and U2429 (N_2429,N_2081,N_2246);
xor U2430 (N_2430,N_2207,N_2242);
or U2431 (N_2431,N_2123,N_2229);
nand U2432 (N_2432,N_2086,N_2211);
nor U2433 (N_2433,N_2073,N_2023);
nor U2434 (N_2434,N_2179,N_2045);
and U2435 (N_2435,N_2178,N_2065);
and U2436 (N_2436,N_2158,N_2006);
nand U2437 (N_2437,N_2204,N_2223);
and U2438 (N_2438,N_2020,N_2245);
nor U2439 (N_2439,N_2099,N_2235);
xor U2440 (N_2440,N_2200,N_2017);
nor U2441 (N_2441,N_2087,N_2038);
or U2442 (N_2442,N_2064,N_2031);
nand U2443 (N_2443,N_2238,N_2049);
or U2444 (N_2444,N_2029,N_2034);
nand U2445 (N_2445,N_2105,N_2119);
nor U2446 (N_2446,N_2102,N_2212);
or U2447 (N_2447,N_2029,N_2069);
and U2448 (N_2448,N_2003,N_2181);
xor U2449 (N_2449,N_2009,N_2079);
nor U2450 (N_2450,N_2125,N_2078);
nor U2451 (N_2451,N_2083,N_2220);
nor U2452 (N_2452,N_2067,N_2224);
nor U2453 (N_2453,N_2113,N_2213);
and U2454 (N_2454,N_2121,N_2145);
nand U2455 (N_2455,N_2124,N_2243);
and U2456 (N_2456,N_2066,N_2231);
or U2457 (N_2457,N_2056,N_2059);
and U2458 (N_2458,N_2068,N_2216);
and U2459 (N_2459,N_2119,N_2180);
or U2460 (N_2460,N_2020,N_2080);
xor U2461 (N_2461,N_2097,N_2061);
nor U2462 (N_2462,N_2081,N_2051);
nand U2463 (N_2463,N_2078,N_2183);
or U2464 (N_2464,N_2090,N_2244);
nand U2465 (N_2465,N_2104,N_2161);
nand U2466 (N_2466,N_2144,N_2216);
nand U2467 (N_2467,N_2091,N_2185);
or U2468 (N_2468,N_2158,N_2178);
nand U2469 (N_2469,N_2121,N_2020);
nor U2470 (N_2470,N_2050,N_2201);
and U2471 (N_2471,N_2090,N_2100);
or U2472 (N_2472,N_2019,N_2117);
or U2473 (N_2473,N_2102,N_2106);
nand U2474 (N_2474,N_2184,N_2161);
and U2475 (N_2475,N_2184,N_2144);
or U2476 (N_2476,N_2129,N_2237);
xnor U2477 (N_2477,N_2175,N_2058);
nand U2478 (N_2478,N_2114,N_2134);
nor U2479 (N_2479,N_2189,N_2234);
nor U2480 (N_2480,N_2030,N_2148);
nor U2481 (N_2481,N_2122,N_2027);
xnor U2482 (N_2482,N_2213,N_2198);
nor U2483 (N_2483,N_2031,N_2188);
nor U2484 (N_2484,N_2194,N_2183);
or U2485 (N_2485,N_2155,N_2186);
and U2486 (N_2486,N_2242,N_2003);
or U2487 (N_2487,N_2170,N_2019);
nand U2488 (N_2488,N_2070,N_2007);
xor U2489 (N_2489,N_2106,N_2171);
xor U2490 (N_2490,N_2082,N_2149);
xor U2491 (N_2491,N_2038,N_2023);
xor U2492 (N_2492,N_2188,N_2200);
xnor U2493 (N_2493,N_2127,N_2190);
or U2494 (N_2494,N_2033,N_2110);
nor U2495 (N_2495,N_2015,N_2200);
xnor U2496 (N_2496,N_2233,N_2078);
or U2497 (N_2497,N_2199,N_2031);
nand U2498 (N_2498,N_2158,N_2179);
nand U2499 (N_2499,N_2124,N_2185);
or U2500 (N_2500,N_2286,N_2485);
nor U2501 (N_2501,N_2493,N_2268);
xor U2502 (N_2502,N_2334,N_2272);
or U2503 (N_2503,N_2435,N_2499);
nand U2504 (N_2504,N_2403,N_2339);
and U2505 (N_2505,N_2322,N_2384);
nor U2506 (N_2506,N_2353,N_2447);
or U2507 (N_2507,N_2423,N_2329);
or U2508 (N_2508,N_2360,N_2488);
nand U2509 (N_2509,N_2266,N_2480);
and U2510 (N_2510,N_2290,N_2377);
or U2511 (N_2511,N_2388,N_2416);
nand U2512 (N_2512,N_2490,N_2291);
or U2513 (N_2513,N_2457,N_2308);
xor U2514 (N_2514,N_2301,N_2252);
nor U2515 (N_2515,N_2316,N_2453);
and U2516 (N_2516,N_2305,N_2309);
xnor U2517 (N_2517,N_2426,N_2477);
nor U2518 (N_2518,N_2469,N_2460);
xor U2519 (N_2519,N_2347,N_2487);
and U2520 (N_2520,N_2415,N_2393);
and U2521 (N_2521,N_2411,N_2313);
nand U2522 (N_2522,N_2276,N_2376);
nand U2523 (N_2523,N_2385,N_2267);
nor U2524 (N_2524,N_2364,N_2307);
or U2525 (N_2525,N_2293,N_2401);
nor U2526 (N_2526,N_2427,N_2408);
and U2527 (N_2527,N_2273,N_2303);
and U2528 (N_2528,N_2369,N_2304);
nor U2529 (N_2529,N_2349,N_2254);
or U2530 (N_2530,N_2310,N_2467);
or U2531 (N_2531,N_2399,N_2440);
or U2532 (N_2532,N_2341,N_2260);
and U2533 (N_2533,N_2358,N_2259);
or U2534 (N_2534,N_2354,N_2294);
nand U2535 (N_2535,N_2483,N_2434);
xnor U2536 (N_2536,N_2263,N_2312);
xor U2537 (N_2537,N_2251,N_2441);
nand U2538 (N_2538,N_2298,N_2466);
nor U2539 (N_2539,N_2470,N_2359);
nor U2540 (N_2540,N_2314,N_2438);
or U2541 (N_2541,N_2336,N_2255);
nand U2542 (N_2542,N_2431,N_2279);
or U2543 (N_2543,N_2278,N_2381);
nor U2544 (N_2544,N_2425,N_2397);
and U2545 (N_2545,N_2253,N_2407);
and U2546 (N_2546,N_2283,N_2287);
xnor U2547 (N_2547,N_2390,N_2482);
nor U2548 (N_2548,N_2264,N_2335);
and U2549 (N_2549,N_2420,N_2437);
xnor U2550 (N_2550,N_2323,N_2451);
or U2551 (N_2551,N_2424,N_2296);
nor U2552 (N_2552,N_2345,N_2495);
or U2553 (N_2553,N_2311,N_2474);
nand U2554 (N_2554,N_2327,N_2449);
or U2555 (N_2555,N_2414,N_2400);
nand U2556 (N_2556,N_2362,N_2321);
and U2557 (N_2557,N_2378,N_2281);
nor U2558 (N_2558,N_2394,N_2465);
and U2559 (N_2559,N_2455,N_2459);
or U2560 (N_2560,N_2475,N_2406);
xor U2561 (N_2561,N_2270,N_2257);
and U2562 (N_2562,N_2444,N_2478);
nand U2563 (N_2563,N_2300,N_2452);
xor U2564 (N_2564,N_2492,N_2256);
nand U2565 (N_2565,N_2484,N_2356);
or U2566 (N_2566,N_2436,N_2413);
nor U2567 (N_2567,N_2328,N_2456);
xnor U2568 (N_2568,N_2285,N_2379);
or U2569 (N_2569,N_2491,N_2396);
nand U2570 (N_2570,N_2315,N_2419);
nor U2571 (N_2571,N_2391,N_2338);
and U2572 (N_2572,N_2386,N_2498);
nand U2573 (N_2573,N_2422,N_2370);
xor U2574 (N_2574,N_2486,N_2258);
nand U2575 (N_2575,N_2325,N_2463);
xnor U2576 (N_2576,N_2383,N_2439);
or U2577 (N_2577,N_2375,N_2371);
xnor U2578 (N_2578,N_2344,N_2412);
or U2579 (N_2579,N_2275,N_2472);
xor U2580 (N_2580,N_2489,N_2332);
xor U2581 (N_2581,N_2404,N_2446);
and U2582 (N_2582,N_2355,N_2350);
nand U2583 (N_2583,N_2357,N_2271);
nand U2584 (N_2584,N_2331,N_2297);
nand U2585 (N_2585,N_2342,N_2481);
xnor U2586 (N_2586,N_2318,N_2269);
nor U2587 (N_2587,N_2330,N_2405);
and U2588 (N_2588,N_2471,N_2433);
or U2589 (N_2589,N_2461,N_2365);
nor U2590 (N_2590,N_2380,N_2250);
nand U2591 (N_2591,N_2429,N_2458);
or U2592 (N_2592,N_2351,N_2346);
nor U2593 (N_2593,N_2348,N_2363);
or U2594 (N_2594,N_2374,N_2421);
nor U2595 (N_2595,N_2366,N_2448);
xnor U2596 (N_2596,N_2450,N_2464);
nor U2597 (N_2597,N_2468,N_2292);
or U2598 (N_2598,N_2274,N_2432);
xnor U2599 (N_2599,N_2295,N_2352);
xnor U2600 (N_2600,N_2382,N_2337);
or U2601 (N_2601,N_2387,N_2299);
nand U2602 (N_2602,N_2430,N_2302);
nor U2603 (N_2603,N_2306,N_2261);
nor U2604 (N_2604,N_2288,N_2284);
nor U2605 (N_2605,N_2410,N_2343);
and U2606 (N_2606,N_2392,N_2454);
nor U2607 (N_2607,N_2417,N_2473);
nand U2608 (N_2608,N_2428,N_2262);
nand U2609 (N_2609,N_2418,N_2333);
nor U2610 (N_2610,N_2367,N_2445);
xor U2611 (N_2611,N_2277,N_2373);
nand U2612 (N_2612,N_2280,N_2324);
or U2613 (N_2613,N_2320,N_2340);
xnor U2614 (N_2614,N_2326,N_2282);
and U2615 (N_2615,N_2479,N_2409);
xor U2616 (N_2616,N_2494,N_2497);
xor U2617 (N_2617,N_2289,N_2402);
and U2618 (N_2618,N_2319,N_2476);
or U2619 (N_2619,N_2368,N_2442);
nor U2620 (N_2620,N_2265,N_2443);
nand U2621 (N_2621,N_2389,N_2361);
nand U2622 (N_2622,N_2317,N_2398);
nand U2623 (N_2623,N_2372,N_2496);
nor U2624 (N_2624,N_2395,N_2462);
and U2625 (N_2625,N_2377,N_2472);
and U2626 (N_2626,N_2280,N_2496);
xnor U2627 (N_2627,N_2302,N_2357);
or U2628 (N_2628,N_2301,N_2473);
nand U2629 (N_2629,N_2364,N_2254);
or U2630 (N_2630,N_2294,N_2482);
nand U2631 (N_2631,N_2460,N_2376);
or U2632 (N_2632,N_2330,N_2347);
or U2633 (N_2633,N_2286,N_2452);
or U2634 (N_2634,N_2395,N_2265);
or U2635 (N_2635,N_2432,N_2317);
nor U2636 (N_2636,N_2492,N_2298);
nor U2637 (N_2637,N_2382,N_2401);
nand U2638 (N_2638,N_2386,N_2256);
and U2639 (N_2639,N_2485,N_2299);
and U2640 (N_2640,N_2376,N_2306);
nand U2641 (N_2641,N_2291,N_2366);
xnor U2642 (N_2642,N_2279,N_2476);
nand U2643 (N_2643,N_2439,N_2271);
nor U2644 (N_2644,N_2370,N_2458);
nor U2645 (N_2645,N_2470,N_2265);
or U2646 (N_2646,N_2488,N_2266);
xor U2647 (N_2647,N_2259,N_2339);
nand U2648 (N_2648,N_2496,N_2314);
or U2649 (N_2649,N_2281,N_2316);
and U2650 (N_2650,N_2330,N_2277);
xnor U2651 (N_2651,N_2477,N_2470);
or U2652 (N_2652,N_2350,N_2284);
and U2653 (N_2653,N_2414,N_2453);
xor U2654 (N_2654,N_2299,N_2428);
xnor U2655 (N_2655,N_2257,N_2440);
nor U2656 (N_2656,N_2473,N_2462);
and U2657 (N_2657,N_2404,N_2283);
and U2658 (N_2658,N_2277,N_2362);
nand U2659 (N_2659,N_2324,N_2391);
nand U2660 (N_2660,N_2306,N_2265);
and U2661 (N_2661,N_2308,N_2498);
or U2662 (N_2662,N_2271,N_2346);
nand U2663 (N_2663,N_2437,N_2337);
and U2664 (N_2664,N_2285,N_2329);
and U2665 (N_2665,N_2333,N_2474);
and U2666 (N_2666,N_2382,N_2482);
and U2667 (N_2667,N_2459,N_2291);
or U2668 (N_2668,N_2266,N_2340);
or U2669 (N_2669,N_2450,N_2369);
or U2670 (N_2670,N_2495,N_2325);
or U2671 (N_2671,N_2322,N_2416);
nand U2672 (N_2672,N_2476,N_2454);
nor U2673 (N_2673,N_2396,N_2330);
or U2674 (N_2674,N_2465,N_2359);
xnor U2675 (N_2675,N_2493,N_2395);
or U2676 (N_2676,N_2381,N_2477);
or U2677 (N_2677,N_2255,N_2411);
xnor U2678 (N_2678,N_2370,N_2250);
nor U2679 (N_2679,N_2298,N_2442);
nand U2680 (N_2680,N_2255,N_2293);
and U2681 (N_2681,N_2331,N_2493);
nand U2682 (N_2682,N_2438,N_2339);
nand U2683 (N_2683,N_2451,N_2291);
nor U2684 (N_2684,N_2279,N_2313);
nor U2685 (N_2685,N_2288,N_2386);
and U2686 (N_2686,N_2465,N_2311);
xor U2687 (N_2687,N_2330,N_2335);
nand U2688 (N_2688,N_2272,N_2492);
nor U2689 (N_2689,N_2383,N_2406);
or U2690 (N_2690,N_2372,N_2394);
and U2691 (N_2691,N_2352,N_2350);
nor U2692 (N_2692,N_2482,N_2254);
nor U2693 (N_2693,N_2439,N_2400);
and U2694 (N_2694,N_2334,N_2250);
xor U2695 (N_2695,N_2468,N_2453);
nand U2696 (N_2696,N_2482,N_2445);
or U2697 (N_2697,N_2456,N_2374);
and U2698 (N_2698,N_2282,N_2389);
nor U2699 (N_2699,N_2403,N_2456);
nand U2700 (N_2700,N_2435,N_2372);
and U2701 (N_2701,N_2341,N_2419);
or U2702 (N_2702,N_2313,N_2287);
nor U2703 (N_2703,N_2472,N_2332);
nand U2704 (N_2704,N_2389,N_2435);
or U2705 (N_2705,N_2309,N_2260);
or U2706 (N_2706,N_2286,N_2379);
nor U2707 (N_2707,N_2368,N_2263);
nand U2708 (N_2708,N_2337,N_2359);
xnor U2709 (N_2709,N_2375,N_2251);
xnor U2710 (N_2710,N_2272,N_2496);
nand U2711 (N_2711,N_2355,N_2349);
xnor U2712 (N_2712,N_2447,N_2495);
nand U2713 (N_2713,N_2266,N_2369);
or U2714 (N_2714,N_2263,N_2496);
and U2715 (N_2715,N_2314,N_2256);
or U2716 (N_2716,N_2402,N_2298);
or U2717 (N_2717,N_2285,N_2312);
nor U2718 (N_2718,N_2382,N_2494);
nand U2719 (N_2719,N_2325,N_2403);
nor U2720 (N_2720,N_2273,N_2411);
xor U2721 (N_2721,N_2435,N_2257);
or U2722 (N_2722,N_2367,N_2495);
nand U2723 (N_2723,N_2467,N_2351);
and U2724 (N_2724,N_2286,N_2475);
xnor U2725 (N_2725,N_2283,N_2349);
or U2726 (N_2726,N_2386,N_2387);
or U2727 (N_2727,N_2415,N_2336);
nor U2728 (N_2728,N_2449,N_2396);
or U2729 (N_2729,N_2400,N_2364);
nor U2730 (N_2730,N_2374,N_2301);
nor U2731 (N_2731,N_2471,N_2469);
or U2732 (N_2732,N_2423,N_2443);
and U2733 (N_2733,N_2467,N_2492);
xor U2734 (N_2734,N_2384,N_2369);
or U2735 (N_2735,N_2493,N_2270);
or U2736 (N_2736,N_2382,N_2443);
nor U2737 (N_2737,N_2259,N_2297);
and U2738 (N_2738,N_2449,N_2318);
or U2739 (N_2739,N_2354,N_2415);
nand U2740 (N_2740,N_2329,N_2337);
nand U2741 (N_2741,N_2323,N_2320);
nand U2742 (N_2742,N_2283,N_2340);
or U2743 (N_2743,N_2449,N_2332);
xor U2744 (N_2744,N_2253,N_2402);
or U2745 (N_2745,N_2278,N_2352);
and U2746 (N_2746,N_2494,N_2489);
xor U2747 (N_2747,N_2321,N_2263);
nor U2748 (N_2748,N_2497,N_2367);
nand U2749 (N_2749,N_2477,N_2441);
nand U2750 (N_2750,N_2735,N_2606);
nor U2751 (N_2751,N_2696,N_2547);
and U2752 (N_2752,N_2635,N_2717);
nor U2753 (N_2753,N_2500,N_2625);
nand U2754 (N_2754,N_2709,N_2670);
nor U2755 (N_2755,N_2680,N_2706);
xnor U2756 (N_2756,N_2702,N_2745);
xor U2757 (N_2757,N_2668,N_2535);
or U2758 (N_2758,N_2640,N_2648);
nand U2759 (N_2759,N_2663,N_2510);
nand U2760 (N_2760,N_2587,N_2669);
nor U2761 (N_2761,N_2691,N_2589);
xor U2762 (N_2762,N_2519,N_2679);
nand U2763 (N_2763,N_2581,N_2624);
xor U2764 (N_2764,N_2666,N_2655);
nor U2765 (N_2765,N_2561,N_2560);
nand U2766 (N_2766,N_2749,N_2503);
and U2767 (N_2767,N_2599,N_2722);
xnor U2768 (N_2768,N_2626,N_2556);
nor U2769 (N_2769,N_2657,N_2682);
xnor U2770 (N_2770,N_2674,N_2572);
nand U2771 (N_2771,N_2737,N_2673);
or U2772 (N_2772,N_2537,N_2574);
xor U2773 (N_2773,N_2747,N_2585);
and U2774 (N_2774,N_2542,N_2645);
nor U2775 (N_2775,N_2598,N_2628);
or U2776 (N_2776,N_2681,N_2522);
or U2777 (N_2777,N_2526,N_2734);
or U2778 (N_2778,N_2569,N_2544);
nand U2779 (N_2779,N_2647,N_2531);
nand U2780 (N_2780,N_2557,N_2662);
xnor U2781 (N_2781,N_2578,N_2653);
nor U2782 (N_2782,N_2550,N_2724);
nand U2783 (N_2783,N_2512,N_2593);
nor U2784 (N_2784,N_2746,N_2584);
and U2785 (N_2785,N_2623,N_2549);
and U2786 (N_2786,N_2558,N_2573);
or U2787 (N_2787,N_2693,N_2509);
or U2788 (N_2788,N_2678,N_2592);
nand U2789 (N_2789,N_2533,N_2721);
nor U2790 (N_2790,N_2636,N_2671);
and U2791 (N_2791,N_2715,N_2646);
nand U2792 (N_2792,N_2534,N_2633);
xor U2793 (N_2793,N_2744,N_2742);
and U2794 (N_2794,N_2540,N_2553);
nor U2795 (N_2795,N_2617,N_2541);
nor U2796 (N_2796,N_2731,N_2527);
xnor U2797 (N_2797,N_2718,N_2652);
nand U2798 (N_2798,N_2729,N_2570);
nor U2799 (N_2799,N_2686,N_2667);
xnor U2800 (N_2800,N_2689,N_2575);
and U2801 (N_2801,N_2629,N_2524);
nand U2802 (N_2802,N_2588,N_2571);
or U2803 (N_2803,N_2739,N_2551);
nand U2804 (N_2804,N_2710,N_2658);
or U2805 (N_2805,N_2621,N_2523);
or U2806 (N_2806,N_2603,N_2529);
and U2807 (N_2807,N_2567,N_2504);
and U2808 (N_2808,N_2580,N_2619);
nand U2809 (N_2809,N_2583,N_2609);
xnor U2810 (N_2810,N_2711,N_2604);
nor U2811 (N_2811,N_2532,N_2695);
nand U2812 (N_2812,N_2545,N_2555);
and U2813 (N_2813,N_2659,N_2607);
nand U2814 (N_2814,N_2521,N_2597);
xnor U2815 (N_2815,N_2697,N_2700);
xor U2816 (N_2816,N_2687,N_2631);
or U2817 (N_2817,N_2602,N_2738);
xor U2818 (N_2818,N_2641,N_2639);
nor U2819 (N_2819,N_2632,N_2643);
or U2820 (N_2820,N_2586,N_2660);
or U2821 (N_2821,N_2610,N_2507);
xor U2822 (N_2822,N_2611,N_2614);
nor U2823 (N_2823,N_2634,N_2683);
nand U2824 (N_2824,N_2726,N_2528);
nand U2825 (N_2825,N_2704,N_2513);
nand U2826 (N_2826,N_2568,N_2720);
nor U2827 (N_2827,N_2741,N_2559);
xor U2828 (N_2828,N_2654,N_2501);
nor U2829 (N_2829,N_2713,N_2506);
and U2830 (N_2830,N_2705,N_2516);
nor U2831 (N_2831,N_2725,N_2590);
nand U2832 (N_2832,N_2664,N_2642);
or U2833 (N_2833,N_2656,N_2638);
nor U2834 (N_2834,N_2618,N_2591);
xor U2835 (N_2835,N_2620,N_2605);
or U2836 (N_2836,N_2615,N_2723);
nand U2837 (N_2837,N_2665,N_2736);
nand U2838 (N_2838,N_2613,N_2566);
or U2839 (N_2839,N_2719,N_2596);
xor U2840 (N_2840,N_2546,N_2685);
or U2841 (N_2841,N_2714,N_2514);
nor U2842 (N_2842,N_2577,N_2703);
xnor U2843 (N_2843,N_2672,N_2552);
nor U2844 (N_2844,N_2508,N_2743);
or U2845 (N_2845,N_2601,N_2716);
xnor U2846 (N_2846,N_2684,N_2539);
nand U2847 (N_2847,N_2576,N_2538);
nor U2848 (N_2848,N_2651,N_2690);
nand U2849 (N_2849,N_2548,N_2525);
or U2850 (N_2850,N_2694,N_2728);
nor U2851 (N_2851,N_2650,N_2612);
nor U2852 (N_2852,N_2565,N_2707);
nand U2853 (N_2853,N_2732,N_2644);
and U2854 (N_2854,N_2622,N_2530);
xor U2855 (N_2855,N_2733,N_2701);
xor U2856 (N_2856,N_2637,N_2536);
nor U2857 (N_2857,N_2676,N_2579);
and U2858 (N_2858,N_2727,N_2708);
and U2859 (N_2859,N_2630,N_2517);
and U2860 (N_2860,N_2594,N_2740);
or U2861 (N_2861,N_2692,N_2748);
and U2862 (N_2862,N_2608,N_2730);
and U2863 (N_2863,N_2505,N_2688);
nand U2864 (N_2864,N_2677,N_2518);
nor U2865 (N_2865,N_2675,N_2627);
nand U2866 (N_2866,N_2511,N_2595);
and U2867 (N_2867,N_2564,N_2554);
and U2868 (N_2868,N_2698,N_2502);
nor U2869 (N_2869,N_2562,N_2582);
or U2870 (N_2870,N_2520,N_2699);
and U2871 (N_2871,N_2543,N_2649);
nand U2872 (N_2872,N_2616,N_2515);
or U2873 (N_2873,N_2712,N_2661);
nor U2874 (N_2874,N_2563,N_2600);
nor U2875 (N_2875,N_2554,N_2613);
and U2876 (N_2876,N_2515,N_2576);
and U2877 (N_2877,N_2711,N_2609);
nor U2878 (N_2878,N_2684,N_2700);
xnor U2879 (N_2879,N_2553,N_2532);
and U2880 (N_2880,N_2697,N_2603);
nor U2881 (N_2881,N_2625,N_2605);
or U2882 (N_2882,N_2590,N_2686);
and U2883 (N_2883,N_2692,N_2689);
nand U2884 (N_2884,N_2702,N_2675);
nand U2885 (N_2885,N_2589,N_2650);
nand U2886 (N_2886,N_2628,N_2518);
xor U2887 (N_2887,N_2571,N_2627);
or U2888 (N_2888,N_2524,N_2699);
xor U2889 (N_2889,N_2707,N_2627);
and U2890 (N_2890,N_2687,N_2664);
or U2891 (N_2891,N_2623,N_2724);
or U2892 (N_2892,N_2679,N_2527);
nand U2893 (N_2893,N_2622,N_2510);
and U2894 (N_2894,N_2540,N_2657);
xnor U2895 (N_2895,N_2567,N_2712);
xor U2896 (N_2896,N_2619,N_2626);
or U2897 (N_2897,N_2545,N_2599);
nor U2898 (N_2898,N_2609,N_2658);
nor U2899 (N_2899,N_2674,N_2543);
xor U2900 (N_2900,N_2591,N_2518);
nand U2901 (N_2901,N_2612,N_2698);
and U2902 (N_2902,N_2638,N_2685);
nand U2903 (N_2903,N_2559,N_2650);
or U2904 (N_2904,N_2667,N_2532);
nand U2905 (N_2905,N_2691,N_2709);
nand U2906 (N_2906,N_2542,N_2667);
and U2907 (N_2907,N_2668,N_2619);
and U2908 (N_2908,N_2672,N_2700);
nor U2909 (N_2909,N_2748,N_2614);
and U2910 (N_2910,N_2553,N_2637);
or U2911 (N_2911,N_2739,N_2545);
nor U2912 (N_2912,N_2734,N_2611);
nor U2913 (N_2913,N_2670,N_2701);
and U2914 (N_2914,N_2622,N_2543);
xnor U2915 (N_2915,N_2568,N_2599);
and U2916 (N_2916,N_2674,N_2584);
or U2917 (N_2917,N_2543,N_2732);
nor U2918 (N_2918,N_2716,N_2532);
nor U2919 (N_2919,N_2653,N_2734);
or U2920 (N_2920,N_2502,N_2598);
xor U2921 (N_2921,N_2605,N_2589);
xor U2922 (N_2922,N_2733,N_2705);
or U2923 (N_2923,N_2648,N_2573);
and U2924 (N_2924,N_2722,N_2564);
nor U2925 (N_2925,N_2598,N_2541);
nand U2926 (N_2926,N_2522,N_2636);
or U2927 (N_2927,N_2616,N_2632);
or U2928 (N_2928,N_2538,N_2670);
and U2929 (N_2929,N_2579,N_2508);
nand U2930 (N_2930,N_2667,N_2643);
nor U2931 (N_2931,N_2748,N_2642);
and U2932 (N_2932,N_2610,N_2590);
or U2933 (N_2933,N_2647,N_2525);
nand U2934 (N_2934,N_2739,N_2690);
nor U2935 (N_2935,N_2583,N_2530);
and U2936 (N_2936,N_2675,N_2648);
or U2937 (N_2937,N_2588,N_2569);
and U2938 (N_2938,N_2692,N_2664);
xnor U2939 (N_2939,N_2625,N_2676);
nor U2940 (N_2940,N_2545,N_2699);
and U2941 (N_2941,N_2599,N_2584);
nor U2942 (N_2942,N_2580,N_2552);
xnor U2943 (N_2943,N_2664,N_2576);
nand U2944 (N_2944,N_2579,N_2636);
nor U2945 (N_2945,N_2568,N_2575);
or U2946 (N_2946,N_2588,N_2511);
xnor U2947 (N_2947,N_2618,N_2585);
and U2948 (N_2948,N_2649,N_2555);
xnor U2949 (N_2949,N_2726,N_2650);
nor U2950 (N_2950,N_2509,N_2616);
nand U2951 (N_2951,N_2621,N_2677);
nand U2952 (N_2952,N_2567,N_2609);
nor U2953 (N_2953,N_2603,N_2594);
or U2954 (N_2954,N_2635,N_2718);
xnor U2955 (N_2955,N_2686,N_2735);
nand U2956 (N_2956,N_2576,N_2500);
and U2957 (N_2957,N_2659,N_2685);
and U2958 (N_2958,N_2728,N_2708);
nand U2959 (N_2959,N_2705,N_2680);
or U2960 (N_2960,N_2577,N_2628);
nor U2961 (N_2961,N_2580,N_2616);
nor U2962 (N_2962,N_2626,N_2560);
nand U2963 (N_2963,N_2531,N_2545);
nor U2964 (N_2964,N_2503,N_2679);
nor U2965 (N_2965,N_2584,N_2724);
or U2966 (N_2966,N_2688,N_2503);
xnor U2967 (N_2967,N_2613,N_2672);
or U2968 (N_2968,N_2535,N_2677);
xor U2969 (N_2969,N_2608,N_2745);
and U2970 (N_2970,N_2735,N_2592);
and U2971 (N_2971,N_2558,N_2749);
and U2972 (N_2972,N_2742,N_2723);
nor U2973 (N_2973,N_2643,N_2700);
and U2974 (N_2974,N_2563,N_2547);
and U2975 (N_2975,N_2621,N_2617);
and U2976 (N_2976,N_2672,N_2679);
or U2977 (N_2977,N_2503,N_2528);
xnor U2978 (N_2978,N_2520,N_2713);
or U2979 (N_2979,N_2743,N_2542);
nor U2980 (N_2980,N_2548,N_2524);
nor U2981 (N_2981,N_2579,N_2537);
and U2982 (N_2982,N_2655,N_2615);
nand U2983 (N_2983,N_2635,N_2533);
xnor U2984 (N_2984,N_2704,N_2601);
nor U2985 (N_2985,N_2577,N_2606);
xnor U2986 (N_2986,N_2508,N_2514);
nor U2987 (N_2987,N_2543,N_2688);
xnor U2988 (N_2988,N_2704,N_2694);
xnor U2989 (N_2989,N_2611,N_2657);
nand U2990 (N_2990,N_2518,N_2740);
nor U2991 (N_2991,N_2589,N_2659);
xnor U2992 (N_2992,N_2687,N_2690);
and U2993 (N_2993,N_2569,N_2584);
or U2994 (N_2994,N_2724,N_2632);
nor U2995 (N_2995,N_2674,N_2735);
nor U2996 (N_2996,N_2696,N_2530);
nor U2997 (N_2997,N_2594,N_2621);
and U2998 (N_2998,N_2636,N_2525);
xnor U2999 (N_2999,N_2745,N_2616);
nand U3000 (N_3000,N_2816,N_2853);
nor U3001 (N_3001,N_2989,N_2900);
nor U3002 (N_3002,N_2895,N_2946);
nor U3003 (N_3003,N_2997,N_2775);
or U3004 (N_3004,N_2805,N_2920);
xnor U3005 (N_3005,N_2792,N_2758);
nor U3006 (N_3006,N_2810,N_2784);
xnor U3007 (N_3007,N_2926,N_2832);
nor U3008 (N_3008,N_2872,N_2907);
or U3009 (N_3009,N_2849,N_2873);
nor U3010 (N_3010,N_2906,N_2923);
xor U3011 (N_3011,N_2899,N_2870);
or U3012 (N_3012,N_2842,N_2803);
nor U3013 (N_3013,N_2931,N_2839);
nor U3014 (N_3014,N_2903,N_2773);
or U3015 (N_3015,N_2761,N_2878);
nor U3016 (N_3016,N_2894,N_2859);
and U3017 (N_3017,N_2986,N_2861);
nand U3018 (N_3018,N_2765,N_2959);
or U3019 (N_3019,N_2774,N_2974);
nor U3020 (N_3020,N_2979,N_2807);
nor U3021 (N_3021,N_2957,N_2898);
nor U3022 (N_3022,N_2996,N_2954);
and U3023 (N_3023,N_2818,N_2821);
nor U3024 (N_3024,N_2967,N_2794);
xor U3025 (N_3025,N_2965,N_2752);
nand U3026 (N_3026,N_2831,N_2790);
nor U3027 (N_3027,N_2828,N_2953);
nor U3028 (N_3028,N_2940,N_2933);
or U3029 (N_3029,N_2934,N_2779);
and U3030 (N_3030,N_2945,N_2795);
or U3031 (N_3031,N_2837,N_2801);
nand U3032 (N_3032,N_2776,N_2797);
nand U3033 (N_3033,N_2763,N_2796);
nand U3034 (N_3034,N_2958,N_2885);
xor U3035 (N_3035,N_2988,N_2834);
or U3036 (N_3036,N_2772,N_2938);
nor U3037 (N_3037,N_2982,N_2833);
nor U3038 (N_3038,N_2917,N_2830);
nor U3039 (N_3039,N_2896,N_2860);
nor U3040 (N_3040,N_2864,N_2751);
and U3041 (N_3041,N_2985,N_2890);
nand U3042 (N_3042,N_2835,N_2913);
or U3043 (N_3043,N_2983,N_2962);
and U3044 (N_3044,N_2846,N_2888);
nor U3045 (N_3045,N_2924,N_2754);
nor U3046 (N_3046,N_2882,N_2783);
or U3047 (N_3047,N_2994,N_2929);
and U3048 (N_3048,N_2777,N_2951);
or U3049 (N_3049,N_2867,N_2781);
and U3050 (N_3050,N_2762,N_2936);
or U3051 (N_3051,N_2881,N_2935);
nor U3052 (N_3052,N_2787,N_2876);
nor U3053 (N_3053,N_2961,N_2925);
nand U3054 (N_3054,N_2921,N_2866);
nand U3055 (N_3055,N_2802,N_2939);
or U3056 (N_3056,N_2757,N_2850);
and U3057 (N_3057,N_2844,N_2852);
or U3058 (N_3058,N_2785,N_2897);
xor U3059 (N_3059,N_2756,N_2914);
nand U3060 (N_3060,N_2915,N_2856);
xnor U3061 (N_3061,N_2991,N_2995);
or U3062 (N_3062,N_2868,N_2877);
and U3063 (N_3063,N_2799,N_2966);
and U3064 (N_3064,N_2909,N_2874);
xnor U3065 (N_3065,N_2884,N_2791);
and U3066 (N_3066,N_2817,N_2952);
nand U3067 (N_3067,N_2944,N_2960);
xor U3068 (N_3068,N_2788,N_2889);
nor U3069 (N_3069,N_2863,N_2971);
xnor U3070 (N_3070,N_2911,N_2869);
and U3071 (N_3071,N_2969,N_2922);
or U3072 (N_3072,N_2941,N_2822);
or U3073 (N_3073,N_2750,N_2841);
nor U3074 (N_3074,N_2887,N_2968);
nand U3075 (N_3075,N_2893,N_2764);
or U3076 (N_3076,N_2919,N_2786);
or U3077 (N_3077,N_2981,N_2829);
nand U3078 (N_3078,N_2780,N_2854);
xnor U3079 (N_3079,N_2825,N_2937);
or U3080 (N_3080,N_2843,N_2800);
nand U3081 (N_3081,N_2782,N_2820);
or U3082 (N_3082,N_2767,N_2793);
or U3083 (N_3083,N_2815,N_2766);
or U3084 (N_3084,N_2977,N_2928);
and U3085 (N_3085,N_2814,N_2984);
nor U3086 (N_3086,N_2838,N_2902);
nand U3087 (N_3087,N_2824,N_2886);
and U3088 (N_3088,N_2769,N_2809);
or U3089 (N_3089,N_2949,N_2908);
xnor U3090 (N_3090,N_2845,N_2932);
nand U3091 (N_3091,N_2806,N_2813);
nor U3092 (N_3092,N_2760,N_2771);
xor U3093 (N_3093,N_2858,N_2789);
and U3094 (N_3094,N_2812,N_2865);
nor U3095 (N_3095,N_2955,N_2823);
and U3096 (N_3096,N_2836,N_2892);
nor U3097 (N_3097,N_2950,N_2862);
nor U3098 (N_3098,N_2987,N_2956);
xor U3099 (N_3099,N_2930,N_2755);
nand U3100 (N_3100,N_2847,N_2879);
nand U3101 (N_3101,N_2963,N_2904);
xnor U3102 (N_3102,N_2901,N_2918);
or U3103 (N_3103,N_2993,N_2804);
nor U3104 (N_3104,N_2851,N_2753);
xor U3105 (N_3105,N_2840,N_2770);
xnor U3106 (N_3106,N_2905,N_2916);
nand U3107 (N_3107,N_2964,N_2883);
nand U3108 (N_3108,N_2998,N_2912);
nor U3109 (N_3109,N_2947,N_2857);
or U3110 (N_3110,N_2827,N_2811);
xnor U3111 (N_3111,N_2976,N_2848);
and U3112 (N_3112,N_2819,N_2875);
xnor U3113 (N_3113,N_2871,N_2808);
nand U3114 (N_3114,N_2826,N_2759);
nand U3115 (N_3115,N_2970,N_2942);
nor U3116 (N_3116,N_2798,N_2927);
and U3117 (N_3117,N_2910,N_2948);
nor U3118 (N_3118,N_2975,N_2973);
or U3119 (N_3119,N_2980,N_2972);
and U3120 (N_3120,N_2778,N_2990);
nor U3121 (N_3121,N_2768,N_2891);
or U3122 (N_3122,N_2855,N_2999);
or U3123 (N_3123,N_2880,N_2992);
nor U3124 (N_3124,N_2943,N_2978);
and U3125 (N_3125,N_2963,N_2912);
or U3126 (N_3126,N_2834,N_2958);
and U3127 (N_3127,N_2915,N_2863);
nor U3128 (N_3128,N_2989,N_2912);
xor U3129 (N_3129,N_2997,N_2810);
or U3130 (N_3130,N_2758,N_2801);
nor U3131 (N_3131,N_2887,N_2978);
and U3132 (N_3132,N_2912,N_2806);
and U3133 (N_3133,N_2829,N_2911);
nand U3134 (N_3134,N_2970,N_2861);
or U3135 (N_3135,N_2951,N_2915);
or U3136 (N_3136,N_2956,N_2965);
or U3137 (N_3137,N_2955,N_2827);
xnor U3138 (N_3138,N_2831,N_2899);
nor U3139 (N_3139,N_2752,N_2860);
and U3140 (N_3140,N_2978,N_2966);
and U3141 (N_3141,N_2847,N_2903);
nor U3142 (N_3142,N_2967,N_2946);
or U3143 (N_3143,N_2962,N_2800);
nor U3144 (N_3144,N_2830,N_2954);
and U3145 (N_3145,N_2974,N_2924);
nor U3146 (N_3146,N_2894,N_2917);
nor U3147 (N_3147,N_2917,N_2763);
nand U3148 (N_3148,N_2954,N_2892);
nor U3149 (N_3149,N_2801,N_2779);
and U3150 (N_3150,N_2910,N_2924);
or U3151 (N_3151,N_2886,N_2841);
nor U3152 (N_3152,N_2965,N_2931);
nand U3153 (N_3153,N_2992,N_2910);
or U3154 (N_3154,N_2930,N_2810);
and U3155 (N_3155,N_2793,N_2850);
and U3156 (N_3156,N_2995,N_2938);
nor U3157 (N_3157,N_2775,N_2853);
nor U3158 (N_3158,N_2971,N_2793);
and U3159 (N_3159,N_2967,N_2792);
nor U3160 (N_3160,N_2950,N_2768);
or U3161 (N_3161,N_2800,N_2879);
nor U3162 (N_3162,N_2948,N_2896);
and U3163 (N_3163,N_2966,N_2979);
xnor U3164 (N_3164,N_2963,N_2859);
nor U3165 (N_3165,N_2811,N_2866);
xor U3166 (N_3166,N_2771,N_2862);
xnor U3167 (N_3167,N_2957,N_2788);
xor U3168 (N_3168,N_2798,N_2969);
and U3169 (N_3169,N_2909,N_2890);
nor U3170 (N_3170,N_2805,N_2775);
xor U3171 (N_3171,N_2982,N_2768);
nor U3172 (N_3172,N_2862,N_2772);
xnor U3173 (N_3173,N_2845,N_2825);
nor U3174 (N_3174,N_2833,N_2790);
and U3175 (N_3175,N_2973,N_2988);
and U3176 (N_3176,N_2791,N_2836);
and U3177 (N_3177,N_2958,N_2918);
xnor U3178 (N_3178,N_2752,N_2808);
xor U3179 (N_3179,N_2966,N_2783);
nand U3180 (N_3180,N_2898,N_2881);
and U3181 (N_3181,N_2852,N_2853);
xnor U3182 (N_3182,N_2872,N_2814);
nand U3183 (N_3183,N_2913,N_2906);
xor U3184 (N_3184,N_2983,N_2762);
nand U3185 (N_3185,N_2977,N_2850);
or U3186 (N_3186,N_2752,N_2984);
nand U3187 (N_3187,N_2761,N_2776);
nand U3188 (N_3188,N_2904,N_2790);
and U3189 (N_3189,N_2971,N_2876);
xor U3190 (N_3190,N_2768,N_2760);
and U3191 (N_3191,N_2770,N_2829);
nor U3192 (N_3192,N_2984,N_2807);
and U3193 (N_3193,N_2921,N_2797);
nand U3194 (N_3194,N_2897,N_2834);
and U3195 (N_3195,N_2984,N_2905);
or U3196 (N_3196,N_2853,N_2810);
nand U3197 (N_3197,N_2788,N_2887);
xnor U3198 (N_3198,N_2928,N_2836);
xor U3199 (N_3199,N_2927,N_2914);
nor U3200 (N_3200,N_2766,N_2871);
nor U3201 (N_3201,N_2955,N_2822);
xnor U3202 (N_3202,N_2884,N_2820);
nand U3203 (N_3203,N_2825,N_2842);
xor U3204 (N_3204,N_2967,N_2815);
or U3205 (N_3205,N_2841,N_2776);
nor U3206 (N_3206,N_2911,N_2973);
and U3207 (N_3207,N_2769,N_2885);
nor U3208 (N_3208,N_2839,N_2772);
nor U3209 (N_3209,N_2913,N_2922);
or U3210 (N_3210,N_2945,N_2819);
or U3211 (N_3211,N_2932,N_2784);
nand U3212 (N_3212,N_2774,N_2800);
nor U3213 (N_3213,N_2873,N_2764);
or U3214 (N_3214,N_2756,N_2878);
xnor U3215 (N_3215,N_2795,N_2855);
nor U3216 (N_3216,N_2798,N_2903);
nand U3217 (N_3217,N_2854,N_2775);
nor U3218 (N_3218,N_2920,N_2861);
nand U3219 (N_3219,N_2995,N_2823);
and U3220 (N_3220,N_2930,N_2947);
nand U3221 (N_3221,N_2931,N_2872);
nor U3222 (N_3222,N_2926,N_2901);
nor U3223 (N_3223,N_2804,N_2843);
or U3224 (N_3224,N_2968,N_2977);
nand U3225 (N_3225,N_2899,N_2843);
or U3226 (N_3226,N_2836,N_2886);
or U3227 (N_3227,N_2758,N_2944);
nor U3228 (N_3228,N_2983,N_2767);
nor U3229 (N_3229,N_2910,N_2868);
xnor U3230 (N_3230,N_2822,N_2843);
nand U3231 (N_3231,N_2851,N_2896);
or U3232 (N_3232,N_2953,N_2763);
or U3233 (N_3233,N_2770,N_2824);
and U3234 (N_3234,N_2911,N_2800);
or U3235 (N_3235,N_2945,N_2994);
xor U3236 (N_3236,N_2832,N_2911);
and U3237 (N_3237,N_2877,N_2784);
and U3238 (N_3238,N_2832,N_2943);
nor U3239 (N_3239,N_2934,N_2939);
or U3240 (N_3240,N_2873,N_2821);
or U3241 (N_3241,N_2982,N_2869);
nand U3242 (N_3242,N_2781,N_2844);
nand U3243 (N_3243,N_2854,N_2817);
nor U3244 (N_3244,N_2943,N_2827);
and U3245 (N_3245,N_2936,N_2905);
xor U3246 (N_3246,N_2785,N_2787);
or U3247 (N_3247,N_2872,N_2866);
xor U3248 (N_3248,N_2820,N_2920);
xnor U3249 (N_3249,N_2914,N_2903);
nor U3250 (N_3250,N_3102,N_3192);
or U3251 (N_3251,N_3071,N_3157);
and U3252 (N_3252,N_3015,N_3160);
nor U3253 (N_3253,N_3155,N_3182);
and U3254 (N_3254,N_3083,N_3154);
and U3255 (N_3255,N_3218,N_3189);
nor U3256 (N_3256,N_3111,N_3206);
or U3257 (N_3257,N_3141,N_3005);
nand U3258 (N_3258,N_3235,N_3142);
and U3259 (N_3259,N_3122,N_3038);
nand U3260 (N_3260,N_3242,N_3248);
and U3261 (N_3261,N_3205,N_3069);
and U3262 (N_3262,N_3183,N_3136);
xnor U3263 (N_3263,N_3024,N_3020);
and U3264 (N_3264,N_3135,N_3151);
xor U3265 (N_3265,N_3233,N_3029);
nand U3266 (N_3266,N_3174,N_3078);
nor U3267 (N_3267,N_3149,N_3240);
xnor U3268 (N_3268,N_3224,N_3193);
and U3269 (N_3269,N_3161,N_3067);
nor U3270 (N_3270,N_3030,N_3162);
nand U3271 (N_3271,N_3026,N_3231);
and U3272 (N_3272,N_3222,N_3041);
nor U3273 (N_3273,N_3043,N_3018);
or U3274 (N_3274,N_3239,N_3146);
xor U3275 (N_3275,N_3112,N_3166);
or U3276 (N_3276,N_3040,N_3246);
or U3277 (N_3277,N_3035,N_3191);
xor U3278 (N_3278,N_3089,N_3108);
nand U3279 (N_3279,N_3128,N_3063);
nor U3280 (N_3280,N_3120,N_3131);
xor U3281 (N_3281,N_3060,N_3055);
xor U3282 (N_3282,N_3227,N_3203);
xnor U3283 (N_3283,N_3175,N_3190);
nand U3284 (N_3284,N_3225,N_3057);
nor U3285 (N_3285,N_3168,N_3095);
xnor U3286 (N_3286,N_3051,N_3199);
and U3287 (N_3287,N_3092,N_3046);
xnor U3288 (N_3288,N_3173,N_3000);
xor U3289 (N_3289,N_3186,N_3234);
or U3290 (N_3290,N_3096,N_3232);
nor U3291 (N_3291,N_3008,N_3212);
xor U3292 (N_3292,N_3021,N_3049);
nand U3293 (N_3293,N_3167,N_3153);
xnor U3294 (N_3294,N_3197,N_3126);
and U3295 (N_3295,N_3022,N_3223);
xnor U3296 (N_3296,N_3084,N_3007);
and U3297 (N_3297,N_3130,N_3165);
xor U3298 (N_3298,N_3115,N_3123);
nor U3299 (N_3299,N_3159,N_3214);
nor U3300 (N_3300,N_3068,N_3119);
nand U3301 (N_3301,N_3170,N_3140);
and U3302 (N_3302,N_3150,N_3127);
nand U3303 (N_3303,N_3176,N_3042);
xnor U3304 (N_3304,N_3058,N_3204);
nor U3305 (N_3305,N_3187,N_3039);
and U3306 (N_3306,N_3110,N_3073);
nand U3307 (N_3307,N_3185,N_3062);
xor U3308 (N_3308,N_3098,N_3082);
or U3309 (N_3309,N_3101,N_3181);
or U3310 (N_3310,N_3006,N_3236);
nand U3311 (N_3311,N_3147,N_3072);
xor U3312 (N_3312,N_3001,N_3080);
and U3313 (N_3313,N_3249,N_3109);
or U3314 (N_3314,N_3143,N_3054);
nor U3315 (N_3315,N_3201,N_3211);
or U3316 (N_3316,N_3177,N_3025);
xor U3317 (N_3317,N_3014,N_3180);
or U3318 (N_3318,N_3243,N_3179);
nand U3319 (N_3319,N_3133,N_3106);
xnor U3320 (N_3320,N_3097,N_3134);
nand U3321 (N_3321,N_3105,N_3059);
nand U3322 (N_3322,N_3210,N_3196);
or U3323 (N_3323,N_3081,N_3230);
and U3324 (N_3324,N_3016,N_3028);
nand U3325 (N_3325,N_3076,N_3216);
nor U3326 (N_3326,N_3164,N_3103);
nand U3327 (N_3327,N_3079,N_3221);
or U3328 (N_3328,N_3152,N_3037);
xor U3329 (N_3329,N_3002,N_3163);
nand U3330 (N_3330,N_3229,N_3066);
and U3331 (N_3331,N_3156,N_3023);
nand U3332 (N_3332,N_3032,N_3100);
and U3333 (N_3333,N_3129,N_3117);
nor U3334 (N_3334,N_3172,N_3070);
or U3335 (N_3335,N_3208,N_3009);
nand U3336 (N_3336,N_3019,N_3144);
or U3337 (N_3337,N_3148,N_3226);
and U3338 (N_3338,N_3138,N_3116);
nand U3339 (N_3339,N_3031,N_3075);
nand U3340 (N_3340,N_3200,N_3033);
nand U3341 (N_3341,N_3050,N_3013);
and U3342 (N_3342,N_3132,N_3012);
or U3343 (N_3343,N_3094,N_3053);
or U3344 (N_3344,N_3184,N_3048);
or U3345 (N_3345,N_3195,N_3158);
nand U3346 (N_3346,N_3171,N_3085);
and U3347 (N_3347,N_3027,N_3064);
nand U3348 (N_3348,N_3099,N_3034);
nor U3349 (N_3349,N_3074,N_3125);
nor U3350 (N_3350,N_3217,N_3220);
and U3351 (N_3351,N_3036,N_3114);
nand U3352 (N_3352,N_3202,N_3241);
nand U3353 (N_3353,N_3086,N_3118);
nand U3354 (N_3354,N_3004,N_3245);
or U3355 (N_3355,N_3169,N_3090);
nor U3356 (N_3356,N_3137,N_3188);
and U3357 (N_3357,N_3104,N_3091);
xor U3358 (N_3358,N_3061,N_3087);
and U3359 (N_3359,N_3121,N_3065);
xor U3360 (N_3360,N_3011,N_3194);
nand U3361 (N_3361,N_3107,N_3113);
and U3362 (N_3362,N_3017,N_3056);
or U3363 (N_3363,N_3145,N_3213);
and U3364 (N_3364,N_3237,N_3124);
xor U3365 (N_3365,N_3139,N_3209);
nor U3366 (N_3366,N_3010,N_3093);
or U3367 (N_3367,N_3215,N_3003);
or U3368 (N_3368,N_3198,N_3244);
or U3369 (N_3369,N_3077,N_3047);
and U3370 (N_3370,N_3088,N_3247);
nand U3371 (N_3371,N_3207,N_3228);
and U3372 (N_3372,N_3045,N_3052);
or U3373 (N_3373,N_3238,N_3219);
xnor U3374 (N_3374,N_3044,N_3178);
and U3375 (N_3375,N_3094,N_3201);
or U3376 (N_3376,N_3120,N_3004);
and U3377 (N_3377,N_3029,N_3085);
nor U3378 (N_3378,N_3182,N_3228);
xor U3379 (N_3379,N_3161,N_3116);
nand U3380 (N_3380,N_3092,N_3008);
or U3381 (N_3381,N_3193,N_3074);
and U3382 (N_3382,N_3184,N_3237);
xor U3383 (N_3383,N_3089,N_3226);
nor U3384 (N_3384,N_3169,N_3009);
xor U3385 (N_3385,N_3021,N_3151);
nor U3386 (N_3386,N_3075,N_3198);
nor U3387 (N_3387,N_3051,N_3223);
or U3388 (N_3388,N_3186,N_3154);
nand U3389 (N_3389,N_3164,N_3149);
nand U3390 (N_3390,N_3006,N_3088);
or U3391 (N_3391,N_3065,N_3221);
xnor U3392 (N_3392,N_3016,N_3022);
or U3393 (N_3393,N_3097,N_3198);
and U3394 (N_3394,N_3089,N_3027);
nand U3395 (N_3395,N_3084,N_3155);
nand U3396 (N_3396,N_3028,N_3249);
xor U3397 (N_3397,N_3056,N_3129);
and U3398 (N_3398,N_3017,N_3239);
nor U3399 (N_3399,N_3113,N_3178);
nand U3400 (N_3400,N_3190,N_3131);
or U3401 (N_3401,N_3123,N_3053);
nand U3402 (N_3402,N_3063,N_3207);
or U3403 (N_3403,N_3215,N_3199);
xnor U3404 (N_3404,N_3120,N_3171);
or U3405 (N_3405,N_3247,N_3146);
xnor U3406 (N_3406,N_3013,N_3243);
or U3407 (N_3407,N_3072,N_3098);
and U3408 (N_3408,N_3202,N_3021);
or U3409 (N_3409,N_3104,N_3120);
nor U3410 (N_3410,N_3106,N_3239);
and U3411 (N_3411,N_3222,N_3082);
and U3412 (N_3412,N_3208,N_3162);
nand U3413 (N_3413,N_3062,N_3021);
nor U3414 (N_3414,N_3248,N_3094);
xor U3415 (N_3415,N_3235,N_3219);
nand U3416 (N_3416,N_3193,N_3114);
and U3417 (N_3417,N_3116,N_3240);
or U3418 (N_3418,N_3127,N_3241);
nor U3419 (N_3419,N_3191,N_3137);
nor U3420 (N_3420,N_3236,N_3137);
nor U3421 (N_3421,N_3228,N_3072);
and U3422 (N_3422,N_3105,N_3093);
nor U3423 (N_3423,N_3152,N_3088);
nor U3424 (N_3424,N_3138,N_3180);
xor U3425 (N_3425,N_3039,N_3007);
nor U3426 (N_3426,N_3201,N_3182);
xnor U3427 (N_3427,N_3168,N_3244);
xnor U3428 (N_3428,N_3207,N_3072);
nor U3429 (N_3429,N_3067,N_3235);
nor U3430 (N_3430,N_3193,N_3064);
and U3431 (N_3431,N_3177,N_3137);
and U3432 (N_3432,N_3058,N_3036);
nand U3433 (N_3433,N_3168,N_3059);
or U3434 (N_3434,N_3030,N_3077);
nand U3435 (N_3435,N_3245,N_3193);
nand U3436 (N_3436,N_3056,N_3176);
xnor U3437 (N_3437,N_3006,N_3193);
and U3438 (N_3438,N_3203,N_3008);
nand U3439 (N_3439,N_3185,N_3139);
and U3440 (N_3440,N_3169,N_3039);
and U3441 (N_3441,N_3192,N_3160);
nand U3442 (N_3442,N_3136,N_3021);
and U3443 (N_3443,N_3013,N_3125);
and U3444 (N_3444,N_3209,N_3117);
xnor U3445 (N_3445,N_3210,N_3071);
xnor U3446 (N_3446,N_3075,N_3135);
and U3447 (N_3447,N_3189,N_3047);
nor U3448 (N_3448,N_3009,N_3163);
nor U3449 (N_3449,N_3216,N_3030);
nor U3450 (N_3450,N_3246,N_3003);
nand U3451 (N_3451,N_3073,N_3040);
or U3452 (N_3452,N_3028,N_3166);
xor U3453 (N_3453,N_3198,N_3148);
nand U3454 (N_3454,N_3208,N_3100);
nor U3455 (N_3455,N_3000,N_3014);
xor U3456 (N_3456,N_3125,N_3174);
or U3457 (N_3457,N_3187,N_3030);
xnor U3458 (N_3458,N_3178,N_3007);
nor U3459 (N_3459,N_3099,N_3234);
or U3460 (N_3460,N_3064,N_3247);
xnor U3461 (N_3461,N_3012,N_3016);
and U3462 (N_3462,N_3053,N_3114);
nand U3463 (N_3463,N_3147,N_3218);
or U3464 (N_3464,N_3120,N_3122);
nand U3465 (N_3465,N_3091,N_3182);
or U3466 (N_3466,N_3127,N_3088);
nand U3467 (N_3467,N_3167,N_3020);
or U3468 (N_3468,N_3167,N_3083);
xnor U3469 (N_3469,N_3132,N_3003);
or U3470 (N_3470,N_3244,N_3201);
and U3471 (N_3471,N_3130,N_3081);
nand U3472 (N_3472,N_3072,N_3215);
nand U3473 (N_3473,N_3226,N_3209);
and U3474 (N_3474,N_3140,N_3032);
nand U3475 (N_3475,N_3085,N_3222);
nand U3476 (N_3476,N_3165,N_3098);
nand U3477 (N_3477,N_3232,N_3043);
and U3478 (N_3478,N_3207,N_3178);
nand U3479 (N_3479,N_3029,N_3015);
nand U3480 (N_3480,N_3062,N_3234);
nand U3481 (N_3481,N_3083,N_3113);
xnor U3482 (N_3482,N_3206,N_3197);
and U3483 (N_3483,N_3229,N_3065);
xor U3484 (N_3484,N_3134,N_3059);
xnor U3485 (N_3485,N_3028,N_3136);
nand U3486 (N_3486,N_3096,N_3091);
or U3487 (N_3487,N_3041,N_3000);
or U3488 (N_3488,N_3215,N_3034);
xor U3489 (N_3489,N_3142,N_3073);
xor U3490 (N_3490,N_3046,N_3040);
and U3491 (N_3491,N_3229,N_3115);
or U3492 (N_3492,N_3210,N_3171);
or U3493 (N_3493,N_3107,N_3130);
and U3494 (N_3494,N_3107,N_3041);
or U3495 (N_3495,N_3179,N_3022);
xnor U3496 (N_3496,N_3007,N_3041);
nor U3497 (N_3497,N_3023,N_3189);
nor U3498 (N_3498,N_3183,N_3188);
nand U3499 (N_3499,N_3125,N_3051);
xor U3500 (N_3500,N_3258,N_3420);
or U3501 (N_3501,N_3374,N_3383);
or U3502 (N_3502,N_3373,N_3405);
nor U3503 (N_3503,N_3351,N_3350);
nand U3504 (N_3504,N_3365,N_3317);
and U3505 (N_3505,N_3320,N_3397);
nor U3506 (N_3506,N_3311,N_3443);
nor U3507 (N_3507,N_3380,N_3424);
and U3508 (N_3508,N_3256,N_3461);
nand U3509 (N_3509,N_3483,N_3484);
or U3510 (N_3510,N_3411,N_3299);
nand U3511 (N_3511,N_3451,N_3328);
xor U3512 (N_3512,N_3291,N_3340);
xor U3513 (N_3513,N_3498,N_3488);
xnor U3514 (N_3514,N_3415,N_3279);
or U3515 (N_3515,N_3339,N_3416);
nand U3516 (N_3516,N_3422,N_3321);
nand U3517 (N_3517,N_3470,N_3438);
nand U3518 (N_3518,N_3252,N_3342);
nand U3519 (N_3519,N_3436,N_3277);
nand U3520 (N_3520,N_3421,N_3362);
xnor U3521 (N_3521,N_3458,N_3306);
nor U3522 (N_3522,N_3437,N_3396);
xnor U3523 (N_3523,N_3278,N_3301);
nor U3524 (N_3524,N_3469,N_3381);
nand U3525 (N_3525,N_3474,N_3480);
nor U3526 (N_3526,N_3329,N_3456);
xor U3527 (N_3527,N_3442,N_3280);
and U3528 (N_3528,N_3463,N_3444);
xor U3529 (N_3529,N_3270,N_3375);
nor U3530 (N_3530,N_3254,N_3305);
xor U3531 (N_3531,N_3445,N_3401);
or U3532 (N_3532,N_3486,N_3314);
nand U3533 (N_3533,N_3429,N_3347);
or U3534 (N_3534,N_3313,N_3287);
nor U3535 (N_3535,N_3322,N_3410);
xnor U3536 (N_3536,N_3377,N_3435);
and U3537 (N_3537,N_3260,N_3356);
nor U3538 (N_3538,N_3448,N_3478);
nand U3539 (N_3539,N_3457,N_3326);
or U3540 (N_3540,N_3330,N_3315);
nor U3541 (N_3541,N_3338,N_3433);
nor U3542 (N_3542,N_3376,N_3496);
nand U3543 (N_3543,N_3386,N_3434);
or U3544 (N_3544,N_3495,N_3465);
nor U3545 (N_3545,N_3349,N_3364);
nand U3546 (N_3546,N_3359,N_3354);
and U3547 (N_3547,N_3316,N_3454);
and U3548 (N_3548,N_3450,N_3423);
nor U3549 (N_3549,N_3358,N_3263);
nor U3550 (N_3550,N_3440,N_3269);
nor U3551 (N_3551,N_3323,N_3363);
nand U3552 (N_3552,N_3335,N_3418);
nand U3553 (N_3553,N_3459,N_3259);
nor U3554 (N_3554,N_3353,N_3392);
xor U3555 (N_3555,N_3294,N_3309);
xnor U3556 (N_3556,N_3348,N_3327);
and U3557 (N_3557,N_3274,N_3334);
nor U3558 (N_3558,N_3490,N_3406);
xnor U3559 (N_3559,N_3404,N_3408);
nor U3560 (N_3560,N_3303,N_3453);
xor U3561 (N_3561,N_3345,N_3388);
or U3562 (N_3562,N_3462,N_3267);
xor U3563 (N_3563,N_3307,N_3476);
and U3564 (N_3564,N_3394,N_3355);
or U3565 (N_3565,N_3412,N_3419);
or U3566 (N_3566,N_3369,N_3302);
nand U3567 (N_3567,N_3293,N_3281);
nor U3568 (N_3568,N_3393,N_3425);
or U3569 (N_3569,N_3265,N_3288);
xnor U3570 (N_3570,N_3409,N_3471);
xor U3571 (N_3571,N_3489,N_3285);
xor U3572 (N_3572,N_3331,N_3446);
nand U3573 (N_3573,N_3266,N_3497);
nand U3574 (N_3574,N_3477,N_3325);
nor U3575 (N_3575,N_3466,N_3426);
and U3576 (N_3576,N_3282,N_3275);
and U3577 (N_3577,N_3297,N_3271);
nand U3578 (N_3578,N_3413,N_3402);
nand U3579 (N_3579,N_3475,N_3487);
nor U3580 (N_3580,N_3391,N_3439);
nor U3581 (N_3581,N_3343,N_3468);
or U3582 (N_3582,N_3398,N_3361);
xor U3583 (N_3583,N_3352,N_3414);
nand U3584 (N_3584,N_3492,N_3276);
nor U3585 (N_3585,N_3289,N_3472);
nand U3586 (N_3586,N_3455,N_3296);
xor U3587 (N_3587,N_3399,N_3253);
nor U3588 (N_3588,N_3449,N_3372);
nor U3589 (N_3589,N_3336,N_3333);
and U3590 (N_3590,N_3379,N_3264);
nand U3591 (N_3591,N_3382,N_3417);
and U3592 (N_3592,N_3344,N_3499);
or U3593 (N_3593,N_3257,N_3395);
xor U3594 (N_3594,N_3251,N_3360);
xor U3595 (N_3595,N_3272,N_3368);
or U3596 (N_3596,N_3284,N_3273);
xnor U3597 (N_3597,N_3310,N_3400);
nor U3598 (N_3598,N_3366,N_3371);
xnor U3599 (N_3599,N_3493,N_3290);
and U3600 (N_3600,N_3387,N_3268);
nor U3601 (N_3601,N_3431,N_3407);
nand U3602 (N_3602,N_3385,N_3357);
nor U3603 (N_3603,N_3286,N_3447);
and U3604 (N_3604,N_3432,N_3460);
nor U3605 (N_3605,N_3473,N_3261);
nor U3606 (N_3606,N_3295,N_3292);
nor U3607 (N_3607,N_3452,N_3491);
nor U3608 (N_3608,N_3283,N_3384);
or U3609 (N_3609,N_3250,N_3341);
nor U3610 (N_3610,N_3312,N_3485);
and U3611 (N_3611,N_3262,N_3427);
nand U3612 (N_3612,N_3255,N_3403);
and U3613 (N_3613,N_3479,N_3464);
and U3614 (N_3614,N_3298,N_3337);
xnor U3615 (N_3615,N_3494,N_3389);
and U3616 (N_3616,N_3308,N_3319);
nand U3617 (N_3617,N_3441,N_3378);
or U3618 (N_3618,N_3332,N_3324);
nand U3619 (N_3619,N_3370,N_3482);
xor U3620 (N_3620,N_3467,N_3481);
or U3621 (N_3621,N_3430,N_3318);
xnor U3622 (N_3622,N_3390,N_3428);
nor U3623 (N_3623,N_3346,N_3367);
nand U3624 (N_3624,N_3304,N_3300);
or U3625 (N_3625,N_3271,N_3387);
xnor U3626 (N_3626,N_3394,N_3485);
and U3627 (N_3627,N_3491,N_3299);
or U3628 (N_3628,N_3326,N_3483);
nand U3629 (N_3629,N_3394,N_3335);
and U3630 (N_3630,N_3439,N_3498);
and U3631 (N_3631,N_3445,N_3400);
xnor U3632 (N_3632,N_3328,N_3473);
or U3633 (N_3633,N_3340,N_3447);
xor U3634 (N_3634,N_3250,N_3467);
and U3635 (N_3635,N_3473,N_3343);
and U3636 (N_3636,N_3451,N_3426);
and U3637 (N_3637,N_3329,N_3326);
or U3638 (N_3638,N_3461,N_3298);
nand U3639 (N_3639,N_3256,N_3398);
xnor U3640 (N_3640,N_3485,N_3287);
nor U3641 (N_3641,N_3399,N_3430);
nor U3642 (N_3642,N_3383,N_3342);
and U3643 (N_3643,N_3415,N_3296);
and U3644 (N_3644,N_3337,N_3467);
and U3645 (N_3645,N_3489,N_3379);
nor U3646 (N_3646,N_3388,N_3316);
or U3647 (N_3647,N_3414,N_3323);
nand U3648 (N_3648,N_3348,N_3330);
nor U3649 (N_3649,N_3487,N_3297);
or U3650 (N_3650,N_3326,N_3461);
or U3651 (N_3651,N_3482,N_3449);
nor U3652 (N_3652,N_3400,N_3408);
xor U3653 (N_3653,N_3321,N_3427);
nand U3654 (N_3654,N_3495,N_3307);
nor U3655 (N_3655,N_3449,N_3431);
nor U3656 (N_3656,N_3395,N_3377);
or U3657 (N_3657,N_3271,N_3296);
and U3658 (N_3658,N_3370,N_3306);
and U3659 (N_3659,N_3442,N_3298);
xor U3660 (N_3660,N_3310,N_3366);
xnor U3661 (N_3661,N_3498,N_3316);
xnor U3662 (N_3662,N_3292,N_3445);
nor U3663 (N_3663,N_3287,N_3269);
xor U3664 (N_3664,N_3264,N_3448);
and U3665 (N_3665,N_3262,N_3423);
xor U3666 (N_3666,N_3272,N_3495);
and U3667 (N_3667,N_3297,N_3356);
xor U3668 (N_3668,N_3354,N_3268);
xnor U3669 (N_3669,N_3396,N_3467);
and U3670 (N_3670,N_3373,N_3287);
or U3671 (N_3671,N_3418,N_3477);
nand U3672 (N_3672,N_3304,N_3294);
nor U3673 (N_3673,N_3359,N_3337);
nand U3674 (N_3674,N_3267,N_3260);
or U3675 (N_3675,N_3356,N_3445);
nand U3676 (N_3676,N_3360,N_3475);
nand U3677 (N_3677,N_3429,N_3415);
nor U3678 (N_3678,N_3352,N_3315);
and U3679 (N_3679,N_3257,N_3408);
xnor U3680 (N_3680,N_3345,N_3423);
xnor U3681 (N_3681,N_3488,N_3445);
nand U3682 (N_3682,N_3310,N_3335);
xnor U3683 (N_3683,N_3344,N_3448);
or U3684 (N_3684,N_3304,N_3440);
or U3685 (N_3685,N_3309,N_3482);
or U3686 (N_3686,N_3351,N_3412);
nor U3687 (N_3687,N_3256,N_3462);
nand U3688 (N_3688,N_3331,N_3487);
xor U3689 (N_3689,N_3375,N_3473);
and U3690 (N_3690,N_3386,N_3307);
xnor U3691 (N_3691,N_3320,N_3499);
or U3692 (N_3692,N_3416,N_3480);
nor U3693 (N_3693,N_3446,N_3314);
or U3694 (N_3694,N_3406,N_3269);
nand U3695 (N_3695,N_3366,N_3260);
xor U3696 (N_3696,N_3424,N_3385);
nand U3697 (N_3697,N_3371,N_3454);
or U3698 (N_3698,N_3486,N_3459);
xnor U3699 (N_3699,N_3413,N_3272);
xnor U3700 (N_3700,N_3359,N_3437);
and U3701 (N_3701,N_3436,N_3265);
xnor U3702 (N_3702,N_3301,N_3431);
or U3703 (N_3703,N_3306,N_3285);
nor U3704 (N_3704,N_3272,N_3260);
xnor U3705 (N_3705,N_3414,N_3468);
nand U3706 (N_3706,N_3335,N_3318);
and U3707 (N_3707,N_3410,N_3414);
nor U3708 (N_3708,N_3448,N_3261);
nor U3709 (N_3709,N_3282,N_3369);
nand U3710 (N_3710,N_3494,N_3294);
nor U3711 (N_3711,N_3253,N_3428);
nand U3712 (N_3712,N_3445,N_3489);
xnor U3713 (N_3713,N_3413,N_3305);
nand U3714 (N_3714,N_3436,N_3332);
or U3715 (N_3715,N_3432,N_3412);
and U3716 (N_3716,N_3470,N_3411);
nand U3717 (N_3717,N_3254,N_3314);
nand U3718 (N_3718,N_3308,N_3460);
nor U3719 (N_3719,N_3267,N_3456);
and U3720 (N_3720,N_3310,N_3439);
nand U3721 (N_3721,N_3417,N_3315);
or U3722 (N_3722,N_3447,N_3417);
xnor U3723 (N_3723,N_3250,N_3447);
nor U3724 (N_3724,N_3327,N_3446);
xor U3725 (N_3725,N_3331,N_3440);
nand U3726 (N_3726,N_3294,N_3263);
nand U3727 (N_3727,N_3365,N_3489);
xnor U3728 (N_3728,N_3393,N_3330);
nor U3729 (N_3729,N_3468,N_3342);
xnor U3730 (N_3730,N_3499,N_3455);
xor U3731 (N_3731,N_3274,N_3313);
nor U3732 (N_3732,N_3497,N_3433);
nand U3733 (N_3733,N_3425,N_3385);
or U3734 (N_3734,N_3370,N_3342);
xor U3735 (N_3735,N_3367,N_3311);
nor U3736 (N_3736,N_3366,N_3309);
nand U3737 (N_3737,N_3326,N_3492);
xnor U3738 (N_3738,N_3262,N_3451);
nor U3739 (N_3739,N_3375,N_3338);
and U3740 (N_3740,N_3290,N_3477);
or U3741 (N_3741,N_3352,N_3474);
and U3742 (N_3742,N_3387,N_3287);
xor U3743 (N_3743,N_3342,N_3260);
nand U3744 (N_3744,N_3474,N_3435);
and U3745 (N_3745,N_3393,N_3381);
or U3746 (N_3746,N_3291,N_3456);
nor U3747 (N_3747,N_3273,N_3362);
nand U3748 (N_3748,N_3293,N_3344);
xnor U3749 (N_3749,N_3446,N_3389);
and U3750 (N_3750,N_3744,N_3626);
or U3751 (N_3751,N_3691,N_3531);
or U3752 (N_3752,N_3747,N_3679);
xnor U3753 (N_3753,N_3632,N_3578);
xnor U3754 (N_3754,N_3646,N_3650);
nand U3755 (N_3755,N_3611,N_3584);
nor U3756 (N_3756,N_3715,N_3535);
xor U3757 (N_3757,N_3690,N_3716);
nand U3758 (N_3758,N_3558,N_3540);
or U3759 (N_3759,N_3649,N_3731);
or U3760 (N_3760,N_3534,N_3500);
nor U3761 (N_3761,N_3682,N_3645);
or U3762 (N_3762,N_3594,N_3520);
nor U3763 (N_3763,N_3681,N_3568);
and U3764 (N_3764,N_3538,N_3669);
and U3765 (N_3765,N_3614,N_3724);
nand U3766 (N_3766,N_3709,N_3729);
nand U3767 (N_3767,N_3642,N_3551);
nor U3768 (N_3768,N_3530,N_3554);
nand U3769 (N_3769,N_3593,N_3583);
or U3770 (N_3770,N_3548,N_3563);
nand U3771 (N_3771,N_3562,N_3510);
nor U3772 (N_3772,N_3565,N_3630);
and U3773 (N_3773,N_3671,N_3670);
and U3774 (N_3774,N_3532,N_3730);
xnor U3775 (N_3775,N_3678,N_3580);
or U3776 (N_3776,N_3528,N_3739);
nor U3777 (N_3777,N_3576,N_3597);
xnor U3778 (N_3778,N_3640,N_3648);
nor U3779 (N_3779,N_3717,N_3564);
nand U3780 (N_3780,N_3543,N_3738);
nand U3781 (N_3781,N_3725,N_3522);
xor U3782 (N_3782,N_3675,N_3608);
or U3783 (N_3783,N_3695,N_3708);
xnor U3784 (N_3784,N_3634,N_3697);
nand U3785 (N_3785,N_3514,N_3566);
nor U3786 (N_3786,N_3592,N_3742);
or U3787 (N_3787,N_3736,N_3647);
nor U3788 (N_3788,N_3735,N_3589);
nor U3789 (N_3789,N_3602,N_3655);
xnor U3790 (N_3790,N_3627,N_3526);
nand U3791 (N_3791,N_3667,N_3687);
xor U3792 (N_3792,N_3605,N_3559);
nor U3793 (N_3793,N_3550,N_3711);
nor U3794 (N_3794,N_3686,N_3633);
nand U3795 (N_3795,N_3518,N_3672);
xnor U3796 (N_3796,N_3643,N_3707);
and U3797 (N_3797,N_3749,N_3572);
nor U3798 (N_3798,N_3521,N_3631);
nor U3799 (N_3799,N_3547,N_3620);
xor U3800 (N_3800,N_3657,N_3609);
or U3801 (N_3801,N_3513,N_3629);
xnor U3802 (N_3802,N_3665,N_3727);
and U3803 (N_3803,N_3516,N_3740);
and U3804 (N_3804,N_3601,N_3734);
and U3805 (N_3805,N_3636,N_3689);
nand U3806 (N_3806,N_3698,N_3737);
xnor U3807 (N_3807,N_3658,N_3660);
nand U3808 (N_3808,N_3654,N_3573);
xnor U3809 (N_3809,N_3668,N_3503);
and U3810 (N_3810,N_3666,N_3718);
nor U3811 (N_3811,N_3639,N_3577);
xnor U3812 (N_3812,N_3508,N_3635);
nand U3813 (N_3813,N_3515,N_3509);
xnor U3814 (N_3814,N_3536,N_3546);
nor U3815 (N_3815,N_3652,N_3641);
and U3816 (N_3816,N_3527,N_3603);
xnor U3817 (N_3817,N_3651,N_3502);
nor U3818 (N_3818,N_3507,N_3741);
nor U3819 (N_3819,N_3714,N_3539);
nand U3820 (N_3820,N_3524,N_3748);
or U3821 (N_3821,N_3719,N_3713);
nand U3822 (N_3822,N_3595,N_3553);
nand U3823 (N_3823,N_3541,N_3512);
or U3824 (N_3824,N_3533,N_3720);
nand U3825 (N_3825,N_3560,N_3732);
nand U3826 (N_3826,N_3506,N_3612);
nand U3827 (N_3827,N_3569,N_3517);
and U3828 (N_3828,N_3557,N_3574);
xor U3829 (N_3829,N_3680,N_3616);
nand U3830 (N_3830,N_3549,N_3607);
and U3831 (N_3831,N_3590,N_3706);
and U3832 (N_3832,N_3505,N_3542);
nand U3833 (N_3833,N_3705,N_3700);
nor U3834 (N_3834,N_3610,N_3677);
xor U3835 (N_3835,N_3617,N_3653);
nor U3836 (N_3836,N_3519,N_3674);
or U3837 (N_3837,N_3661,N_3637);
or U3838 (N_3838,N_3659,N_3663);
nand U3839 (N_3839,N_3523,N_3723);
nor U3840 (N_3840,N_3571,N_3575);
xor U3841 (N_3841,N_3644,N_3555);
nor U3842 (N_3842,N_3685,N_3693);
or U3843 (N_3843,N_3694,N_3701);
nand U3844 (N_3844,N_3544,N_3537);
and U3845 (N_3845,N_3664,N_3622);
xnor U3846 (N_3846,N_3606,N_3628);
xnor U3847 (N_3847,N_3545,N_3746);
and U3848 (N_3848,N_3704,N_3529);
xnor U3849 (N_3849,N_3623,N_3587);
nor U3850 (N_3850,N_3710,N_3501);
xnor U3851 (N_3851,N_3702,N_3656);
nor U3852 (N_3852,N_3688,N_3638);
or U3853 (N_3853,N_3621,N_3722);
or U3854 (N_3854,N_3683,N_3581);
nand U3855 (N_3855,N_3570,N_3599);
and U3856 (N_3856,N_3556,N_3721);
and U3857 (N_3857,N_3588,N_3615);
and U3858 (N_3858,N_3586,N_3745);
or U3859 (N_3859,N_3726,N_3684);
nor U3860 (N_3860,N_3703,N_3673);
nor U3861 (N_3861,N_3598,N_3525);
xor U3862 (N_3862,N_3567,N_3696);
and U3863 (N_3863,N_3728,N_3582);
xor U3864 (N_3864,N_3585,N_3579);
or U3865 (N_3865,N_3619,N_3676);
xnor U3866 (N_3866,N_3692,N_3561);
nand U3867 (N_3867,N_3733,N_3613);
nand U3868 (N_3868,N_3552,N_3504);
and U3869 (N_3869,N_3662,N_3591);
and U3870 (N_3870,N_3511,N_3604);
and U3871 (N_3871,N_3596,N_3618);
xor U3872 (N_3872,N_3600,N_3743);
xnor U3873 (N_3873,N_3625,N_3712);
xor U3874 (N_3874,N_3624,N_3699);
xor U3875 (N_3875,N_3512,N_3574);
or U3876 (N_3876,N_3534,N_3627);
or U3877 (N_3877,N_3701,N_3610);
xor U3878 (N_3878,N_3632,N_3543);
nor U3879 (N_3879,N_3628,N_3704);
or U3880 (N_3880,N_3503,N_3596);
or U3881 (N_3881,N_3579,N_3588);
nand U3882 (N_3882,N_3600,N_3702);
nor U3883 (N_3883,N_3534,N_3739);
or U3884 (N_3884,N_3652,N_3518);
nor U3885 (N_3885,N_3665,N_3658);
nand U3886 (N_3886,N_3625,N_3517);
or U3887 (N_3887,N_3710,N_3683);
nor U3888 (N_3888,N_3564,N_3735);
nand U3889 (N_3889,N_3588,N_3594);
and U3890 (N_3890,N_3692,N_3570);
and U3891 (N_3891,N_3721,N_3652);
xor U3892 (N_3892,N_3591,N_3697);
and U3893 (N_3893,N_3517,N_3614);
nor U3894 (N_3894,N_3749,N_3744);
and U3895 (N_3895,N_3619,N_3710);
xnor U3896 (N_3896,N_3726,N_3581);
nor U3897 (N_3897,N_3510,N_3656);
or U3898 (N_3898,N_3588,N_3677);
nor U3899 (N_3899,N_3551,N_3618);
nor U3900 (N_3900,N_3612,N_3746);
nor U3901 (N_3901,N_3657,N_3505);
or U3902 (N_3902,N_3709,N_3622);
xnor U3903 (N_3903,N_3718,N_3716);
nor U3904 (N_3904,N_3596,N_3646);
or U3905 (N_3905,N_3619,N_3633);
nand U3906 (N_3906,N_3593,N_3616);
nand U3907 (N_3907,N_3619,N_3540);
or U3908 (N_3908,N_3705,N_3540);
nor U3909 (N_3909,N_3731,N_3664);
xnor U3910 (N_3910,N_3696,N_3677);
or U3911 (N_3911,N_3709,N_3605);
or U3912 (N_3912,N_3676,N_3701);
xor U3913 (N_3913,N_3689,N_3627);
nand U3914 (N_3914,N_3513,N_3663);
or U3915 (N_3915,N_3688,N_3563);
and U3916 (N_3916,N_3699,N_3553);
nand U3917 (N_3917,N_3739,N_3617);
nand U3918 (N_3918,N_3672,N_3687);
xor U3919 (N_3919,N_3715,N_3613);
nand U3920 (N_3920,N_3721,N_3541);
and U3921 (N_3921,N_3554,N_3611);
or U3922 (N_3922,N_3604,N_3624);
nand U3923 (N_3923,N_3555,N_3628);
xor U3924 (N_3924,N_3558,N_3515);
or U3925 (N_3925,N_3700,N_3558);
nor U3926 (N_3926,N_3540,N_3531);
or U3927 (N_3927,N_3586,N_3660);
nor U3928 (N_3928,N_3716,N_3629);
xor U3929 (N_3929,N_3682,N_3709);
nand U3930 (N_3930,N_3611,N_3709);
xnor U3931 (N_3931,N_3701,N_3625);
xor U3932 (N_3932,N_3611,N_3632);
nand U3933 (N_3933,N_3617,N_3643);
nor U3934 (N_3934,N_3625,N_3530);
xnor U3935 (N_3935,N_3536,N_3575);
xnor U3936 (N_3936,N_3658,N_3608);
xnor U3937 (N_3937,N_3586,N_3563);
and U3938 (N_3938,N_3620,N_3690);
nor U3939 (N_3939,N_3500,N_3613);
or U3940 (N_3940,N_3528,N_3652);
xor U3941 (N_3941,N_3599,N_3502);
and U3942 (N_3942,N_3668,N_3621);
nor U3943 (N_3943,N_3675,N_3567);
xor U3944 (N_3944,N_3580,N_3598);
nand U3945 (N_3945,N_3747,N_3705);
nand U3946 (N_3946,N_3715,N_3634);
nand U3947 (N_3947,N_3602,N_3727);
xor U3948 (N_3948,N_3716,N_3722);
xnor U3949 (N_3949,N_3670,N_3532);
or U3950 (N_3950,N_3715,N_3661);
nor U3951 (N_3951,N_3651,N_3592);
and U3952 (N_3952,N_3511,N_3699);
and U3953 (N_3953,N_3689,N_3632);
and U3954 (N_3954,N_3704,N_3647);
xnor U3955 (N_3955,N_3642,N_3667);
nand U3956 (N_3956,N_3664,N_3617);
nor U3957 (N_3957,N_3690,N_3660);
nand U3958 (N_3958,N_3513,N_3745);
nor U3959 (N_3959,N_3509,N_3663);
nor U3960 (N_3960,N_3580,N_3566);
or U3961 (N_3961,N_3562,N_3600);
xor U3962 (N_3962,N_3589,N_3667);
nor U3963 (N_3963,N_3601,N_3591);
nand U3964 (N_3964,N_3746,N_3700);
xnor U3965 (N_3965,N_3607,N_3526);
or U3966 (N_3966,N_3532,N_3622);
nand U3967 (N_3967,N_3705,N_3541);
or U3968 (N_3968,N_3715,N_3592);
xor U3969 (N_3969,N_3691,N_3720);
or U3970 (N_3970,N_3547,N_3529);
nand U3971 (N_3971,N_3523,N_3641);
and U3972 (N_3972,N_3567,N_3585);
nand U3973 (N_3973,N_3706,N_3748);
xnor U3974 (N_3974,N_3706,N_3638);
nor U3975 (N_3975,N_3630,N_3689);
xnor U3976 (N_3976,N_3654,N_3538);
xor U3977 (N_3977,N_3714,N_3602);
or U3978 (N_3978,N_3573,N_3689);
and U3979 (N_3979,N_3518,N_3725);
nor U3980 (N_3980,N_3684,N_3523);
or U3981 (N_3981,N_3722,N_3685);
or U3982 (N_3982,N_3534,N_3576);
or U3983 (N_3983,N_3636,N_3719);
xnor U3984 (N_3984,N_3672,N_3554);
nor U3985 (N_3985,N_3729,N_3505);
and U3986 (N_3986,N_3726,N_3660);
nor U3987 (N_3987,N_3570,N_3730);
or U3988 (N_3988,N_3659,N_3655);
nor U3989 (N_3989,N_3518,N_3548);
xor U3990 (N_3990,N_3525,N_3736);
and U3991 (N_3991,N_3684,N_3671);
nand U3992 (N_3992,N_3577,N_3594);
and U3993 (N_3993,N_3643,N_3647);
and U3994 (N_3994,N_3726,N_3566);
and U3995 (N_3995,N_3684,N_3664);
or U3996 (N_3996,N_3708,N_3673);
nand U3997 (N_3997,N_3616,N_3518);
or U3998 (N_3998,N_3524,N_3740);
and U3999 (N_3999,N_3709,N_3510);
nand U4000 (N_4000,N_3944,N_3870);
nand U4001 (N_4001,N_3958,N_3946);
xnor U4002 (N_4002,N_3804,N_3873);
and U4003 (N_4003,N_3831,N_3939);
and U4004 (N_4004,N_3762,N_3924);
nor U4005 (N_4005,N_3895,N_3844);
xor U4006 (N_4006,N_3894,N_3927);
or U4007 (N_4007,N_3820,N_3971);
xnor U4008 (N_4008,N_3891,N_3876);
nor U4009 (N_4009,N_3918,N_3845);
and U4010 (N_4010,N_3818,N_3886);
and U4011 (N_4011,N_3902,N_3771);
and U4012 (N_4012,N_3840,N_3814);
and U4013 (N_4013,N_3772,N_3950);
nand U4014 (N_4014,N_3775,N_3853);
xor U4015 (N_4015,N_3789,N_3782);
nor U4016 (N_4016,N_3882,N_3878);
nand U4017 (N_4017,N_3833,N_3903);
and U4018 (N_4018,N_3969,N_3807);
and U4019 (N_4019,N_3995,N_3795);
nand U4020 (N_4020,N_3864,N_3994);
nor U4021 (N_4021,N_3884,N_3913);
nor U4022 (N_4022,N_3912,N_3761);
and U4023 (N_4023,N_3999,N_3955);
and U4024 (N_4024,N_3824,N_3809);
xor U4025 (N_4025,N_3838,N_3869);
and U4026 (N_4026,N_3964,N_3861);
and U4027 (N_4027,N_3900,N_3921);
and U4028 (N_4028,N_3909,N_3816);
or U4029 (N_4029,N_3863,N_3951);
or U4030 (N_4030,N_3888,N_3952);
xor U4031 (N_4031,N_3908,N_3826);
nand U4032 (N_4032,N_3843,N_3925);
nand U4033 (N_4033,N_3957,N_3791);
xnor U4034 (N_4034,N_3779,N_3752);
xnor U4035 (N_4035,N_3874,N_3788);
or U4036 (N_4036,N_3758,N_3937);
xnor U4037 (N_4037,N_3941,N_3811);
nor U4038 (N_4038,N_3839,N_3947);
and U4039 (N_4039,N_3805,N_3897);
or U4040 (N_4040,N_3865,N_3892);
xor U4041 (N_4041,N_3926,N_3773);
nor U4042 (N_4042,N_3883,N_3760);
or U4043 (N_4043,N_3851,N_3750);
and U4044 (N_4044,N_3783,N_3956);
nand U4045 (N_4045,N_3769,N_3846);
nor U4046 (N_4046,N_3875,N_3754);
nand U4047 (N_4047,N_3922,N_3827);
nor U4048 (N_4048,N_3765,N_3972);
nand U4049 (N_4049,N_3860,N_3932);
nor U4050 (N_4050,N_3978,N_3755);
and U4051 (N_4051,N_3810,N_3756);
nor U4052 (N_4052,N_3928,N_3934);
or U4053 (N_4053,N_3935,N_3793);
xor U4054 (N_4054,N_3989,N_3829);
xor U4055 (N_4055,N_3796,N_3974);
or U4056 (N_4056,N_3830,N_3889);
and U4057 (N_4057,N_3966,N_3848);
nor U4058 (N_4058,N_3753,N_3907);
and U4059 (N_4059,N_3915,N_3806);
and U4060 (N_4060,N_3898,N_3901);
or U4061 (N_4061,N_3914,N_3817);
or U4062 (N_4062,N_3837,N_3973);
nor U4063 (N_4063,N_3786,N_3970);
nor U4064 (N_4064,N_3866,N_3929);
xor U4065 (N_4065,N_3906,N_3961);
or U4066 (N_4066,N_3792,N_3797);
nor U4067 (N_4067,N_3808,N_3868);
and U4068 (N_4068,N_3780,N_3911);
nand U4069 (N_4069,N_3859,N_3784);
nor U4070 (N_4070,N_3832,N_3962);
nor U4071 (N_4071,N_3977,N_3990);
and U4072 (N_4072,N_3953,N_3858);
nor U4073 (N_4073,N_3942,N_3813);
or U4074 (N_4074,N_3896,N_3904);
nand U4075 (N_4075,N_3800,N_3770);
or U4076 (N_4076,N_3879,N_3967);
xnor U4077 (N_4077,N_3790,N_3917);
nand U4078 (N_4078,N_3949,N_3959);
and U4079 (N_4079,N_3857,N_3986);
nor U4080 (N_4080,N_3825,N_3774);
and U4081 (N_4081,N_3976,N_3812);
and U4082 (N_4082,N_3768,N_3842);
or U4083 (N_4083,N_3777,N_3887);
xor U4084 (N_4084,N_3930,N_3751);
nor U4085 (N_4085,N_3759,N_3763);
nand U4086 (N_4086,N_3821,N_3822);
nand U4087 (N_4087,N_3938,N_3785);
xnor U4088 (N_4088,N_3867,N_3880);
nand U4089 (N_4089,N_3778,N_3787);
or U4090 (N_4090,N_3852,N_3945);
nand U4091 (N_4091,N_3931,N_3854);
and U4092 (N_4092,N_3980,N_3943);
or U4093 (N_4093,N_3998,N_3987);
and U4094 (N_4094,N_3910,N_3920);
nand U4095 (N_4095,N_3996,N_3948);
nor U4096 (N_4096,N_3871,N_3819);
xnor U4097 (N_4097,N_3899,N_3802);
and U4098 (N_4098,N_3799,N_3988);
nor U4099 (N_4099,N_3836,N_3997);
and U4100 (N_4100,N_3936,N_3835);
xor U4101 (N_4101,N_3828,N_3933);
and U4102 (N_4102,N_3834,N_3965);
and U4103 (N_4103,N_3803,N_3981);
xnor U4104 (N_4104,N_3798,N_3992);
nand U4105 (N_4105,N_3781,N_3975);
and U4106 (N_4106,N_3776,N_3757);
nand U4107 (N_4107,N_3968,N_3872);
or U4108 (N_4108,N_3985,N_3982);
nor U4109 (N_4109,N_3979,N_3923);
xnor U4110 (N_4110,N_3850,N_3963);
or U4111 (N_4111,N_3815,N_3960);
nand U4112 (N_4112,N_3940,N_3856);
xnor U4113 (N_4113,N_3954,N_3766);
or U4114 (N_4114,N_3984,N_3890);
nand U4115 (N_4115,N_3841,N_3823);
nand U4116 (N_4116,N_3893,N_3801);
nand U4117 (N_4117,N_3764,N_3847);
xnor U4118 (N_4118,N_3862,N_3916);
or U4119 (N_4119,N_3849,N_3919);
xor U4120 (N_4120,N_3877,N_3881);
and U4121 (N_4121,N_3993,N_3905);
nor U4122 (N_4122,N_3885,N_3855);
or U4123 (N_4123,N_3991,N_3767);
nor U4124 (N_4124,N_3983,N_3794);
or U4125 (N_4125,N_3767,N_3896);
nand U4126 (N_4126,N_3875,N_3838);
or U4127 (N_4127,N_3903,N_3993);
or U4128 (N_4128,N_3794,N_3896);
nand U4129 (N_4129,N_3903,N_3870);
xnor U4130 (N_4130,N_3994,N_3876);
and U4131 (N_4131,N_3790,N_3768);
or U4132 (N_4132,N_3973,N_3912);
and U4133 (N_4133,N_3912,N_3840);
and U4134 (N_4134,N_3833,N_3842);
nand U4135 (N_4135,N_3930,N_3858);
xnor U4136 (N_4136,N_3779,N_3866);
and U4137 (N_4137,N_3876,N_3809);
nor U4138 (N_4138,N_3760,N_3859);
and U4139 (N_4139,N_3893,N_3881);
nor U4140 (N_4140,N_3751,N_3898);
nand U4141 (N_4141,N_3884,N_3843);
or U4142 (N_4142,N_3974,N_3868);
nand U4143 (N_4143,N_3750,N_3862);
nor U4144 (N_4144,N_3930,N_3818);
and U4145 (N_4145,N_3873,N_3941);
or U4146 (N_4146,N_3774,N_3757);
or U4147 (N_4147,N_3940,N_3764);
nand U4148 (N_4148,N_3812,N_3960);
xnor U4149 (N_4149,N_3987,N_3932);
or U4150 (N_4150,N_3773,N_3820);
or U4151 (N_4151,N_3925,N_3770);
nor U4152 (N_4152,N_3784,N_3770);
or U4153 (N_4153,N_3913,N_3987);
nor U4154 (N_4154,N_3968,N_3990);
nand U4155 (N_4155,N_3912,N_3978);
or U4156 (N_4156,N_3881,N_3820);
nor U4157 (N_4157,N_3864,N_3813);
xor U4158 (N_4158,N_3953,N_3867);
nor U4159 (N_4159,N_3982,N_3954);
nor U4160 (N_4160,N_3958,N_3862);
or U4161 (N_4161,N_3922,N_3858);
xor U4162 (N_4162,N_3940,N_3914);
xnor U4163 (N_4163,N_3941,N_3904);
xnor U4164 (N_4164,N_3805,N_3823);
and U4165 (N_4165,N_3811,N_3977);
or U4166 (N_4166,N_3899,N_3932);
xor U4167 (N_4167,N_3888,N_3795);
nor U4168 (N_4168,N_3978,N_3990);
xor U4169 (N_4169,N_3815,N_3798);
xor U4170 (N_4170,N_3826,N_3927);
nor U4171 (N_4171,N_3785,N_3751);
or U4172 (N_4172,N_3884,N_3769);
xor U4173 (N_4173,N_3757,N_3752);
and U4174 (N_4174,N_3972,N_3911);
or U4175 (N_4175,N_3765,N_3815);
and U4176 (N_4176,N_3786,N_3768);
nand U4177 (N_4177,N_3841,N_3810);
xor U4178 (N_4178,N_3859,N_3770);
xnor U4179 (N_4179,N_3848,N_3761);
nand U4180 (N_4180,N_3850,N_3794);
or U4181 (N_4181,N_3973,N_3776);
or U4182 (N_4182,N_3847,N_3911);
or U4183 (N_4183,N_3840,N_3905);
nor U4184 (N_4184,N_3871,N_3833);
xnor U4185 (N_4185,N_3759,N_3926);
nor U4186 (N_4186,N_3806,N_3773);
nor U4187 (N_4187,N_3903,N_3992);
xnor U4188 (N_4188,N_3931,N_3807);
and U4189 (N_4189,N_3800,N_3889);
nor U4190 (N_4190,N_3943,N_3852);
or U4191 (N_4191,N_3896,N_3977);
and U4192 (N_4192,N_3855,N_3909);
nand U4193 (N_4193,N_3977,N_3830);
xnor U4194 (N_4194,N_3961,N_3797);
or U4195 (N_4195,N_3998,N_3781);
or U4196 (N_4196,N_3933,N_3837);
nand U4197 (N_4197,N_3926,N_3863);
nand U4198 (N_4198,N_3752,N_3885);
nand U4199 (N_4199,N_3842,N_3836);
xor U4200 (N_4200,N_3939,N_3934);
xor U4201 (N_4201,N_3909,N_3815);
xor U4202 (N_4202,N_3933,N_3959);
or U4203 (N_4203,N_3803,N_3807);
nand U4204 (N_4204,N_3845,N_3904);
xnor U4205 (N_4205,N_3847,N_3790);
or U4206 (N_4206,N_3791,N_3968);
xnor U4207 (N_4207,N_3841,N_3996);
nor U4208 (N_4208,N_3808,N_3864);
nor U4209 (N_4209,N_3840,N_3771);
xor U4210 (N_4210,N_3988,N_3992);
nand U4211 (N_4211,N_3764,N_3757);
nand U4212 (N_4212,N_3791,N_3830);
or U4213 (N_4213,N_3788,N_3797);
or U4214 (N_4214,N_3853,N_3951);
or U4215 (N_4215,N_3944,N_3840);
xnor U4216 (N_4216,N_3790,N_3937);
nand U4217 (N_4217,N_3892,N_3931);
xor U4218 (N_4218,N_3771,N_3839);
nor U4219 (N_4219,N_3886,N_3838);
nor U4220 (N_4220,N_3895,N_3878);
xnor U4221 (N_4221,N_3978,N_3945);
xor U4222 (N_4222,N_3790,N_3888);
and U4223 (N_4223,N_3942,N_3986);
or U4224 (N_4224,N_3892,N_3869);
xor U4225 (N_4225,N_3950,N_3829);
nand U4226 (N_4226,N_3916,N_3865);
nor U4227 (N_4227,N_3777,N_3889);
xor U4228 (N_4228,N_3958,N_3974);
or U4229 (N_4229,N_3913,N_3849);
nand U4230 (N_4230,N_3767,N_3843);
xnor U4231 (N_4231,N_3940,N_3965);
or U4232 (N_4232,N_3832,N_3952);
nor U4233 (N_4233,N_3996,N_3873);
and U4234 (N_4234,N_3840,N_3824);
nand U4235 (N_4235,N_3974,N_3756);
nand U4236 (N_4236,N_3971,N_3845);
nand U4237 (N_4237,N_3828,N_3797);
xor U4238 (N_4238,N_3768,N_3801);
and U4239 (N_4239,N_3942,N_3885);
or U4240 (N_4240,N_3765,N_3839);
nor U4241 (N_4241,N_3793,N_3917);
or U4242 (N_4242,N_3974,N_3776);
or U4243 (N_4243,N_3880,N_3946);
and U4244 (N_4244,N_3794,N_3829);
nor U4245 (N_4245,N_3966,N_3866);
or U4246 (N_4246,N_3841,N_3974);
nor U4247 (N_4247,N_3965,N_3933);
xor U4248 (N_4248,N_3788,N_3976);
xor U4249 (N_4249,N_3944,N_3777);
xor U4250 (N_4250,N_4234,N_4039);
xor U4251 (N_4251,N_4081,N_4242);
or U4252 (N_4252,N_4046,N_4137);
nor U4253 (N_4253,N_4052,N_4105);
or U4254 (N_4254,N_4027,N_4021);
or U4255 (N_4255,N_4016,N_4131);
xor U4256 (N_4256,N_4152,N_4116);
and U4257 (N_4257,N_4043,N_4031);
xor U4258 (N_4258,N_4051,N_4214);
and U4259 (N_4259,N_4066,N_4202);
xnor U4260 (N_4260,N_4068,N_4171);
nand U4261 (N_4261,N_4036,N_4084);
nand U4262 (N_4262,N_4118,N_4246);
and U4263 (N_4263,N_4080,N_4102);
nand U4264 (N_4264,N_4247,N_4008);
nand U4265 (N_4265,N_4147,N_4101);
or U4266 (N_4266,N_4162,N_4187);
xnor U4267 (N_4267,N_4138,N_4153);
nand U4268 (N_4268,N_4075,N_4204);
and U4269 (N_4269,N_4061,N_4127);
or U4270 (N_4270,N_4073,N_4164);
xnor U4271 (N_4271,N_4042,N_4109);
xor U4272 (N_4272,N_4169,N_4132);
or U4273 (N_4273,N_4064,N_4041);
xnor U4274 (N_4274,N_4123,N_4212);
xor U4275 (N_4275,N_4026,N_4136);
and U4276 (N_4276,N_4158,N_4056);
nand U4277 (N_4277,N_4062,N_4044);
nor U4278 (N_4278,N_4049,N_4078);
nor U4279 (N_4279,N_4150,N_4037);
or U4280 (N_4280,N_4085,N_4151);
or U4281 (N_4281,N_4103,N_4025);
xnor U4282 (N_4282,N_4106,N_4217);
nor U4283 (N_4283,N_4114,N_4201);
nand U4284 (N_4284,N_4122,N_4054);
xnor U4285 (N_4285,N_4249,N_4094);
xor U4286 (N_4286,N_4199,N_4216);
nor U4287 (N_4287,N_4172,N_4191);
xnor U4288 (N_4288,N_4226,N_4221);
xor U4289 (N_4289,N_4163,N_4227);
or U4290 (N_4290,N_4135,N_4010);
nor U4291 (N_4291,N_4072,N_4230);
nand U4292 (N_4292,N_4090,N_4190);
and U4293 (N_4293,N_4192,N_4117);
nor U4294 (N_4294,N_4086,N_4184);
or U4295 (N_4295,N_4240,N_4140);
nor U4296 (N_4296,N_4003,N_4071);
nor U4297 (N_4297,N_4166,N_4015);
and U4298 (N_4298,N_4093,N_4097);
nand U4299 (N_4299,N_4239,N_4165);
nand U4300 (N_4300,N_4023,N_4007);
and U4301 (N_4301,N_4012,N_4148);
nor U4302 (N_4302,N_4092,N_4188);
and U4303 (N_4303,N_4045,N_4218);
nand U4304 (N_4304,N_4047,N_4161);
xor U4305 (N_4305,N_4119,N_4206);
or U4306 (N_4306,N_4142,N_4124);
xnor U4307 (N_4307,N_4223,N_4149);
nand U4308 (N_4308,N_4197,N_4168);
or U4309 (N_4309,N_4112,N_4076);
xnor U4310 (N_4310,N_4180,N_4098);
nand U4311 (N_4311,N_4111,N_4213);
xnor U4312 (N_4312,N_4243,N_4175);
xnor U4313 (N_4313,N_4057,N_4013);
nand U4314 (N_4314,N_4174,N_4205);
xnor U4315 (N_4315,N_4233,N_4034);
and U4316 (N_4316,N_4079,N_4203);
or U4317 (N_4317,N_4182,N_4096);
and U4318 (N_4318,N_4110,N_4053);
or U4319 (N_4319,N_4095,N_4225);
xor U4320 (N_4320,N_4228,N_4024);
nand U4321 (N_4321,N_4130,N_4077);
nor U4322 (N_4322,N_4219,N_4173);
nor U4323 (N_4323,N_4040,N_4156);
nand U4324 (N_4324,N_4198,N_4139);
nand U4325 (N_4325,N_4038,N_4006);
and U4326 (N_4326,N_4179,N_4170);
xor U4327 (N_4327,N_4238,N_4210);
and U4328 (N_4328,N_4146,N_4215);
nor U4329 (N_4329,N_4019,N_4222);
and U4330 (N_4330,N_4104,N_4209);
and U4331 (N_4331,N_4145,N_4089);
nor U4332 (N_4332,N_4108,N_4065);
or U4333 (N_4333,N_4129,N_4014);
xnor U4334 (N_4334,N_4196,N_4121);
xnor U4335 (N_4335,N_4126,N_4004);
and U4336 (N_4336,N_4082,N_4113);
xor U4337 (N_4337,N_4176,N_4028);
nor U4338 (N_4338,N_4100,N_4177);
nor U4339 (N_4339,N_4193,N_4125);
nand U4340 (N_4340,N_4241,N_4059);
nand U4341 (N_4341,N_4224,N_4185);
nand U4342 (N_4342,N_4133,N_4211);
nand U4343 (N_4343,N_4134,N_4115);
and U4344 (N_4344,N_4181,N_4144);
nor U4345 (N_4345,N_4002,N_4245);
or U4346 (N_4346,N_4033,N_4030);
and U4347 (N_4347,N_4237,N_4020);
nand U4348 (N_4348,N_4159,N_4074);
nor U4349 (N_4349,N_4099,N_4154);
and U4350 (N_4350,N_4000,N_4005);
nand U4351 (N_4351,N_4069,N_4220);
and U4352 (N_4352,N_4178,N_4060);
or U4353 (N_4353,N_4141,N_4029);
nor U4354 (N_4354,N_4001,N_4231);
nand U4355 (N_4355,N_4194,N_4058);
xor U4356 (N_4356,N_4070,N_4107);
nor U4357 (N_4357,N_4189,N_4088);
nand U4358 (N_4358,N_4050,N_4244);
or U4359 (N_4359,N_4022,N_4183);
xnor U4360 (N_4360,N_4160,N_4120);
or U4361 (N_4361,N_4195,N_4235);
xnor U4362 (N_4362,N_4167,N_4128);
nand U4363 (N_4363,N_4248,N_4035);
or U4364 (N_4364,N_4091,N_4236);
xnor U4365 (N_4365,N_4207,N_4229);
nor U4366 (N_4366,N_4011,N_4200);
xnor U4367 (N_4367,N_4155,N_4186);
xnor U4368 (N_4368,N_4157,N_4018);
nand U4369 (N_4369,N_4232,N_4063);
nor U4370 (N_4370,N_4083,N_4067);
nand U4371 (N_4371,N_4087,N_4032);
nand U4372 (N_4372,N_4017,N_4048);
xor U4373 (N_4373,N_4208,N_4055);
nand U4374 (N_4374,N_4009,N_4143);
nand U4375 (N_4375,N_4134,N_4075);
or U4376 (N_4376,N_4115,N_4038);
nand U4377 (N_4377,N_4113,N_4167);
nand U4378 (N_4378,N_4127,N_4140);
nor U4379 (N_4379,N_4051,N_4141);
and U4380 (N_4380,N_4190,N_4155);
nor U4381 (N_4381,N_4198,N_4066);
nand U4382 (N_4382,N_4187,N_4016);
and U4383 (N_4383,N_4023,N_4058);
nor U4384 (N_4384,N_4235,N_4152);
nand U4385 (N_4385,N_4109,N_4087);
or U4386 (N_4386,N_4182,N_4106);
nand U4387 (N_4387,N_4206,N_4006);
nand U4388 (N_4388,N_4055,N_4150);
xnor U4389 (N_4389,N_4097,N_4115);
or U4390 (N_4390,N_4140,N_4026);
and U4391 (N_4391,N_4027,N_4097);
or U4392 (N_4392,N_4012,N_4084);
nand U4393 (N_4393,N_4038,N_4176);
or U4394 (N_4394,N_4125,N_4167);
nor U4395 (N_4395,N_4046,N_4017);
xor U4396 (N_4396,N_4143,N_4088);
and U4397 (N_4397,N_4222,N_4059);
xnor U4398 (N_4398,N_4078,N_4150);
nand U4399 (N_4399,N_4123,N_4119);
or U4400 (N_4400,N_4185,N_4242);
xnor U4401 (N_4401,N_4177,N_4245);
xor U4402 (N_4402,N_4183,N_4245);
and U4403 (N_4403,N_4081,N_4230);
xnor U4404 (N_4404,N_4002,N_4215);
nor U4405 (N_4405,N_4049,N_4212);
xor U4406 (N_4406,N_4201,N_4014);
nand U4407 (N_4407,N_4000,N_4087);
nor U4408 (N_4408,N_4003,N_4133);
and U4409 (N_4409,N_4174,N_4046);
xor U4410 (N_4410,N_4076,N_4098);
and U4411 (N_4411,N_4000,N_4019);
and U4412 (N_4412,N_4003,N_4012);
nor U4413 (N_4413,N_4043,N_4054);
and U4414 (N_4414,N_4131,N_4018);
xor U4415 (N_4415,N_4226,N_4117);
and U4416 (N_4416,N_4201,N_4140);
xor U4417 (N_4417,N_4004,N_4192);
nor U4418 (N_4418,N_4136,N_4064);
nor U4419 (N_4419,N_4135,N_4144);
xnor U4420 (N_4420,N_4135,N_4155);
or U4421 (N_4421,N_4001,N_4150);
and U4422 (N_4422,N_4183,N_4041);
xnor U4423 (N_4423,N_4179,N_4216);
nor U4424 (N_4424,N_4215,N_4206);
xnor U4425 (N_4425,N_4207,N_4180);
nor U4426 (N_4426,N_4185,N_4121);
nand U4427 (N_4427,N_4066,N_4002);
and U4428 (N_4428,N_4028,N_4063);
nor U4429 (N_4429,N_4242,N_4039);
xor U4430 (N_4430,N_4028,N_4213);
and U4431 (N_4431,N_4212,N_4000);
nor U4432 (N_4432,N_4002,N_4082);
nor U4433 (N_4433,N_4090,N_4008);
nor U4434 (N_4434,N_4122,N_4186);
or U4435 (N_4435,N_4065,N_4100);
and U4436 (N_4436,N_4172,N_4234);
and U4437 (N_4437,N_4021,N_4221);
nor U4438 (N_4438,N_4113,N_4066);
xnor U4439 (N_4439,N_4019,N_4108);
xor U4440 (N_4440,N_4104,N_4206);
or U4441 (N_4441,N_4111,N_4168);
and U4442 (N_4442,N_4037,N_4200);
nand U4443 (N_4443,N_4084,N_4144);
and U4444 (N_4444,N_4221,N_4084);
nor U4445 (N_4445,N_4016,N_4132);
nor U4446 (N_4446,N_4110,N_4094);
xor U4447 (N_4447,N_4137,N_4213);
xor U4448 (N_4448,N_4062,N_4120);
nor U4449 (N_4449,N_4247,N_4034);
or U4450 (N_4450,N_4129,N_4162);
and U4451 (N_4451,N_4182,N_4214);
nor U4452 (N_4452,N_4128,N_4160);
and U4453 (N_4453,N_4225,N_4031);
xor U4454 (N_4454,N_4211,N_4007);
and U4455 (N_4455,N_4002,N_4045);
or U4456 (N_4456,N_4097,N_4201);
nor U4457 (N_4457,N_4168,N_4138);
or U4458 (N_4458,N_4041,N_4246);
nand U4459 (N_4459,N_4137,N_4187);
and U4460 (N_4460,N_4062,N_4134);
nand U4461 (N_4461,N_4144,N_4097);
xor U4462 (N_4462,N_4226,N_4101);
and U4463 (N_4463,N_4201,N_4207);
or U4464 (N_4464,N_4028,N_4140);
and U4465 (N_4465,N_4151,N_4202);
xnor U4466 (N_4466,N_4101,N_4185);
xnor U4467 (N_4467,N_4068,N_4041);
and U4468 (N_4468,N_4012,N_4240);
nand U4469 (N_4469,N_4160,N_4130);
xnor U4470 (N_4470,N_4148,N_4139);
nand U4471 (N_4471,N_4213,N_4154);
and U4472 (N_4472,N_4124,N_4046);
nor U4473 (N_4473,N_4146,N_4209);
nand U4474 (N_4474,N_4050,N_4049);
and U4475 (N_4475,N_4135,N_4085);
xnor U4476 (N_4476,N_4125,N_4103);
nand U4477 (N_4477,N_4091,N_4023);
nand U4478 (N_4478,N_4235,N_4094);
or U4479 (N_4479,N_4065,N_4163);
or U4480 (N_4480,N_4210,N_4203);
and U4481 (N_4481,N_4063,N_4219);
xnor U4482 (N_4482,N_4109,N_4131);
nor U4483 (N_4483,N_4196,N_4069);
nor U4484 (N_4484,N_4180,N_4201);
xnor U4485 (N_4485,N_4058,N_4218);
xnor U4486 (N_4486,N_4115,N_4218);
and U4487 (N_4487,N_4134,N_4164);
nand U4488 (N_4488,N_4139,N_4049);
or U4489 (N_4489,N_4089,N_4036);
xor U4490 (N_4490,N_4243,N_4114);
xnor U4491 (N_4491,N_4062,N_4220);
xor U4492 (N_4492,N_4120,N_4048);
nor U4493 (N_4493,N_4022,N_4219);
xnor U4494 (N_4494,N_4109,N_4066);
and U4495 (N_4495,N_4013,N_4045);
nor U4496 (N_4496,N_4044,N_4055);
or U4497 (N_4497,N_4089,N_4070);
xor U4498 (N_4498,N_4179,N_4100);
and U4499 (N_4499,N_4041,N_4227);
xor U4500 (N_4500,N_4350,N_4420);
and U4501 (N_4501,N_4366,N_4330);
nor U4502 (N_4502,N_4468,N_4379);
nor U4503 (N_4503,N_4298,N_4260);
xor U4504 (N_4504,N_4336,N_4266);
nand U4505 (N_4505,N_4281,N_4452);
nor U4506 (N_4506,N_4325,N_4255);
and U4507 (N_4507,N_4317,N_4465);
xnor U4508 (N_4508,N_4416,N_4490);
nand U4509 (N_4509,N_4347,N_4444);
nor U4510 (N_4510,N_4495,N_4426);
nor U4511 (N_4511,N_4349,N_4391);
nor U4512 (N_4512,N_4436,N_4384);
and U4513 (N_4513,N_4457,N_4389);
nand U4514 (N_4514,N_4378,N_4311);
xor U4515 (N_4515,N_4337,N_4334);
nor U4516 (N_4516,N_4482,N_4252);
xor U4517 (N_4517,N_4333,N_4306);
nor U4518 (N_4518,N_4327,N_4332);
xnor U4519 (N_4519,N_4491,N_4446);
xor U4520 (N_4520,N_4447,N_4424);
or U4521 (N_4521,N_4361,N_4450);
nor U4522 (N_4522,N_4319,N_4386);
and U4523 (N_4523,N_4274,N_4323);
nor U4524 (N_4524,N_4415,N_4371);
or U4525 (N_4525,N_4394,N_4487);
or U4526 (N_4526,N_4357,N_4368);
and U4527 (N_4527,N_4278,N_4393);
or U4528 (N_4528,N_4477,N_4429);
or U4529 (N_4529,N_4380,N_4381);
or U4530 (N_4530,N_4408,N_4438);
nand U4531 (N_4531,N_4483,N_4418);
and U4532 (N_4532,N_4304,N_4251);
nor U4533 (N_4533,N_4356,N_4462);
nor U4534 (N_4534,N_4360,N_4432);
xor U4535 (N_4535,N_4470,N_4484);
or U4536 (N_4536,N_4433,N_4466);
and U4537 (N_4537,N_4414,N_4346);
xor U4538 (N_4538,N_4498,N_4390);
nor U4539 (N_4539,N_4258,N_4285);
nand U4540 (N_4540,N_4308,N_4267);
and U4541 (N_4541,N_4279,N_4343);
nand U4542 (N_4542,N_4339,N_4291);
nor U4543 (N_4543,N_4413,N_4352);
and U4544 (N_4544,N_4376,N_4388);
or U4545 (N_4545,N_4448,N_4312);
xnor U4546 (N_4546,N_4476,N_4276);
nand U4547 (N_4547,N_4454,N_4481);
nand U4548 (N_4548,N_4397,N_4303);
nor U4549 (N_4549,N_4421,N_4265);
nor U4550 (N_4550,N_4459,N_4348);
and U4551 (N_4551,N_4375,N_4427);
nand U4552 (N_4552,N_4492,N_4461);
xor U4553 (N_4553,N_4353,N_4417);
or U4554 (N_4554,N_4485,N_4321);
nand U4555 (N_4555,N_4363,N_4269);
xor U4556 (N_4556,N_4309,N_4369);
nor U4557 (N_4557,N_4342,N_4340);
nand U4558 (N_4558,N_4404,N_4439);
and U4559 (N_4559,N_4268,N_4445);
or U4560 (N_4560,N_4440,N_4316);
and U4561 (N_4561,N_4292,N_4354);
nand U4562 (N_4562,N_4314,N_4405);
and U4563 (N_4563,N_4295,N_4344);
xor U4564 (N_4564,N_4437,N_4254);
and U4565 (N_4565,N_4296,N_4443);
and U4566 (N_4566,N_4335,N_4403);
and U4567 (N_4567,N_4367,N_4358);
xor U4568 (N_4568,N_4474,N_4257);
and U4569 (N_4569,N_4401,N_4469);
xnor U4570 (N_4570,N_4402,N_4256);
and U4571 (N_4571,N_4382,N_4277);
nand U4572 (N_4572,N_4434,N_4451);
xnor U4573 (N_4573,N_4494,N_4280);
nand U4574 (N_4574,N_4262,N_4387);
xor U4575 (N_4575,N_4407,N_4430);
nand U4576 (N_4576,N_4250,N_4423);
xnor U4577 (N_4577,N_4275,N_4288);
nand U4578 (N_4578,N_4324,N_4273);
or U4579 (N_4579,N_4431,N_4253);
nand U4580 (N_4580,N_4270,N_4345);
nand U4581 (N_4581,N_4372,N_4460);
nor U4582 (N_4582,N_4489,N_4486);
or U4583 (N_4583,N_4294,N_4458);
nand U4584 (N_4584,N_4287,N_4264);
and U4585 (N_4585,N_4331,N_4315);
nand U4586 (N_4586,N_4326,N_4441);
or U4587 (N_4587,N_4374,N_4307);
and U4588 (N_4588,N_4272,N_4320);
nor U4589 (N_4589,N_4463,N_4364);
and U4590 (N_4590,N_4392,N_4456);
and U4591 (N_4591,N_4377,N_4385);
nand U4592 (N_4592,N_4467,N_4496);
or U4593 (N_4593,N_4290,N_4322);
and U4594 (N_4594,N_4411,N_4302);
xor U4595 (N_4595,N_4488,N_4355);
or U4596 (N_4596,N_4478,N_4299);
or U4597 (N_4597,N_4283,N_4455);
xor U4598 (N_4598,N_4383,N_4400);
nand U4599 (N_4599,N_4425,N_4422);
nand U4600 (N_4600,N_4373,N_4329);
nor U4601 (N_4601,N_4341,N_4442);
nor U4602 (N_4602,N_4286,N_4365);
xnor U4603 (N_4603,N_4471,N_4300);
and U4604 (N_4604,N_4435,N_4351);
or U4605 (N_4605,N_4419,N_4472);
xor U4606 (N_4606,N_4428,N_4493);
or U4607 (N_4607,N_4406,N_4362);
nand U4608 (N_4608,N_4259,N_4282);
nand U4609 (N_4609,N_4395,N_4305);
or U4610 (N_4610,N_4338,N_4464);
nor U4611 (N_4611,N_4480,N_4499);
xor U4612 (N_4612,N_4328,N_4318);
or U4613 (N_4613,N_4497,N_4398);
nor U4614 (N_4614,N_4370,N_4271);
nand U4615 (N_4615,N_4412,N_4396);
nand U4616 (N_4616,N_4293,N_4359);
xnor U4617 (N_4617,N_4261,N_4409);
nand U4618 (N_4618,N_4399,N_4313);
and U4619 (N_4619,N_4479,N_4473);
nand U4620 (N_4620,N_4301,N_4475);
nand U4621 (N_4621,N_4453,N_4263);
xor U4622 (N_4622,N_4410,N_4284);
xnor U4623 (N_4623,N_4310,N_4297);
or U4624 (N_4624,N_4289,N_4449);
and U4625 (N_4625,N_4492,N_4254);
nor U4626 (N_4626,N_4498,N_4369);
and U4627 (N_4627,N_4377,N_4430);
and U4628 (N_4628,N_4331,N_4417);
or U4629 (N_4629,N_4392,N_4291);
nor U4630 (N_4630,N_4339,N_4461);
nand U4631 (N_4631,N_4275,N_4355);
and U4632 (N_4632,N_4391,N_4347);
or U4633 (N_4633,N_4270,N_4476);
nor U4634 (N_4634,N_4433,N_4420);
nand U4635 (N_4635,N_4275,N_4498);
or U4636 (N_4636,N_4443,N_4459);
or U4637 (N_4637,N_4357,N_4477);
and U4638 (N_4638,N_4479,N_4332);
nand U4639 (N_4639,N_4349,N_4472);
nor U4640 (N_4640,N_4438,N_4416);
or U4641 (N_4641,N_4256,N_4297);
or U4642 (N_4642,N_4318,N_4447);
or U4643 (N_4643,N_4250,N_4384);
or U4644 (N_4644,N_4333,N_4283);
and U4645 (N_4645,N_4301,N_4491);
nor U4646 (N_4646,N_4385,N_4499);
nor U4647 (N_4647,N_4293,N_4356);
or U4648 (N_4648,N_4383,N_4270);
nand U4649 (N_4649,N_4374,N_4257);
xnor U4650 (N_4650,N_4448,N_4481);
or U4651 (N_4651,N_4416,N_4257);
nor U4652 (N_4652,N_4396,N_4269);
nor U4653 (N_4653,N_4271,N_4253);
nand U4654 (N_4654,N_4470,N_4458);
xnor U4655 (N_4655,N_4339,N_4332);
nor U4656 (N_4656,N_4343,N_4497);
xor U4657 (N_4657,N_4253,N_4470);
and U4658 (N_4658,N_4436,N_4403);
nor U4659 (N_4659,N_4410,N_4277);
and U4660 (N_4660,N_4270,N_4382);
and U4661 (N_4661,N_4380,N_4366);
xor U4662 (N_4662,N_4381,N_4314);
nand U4663 (N_4663,N_4351,N_4258);
and U4664 (N_4664,N_4296,N_4398);
nand U4665 (N_4665,N_4272,N_4386);
nand U4666 (N_4666,N_4318,N_4267);
or U4667 (N_4667,N_4384,N_4397);
xnor U4668 (N_4668,N_4379,N_4393);
nand U4669 (N_4669,N_4384,N_4333);
or U4670 (N_4670,N_4377,N_4305);
and U4671 (N_4671,N_4272,N_4495);
or U4672 (N_4672,N_4397,N_4321);
nand U4673 (N_4673,N_4368,N_4468);
and U4674 (N_4674,N_4374,N_4274);
nand U4675 (N_4675,N_4496,N_4493);
nand U4676 (N_4676,N_4403,N_4386);
and U4677 (N_4677,N_4409,N_4285);
xnor U4678 (N_4678,N_4469,N_4376);
nor U4679 (N_4679,N_4349,N_4345);
xor U4680 (N_4680,N_4491,N_4440);
nand U4681 (N_4681,N_4363,N_4281);
xor U4682 (N_4682,N_4370,N_4307);
and U4683 (N_4683,N_4498,N_4325);
and U4684 (N_4684,N_4286,N_4379);
xnor U4685 (N_4685,N_4390,N_4304);
or U4686 (N_4686,N_4484,N_4279);
and U4687 (N_4687,N_4330,N_4499);
nand U4688 (N_4688,N_4317,N_4441);
nand U4689 (N_4689,N_4255,N_4488);
nand U4690 (N_4690,N_4358,N_4432);
and U4691 (N_4691,N_4421,N_4274);
nor U4692 (N_4692,N_4473,N_4316);
and U4693 (N_4693,N_4440,N_4422);
and U4694 (N_4694,N_4384,N_4381);
xor U4695 (N_4695,N_4478,N_4328);
nor U4696 (N_4696,N_4395,N_4277);
or U4697 (N_4697,N_4411,N_4310);
nand U4698 (N_4698,N_4398,N_4383);
xor U4699 (N_4699,N_4317,N_4438);
nand U4700 (N_4700,N_4445,N_4490);
or U4701 (N_4701,N_4483,N_4303);
nand U4702 (N_4702,N_4258,N_4430);
nand U4703 (N_4703,N_4485,N_4438);
nand U4704 (N_4704,N_4454,N_4275);
or U4705 (N_4705,N_4335,N_4275);
xor U4706 (N_4706,N_4442,N_4453);
nand U4707 (N_4707,N_4436,N_4495);
nand U4708 (N_4708,N_4491,N_4311);
xnor U4709 (N_4709,N_4480,N_4488);
or U4710 (N_4710,N_4267,N_4382);
nand U4711 (N_4711,N_4446,N_4498);
nand U4712 (N_4712,N_4291,N_4278);
and U4713 (N_4713,N_4362,N_4432);
nor U4714 (N_4714,N_4435,N_4387);
nand U4715 (N_4715,N_4496,N_4262);
nor U4716 (N_4716,N_4282,N_4276);
nand U4717 (N_4717,N_4332,N_4371);
nor U4718 (N_4718,N_4397,N_4329);
nand U4719 (N_4719,N_4343,N_4308);
xor U4720 (N_4720,N_4451,N_4319);
or U4721 (N_4721,N_4277,N_4475);
nand U4722 (N_4722,N_4425,N_4434);
nand U4723 (N_4723,N_4301,N_4453);
xnor U4724 (N_4724,N_4335,N_4299);
xnor U4725 (N_4725,N_4438,N_4355);
nor U4726 (N_4726,N_4483,N_4426);
or U4727 (N_4727,N_4468,N_4367);
nand U4728 (N_4728,N_4272,N_4305);
xor U4729 (N_4729,N_4394,N_4483);
or U4730 (N_4730,N_4425,N_4430);
nand U4731 (N_4731,N_4304,N_4438);
or U4732 (N_4732,N_4466,N_4271);
nand U4733 (N_4733,N_4279,N_4396);
and U4734 (N_4734,N_4430,N_4332);
nand U4735 (N_4735,N_4462,N_4397);
nand U4736 (N_4736,N_4372,N_4287);
nor U4737 (N_4737,N_4344,N_4339);
xnor U4738 (N_4738,N_4359,N_4479);
or U4739 (N_4739,N_4379,N_4258);
or U4740 (N_4740,N_4286,N_4461);
nor U4741 (N_4741,N_4253,N_4489);
nand U4742 (N_4742,N_4363,N_4407);
or U4743 (N_4743,N_4254,N_4450);
or U4744 (N_4744,N_4358,N_4370);
and U4745 (N_4745,N_4418,N_4364);
nor U4746 (N_4746,N_4356,N_4461);
and U4747 (N_4747,N_4256,N_4327);
nand U4748 (N_4748,N_4297,N_4459);
or U4749 (N_4749,N_4379,N_4278);
and U4750 (N_4750,N_4621,N_4571);
or U4751 (N_4751,N_4720,N_4664);
nor U4752 (N_4752,N_4557,N_4543);
nor U4753 (N_4753,N_4548,N_4577);
and U4754 (N_4754,N_4511,N_4653);
and U4755 (N_4755,N_4615,N_4510);
xor U4756 (N_4756,N_4643,N_4675);
xor U4757 (N_4757,N_4626,N_4724);
and U4758 (N_4758,N_4561,N_4657);
nand U4759 (N_4759,N_4665,N_4678);
xor U4760 (N_4760,N_4682,N_4674);
or U4761 (N_4761,N_4722,N_4690);
xor U4762 (N_4762,N_4546,N_4651);
nor U4763 (N_4763,N_4705,N_4687);
nand U4764 (N_4764,N_4628,N_4619);
nand U4765 (N_4765,N_4707,N_4679);
nor U4766 (N_4766,N_4627,N_4594);
nand U4767 (N_4767,N_4701,N_4620);
nor U4768 (N_4768,N_4728,N_4648);
nand U4769 (N_4769,N_4566,N_4520);
xnor U4770 (N_4770,N_4662,N_4733);
nor U4771 (N_4771,N_4528,N_4578);
xor U4772 (N_4772,N_4590,N_4505);
nor U4773 (N_4773,N_4740,N_4535);
and U4774 (N_4774,N_4506,N_4656);
nand U4775 (N_4775,N_4743,N_4522);
nor U4776 (N_4776,N_4671,N_4610);
and U4777 (N_4777,N_4727,N_4599);
nor U4778 (N_4778,N_4638,N_4518);
or U4779 (N_4779,N_4581,N_4604);
or U4780 (N_4780,N_4725,N_4647);
and U4781 (N_4781,N_4541,N_4650);
or U4782 (N_4782,N_4613,N_4689);
or U4783 (N_4783,N_4715,N_4663);
nand U4784 (N_4784,N_4684,N_4532);
nor U4785 (N_4785,N_4645,N_4609);
or U4786 (N_4786,N_4642,N_4596);
nand U4787 (N_4787,N_4616,N_4508);
xnor U4788 (N_4788,N_4726,N_4691);
or U4789 (N_4789,N_4635,N_4608);
and U4790 (N_4790,N_4661,N_4529);
xnor U4791 (N_4791,N_4533,N_4730);
nor U4792 (N_4792,N_4629,N_4592);
xnor U4793 (N_4793,N_4617,N_4563);
or U4794 (N_4794,N_4560,N_4589);
nand U4795 (N_4795,N_4697,N_4696);
or U4796 (N_4796,N_4591,N_4503);
and U4797 (N_4797,N_4554,N_4540);
and U4798 (N_4798,N_4717,N_4695);
nor U4799 (N_4799,N_4637,N_4639);
xor U4800 (N_4800,N_4585,N_4747);
xnor U4801 (N_4801,N_4716,N_4685);
and U4802 (N_4802,N_4746,N_4739);
xor U4803 (N_4803,N_4744,N_4545);
or U4804 (N_4804,N_4600,N_4501);
xnor U4805 (N_4805,N_4527,N_4605);
nor U4806 (N_4806,N_4693,N_4521);
nor U4807 (N_4807,N_4700,N_4660);
xnor U4808 (N_4808,N_4672,N_4668);
and U4809 (N_4809,N_4514,N_4516);
nor U4810 (N_4810,N_4593,N_4749);
or U4811 (N_4811,N_4573,N_4513);
nand U4812 (N_4812,N_4745,N_4688);
or U4813 (N_4813,N_4658,N_4704);
xnor U4814 (N_4814,N_4703,N_4547);
nand U4815 (N_4815,N_4719,N_4748);
xnor U4816 (N_4816,N_4569,N_4711);
nand U4817 (N_4817,N_4710,N_4504);
xor U4818 (N_4818,N_4699,N_4702);
and U4819 (N_4819,N_4713,N_4595);
and U4820 (N_4820,N_4732,N_4630);
or U4821 (N_4821,N_4572,N_4666);
and U4822 (N_4822,N_4586,N_4706);
nand U4823 (N_4823,N_4574,N_4537);
nand U4824 (N_4824,N_4550,N_4526);
or U4825 (N_4825,N_4644,N_4597);
or U4826 (N_4826,N_4502,N_4525);
or U4827 (N_4827,N_4539,N_4680);
nor U4828 (N_4828,N_4735,N_4524);
xnor U4829 (N_4829,N_4623,N_4742);
nand U4830 (N_4830,N_4721,N_4555);
nor U4831 (N_4831,N_4737,N_4576);
xnor U4832 (N_4832,N_4714,N_4587);
nand U4833 (N_4833,N_4552,N_4512);
nor U4834 (N_4834,N_4530,N_4712);
and U4835 (N_4835,N_4729,N_4708);
and U4836 (N_4836,N_4632,N_4633);
nand U4837 (N_4837,N_4558,N_4567);
and U4838 (N_4838,N_4709,N_4659);
or U4839 (N_4839,N_4618,N_4575);
and U4840 (N_4840,N_4523,N_4614);
xnor U4841 (N_4841,N_4584,N_4652);
xor U4842 (N_4842,N_4683,N_4519);
or U4843 (N_4843,N_4669,N_4692);
xor U4844 (N_4844,N_4736,N_4667);
xor U4845 (N_4845,N_4741,N_4579);
xnor U4846 (N_4846,N_4636,N_4515);
or U4847 (N_4847,N_4718,N_4602);
or U4848 (N_4848,N_4698,N_4606);
and U4849 (N_4849,N_4583,N_4549);
nor U4850 (N_4850,N_4603,N_4723);
nand U4851 (N_4851,N_4676,N_4564);
and U4852 (N_4852,N_4588,N_4568);
or U4853 (N_4853,N_4565,N_4556);
xnor U4854 (N_4854,N_4598,N_4673);
and U4855 (N_4855,N_4509,N_4536);
xor U4856 (N_4856,N_4542,N_4611);
xor U4857 (N_4857,N_4500,N_4734);
xor U4858 (N_4858,N_4544,N_4607);
nor U4859 (N_4859,N_4531,N_4562);
xnor U4860 (N_4860,N_4601,N_4634);
or U4861 (N_4861,N_4570,N_4625);
or U4862 (N_4862,N_4517,N_4640);
xnor U4863 (N_4863,N_4686,N_4649);
nand U4864 (N_4864,N_4738,N_4559);
or U4865 (N_4865,N_4553,N_4681);
and U4866 (N_4866,N_4670,N_4694);
and U4867 (N_4867,N_4534,N_4507);
nand U4868 (N_4868,N_4622,N_4655);
and U4869 (N_4869,N_4646,N_4538);
xor U4870 (N_4870,N_4582,N_4631);
xor U4871 (N_4871,N_4624,N_4641);
xor U4872 (N_4872,N_4551,N_4580);
nand U4873 (N_4873,N_4612,N_4731);
nor U4874 (N_4874,N_4654,N_4677);
or U4875 (N_4875,N_4608,N_4688);
xor U4876 (N_4876,N_4725,N_4700);
xor U4877 (N_4877,N_4598,N_4744);
xnor U4878 (N_4878,N_4635,N_4715);
nand U4879 (N_4879,N_4590,N_4718);
nor U4880 (N_4880,N_4748,N_4676);
xnor U4881 (N_4881,N_4539,N_4730);
or U4882 (N_4882,N_4616,N_4525);
nand U4883 (N_4883,N_4710,N_4548);
and U4884 (N_4884,N_4689,N_4530);
xnor U4885 (N_4885,N_4594,N_4604);
and U4886 (N_4886,N_4547,N_4560);
xnor U4887 (N_4887,N_4632,N_4615);
nor U4888 (N_4888,N_4710,N_4713);
and U4889 (N_4889,N_4733,N_4702);
nor U4890 (N_4890,N_4610,N_4527);
xor U4891 (N_4891,N_4592,N_4707);
or U4892 (N_4892,N_4642,N_4649);
nand U4893 (N_4893,N_4740,N_4551);
xor U4894 (N_4894,N_4671,N_4547);
nand U4895 (N_4895,N_4743,N_4687);
nor U4896 (N_4896,N_4584,N_4575);
nand U4897 (N_4897,N_4706,N_4562);
xnor U4898 (N_4898,N_4505,N_4593);
and U4899 (N_4899,N_4730,N_4524);
nand U4900 (N_4900,N_4614,N_4647);
or U4901 (N_4901,N_4581,N_4629);
xor U4902 (N_4902,N_4584,N_4736);
or U4903 (N_4903,N_4501,N_4535);
xor U4904 (N_4904,N_4628,N_4698);
or U4905 (N_4905,N_4567,N_4576);
and U4906 (N_4906,N_4670,N_4672);
and U4907 (N_4907,N_4635,N_4678);
and U4908 (N_4908,N_4573,N_4732);
nor U4909 (N_4909,N_4514,N_4649);
nand U4910 (N_4910,N_4676,N_4710);
or U4911 (N_4911,N_4601,N_4580);
xnor U4912 (N_4912,N_4501,N_4646);
nor U4913 (N_4913,N_4722,N_4528);
nor U4914 (N_4914,N_4588,N_4650);
nand U4915 (N_4915,N_4647,N_4728);
xnor U4916 (N_4916,N_4663,N_4523);
xnor U4917 (N_4917,N_4617,N_4722);
nor U4918 (N_4918,N_4612,N_4595);
xor U4919 (N_4919,N_4591,N_4648);
nor U4920 (N_4920,N_4690,N_4607);
or U4921 (N_4921,N_4547,N_4552);
or U4922 (N_4922,N_4547,N_4621);
xor U4923 (N_4923,N_4524,N_4627);
nor U4924 (N_4924,N_4514,N_4682);
and U4925 (N_4925,N_4665,N_4587);
and U4926 (N_4926,N_4507,N_4630);
xnor U4927 (N_4927,N_4711,N_4681);
nand U4928 (N_4928,N_4642,N_4631);
xnor U4929 (N_4929,N_4640,N_4588);
nor U4930 (N_4930,N_4607,N_4571);
nor U4931 (N_4931,N_4700,N_4545);
or U4932 (N_4932,N_4747,N_4648);
or U4933 (N_4933,N_4629,N_4719);
xor U4934 (N_4934,N_4559,N_4512);
or U4935 (N_4935,N_4645,N_4707);
or U4936 (N_4936,N_4545,N_4573);
and U4937 (N_4937,N_4640,N_4697);
nor U4938 (N_4938,N_4748,N_4651);
or U4939 (N_4939,N_4591,N_4621);
nor U4940 (N_4940,N_4572,N_4662);
nor U4941 (N_4941,N_4624,N_4716);
xor U4942 (N_4942,N_4591,N_4541);
xor U4943 (N_4943,N_4618,N_4530);
xnor U4944 (N_4944,N_4657,N_4535);
or U4945 (N_4945,N_4515,N_4637);
or U4946 (N_4946,N_4618,N_4718);
xor U4947 (N_4947,N_4664,N_4622);
and U4948 (N_4948,N_4662,N_4684);
and U4949 (N_4949,N_4502,N_4503);
nor U4950 (N_4950,N_4605,N_4682);
or U4951 (N_4951,N_4676,N_4737);
xor U4952 (N_4952,N_4735,N_4513);
xor U4953 (N_4953,N_4646,N_4508);
or U4954 (N_4954,N_4573,N_4544);
and U4955 (N_4955,N_4731,N_4734);
and U4956 (N_4956,N_4725,N_4681);
xnor U4957 (N_4957,N_4728,N_4567);
xor U4958 (N_4958,N_4696,N_4702);
nand U4959 (N_4959,N_4745,N_4568);
or U4960 (N_4960,N_4536,N_4669);
or U4961 (N_4961,N_4569,N_4628);
or U4962 (N_4962,N_4703,N_4685);
nor U4963 (N_4963,N_4666,N_4667);
and U4964 (N_4964,N_4574,N_4725);
nand U4965 (N_4965,N_4736,N_4568);
nand U4966 (N_4966,N_4547,N_4726);
xor U4967 (N_4967,N_4525,N_4592);
and U4968 (N_4968,N_4585,N_4582);
or U4969 (N_4969,N_4744,N_4730);
nor U4970 (N_4970,N_4719,N_4616);
xnor U4971 (N_4971,N_4689,N_4705);
xor U4972 (N_4972,N_4665,N_4567);
nor U4973 (N_4973,N_4705,N_4640);
or U4974 (N_4974,N_4533,N_4581);
and U4975 (N_4975,N_4699,N_4634);
xnor U4976 (N_4976,N_4690,N_4515);
nor U4977 (N_4977,N_4654,N_4671);
xnor U4978 (N_4978,N_4657,N_4523);
xnor U4979 (N_4979,N_4628,N_4530);
xor U4980 (N_4980,N_4591,N_4547);
xor U4981 (N_4981,N_4576,N_4674);
and U4982 (N_4982,N_4612,N_4553);
or U4983 (N_4983,N_4731,N_4523);
nor U4984 (N_4984,N_4549,N_4680);
nand U4985 (N_4985,N_4732,N_4521);
or U4986 (N_4986,N_4515,N_4716);
or U4987 (N_4987,N_4694,N_4677);
nand U4988 (N_4988,N_4516,N_4705);
nand U4989 (N_4989,N_4733,N_4610);
and U4990 (N_4990,N_4529,N_4679);
xnor U4991 (N_4991,N_4580,N_4664);
and U4992 (N_4992,N_4569,N_4693);
nand U4993 (N_4993,N_4744,N_4674);
xnor U4994 (N_4994,N_4687,N_4500);
nor U4995 (N_4995,N_4553,N_4547);
or U4996 (N_4996,N_4549,N_4581);
or U4997 (N_4997,N_4521,N_4544);
nand U4998 (N_4998,N_4662,N_4504);
xnor U4999 (N_4999,N_4732,N_4586);
or U5000 (N_5000,N_4768,N_4775);
xor U5001 (N_5001,N_4864,N_4952);
or U5002 (N_5002,N_4854,N_4946);
xnor U5003 (N_5003,N_4836,N_4944);
or U5004 (N_5004,N_4782,N_4758);
nand U5005 (N_5005,N_4874,N_4898);
or U5006 (N_5006,N_4842,N_4839);
nor U5007 (N_5007,N_4915,N_4823);
nand U5008 (N_5008,N_4967,N_4986);
or U5009 (N_5009,N_4834,N_4963);
or U5010 (N_5010,N_4762,N_4935);
nand U5011 (N_5011,N_4752,N_4883);
nand U5012 (N_5012,N_4811,N_4943);
or U5013 (N_5013,N_4779,N_4895);
and U5014 (N_5014,N_4793,N_4896);
xnor U5015 (N_5015,N_4973,N_4994);
and U5016 (N_5016,N_4800,N_4786);
nor U5017 (N_5017,N_4788,N_4947);
nor U5018 (N_5018,N_4783,N_4919);
nor U5019 (N_5019,N_4987,N_4849);
or U5020 (N_5020,N_4795,N_4778);
and U5021 (N_5021,N_4867,N_4803);
or U5022 (N_5022,N_4798,N_4766);
and U5023 (N_5023,N_4911,N_4923);
or U5024 (N_5024,N_4859,N_4807);
nand U5025 (N_5025,N_4890,N_4908);
and U5026 (N_5026,N_4785,N_4948);
nand U5027 (N_5027,N_4759,N_4830);
nor U5028 (N_5028,N_4950,N_4875);
xor U5029 (N_5029,N_4824,N_4945);
or U5030 (N_5030,N_4953,N_4951);
xor U5031 (N_5031,N_4750,N_4767);
or U5032 (N_5032,N_4906,N_4774);
nor U5033 (N_5033,N_4940,N_4927);
nand U5034 (N_5034,N_4949,N_4843);
xor U5035 (N_5035,N_4847,N_4769);
or U5036 (N_5036,N_4932,N_4799);
or U5037 (N_5037,N_4812,N_4837);
xnor U5038 (N_5038,N_4855,N_4869);
or U5039 (N_5039,N_4876,N_4910);
or U5040 (N_5040,N_4970,N_4805);
nand U5041 (N_5041,N_4791,N_4770);
nor U5042 (N_5042,N_4790,N_4870);
xor U5043 (N_5043,N_4931,N_4872);
xor U5044 (N_5044,N_4954,N_4968);
or U5045 (N_5045,N_4825,N_4801);
xor U5046 (N_5046,N_4974,N_4865);
nand U5047 (N_5047,N_4903,N_4886);
nor U5048 (N_5048,N_4871,N_4818);
xnor U5049 (N_5049,N_4754,N_4833);
and U5050 (N_5050,N_4985,N_4936);
nand U5051 (N_5051,N_4901,N_4827);
nor U5052 (N_5052,N_4921,N_4913);
or U5053 (N_5053,N_4857,N_4815);
or U5054 (N_5054,N_4992,N_4982);
nor U5055 (N_5055,N_4980,N_4930);
and U5056 (N_5056,N_4848,N_4941);
nand U5057 (N_5057,N_4862,N_4844);
and U5058 (N_5058,N_4971,N_4972);
xor U5059 (N_5059,N_4822,N_4899);
and U5060 (N_5060,N_4764,N_4958);
nand U5061 (N_5061,N_4981,N_4991);
or U5062 (N_5062,N_4780,N_4956);
and U5063 (N_5063,N_4802,N_4888);
or U5064 (N_5064,N_4960,N_4893);
or U5065 (N_5065,N_4853,N_4897);
nor U5066 (N_5066,N_4832,N_4850);
xnor U5067 (N_5067,N_4957,N_4892);
xnor U5068 (N_5068,N_4784,N_4858);
or U5069 (N_5069,N_4751,N_4926);
xnor U5070 (N_5070,N_4878,N_4877);
or U5071 (N_5071,N_4776,N_4763);
nand U5072 (N_5072,N_4959,N_4757);
xnor U5073 (N_5073,N_4942,N_4755);
and U5074 (N_5074,N_4835,N_4765);
nor U5075 (N_5075,N_4852,N_4975);
or U5076 (N_5076,N_4846,N_4821);
nor U5077 (N_5077,N_4868,N_4756);
nor U5078 (N_5078,N_4965,N_4841);
nand U5079 (N_5079,N_4900,N_4820);
or U5080 (N_5080,N_4796,N_4797);
xor U5081 (N_5081,N_4760,N_4920);
nor U5082 (N_5082,N_4845,N_4983);
and U5083 (N_5083,N_4933,N_4912);
xor U5084 (N_5084,N_4929,N_4996);
and U5085 (N_5085,N_4977,N_4819);
nand U5086 (N_5086,N_4990,N_4840);
or U5087 (N_5087,N_4997,N_4863);
xor U5088 (N_5088,N_4884,N_4814);
or U5089 (N_5089,N_4804,N_4925);
or U5090 (N_5090,N_4998,N_4969);
and U5091 (N_5091,N_4961,N_4831);
nand U5092 (N_5092,N_4993,N_4772);
and U5093 (N_5093,N_4777,N_4794);
and U5094 (N_5094,N_4966,N_4808);
nand U5095 (N_5095,N_4909,N_4889);
nor U5096 (N_5096,N_4976,N_4904);
nand U5097 (N_5097,N_4873,N_4826);
nand U5098 (N_5098,N_4771,N_4964);
xor U5099 (N_5099,N_4894,N_4891);
or U5100 (N_5100,N_4813,N_4934);
xor U5101 (N_5101,N_4816,N_4817);
nor U5102 (N_5102,N_4881,N_4838);
xor U5103 (N_5103,N_4810,N_4999);
or U5104 (N_5104,N_4789,N_4753);
and U5105 (N_5105,N_4922,N_4984);
or U5106 (N_5106,N_4866,N_4995);
or U5107 (N_5107,N_4955,N_4828);
xnor U5108 (N_5108,N_4851,N_4887);
nor U5109 (N_5109,N_4918,N_4829);
nor U5110 (N_5110,N_4962,N_4905);
nor U5111 (N_5111,N_4924,N_4916);
or U5112 (N_5112,N_4882,N_4978);
nor U5113 (N_5113,N_4885,N_4787);
and U5114 (N_5114,N_4806,N_4917);
nor U5115 (N_5115,N_4861,N_4879);
nand U5116 (N_5116,N_4773,N_4937);
nor U5117 (N_5117,N_4792,N_4914);
nor U5118 (N_5118,N_4761,N_4928);
nor U5119 (N_5119,N_4809,N_4938);
nand U5120 (N_5120,N_4856,N_4902);
or U5121 (N_5121,N_4988,N_4781);
xor U5122 (N_5122,N_4907,N_4939);
and U5123 (N_5123,N_4979,N_4989);
nand U5124 (N_5124,N_4880,N_4860);
nor U5125 (N_5125,N_4829,N_4881);
xnor U5126 (N_5126,N_4830,N_4838);
nand U5127 (N_5127,N_4975,N_4805);
and U5128 (N_5128,N_4859,N_4858);
or U5129 (N_5129,N_4754,N_4931);
xnor U5130 (N_5130,N_4915,N_4859);
or U5131 (N_5131,N_4848,N_4939);
nor U5132 (N_5132,N_4938,N_4774);
and U5133 (N_5133,N_4758,N_4872);
xor U5134 (N_5134,N_4894,N_4954);
and U5135 (N_5135,N_4942,N_4827);
nand U5136 (N_5136,N_4764,N_4856);
nand U5137 (N_5137,N_4915,N_4901);
and U5138 (N_5138,N_4850,N_4783);
nor U5139 (N_5139,N_4875,N_4789);
xor U5140 (N_5140,N_4964,N_4873);
nand U5141 (N_5141,N_4836,N_4934);
or U5142 (N_5142,N_4983,N_4869);
or U5143 (N_5143,N_4906,N_4756);
xor U5144 (N_5144,N_4993,N_4882);
nand U5145 (N_5145,N_4998,N_4862);
and U5146 (N_5146,N_4808,N_4973);
nand U5147 (N_5147,N_4871,N_4823);
xor U5148 (N_5148,N_4765,N_4815);
and U5149 (N_5149,N_4922,N_4952);
and U5150 (N_5150,N_4869,N_4982);
and U5151 (N_5151,N_4881,N_4880);
and U5152 (N_5152,N_4883,N_4890);
nand U5153 (N_5153,N_4901,N_4929);
or U5154 (N_5154,N_4982,N_4769);
xor U5155 (N_5155,N_4844,N_4834);
xor U5156 (N_5156,N_4893,N_4913);
nand U5157 (N_5157,N_4872,N_4762);
nor U5158 (N_5158,N_4798,N_4985);
xor U5159 (N_5159,N_4912,N_4849);
xor U5160 (N_5160,N_4896,N_4940);
or U5161 (N_5161,N_4859,N_4795);
xnor U5162 (N_5162,N_4870,N_4807);
and U5163 (N_5163,N_4938,N_4799);
xor U5164 (N_5164,N_4752,N_4881);
or U5165 (N_5165,N_4853,N_4756);
nand U5166 (N_5166,N_4983,N_4837);
nor U5167 (N_5167,N_4951,N_4976);
and U5168 (N_5168,N_4752,N_4931);
xnor U5169 (N_5169,N_4927,N_4786);
nor U5170 (N_5170,N_4908,N_4811);
nor U5171 (N_5171,N_4953,N_4764);
nand U5172 (N_5172,N_4751,N_4990);
or U5173 (N_5173,N_4937,N_4751);
nor U5174 (N_5174,N_4881,N_4856);
xnor U5175 (N_5175,N_4875,N_4869);
nand U5176 (N_5176,N_4900,N_4997);
or U5177 (N_5177,N_4808,N_4977);
and U5178 (N_5178,N_4923,N_4988);
or U5179 (N_5179,N_4832,N_4978);
or U5180 (N_5180,N_4823,N_4752);
nand U5181 (N_5181,N_4750,N_4775);
or U5182 (N_5182,N_4899,N_4872);
nor U5183 (N_5183,N_4868,N_4985);
xnor U5184 (N_5184,N_4982,N_4861);
and U5185 (N_5185,N_4849,N_4755);
nand U5186 (N_5186,N_4775,N_4829);
nand U5187 (N_5187,N_4767,N_4963);
nand U5188 (N_5188,N_4924,N_4841);
xnor U5189 (N_5189,N_4774,N_4963);
nor U5190 (N_5190,N_4894,N_4871);
or U5191 (N_5191,N_4786,N_4922);
nor U5192 (N_5192,N_4981,N_4840);
and U5193 (N_5193,N_4984,N_4964);
nand U5194 (N_5194,N_4872,N_4795);
nor U5195 (N_5195,N_4870,N_4888);
or U5196 (N_5196,N_4909,N_4796);
xnor U5197 (N_5197,N_4828,N_4984);
nand U5198 (N_5198,N_4854,N_4984);
nor U5199 (N_5199,N_4793,N_4893);
xnor U5200 (N_5200,N_4904,N_4830);
and U5201 (N_5201,N_4789,N_4843);
nor U5202 (N_5202,N_4858,N_4866);
xor U5203 (N_5203,N_4929,N_4847);
xor U5204 (N_5204,N_4814,N_4833);
nand U5205 (N_5205,N_4781,N_4810);
xor U5206 (N_5206,N_4781,N_4809);
or U5207 (N_5207,N_4889,N_4911);
or U5208 (N_5208,N_4922,N_4785);
nand U5209 (N_5209,N_4998,N_4939);
and U5210 (N_5210,N_4846,N_4862);
nor U5211 (N_5211,N_4898,N_4799);
xnor U5212 (N_5212,N_4987,N_4904);
or U5213 (N_5213,N_4962,N_4864);
or U5214 (N_5214,N_4970,N_4848);
nand U5215 (N_5215,N_4900,N_4829);
nand U5216 (N_5216,N_4858,N_4843);
nand U5217 (N_5217,N_4993,N_4757);
xnor U5218 (N_5218,N_4872,N_4798);
and U5219 (N_5219,N_4866,N_4778);
and U5220 (N_5220,N_4858,N_4770);
nand U5221 (N_5221,N_4949,N_4847);
nor U5222 (N_5222,N_4875,N_4888);
nand U5223 (N_5223,N_4817,N_4896);
xor U5224 (N_5224,N_4827,N_4889);
nor U5225 (N_5225,N_4764,N_4952);
xnor U5226 (N_5226,N_4865,N_4790);
or U5227 (N_5227,N_4860,N_4870);
xnor U5228 (N_5228,N_4968,N_4752);
nand U5229 (N_5229,N_4950,N_4991);
nand U5230 (N_5230,N_4801,N_4819);
nor U5231 (N_5231,N_4857,N_4792);
or U5232 (N_5232,N_4850,N_4813);
nor U5233 (N_5233,N_4998,N_4970);
and U5234 (N_5234,N_4921,N_4934);
and U5235 (N_5235,N_4901,N_4795);
and U5236 (N_5236,N_4767,N_4978);
and U5237 (N_5237,N_4936,N_4973);
xnor U5238 (N_5238,N_4821,N_4986);
xor U5239 (N_5239,N_4981,N_4919);
nand U5240 (N_5240,N_4946,N_4791);
xor U5241 (N_5241,N_4931,N_4844);
nor U5242 (N_5242,N_4974,N_4954);
and U5243 (N_5243,N_4859,N_4957);
xor U5244 (N_5244,N_4843,N_4923);
or U5245 (N_5245,N_4921,N_4839);
or U5246 (N_5246,N_4867,N_4970);
and U5247 (N_5247,N_4888,N_4882);
nand U5248 (N_5248,N_4867,N_4922);
or U5249 (N_5249,N_4905,N_4796);
nor U5250 (N_5250,N_5051,N_5101);
and U5251 (N_5251,N_5159,N_5153);
and U5252 (N_5252,N_5194,N_5208);
nor U5253 (N_5253,N_5002,N_5138);
and U5254 (N_5254,N_5158,N_5136);
and U5255 (N_5255,N_5045,N_5007);
xor U5256 (N_5256,N_5084,N_5247);
nand U5257 (N_5257,N_5106,N_5026);
or U5258 (N_5258,N_5086,N_5048);
or U5259 (N_5259,N_5050,N_5028);
or U5260 (N_5260,N_5019,N_5183);
nor U5261 (N_5261,N_5146,N_5065);
and U5262 (N_5262,N_5118,N_5020);
nand U5263 (N_5263,N_5066,N_5054);
and U5264 (N_5264,N_5221,N_5189);
and U5265 (N_5265,N_5003,N_5175);
xor U5266 (N_5266,N_5190,N_5052);
xnor U5267 (N_5267,N_5214,N_5133);
or U5268 (N_5268,N_5041,N_5017);
xor U5269 (N_5269,N_5234,N_5244);
or U5270 (N_5270,N_5070,N_5197);
or U5271 (N_5271,N_5248,N_5218);
nor U5272 (N_5272,N_5043,N_5167);
nand U5273 (N_5273,N_5223,N_5035);
nand U5274 (N_5274,N_5130,N_5098);
xor U5275 (N_5275,N_5195,N_5077);
and U5276 (N_5276,N_5231,N_5014);
nor U5277 (N_5277,N_5230,N_5210);
and U5278 (N_5278,N_5091,N_5193);
nor U5279 (N_5279,N_5036,N_5216);
nor U5280 (N_5280,N_5022,N_5220);
or U5281 (N_5281,N_5088,N_5137);
xnor U5282 (N_5282,N_5010,N_5225);
nand U5283 (N_5283,N_5192,N_5170);
or U5284 (N_5284,N_5038,N_5173);
nor U5285 (N_5285,N_5085,N_5081);
or U5286 (N_5286,N_5152,N_5059);
and U5287 (N_5287,N_5200,N_5163);
or U5288 (N_5288,N_5129,N_5040);
or U5289 (N_5289,N_5114,N_5068);
nor U5290 (N_5290,N_5187,N_5232);
nand U5291 (N_5291,N_5061,N_5171);
and U5292 (N_5292,N_5083,N_5094);
nor U5293 (N_5293,N_5157,N_5009);
and U5294 (N_5294,N_5119,N_5069);
nand U5295 (N_5295,N_5034,N_5087);
nor U5296 (N_5296,N_5228,N_5080);
or U5297 (N_5297,N_5063,N_5249);
xor U5298 (N_5298,N_5209,N_5179);
and U5299 (N_5299,N_5053,N_5093);
nand U5300 (N_5300,N_5215,N_5046);
and U5301 (N_5301,N_5027,N_5057);
and U5302 (N_5302,N_5031,N_5226);
xnor U5303 (N_5303,N_5033,N_5030);
nor U5304 (N_5304,N_5217,N_5047);
xor U5305 (N_5305,N_5164,N_5201);
nand U5306 (N_5306,N_5161,N_5011);
or U5307 (N_5307,N_5125,N_5240);
nand U5308 (N_5308,N_5202,N_5120);
xnor U5309 (N_5309,N_5102,N_5180);
or U5310 (N_5310,N_5224,N_5141);
or U5311 (N_5311,N_5108,N_5131);
and U5312 (N_5312,N_5188,N_5072);
nand U5313 (N_5313,N_5184,N_5029);
and U5314 (N_5314,N_5090,N_5095);
xnor U5315 (N_5315,N_5203,N_5169);
nor U5316 (N_5316,N_5039,N_5227);
nand U5317 (N_5317,N_5135,N_5073);
or U5318 (N_5318,N_5079,N_5075);
nand U5319 (N_5319,N_5117,N_5100);
xnor U5320 (N_5320,N_5116,N_5018);
xnor U5321 (N_5321,N_5145,N_5055);
or U5322 (N_5322,N_5071,N_5096);
or U5323 (N_5323,N_5186,N_5056);
and U5324 (N_5324,N_5205,N_5185);
nor U5325 (N_5325,N_5115,N_5219);
xnor U5326 (N_5326,N_5013,N_5037);
or U5327 (N_5327,N_5139,N_5113);
xor U5328 (N_5328,N_5241,N_5111);
xnor U5329 (N_5329,N_5123,N_5245);
nand U5330 (N_5330,N_5148,N_5092);
xor U5331 (N_5331,N_5021,N_5032);
nand U5332 (N_5332,N_5182,N_5198);
nor U5333 (N_5333,N_5067,N_5122);
nand U5334 (N_5334,N_5104,N_5229);
or U5335 (N_5335,N_5024,N_5155);
or U5336 (N_5336,N_5156,N_5103);
and U5337 (N_5337,N_5239,N_5023);
xnor U5338 (N_5338,N_5154,N_5207);
nand U5339 (N_5339,N_5177,N_5060);
or U5340 (N_5340,N_5213,N_5049);
or U5341 (N_5341,N_5126,N_5062);
nor U5342 (N_5342,N_5144,N_5121);
and U5343 (N_5343,N_5212,N_5000);
or U5344 (N_5344,N_5140,N_5107);
nand U5345 (N_5345,N_5006,N_5147);
nor U5346 (N_5346,N_5112,N_5099);
nand U5347 (N_5347,N_5165,N_5199);
or U5348 (N_5348,N_5008,N_5015);
xnor U5349 (N_5349,N_5078,N_5110);
nand U5350 (N_5350,N_5236,N_5004);
or U5351 (N_5351,N_5237,N_5076);
or U5352 (N_5352,N_5160,N_5105);
and U5353 (N_5353,N_5162,N_5172);
xnor U5354 (N_5354,N_5064,N_5211);
and U5355 (N_5355,N_5074,N_5181);
and U5356 (N_5356,N_5128,N_5168);
and U5357 (N_5357,N_5001,N_5127);
nor U5358 (N_5358,N_5176,N_5143);
nor U5359 (N_5359,N_5109,N_5178);
nor U5360 (N_5360,N_5042,N_5149);
nand U5361 (N_5361,N_5005,N_5206);
xor U5362 (N_5362,N_5196,N_5166);
xnor U5363 (N_5363,N_5174,N_5142);
nor U5364 (N_5364,N_5246,N_5025);
xor U5365 (N_5365,N_5082,N_5012);
xor U5366 (N_5366,N_5222,N_5235);
nor U5367 (N_5367,N_5204,N_5044);
and U5368 (N_5368,N_5016,N_5134);
nand U5369 (N_5369,N_5191,N_5058);
xor U5370 (N_5370,N_5089,N_5242);
and U5371 (N_5371,N_5238,N_5097);
and U5372 (N_5372,N_5233,N_5132);
nor U5373 (N_5373,N_5150,N_5243);
or U5374 (N_5374,N_5151,N_5124);
nand U5375 (N_5375,N_5021,N_5205);
xor U5376 (N_5376,N_5023,N_5036);
xor U5377 (N_5377,N_5116,N_5166);
nand U5378 (N_5378,N_5014,N_5001);
nor U5379 (N_5379,N_5114,N_5004);
xor U5380 (N_5380,N_5214,N_5131);
nor U5381 (N_5381,N_5230,N_5215);
xnor U5382 (N_5382,N_5110,N_5157);
or U5383 (N_5383,N_5016,N_5084);
and U5384 (N_5384,N_5158,N_5062);
nor U5385 (N_5385,N_5163,N_5125);
nor U5386 (N_5386,N_5246,N_5030);
xor U5387 (N_5387,N_5245,N_5007);
or U5388 (N_5388,N_5221,N_5217);
nand U5389 (N_5389,N_5088,N_5216);
or U5390 (N_5390,N_5040,N_5220);
or U5391 (N_5391,N_5190,N_5108);
nand U5392 (N_5392,N_5172,N_5094);
nor U5393 (N_5393,N_5192,N_5024);
or U5394 (N_5394,N_5035,N_5119);
nor U5395 (N_5395,N_5029,N_5213);
nand U5396 (N_5396,N_5128,N_5058);
nand U5397 (N_5397,N_5246,N_5245);
and U5398 (N_5398,N_5209,N_5154);
and U5399 (N_5399,N_5153,N_5102);
xor U5400 (N_5400,N_5088,N_5038);
and U5401 (N_5401,N_5067,N_5144);
nand U5402 (N_5402,N_5236,N_5083);
nor U5403 (N_5403,N_5007,N_5212);
or U5404 (N_5404,N_5142,N_5008);
or U5405 (N_5405,N_5204,N_5144);
xor U5406 (N_5406,N_5051,N_5116);
nand U5407 (N_5407,N_5147,N_5107);
and U5408 (N_5408,N_5027,N_5134);
or U5409 (N_5409,N_5249,N_5171);
nor U5410 (N_5410,N_5208,N_5110);
nor U5411 (N_5411,N_5107,N_5031);
xnor U5412 (N_5412,N_5151,N_5197);
and U5413 (N_5413,N_5147,N_5099);
xnor U5414 (N_5414,N_5146,N_5131);
and U5415 (N_5415,N_5047,N_5160);
xnor U5416 (N_5416,N_5183,N_5042);
or U5417 (N_5417,N_5141,N_5247);
nand U5418 (N_5418,N_5202,N_5231);
nand U5419 (N_5419,N_5039,N_5120);
or U5420 (N_5420,N_5156,N_5115);
xor U5421 (N_5421,N_5163,N_5054);
or U5422 (N_5422,N_5042,N_5052);
nor U5423 (N_5423,N_5167,N_5155);
nand U5424 (N_5424,N_5220,N_5072);
xnor U5425 (N_5425,N_5003,N_5051);
and U5426 (N_5426,N_5103,N_5099);
and U5427 (N_5427,N_5041,N_5098);
nand U5428 (N_5428,N_5103,N_5166);
nand U5429 (N_5429,N_5060,N_5085);
nor U5430 (N_5430,N_5073,N_5235);
xnor U5431 (N_5431,N_5214,N_5033);
nor U5432 (N_5432,N_5090,N_5118);
nor U5433 (N_5433,N_5063,N_5174);
xnor U5434 (N_5434,N_5072,N_5221);
and U5435 (N_5435,N_5106,N_5044);
nand U5436 (N_5436,N_5204,N_5158);
or U5437 (N_5437,N_5184,N_5016);
or U5438 (N_5438,N_5082,N_5199);
and U5439 (N_5439,N_5116,N_5064);
nor U5440 (N_5440,N_5176,N_5059);
nand U5441 (N_5441,N_5162,N_5083);
nand U5442 (N_5442,N_5026,N_5021);
xnor U5443 (N_5443,N_5010,N_5115);
nor U5444 (N_5444,N_5067,N_5072);
nor U5445 (N_5445,N_5048,N_5096);
xnor U5446 (N_5446,N_5041,N_5093);
and U5447 (N_5447,N_5221,N_5175);
nand U5448 (N_5448,N_5108,N_5221);
nor U5449 (N_5449,N_5098,N_5139);
nor U5450 (N_5450,N_5066,N_5082);
nor U5451 (N_5451,N_5147,N_5247);
and U5452 (N_5452,N_5029,N_5124);
or U5453 (N_5453,N_5161,N_5221);
xor U5454 (N_5454,N_5047,N_5086);
and U5455 (N_5455,N_5055,N_5028);
or U5456 (N_5456,N_5231,N_5229);
nand U5457 (N_5457,N_5146,N_5011);
nand U5458 (N_5458,N_5048,N_5061);
xor U5459 (N_5459,N_5123,N_5136);
xnor U5460 (N_5460,N_5209,N_5056);
or U5461 (N_5461,N_5077,N_5131);
nand U5462 (N_5462,N_5220,N_5013);
and U5463 (N_5463,N_5150,N_5053);
nor U5464 (N_5464,N_5234,N_5197);
or U5465 (N_5465,N_5071,N_5043);
and U5466 (N_5466,N_5003,N_5075);
or U5467 (N_5467,N_5166,N_5163);
or U5468 (N_5468,N_5057,N_5050);
nand U5469 (N_5469,N_5219,N_5027);
and U5470 (N_5470,N_5017,N_5198);
nor U5471 (N_5471,N_5160,N_5060);
nor U5472 (N_5472,N_5021,N_5081);
nand U5473 (N_5473,N_5247,N_5155);
nor U5474 (N_5474,N_5202,N_5179);
or U5475 (N_5475,N_5138,N_5157);
xnor U5476 (N_5476,N_5244,N_5214);
and U5477 (N_5477,N_5140,N_5133);
xor U5478 (N_5478,N_5017,N_5183);
xor U5479 (N_5479,N_5097,N_5158);
xnor U5480 (N_5480,N_5230,N_5171);
nand U5481 (N_5481,N_5047,N_5173);
nand U5482 (N_5482,N_5094,N_5005);
nand U5483 (N_5483,N_5167,N_5136);
or U5484 (N_5484,N_5170,N_5108);
nand U5485 (N_5485,N_5235,N_5175);
nor U5486 (N_5486,N_5103,N_5241);
or U5487 (N_5487,N_5068,N_5098);
nand U5488 (N_5488,N_5064,N_5113);
nor U5489 (N_5489,N_5022,N_5012);
xor U5490 (N_5490,N_5059,N_5064);
xnor U5491 (N_5491,N_5078,N_5117);
nand U5492 (N_5492,N_5203,N_5249);
xnor U5493 (N_5493,N_5045,N_5148);
and U5494 (N_5494,N_5200,N_5000);
or U5495 (N_5495,N_5224,N_5156);
nand U5496 (N_5496,N_5082,N_5085);
nand U5497 (N_5497,N_5089,N_5059);
nor U5498 (N_5498,N_5152,N_5130);
xor U5499 (N_5499,N_5018,N_5220);
nand U5500 (N_5500,N_5417,N_5462);
or U5501 (N_5501,N_5480,N_5348);
nor U5502 (N_5502,N_5264,N_5288);
and U5503 (N_5503,N_5404,N_5250);
or U5504 (N_5504,N_5495,N_5367);
nor U5505 (N_5505,N_5469,N_5328);
nand U5506 (N_5506,N_5483,N_5354);
or U5507 (N_5507,N_5306,N_5361);
nand U5508 (N_5508,N_5323,N_5319);
or U5509 (N_5509,N_5267,N_5254);
nand U5510 (N_5510,N_5358,N_5347);
or U5511 (N_5511,N_5357,N_5396);
nand U5512 (N_5512,N_5496,N_5471);
xnor U5513 (N_5513,N_5460,N_5443);
or U5514 (N_5514,N_5313,N_5437);
and U5515 (N_5515,N_5377,N_5416);
xor U5516 (N_5516,N_5302,N_5286);
or U5517 (N_5517,N_5331,N_5273);
or U5518 (N_5518,N_5397,N_5499);
nor U5519 (N_5519,N_5484,N_5420);
xnor U5520 (N_5520,N_5373,N_5477);
nand U5521 (N_5521,N_5431,N_5285);
and U5522 (N_5522,N_5395,N_5444);
and U5523 (N_5523,N_5493,N_5283);
or U5524 (N_5524,N_5360,N_5301);
xor U5525 (N_5525,N_5317,N_5266);
xor U5526 (N_5526,N_5352,N_5472);
or U5527 (N_5527,N_5439,N_5304);
nand U5528 (N_5528,N_5294,N_5337);
or U5529 (N_5529,N_5277,N_5316);
nor U5530 (N_5530,N_5494,N_5338);
and U5531 (N_5531,N_5315,N_5461);
nor U5532 (N_5532,N_5401,N_5451);
and U5533 (N_5533,N_5255,N_5345);
or U5534 (N_5534,N_5385,N_5275);
nand U5535 (N_5535,N_5473,N_5375);
nor U5536 (N_5536,N_5428,N_5298);
or U5537 (N_5537,N_5307,N_5436);
xnor U5538 (N_5538,N_5262,N_5394);
and U5539 (N_5539,N_5458,N_5498);
xnor U5540 (N_5540,N_5265,N_5445);
xor U5541 (N_5541,N_5467,N_5497);
or U5542 (N_5542,N_5466,N_5336);
nand U5543 (N_5543,N_5435,N_5363);
nor U5544 (N_5544,N_5455,N_5343);
xnor U5545 (N_5545,N_5491,N_5379);
nor U5546 (N_5546,N_5423,N_5413);
nand U5547 (N_5547,N_5274,N_5448);
xor U5548 (N_5548,N_5470,N_5412);
or U5549 (N_5549,N_5297,N_5474);
nand U5550 (N_5550,N_5456,N_5432);
nand U5551 (N_5551,N_5410,N_5415);
or U5552 (N_5552,N_5457,N_5405);
or U5553 (N_5553,N_5406,N_5479);
and U5554 (N_5554,N_5434,N_5369);
nand U5555 (N_5555,N_5291,N_5251);
or U5556 (N_5556,N_5453,N_5409);
or U5557 (N_5557,N_5475,N_5351);
nor U5558 (N_5558,N_5280,N_5365);
and U5559 (N_5559,N_5296,N_5334);
and U5560 (N_5560,N_5468,N_5287);
and U5561 (N_5561,N_5408,N_5449);
nand U5562 (N_5562,N_5447,N_5327);
or U5563 (N_5563,N_5350,N_5344);
and U5564 (N_5564,N_5488,N_5340);
nand U5565 (N_5565,N_5421,N_5402);
nand U5566 (N_5566,N_5368,N_5278);
xnor U5567 (N_5567,N_5333,N_5486);
xor U5568 (N_5568,N_5364,N_5425);
nor U5569 (N_5569,N_5482,N_5299);
or U5570 (N_5570,N_5349,N_5263);
and U5571 (N_5571,N_5381,N_5342);
xor U5572 (N_5572,N_5322,N_5269);
and U5573 (N_5573,N_5355,N_5320);
and U5574 (N_5574,N_5450,N_5332);
or U5575 (N_5575,N_5268,N_5384);
or U5576 (N_5576,N_5300,N_5446);
and U5577 (N_5577,N_5370,N_5330);
and U5578 (N_5578,N_5426,N_5429);
or U5579 (N_5579,N_5492,N_5390);
nand U5580 (N_5580,N_5374,N_5414);
and U5581 (N_5581,N_5292,N_5487);
nor U5582 (N_5582,N_5270,N_5258);
nor U5583 (N_5583,N_5289,N_5438);
xor U5584 (N_5584,N_5485,N_5441);
or U5585 (N_5585,N_5284,N_5389);
nand U5586 (N_5586,N_5276,N_5424);
or U5587 (N_5587,N_5256,N_5372);
nand U5588 (N_5588,N_5309,N_5324);
nand U5589 (N_5589,N_5388,N_5387);
or U5590 (N_5590,N_5359,N_5356);
nor U5591 (N_5591,N_5318,N_5386);
or U5592 (N_5592,N_5454,N_5293);
and U5593 (N_5593,N_5272,N_5489);
nor U5594 (N_5594,N_5392,N_5419);
nor U5595 (N_5595,N_5411,N_5259);
nand U5596 (N_5596,N_5490,N_5311);
and U5597 (N_5597,N_5346,N_5393);
nor U5598 (N_5598,N_5481,N_5391);
and U5599 (N_5599,N_5383,N_5418);
or U5600 (N_5600,N_5335,N_5362);
and U5601 (N_5601,N_5465,N_5400);
xnor U5602 (N_5602,N_5329,N_5326);
or U5603 (N_5603,N_5312,N_5427);
nand U5604 (N_5604,N_5378,N_5398);
or U5605 (N_5605,N_5295,N_5339);
nand U5606 (N_5606,N_5478,N_5407);
or U5607 (N_5607,N_5476,N_5279);
xnor U5608 (N_5608,N_5380,N_5290);
nor U5609 (N_5609,N_5281,N_5308);
and U5610 (N_5610,N_5253,N_5303);
nor U5611 (N_5611,N_5252,N_5366);
nor U5612 (N_5612,N_5310,N_5459);
nand U5613 (N_5613,N_5341,N_5271);
or U5614 (N_5614,N_5261,N_5305);
xnor U5615 (N_5615,N_5403,N_5422);
or U5616 (N_5616,N_5321,N_5282);
nor U5617 (N_5617,N_5464,N_5257);
or U5618 (N_5618,N_5325,N_5260);
xor U5619 (N_5619,N_5376,N_5452);
or U5620 (N_5620,N_5382,N_5399);
and U5621 (N_5621,N_5430,N_5463);
and U5622 (N_5622,N_5353,N_5440);
or U5623 (N_5623,N_5371,N_5314);
or U5624 (N_5624,N_5442,N_5433);
xnor U5625 (N_5625,N_5461,N_5382);
nand U5626 (N_5626,N_5457,N_5473);
xor U5627 (N_5627,N_5459,N_5373);
or U5628 (N_5628,N_5286,N_5464);
and U5629 (N_5629,N_5295,N_5404);
xnor U5630 (N_5630,N_5424,N_5301);
nor U5631 (N_5631,N_5266,N_5362);
and U5632 (N_5632,N_5467,N_5347);
nor U5633 (N_5633,N_5398,N_5400);
and U5634 (N_5634,N_5409,N_5294);
nor U5635 (N_5635,N_5278,N_5258);
and U5636 (N_5636,N_5359,N_5475);
or U5637 (N_5637,N_5385,N_5394);
nand U5638 (N_5638,N_5481,N_5288);
xnor U5639 (N_5639,N_5420,N_5421);
and U5640 (N_5640,N_5406,N_5490);
or U5641 (N_5641,N_5275,N_5483);
nand U5642 (N_5642,N_5285,N_5292);
nor U5643 (N_5643,N_5460,N_5269);
nor U5644 (N_5644,N_5481,N_5329);
or U5645 (N_5645,N_5349,N_5458);
and U5646 (N_5646,N_5362,N_5338);
xnor U5647 (N_5647,N_5255,N_5251);
nand U5648 (N_5648,N_5430,N_5474);
nor U5649 (N_5649,N_5306,N_5381);
nand U5650 (N_5650,N_5385,N_5438);
nand U5651 (N_5651,N_5498,N_5399);
nor U5652 (N_5652,N_5285,N_5256);
or U5653 (N_5653,N_5459,N_5252);
and U5654 (N_5654,N_5430,N_5339);
xor U5655 (N_5655,N_5263,N_5442);
or U5656 (N_5656,N_5407,N_5345);
nand U5657 (N_5657,N_5452,N_5264);
nand U5658 (N_5658,N_5394,N_5431);
nand U5659 (N_5659,N_5402,N_5268);
nand U5660 (N_5660,N_5494,N_5460);
nor U5661 (N_5661,N_5274,N_5313);
and U5662 (N_5662,N_5311,N_5326);
xor U5663 (N_5663,N_5465,N_5324);
xor U5664 (N_5664,N_5280,N_5257);
xor U5665 (N_5665,N_5453,N_5340);
nor U5666 (N_5666,N_5298,N_5376);
nand U5667 (N_5667,N_5273,N_5297);
nand U5668 (N_5668,N_5400,N_5474);
nand U5669 (N_5669,N_5251,N_5365);
and U5670 (N_5670,N_5337,N_5420);
nor U5671 (N_5671,N_5361,N_5263);
nor U5672 (N_5672,N_5269,N_5443);
nand U5673 (N_5673,N_5488,N_5490);
xnor U5674 (N_5674,N_5459,N_5307);
and U5675 (N_5675,N_5268,N_5427);
or U5676 (N_5676,N_5462,N_5270);
xor U5677 (N_5677,N_5369,N_5471);
nand U5678 (N_5678,N_5477,N_5257);
xnor U5679 (N_5679,N_5305,N_5424);
xnor U5680 (N_5680,N_5314,N_5394);
nand U5681 (N_5681,N_5343,N_5321);
and U5682 (N_5682,N_5461,N_5390);
nor U5683 (N_5683,N_5461,N_5448);
nand U5684 (N_5684,N_5369,N_5457);
nand U5685 (N_5685,N_5321,N_5290);
xnor U5686 (N_5686,N_5422,N_5331);
and U5687 (N_5687,N_5392,N_5480);
or U5688 (N_5688,N_5376,N_5463);
xor U5689 (N_5689,N_5270,N_5402);
nand U5690 (N_5690,N_5499,N_5462);
or U5691 (N_5691,N_5498,N_5423);
nand U5692 (N_5692,N_5257,N_5335);
nor U5693 (N_5693,N_5270,N_5371);
and U5694 (N_5694,N_5340,N_5270);
nor U5695 (N_5695,N_5328,N_5314);
and U5696 (N_5696,N_5461,N_5409);
and U5697 (N_5697,N_5460,N_5489);
and U5698 (N_5698,N_5401,N_5266);
and U5699 (N_5699,N_5463,N_5299);
or U5700 (N_5700,N_5307,N_5336);
nor U5701 (N_5701,N_5260,N_5307);
xor U5702 (N_5702,N_5447,N_5392);
and U5703 (N_5703,N_5328,N_5348);
or U5704 (N_5704,N_5475,N_5255);
or U5705 (N_5705,N_5333,N_5497);
xor U5706 (N_5706,N_5259,N_5292);
nor U5707 (N_5707,N_5490,N_5424);
nor U5708 (N_5708,N_5491,N_5421);
or U5709 (N_5709,N_5470,N_5410);
nand U5710 (N_5710,N_5476,N_5267);
or U5711 (N_5711,N_5325,N_5313);
nor U5712 (N_5712,N_5361,N_5372);
or U5713 (N_5713,N_5409,N_5268);
nor U5714 (N_5714,N_5302,N_5320);
and U5715 (N_5715,N_5459,N_5435);
xnor U5716 (N_5716,N_5357,N_5403);
and U5717 (N_5717,N_5474,N_5315);
xnor U5718 (N_5718,N_5476,N_5441);
xnor U5719 (N_5719,N_5497,N_5410);
xnor U5720 (N_5720,N_5314,N_5415);
or U5721 (N_5721,N_5310,N_5363);
and U5722 (N_5722,N_5263,N_5274);
nand U5723 (N_5723,N_5254,N_5357);
nor U5724 (N_5724,N_5423,N_5416);
nor U5725 (N_5725,N_5464,N_5262);
and U5726 (N_5726,N_5368,N_5409);
xnor U5727 (N_5727,N_5288,N_5420);
xor U5728 (N_5728,N_5269,N_5357);
or U5729 (N_5729,N_5427,N_5457);
xnor U5730 (N_5730,N_5485,N_5331);
and U5731 (N_5731,N_5436,N_5327);
and U5732 (N_5732,N_5293,N_5498);
nand U5733 (N_5733,N_5437,N_5307);
and U5734 (N_5734,N_5430,N_5362);
xnor U5735 (N_5735,N_5350,N_5396);
or U5736 (N_5736,N_5283,N_5425);
nor U5737 (N_5737,N_5252,N_5480);
nor U5738 (N_5738,N_5395,N_5456);
nor U5739 (N_5739,N_5305,N_5279);
or U5740 (N_5740,N_5497,N_5308);
xor U5741 (N_5741,N_5336,N_5299);
or U5742 (N_5742,N_5365,N_5443);
nor U5743 (N_5743,N_5406,N_5296);
xnor U5744 (N_5744,N_5308,N_5427);
nor U5745 (N_5745,N_5409,N_5300);
and U5746 (N_5746,N_5457,N_5419);
nand U5747 (N_5747,N_5412,N_5362);
nand U5748 (N_5748,N_5262,N_5497);
xnor U5749 (N_5749,N_5446,N_5428);
nor U5750 (N_5750,N_5563,N_5685);
nor U5751 (N_5751,N_5652,N_5682);
nand U5752 (N_5752,N_5734,N_5641);
nor U5753 (N_5753,N_5599,N_5698);
or U5754 (N_5754,N_5549,N_5586);
and U5755 (N_5755,N_5673,N_5525);
or U5756 (N_5756,N_5645,N_5601);
nand U5757 (N_5757,N_5744,N_5602);
or U5758 (N_5758,N_5657,N_5658);
nor U5759 (N_5759,N_5571,N_5520);
nor U5760 (N_5760,N_5692,N_5527);
and U5761 (N_5761,N_5637,N_5597);
xor U5762 (N_5762,N_5581,N_5731);
nor U5763 (N_5763,N_5509,N_5626);
nand U5764 (N_5764,N_5546,N_5510);
nand U5765 (N_5765,N_5643,N_5655);
xor U5766 (N_5766,N_5729,N_5696);
and U5767 (N_5767,N_5565,N_5539);
and U5768 (N_5768,N_5740,N_5500);
nand U5769 (N_5769,N_5663,N_5543);
nor U5770 (N_5770,N_5676,N_5651);
and U5771 (N_5771,N_5606,N_5735);
nor U5772 (N_5772,N_5512,N_5687);
and U5773 (N_5773,N_5721,N_5552);
xnor U5774 (N_5774,N_5653,N_5580);
nor U5775 (N_5775,N_5679,N_5727);
nor U5776 (N_5776,N_5694,N_5529);
nand U5777 (N_5777,N_5559,N_5741);
xnor U5778 (N_5778,N_5587,N_5714);
or U5779 (N_5779,N_5584,N_5627);
nor U5780 (N_5780,N_5739,N_5569);
xor U5781 (N_5781,N_5554,N_5647);
xnor U5782 (N_5782,N_5594,N_5531);
xor U5783 (N_5783,N_5656,N_5702);
nor U5784 (N_5784,N_5747,N_5621);
or U5785 (N_5785,N_5585,N_5620);
or U5786 (N_5786,N_5650,N_5530);
or U5787 (N_5787,N_5723,N_5590);
nor U5788 (N_5788,N_5556,N_5700);
or U5789 (N_5789,N_5681,N_5607);
xnor U5790 (N_5790,N_5671,N_5522);
or U5791 (N_5791,N_5670,N_5675);
xnor U5792 (N_5792,N_5541,N_5610);
nand U5793 (N_5793,N_5715,N_5557);
nor U5794 (N_5794,N_5718,N_5630);
or U5795 (N_5795,N_5708,N_5664);
and U5796 (N_5796,N_5699,N_5629);
or U5797 (N_5797,N_5667,N_5553);
and U5798 (N_5798,N_5632,N_5619);
xnor U5799 (N_5799,N_5726,N_5506);
nor U5800 (N_5800,N_5591,N_5532);
or U5801 (N_5801,N_5614,N_5697);
or U5802 (N_5802,N_5578,N_5707);
or U5803 (N_5803,N_5745,N_5640);
and U5804 (N_5804,N_5706,N_5513);
nor U5805 (N_5805,N_5633,N_5730);
xor U5806 (N_5806,N_5720,N_5690);
nand U5807 (N_5807,N_5528,N_5518);
nor U5808 (N_5808,N_5574,N_5716);
nor U5809 (N_5809,N_5711,N_5634);
and U5810 (N_5810,N_5540,N_5662);
nor U5811 (N_5811,N_5737,N_5573);
or U5812 (N_5812,N_5588,N_5505);
or U5813 (N_5813,N_5514,N_5649);
or U5814 (N_5814,N_5560,N_5595);
or U5815 (N_5815,N_5547,N_5515);
xnor U5816 (N_5816,N_5644,N_5677);
nor U5817 (N_5817,N_5577,N_5639);
nor U5818 (N_5818,N_5749,N_5542);
and U5819 (N_5819,N_5738,N_5674);
and U5820 (N_5820,N_5558,N_5704);
nand U5821 (N_5821,N_5544,N_5507);
nor U5822 (N_5822,N_5502,N_5576);
or U5823 (N_5823,N_5517,N_5618);
or U5824 (N_5824,N_5736,N_5533);
or U5825 (N_5825,N_5661,N_5669);
xnor U5826 (N_5826,N_5600,N_5659);
and U5827 (N_5827,N_5562,N_5642);
and U5828 (N_5828,N_5603,N_5579);
or U5829 (N_5829,N_5501,N_5617);
and U5830 (N_5830,N_5534,N_5710);
and U5831 (N_5831,N_5713,N_5668);
or U5832 (N_5832,N_5566,N_5508);
and U5833 (N_5833,N_5719,N_5678);
xnor U5834 (N_5834,N_5665,N_5703);
and U5835 (N_5835,N_5688,N_5689);
and U5836 (N_5836,N_5526,N_5561);
nor U5837 (N_5837,N_5538,N_5733);
nand U5838 (N_5838,N_5550,N_5725);
or U5839 (N_5839,N_5609,N_5672);
nand U5840 (N_5840,N_5748,N_5605);
nand U5841 (N_5841,N_5746,N_5516);
or U5842 (N_5842,N_5680,N_5705);
nor U5843 (N_5843,N_5537,N_5615);
or U5844 (N_5844,N_5684,N_5582);
nand U5845 (N_5845,N_5660,N_5598);
and U5846 (N_5846,N_5709,N_5608);
and U5847 (N_5847,N_5548,N_5636);
xor U5848 (N_5848,N_5712,N_5701);
nor U5849 (N_5849,N_5732,N_5613);
xor U5850 (N_5850,N_5519,N_5568);
nor U5851 (N_5851,N_5572,N_5717);
and U5852 (N_5852,N_5524,N_5654);
nor U5853 (N_5853,N_5646,N_5567);
and U5854 (N_5854,N_5691,N_5742);
nor U5855 (N_5855,N_5638,N_5722);
xnor U5856 (N_5856,N_5625,N_5628);
nor U5857 (N_5857,N_5624,N_5593);
nor U5858 (N_5858,N_5575,N_5592);
or U5859 (N_5859,N_5570,N_5631);
and U5860 (N_5860,N_5535,N_5612);
and U5861 (N_5861,N_5596,N_5695);
and U5862 (N_5862,N_5728,N_5551);
or U5863 (N_5863,N_5611,N_5648);
xnor U5864 (N_5864,N_5504,N_5616);
nor U5865 (N_5865,N_5686,N_5724);
and U5866 (N_5866,N_5635,N_5503);
or U5867 (N_5867,N_5583,N_5666);
nor U5868 (N_5868,N_5693,N_5521);
nor U5869 (N_5869,N_5683,N_5545);
xnor U5870 (N_5870,N_5622,N_5523);
xnor U5871 (N_5871,N_5564,N_5623);
and U5872 (N_5872,N_5555,N_5589);
nor U5873 (N_5873,N_5743,N_5604);
or U5874 (N_5874,N_5511,N_5536);
and U5875 (N_5875,N_5692,N_5571);
nor U5876 (N_5876,N_5711,N_5700);
nand U5877 (N_5877,N_5609,N_5725);
and U5878 (N_5878,N_5596,N_5548);
and U5879 (N_5879,N_5503,N_5551);
nand U5880 (N_5880,N_5628,N_5562);
nand U5881 (N_5881,N_5733,N_5611);
or U5882 (N_5882,N_5695,N_5598);
or U5883 (N_5883,N_5545,N_5602);
and U5884 (N_5884,N_5663,N_5590);
xnor U5885 (N_5885,N_5501,N_5591);
nand U5886 (N_5886,N_5648,N_5620);
nor U5887 (N_5887,N_5743,N_5723);
nand U5888 (N_5888,N_5544,N_5696);
and U5889 (N_5889,N_5697,N_5705);
or U5890 (N_5890,N_5659,N_5584);
nand U5891 (N_5891,N_5725,N_5562);
or U5892 (N_5892,N_5614,N_5625);
nand U5893 (N_5893,N_5688,N_5668);
nand U5894 (N_5894,N_5694,N_5667);
or U5895 (N_5895,N_5664,N_5612);
nand U5896 (N_5896,N_5589,N_5585);
and U5897 (N_5897,N_5523,N_5550);
or U5898 (N_5898,N_5602,N_5724);
or U5899 (N_5899,N_5505,N_5747);
or U5900 (N_5900,N_5621,N_5585);
xnor U5901 (N_5901,N_5604,N_5601);
and U5902 (N_5902,N_5527,N_5707);
nor U5903 (N_5903,N_5537,N_5683);
nand U5904 (N_5904,N_5644,N_5692);
xnor U5905 (N_5905,N_5511,N_5543);
and U5906 (N_5906,N_5660,N_5736);
or U5907 (N_5907,N_5691,N_5639);
nor U5908 (N_5908,N_5704,N_5643);
xnor U5909 (N_5909,N_5578,N_5604);
nor U5910 (N_5910,N_5535,N_5736);
nand U5911 (N_5911,N_5524,N_5611);
and U5912 (N_5912,N_5571,N_5720);
nor U5913 (N_5913,N_5728,N_5739);
xnor U5914 (N_5914,N_5591,N_5691);
and U5915 (N_5915,N_5535,N_5688);
nor U5916 (N_5916,N_5601,N_5732);
and U5917 (N_5917,N_5683,N_5716);
xnor U5918 (N_5918,N_5561,N_5620);
xor U5919 (N_5919,N_5722,N_5702);
and U5920 (N_5920,N_5726,N_5670);
or U5921 (N_5921,N_5539,N_5667);
nor U5922 (N_5922,N_5561,N_5580);
xnor U5923 (N_5923,N_5649,N_5737);
nor U5924 (N_5924,N_5512,N_5745);
nand U5925 (N_5925,N_5546,N_5576);
nor U5926 (N_5926,N_5572,N_5741);
nor U5927 (N_5927,N_5649,N_5701);
nand U5928 (N_5928,N_5555,N_5721);
or U5929 (N_5929,N_5673,N_5720);
nor U5930 (N_5930,N_5609,N_5579);
or U5931 (N_5931,N_5508,N_5500);
xor U5932 (N_5932,N_5666,N_5522);
nor U5933 (N_5933,N_5525,N_5567);
xnor U5934 (N_5934,N_5684,N_5658);
xnor U5935 (N_5935,N_5709,N_5696);
xor U5936 (N_5936,N_5690,N_5582);
or U5937 (N_5937,N_5720,N_5573);
xor U5938 (N_5938,N_5649,N_5584);
and U5939 (N_5939,N_5598,N_5645);
nand U5940 (N_5940,N_5586,N_5595);
nor U5941 (N_5941,N_5629,N_5592);
and U5942 (N_5942,N_5640,N_5528);
nand U5943 (N_5943,N_5552,N_5646);
nand U5944 (N_5944,N_5721,N_5541);
nor U5945 (N_5945,N_5649,N_5543);
nor U5946 (N_5946,N_5699,N_5517);
nand U5947 (N_5947,N_5521,N_5661);
xor U5948 (N_5948,N_5651,N_5506);
or U5949 (N_5949,N_5665,N_5633);
nand U5950 (N_5950,N_5510,N_5682);
xnor U5951 (N_5951,N_5537,N_5582);
nor U5952 (N_5952,N_5626,N_5747);
and U5953 (N_5953,N_5716,N_5624);
nand U5954 (N_5954,N_5565,N_5643);
or U5955 (N_5955,N_5629,N_5661);
and U5956 (N_5956,N_5641,N_5726);
xor U5957 (N_5957,N_5567,N_5598);
xnor U5958 (N_5958,N_5543,N_5668);
nor U5959 (N_5959,N_5645,N_5712);
nand U5960 (N_5960,N_5658,N_5682);
nand U5961 (N_5961,N_5567,N_5643);
nand U5962 (N_5962,N_5729,N_5634);
nand U5963 (N_5963,N_5537,N_5662);
nand U5964 (N_5964,N_5599,N_5681);
or U5965 (N_5965,N_5705,N_5706);
nand U5966 (N_5966,N_5573,N_5556);
and U5967 (N_5967,N_5703,N_5648);
and U5968 (N_5968,N_5554,N_5617);
nor U5969 (N_5969,N_5709,N_5629);
xor U5970 (N_5970,N_5544,N_5736);
and U5971 (N_5971,N_5580,N_5712);
and U5972 (N_5972,N_5676,N_5743);
and U5973 (N_5973,N_5504,N_5558);
or U5974 (N_5974,N_5610,N_5614);
xor U5975 (N_5975,N_5727,N_5624);
or U5976 (N_5976,N_5612,N_5731);
and U5977 (N_5977,N_5726,N_5543);
nand U5978 (N_5978,N_5598,N_5748);
nand U5979 (N_5979,N_5566,N_5627);
xnor U5980 (N_5980,N_5504,N_5536);
nor U5981 (N_5981,N_5721,N_5581);
xor U5982 (N_5982,N_5537,N_5740);
nor U5983 (N_5983,N_5625,N_5652);
xnor U5984 (N_5984,N_5589,N_5546);
nand U5985 (N_5985,N_5588,N_5530);
and U5986 (N_5986,N_5566,N_5725);
or U5987 (N_5987,N_5720,N_5612);
nand U5988 (N_5988,N_5717,N_5543);
nand U5989 (N_5989,N_5592,N_5713);
or U5990 (N_5990,N_5710,N_5680);
nand U5991 (N_5991,N_5680,N_5624);
and U5992 (N_5992,N_5581,N_5694);
nand U5993 (N_5993,N_5510,N_5561);
or U5994 (N_5994,N_5708,N_5686);
nor U5995 (N_5995,N_5577,N_5659);
nand U5996 (N_5996,N_5679,N_5500);
nand U5997 (N_5997,N_5533,N_5647);
xor U5998 (N_5998,N_5698,N_5680);
nand U5999 (N_5999,N_5557,N_5742);
or U6000 (N_6000,N_5891,N_5801);
or U6001 (N_6001,N_5792,N_5964);
nor U6002 (N_6002,N_5900,N_5903);
nor U6003 (N_6003,N_5895,N_5876);
nand U6004 (N_6004,N_5928,N_5938);
xnor U6005 (N_6005,N_5944,N_5889);
or U6006 (N_6006,N_5793,N_5858);
and U6007 (N_6007,N_5764,N_5786);
and U6008 (N_6008,N_5892,N_5835);
nand U6009 (N_6009,N_5896,N_5781);
xnor U6010 (N_6010,N_5911,N_5809);
and U6011 (N_6011,N_5804,N_5899);
nand U6012 (N_6012,N_5841,N_5916);
and U6013 (N_6013,N_5963,N_5825);
nand U6014 (N_6014,N_5874,N_5821);
or U6015 (N_6015,N_5890,N_5819);
and U6016 (N_6016,N_5852,N_5850);
xnor U6017 (N_6017,N_5766,N_5935);
xor U6018 (N_6018,N_5957,N_5864);
nor U6019 (N_6019,N_5912,N_5937);
nand U6020 (N_6020,N_5824,N_5770);
nand U6021 (N_6021,N_5844,N_5826);
nand U6022 (N_6022,N_5830,N_5902);
nand U6023 (N_6023,N_5833,N_5757);
or U6024 (N_6024,N_5782,N_5989);
xor U6025 (N_6025,N_5991,N_5842);
or U6026 (N_6026,N_5914,N_5929);
nand U6027 (N_6027,N_5878,N_5897);
or U6028 (N_6028,N_5885,N_5822);
xnor U6029 (N_6029,N_5956,N_5845);
nor U6030 (N_6030,N_5834,N_5931);
nand U6031 (N_6031,N_5777,N_5775);
and U6032 (N_6032,N_5872,N_5949);
nand U6033 (N_6033,N_5769,N_5838);
nand U6034 (N_6034,N_5827,N_5905);
nand U6035 (N_6035,N_5868,N_5977);
nand U6036 (N_6036,N_5979,N_5799);
or U6037 (N_6037,N_5780,N_5814);
xnor U6038 (N_6038,N_5820,N_5856);
nor U6039 (N_6039,N_5970,N_5969);
or U6040 (N_6040,N_5971,N_5754);
or U6041 (N_6041,N_5960,N_5857);
nor U6042 (N_6042,N_5915,N_5761);
xnor U6043 (N_6043,N_5803,N_5869);
and U6044 (N_6044,N_5785,N_5855);
or U6045 (N_6045,N_5788,N_5783);
and U6046 (N_6046,N_5796,N_5866);
nor U6047 (N_6047,N_5829,N_5887);
nand U6048 (N_6048,N_5948,N_5807);
nand U6049 (N_6049,N_5818,N_5906);
or U6050 (N_6050,N_5907,N_5898);
or U6051 (N_6051,N_5945,N_5919);
nor U6052 (N_6052,N_5815,N_5930);
nor U6053 (N_6053,N_5848,N_5883);
nand U6054 (N_6054,N_5973,N_5942);
and U6055 (N_6055,N_5975,N_5943);
and U6056 (N_6056,N_5880,N_5965);
nor U6057 (N_6057,N_5932,N_5918);
or U6058 (N_6058,N_5993,N_5805);
nand U6059 (N_6059,N_5831,N_5972);
and U6060 (N_6060,N_5924,N_5996);
nand U6061 (N_6061,N_5836,N_5771);
xor U6062 (N_6062,N_5952,N_5851);
and U6063 (N_6063,N_5999,N_5910);
and U6064 (N_6064,N_5976,N_5927);
xor U6065 (N_6065,N_5753,N_5756);
nor U6066 (N_6066,N_5961,N_5791);
nor U6067 (N_6067,N_5763,N_5816);
and U6068 (N_6068,N_5794,N_5837);
xnor U6069 (N_6069,N_5789,N_5861);
nor U6070 (N_6070,N_5779,N_5790);
or U6071 (N_6071,N_5940,N_5750);
or U6072 (N_6072,N_5968,N_5995);
nor U6073 (N_6073,N_5980,N_5759);
and U6074 (N_6074,N_5984,N_5920);
xor U6075 (N_6075,N_5894,N_5862);
or U6076 (N_6076,N_5901,N_5859);
nor U6077 (N_6077,N_5797,N_5812);
nor U6078 (N_6078,N_5986,N_5768);
or U6079 (N_6079,N_5879,N_5776);
or U6080 (N_6080,N_5955,N_5823);
nand U6081 (N_6081,N_5994,N_5967);
and U6082 (N_6082,N_5832,N_5959);
nand U6083 (N_6083,N_5925,N_5817);
nor U6084 (N_6084,N_5787,N_5870);
nand U6085 (N_6085,N_5755,N_5987);
xor U6086 (N_6086,N_5947,N_5784);
nor U6087 (N_6087,N_5758,N_5767);
and U6088 (N_6088,N_5908,N_5765);
xnor U6089 (N_6089,N_5941,N_5958);
or U6090 (N_6090,N_5840,N_5988);
or U6091 (N_6091,N_5939,N_5922);
nor U6092 (N_6092,N_5946,N_5985);
and U6093 (N_6093,N_5888,N_5843);
xor U6094 (N_6094,N_5798,N_5795);
and U6095 (N_6095,N_5962,N_5839);
nand U6096 (N_6096,N_5875,N_5998);
and U6097 (N_6097,N_5893,N_5867);
xor U6098 (N_6098,N_5953,N_5863);
nand U6099 (N_6099,N_5828,N_5773);
and U6100 (N_6100,N_5904,N_5992);
and U6101 (N_6101,N_5974,N_5854);
nand U6102 (N_6102,N_5810,N_5936);
nor U6103 (N_6103,N_5997,N_5865);
nor U6104 (N_6104,N_5778,N_5800);
and U6105 (N_6105,N_5751,N_5752);
nand U6106 (N_6106,N_5966,N_5983);
nand U6107 (N_6107,N_5847,N_5913);
xnor U6108 (N_6108,N_5982,N_5950);
nand U6109 (N_6109,N_5881,N_5951);
or U6110 (N_6110,N_5871,N_5808);
nor U6111 (N_6111,N_5762,N_5934);
or U6112 (N_6112,N_5853,N_5990);
nand U6113 (N_6113,N_5909,N_5923);
xnor U6114 (N_6114,N_5860,N_5849);
and U6115 (N_6115,N_5882,N_5917);
or U6116 (N_6116,N_5802,N_5760);
nor U6117 (N_6117,N_5813,N_5954);
nor U6118 (N_6118,N_5877,N_5873);
or U6119 (N_6119,N_5926,N_5978);
and U6120 (N_6120,N_5774,N_5921);
nand U6121 (N_6121,N_5811,N_5884);
nand U6122 (N_6122,N_5886,N_5981);
and U6123 (N_6123,N_5806,N_5772);
xor U6124 (N_6124,N_5933,N_5846);
and U6125 (N_6125,N_5757,N_5887);
nor U6126 (N_6126,N_5757,N_5989);
nand U6127 (N_6127,N_5787,N_5840);
nor U6128 (N_6128,N_5934,N_5926);
and U6129 (N_6129,N_5888,N_5996);
xor U6130 (N_6130,N_5956,N_5836);
nand U6131 (N_6131,N_5810,N_5991);
nand U6132 (N_6132,N_5990,N_5915);
and U6133 (N_6133,N_5933,N_5916);
and U6134 (N_6134,N_5956,N_5768);
and U6135 (N_6135,N_5932,N_5941);
xor U6136 (N_6136,N_5868,N_5961);
nand U6137 (N_6137,N_5752,N_5886);
or U6138 (N_6138,N_5928,N_5888);
xor U6139 (N_6139,N_5966,N_5935);
or U6140 (N_6140,N_5769,N_5984);
and U6141 (N_6141,N_5943,N_5962);
nor U6142 (N_6142,N_5983,N_5890);
and U6143 (N_6143,N_5914,N_5896);
and U6144 (N_6144,N_5767,N_5798);
and U6145 (N_6145,N_5954,N_5928);
or U6146 (N_6146,N_5871,N_5880);
or U6147 (N_6147,N_5959,N_5885);
and U6148 (N_6148,N_5963,N_5886);
nand U6149 (N_6149,N_5814,N_5875);
xor U6150 (N_6150,N_5980,N_5827);
or U6151 (N_6151,N_5996,N_5901);
and U6152 (N_6152,N_5773,N_5774);
nand U6153 (N_6153,N_5983,N_5854);
or U6154 (N_6154,N_5775,N_5841);
xnor U6155 (N_6155,N_5775,N_5854);
nand U6156 (N_6156,N_5791,N_5810);
nor U6157 (N_6157,N_5974,N_5896);
xnor U6158 (N_6158,N_5750,N_5828);
xor U6159 (N_6159,N_5868,N_5942);
nand U6160 (N_6160,N_5908,N_5886);
nand U6161 (N_6161,N_5951,N_5985);
nor U6162 (N_6162,N_5809,N_5930);
or U6163 (N_6163,N_5850,N_5843);
or U6164 (N_6164,N_5773,N_5799);
nand U6165 (N_6165,N_5944,N_5801);
nand U6166 (N_6166,N_5775,N_5963);
and U6167 (N_6167,N_5897,N_5883);
and U6168 (N_6168,N_5808,N_5881);
nor U6169 (N_6169,N_5776,N_5750);
nor U6170 (N_6170,N_5909,N_5932);
nand U6171 (N_6171,N_5886,N_5892);
and U6172 (N_6172,N_5827,N_5911);
and U6173 (N_6173,N_5886,N_5856);
or U6174 (N_6174,N_5882,N_5812);
and U6175 (N_6175,N_5826,N_5913);
nand U6176 (N_6176,N_5753,N_5835);
nor U6177 (N_6177,N_5866,N_5848);
and U6178 (N_6178,N_5922,N_5909);
xnor U6179 (N_6179,N_5766,N_5961);
nor U6180 (N_6180,N_5925,N_5860);
xnor U6181 (N_6181,N_5781,N_5996);
nand U6182 (N_6182,N_5973,N_5773);
and U6183 (N_6183,N_5843,N_5886);
nor U6184 (N_6184,N_5861,N_5786);
nor U6185 (N_6185,N_5840,N_5995);
nand U6186 (N_6186,N_5781,N_5792);
nor U6187 (N_6187,N_5989,N_5987);
and U6188 (N_6188,N_5753,N_5926);
nor U6189 (N_6189,N_5827,N_5935);
and U6190 (N_6190,N_5767,N_5760);
and U6191 (N_6191,N_5907,N_5924);
xnor U6192 (N_6192,N_5811,N_5990);
nor U6193 (N_6193,N_5963,N_5818);
nor U6194 (N_6194,N_5957,N_5758);
nor U6195 (N_6195,N_5928,N_5882);
nand U6196 (N_6196,N_5959,N_5800);
nor U6197 (N_6197,N_5999,N_5996);
xor U6198 (N_6198,N_5827,N_5756);
and U6199 (N_6199,N_5798,N_5846);
or U6200 (N_6200,N_5847,N_5988);
nand U6201 (N_6201,N_5769,N_5958);
or U6202 (N_6202,N_5845,N_5964);
nor U6203 (N_6203,N_5934,N_5754);
and U6204 (N_6204,N_5811,N_5813);
nand U6205 (N_6205,N_5911,N_5891);
and U6206 (N_6206,N_5796,N_5777);
nand U6207 (N_6207,N_5800,N_5886);
nor U6208 (N_6208,N_5778,N_5900);
or U6209 (N_6209,N_5758,N_5845);
nor U6210 (N_6210,N_5765,N_5821);
or U6211 (N_6211,N_5769,N_5869);
xor U6212 (N_6212,N_5783,N_5877);
xor U6213 (N_6213,N_5756,N_5973);
nor U6214 (N_6214,N_5851,N_5949);
xor U6215 (N_6215,N_5963,N_5788);
nor U6216 (N_6216,N_5799,N_5959);
or U6217 (N_6217,N_5977,N_5859);
xor U6218 (N_6218,N_5818,N_5887);
xor U6219 (N_6219,N_5921,N_5804);
nand U6220 (N_6220,N_5923,N_5908);
xor U6221 (N_6221,N_5832,N_5826);
and U6222 (N_6222,N_5883,N_5872);
xor U6223 (N_6223,N_5915,N_5979);
and U6224 (N_6224,N_5849,N_5793);
or U6225 (N_6225,N_5899,N_5909);
nor U6226 (N_6226,N_5874,N_5983);
nor U6227 (N_6227,N_5904,N_5932);
nand U6228 (N_6228,N_5881,N_5789);
or U6229 (N_6229,N_5899,N_5965);
and U6230 (N_6230,N_5897,N_5831);
or U6231 (N_6231,N_5828,N_5817);
xor U6232 (N_6232,N_5857,N_5861);
nand U6233 (N_6233,N_5753,N_5909);
or U6234 (N_6234,N_5822,N_5916);
nand U6235 (N_6235,N_5816,N_5859);
or U6236 (N_6236,N_5768,N_5927);
xnor U6237 (N_6237,N_5908,N_5869);
xor U6238 (N_6238,N_5995,N_5980);
nand U6239 (N_6239,N_5767,N_5773);
xnor U6240 (N_6240,N_5991,N_5985);
xnor U6241 (N_6241,N_5948,N_5958);
nand U6242 (N_6242,N_5905,N_5792);
nor U6243 (N_6243,N_5846,N_5767);
nor U6244 (N_6244,N_5789,N_5755);
xor U6245 (N_6245,N_5893,N_5796);
xor U6246 (N_6246,N_5900,N_5916);
or U6247 (N_6247,N_5753,N_5766);
and U6248 (N_6248,N_5872,N_5847);
xor U6249 (N_6249,N_5774,N_5771);
nor U6250 (N_6250,N_6040,N_6139);
xnor U6251 (N_6251,N_6109,N_6206);
xnor U6252 (N_6252,N_6110,N_6166);
nor U6253 (N_6253,N_6188,N_6158);
and U6254 (N_6254,N_6190,N_6242);
nor U6255 (N_6255,N_6221,N_6087);
and U6256 (N_6256,N_6127,N_6005);
and U6257 (N_6257,N_6006,N_6026);
or U6258 (N_6258,N_6047,N_6069);
nand U6259 (N_6259,N_6182,N_6028);
or U6260 (N_6260,N_6164,N_6238);
or U6261 (N_6261,N_6223,N_6000);
and U6262 (N_6262,N_6219,N_6147);
nand U6263 (N_6263,N_6211,N_6120);
nor U6264 (N_6264,N_6133,N_6093);
nand U6265 (N_6265,N_6151,N_6220);
and U6266 (N_6266,N_6153,N_6117);
nand U6267 (N_6267,N_6099,N_6012);
nor U6268 (N_6268,N_6014,N_6107);
nor U6269 (N_6269,N_6094,N_6171);
and U6270 (N_6270,N_6236,N_6168);
nand U6271 (N_6271,N_6249,N_6024);
nand U6272 (N_6272,N_6111,N_6141);
or U6273 (N_6273,N_6149,N_6010);
and U6274 (N_6274,N_6072,N_6246);
nand U6275 (N_6275,N_6082,N_6064);
nor U6276 (N_6276,N_6029,N_6144);
nor U6277 (N_6277,N_6131,N_6180);
xor U6278 (N_6278,N_6178,N_6034);
nor U6279 (N_6279,N_6090,N_6142);
xnor U6280 (N_6280,N_6212,N_6112);
or U6281 (N_6281,N_6031,N_6032);
xor U6282 (N_6282,N_6247,N_6183);
nand U6283 (N_6283,N_6136,N_6085);
nand U6284 (N_6284,N_6067,N_6020);
nor U6285 (N_6285,N_6083,N_6209);
nand U6286 (N_6286,N_6013,N_6145);
xnor U6287 (N_6287,N_6123,N_6002);
and U6288 (N_6288,N_6042,N_6074);
xnor U6289 (N_6289,N_6025,N_6222);
nand U6290 (N_6290,N_6003,N_6241);
xor U6291 (N_6291,N_6038,N_6102);
or U6292 (N_6292,N_6049,N_6231);
xnor U6293 (N_6293,N_6077,N_6174);
nor U6294 (N_6294,N_6179,N_6098);
and U6295 (N_6295,N_6134,N_6041);
nand U6296 (N_6296,N_6050,N_6185);
nand U6297 (N_6297,N_6066,N_6137);
nand U6298 (N_6298,N_6015,N_6202);
nand U6299 (N_6299,N_6103,N_6161);
nor U6300 (N_6300,N_6073,N_6106);
xnor U6301 (N_6301,N_6167,N_6101);
nand U6302 (N_6302,N_6229,N_6104);
xnor U6303 (N_6303,N_6157,N_6227);
nor U6304 (N_6304,N_6060,N_6243);
nand U6305 (N_6305,N_6114,N_6004);
or U6306 (N_6306,N_6030,N_6019);
nor U6307 (N_6307,N_6172,N_6045);
nor U6308 (N_6308,N_6197,N_6080);
xnor U6309 (N_6309,N_6065,N_6175);
nor U6310 (N_6310,N_6037,N_6070);
and U6311 (N_6311,N_6048,N_6152);
nand U6312 (N_6312,N_6226,N_6196);
nand U6313 (N_6313,N_6043,N_6105);
nor U6314 (N_6314,N_6135,N_6011);
nor U6315 (N_6315,N_6095,N_6063);
and U6316 (N_6316,N_6071,N_6100);
or U6317 (N_6317,N_6201,N_6078);
or U6318 (N_6318,N_6176,N_6009);
nor U6319 (N_6319,N_6075,N_6205);
or U6320 (N_6320,N_6181,N_6208);
or U6321 (N_6321,N_6035,N_6097);
nor U6322 (N_6322,N_6195,N_6173);
nor U6323 (N_6323,N_6210,N_6194);
nor U6324 (N_6324,N_6232,N_6129);
or U6325 (N_6325,N_6001,N_6160);
nor U6326 (N_6326,N_6079,N_6027);
or U6327 (N_6327,N_6008,N_6096);
and U6328 (N_6328,N_6051,N_6061);
or U6329 (N_6329,N_6039,N_6062);
and U6330 (N_6330,N_6216,N_6125);
nor U6331 (N_6331,N_6213,N_6113);
nor U6332 (N_6332,N_6245,N_6054);
nor U6333 (N_6333,N_6122,N_6156);
or U6334 (N_6334,N_6022,N_6148);
xor U6335 (N_6335,N_6116,N_6233);
nand U6336 (N_6336,N_6186,N_6244);
or U6337 (N_6337,N_6053,N_6132);
xor U6338 (N_6338,N_6184,N_6052);
xor U6339 (N_6339,N_6187,N_6169);
and U6340 (N_6340,N_6046,N_6198);
and U6341 (N_6341,N_6215,N_6128);
and U6342 (N_6342,N_6217,N_6057);
and U6343 (N_6343,N_6119,N_6155);
xnor U6344 (N_6344,N_6191,N_6214);
xor U6345 (N_6345,N_6193,N_6089);
nor U6346 (N_6346,N_6007,N_6055);
nand U6347 (N_6347,N_6235,N_6189);
xnor U6348 (N_6348,N_6162,N_6084);
nand U6349 (N_6349,N_6121,N_6023);
or U6350 (N_6350,N_6138,N_6203);
or U6351 (N_6351,N_6154,N_6115);
nand U6352 (N_6352,N_6159,N_6248);
nor U6353 (N_6353,N_6200,N_6225);
or U6354 (N_6354,N_6068,N_6228);
nor U6355 (N_6355,N_6033,N_6036);
xnor U6356 (N_6356,N_6170,N_6021);
nor U6357 (N_6357,N_6143,N_6081);
nor U6358 (N_6358,N_6199,N_6058);
nand U6359 (N_6359,N_6018,N_6118);
nand U6360 (N_6360,N_6091,N_6237);
xnor U6361 (N_6361,N_6146,N_6108);
nor U6362 (N_6362,N_6207,N_6224);
or U6363 (N_6363,N_6140,N_6234);
xor U6364 (N_6364,N_6017,N_6124);
and U6365 (N_6365,N_6150,N_6088);
or U6366 (N_6366,N_6240,N_6056);
xor U6367 (N_6367,N_6044,N_6239);
xnor U6368 (N_6368,N_6086,N_6204);
nor U6369 (N_6369,N_6059,N_6163);
nand U6370 (N_6370,N_6218,N_6130);
or U6371 (N_6371,N_6177,N_6192);
and U6372 (N_6372,N_6230,N_6016);
nand U6373 (N_6373,N_6126,N_6165);
or U6374 (N_6374,N_6076,N_6092);
nand U6375 (N_6375,N_6038,N_6190);
or U6376 (N_6376,N_6015,N_6216);
nor U6377 (N_6377,N_6020,N_6235);
or U6378 (N_6378,N_6161,N_6182);
xor U6379 (N_6379,N_6247,N_6063);
nor U6380 (N_6380,N_6234,N_6001);
nor U6381 (N_6381,N_6009,N_6166);
and U6382 (N_6382,N_6043,N_6144);
or U6383 (N_6383,N_6178,N_6033);
xor U6384 (N_6384,N_6002,N_6120);
or U6385 (N_6385,N_6095,N_6128);
xor U6386 (N_6386,N_6060,N_6202);
xor U6387 (N_6387,N_6228,N_6202);
xnor U6388 (N_6388,N_6204,N_6178);
nor U6389 (N_6389,N_6084,N_6189);
or U6390 (N_6390,N_6083,N_6162);
or U6391 (N_6391,N_6124,N_6201);
xor U6392 (N_6392,N_6155,N_6175);
and U6393 (N_6393,N_6087,N_6234);
or U6394 (N_6394,N_6030,N_6163);
or U6395 (N_6395,N_6223,N_6045);
or U6396 (N_6396,N_6071,N_6176);
or U6397 (N_6397,N_6132,N_6134);
nand U6398 (N_6398,N_6193,N_6011);
or U6399 (N_6399,N_6068,N_6039);
or U6400 (N_6400,N_6148,N_6169);
nand U6401 (N_6401,N_6092,N_6067);
or U6402 (N_6402,N_6077,N_6121);
xor U6403 (N_6403,N_6046,N_6242);
or U6404 (N_6404,N_6211,N_6115);
nor U6405 (N_6405,N_6243,N_6103);
nor U6406 (N_6406,N_6211,N_6034);
and U6407 (N_6407,N_6057,N_6179);
or U6408 (N_6408,N_6089,N_6048);
and U6409 (N_6409,N_6142,N_6153);
or U6410 (N_6410,N_6111,N_6085);
nand U6411 (N_6411,N_6076,N_6097);
nor U6412 (N_6412,N_6236,N_6104);
xor U6413 (N_6413,N_6102,N_6175);
and U6414 (N_6414,N_6015,N_6039);
nand U6415 (N_6415,N_6109,N_6081);
nand U6416 (N_6416,N_6093,N_6143);
and U6417 (N_6417,N_6119,N_6042);
nand U6418 (N_6418,N_6220,N_6204);
or U6419 (N_6419,N_6219,N_6180);
xnor U6420 (N_6420,N_6143,N_6088);
nand U6421 (N_6421,N_6214,N_6081);
or U6422 (N_6422,N_6081,N_6127);
nor U6423 (N_6423,N_6175,N_6050);
and U6424 (N_6424,N_6078,N_6075);
and U6425 (N_6425,N_6127,N_6032);
nor U6426 (N_6426,N_6184,N_6100);
or U6427 (N_6427,N_6209,N_6103);
nor U6428 (N_6428,N_6065,N_6230);
or U6429 (N_6429,N_6225,N_6197);
nand U6430 (N_6430,N_6216,N_6105);
xnor U6431 (N_6431,N_6130,N_6141);
nand U6432 (N_6432,N_6146,N_6064);
nor U6433 (N_6433,N_6152,N_6222);
and U6434 (N_6434,N_6203,N_6238);
or U6435 (N_6435,N_6158,N_6234);
nor U6436 (N_6436,N_6231,N_6050);
nand U6437 (N_6437,N_6076,N_6043);
xnor U6438 (N_6438,N_6214,N_6069);
nand U6439 (N_6439,N_6170,N_6204);
or U6440 (N_6440,N_6242,N_6078);
nand U6441 (N_6441,N_6046,N_6008);
nand U6442 (N_6442,N_6020,N_6025);
nand U6443 (N_6443,N_6130,N_6043);
nor U6444 (N_6444,N_6245,N_6181);
nor U6445 (N_6445,N_6080,N_6231);
or U6446 (N_6446,N_6004,N_6148);
or U6447 (N_6447,N_6077,N_6221);
nor U6448 (N_6448,N_6099,N_6152);
or U6449 (N_6449,N_6146,N_6202);
or U6450 (N_6450,N_6084,N_6202);
or U6451 (N_6451,N_6097,N_6138);
and U6452 (N_6452,N_6187,N_6027);
and U6453 (N_6453,N_6171,N_6154);
nor U6454 (N_6454,N_6087,N_6132);
xnor U6455 (N_6455,N_6059,N_6120);
nor U6456 (N_6456,N_6226,N_6128);
and U6457 (N_6457,N_6129,N_6155);
and U6458 (N_6458,N_6208,N_6121);
xnor U6459 (N_6459,N_6203,N_6003);
or U6460 (N_6460,N_6249,N_6212);
or U6461 (N_6461,N_6045,N_6195);
nor U6462 (N_6462,N_6207,N_6220);
nand U6463 (N_6463,N_6038,N_6216);
and U6464 (N_6464,N_6008,N_6036);
and U6465 (N_6465,N_6229,N_6202);
xor U6466 (N_6466,N_6207,N_6116);
nor U6467 (N_6467,N_6132,N_6191);
or U6468 (N_6468,N_6241,N_6022);
or U6469 (N_6469,N_6116,N_6245);
nand U6470 (N_6470,N_6122,N_6172);
and U6471 (N_6471,N_6126,N_6007);
nor U6472 (N_6472,N_6000,N_6073);
nor U6473 (N_6473,N_6205,N_6120);
xnor U6474 (N_6474,N_6041,N_6066);
and U6475 (N_6475,N_6003,N_6053);
xor U6476 (N_6476,N_6115,N_6079);
and U6477 (N_6477,N_6123,N_6111);
and U6478 (N_6478,N_6190,N_6049);
or U6479 (N_6479,N_6199,N_6013);
and U6480 (N_6480,N_6105,N_6052);
or U6481 (N_6481,N_6096,N_6025);
nor U6482 (N_6482,N_6176,N_6098);
xnor U6483 (N_6483,N_6220,N_6185);
and U6484 (N_6484,N_6216,N_6052);
xor U6485 (N_6485,N_6186,N_6183);
nor U6486 (N_6486,N_6112,N_6163);
or U6487 (N_6487,N_6177,N_6016);
nand U6488 (N_6488,N_6237,N_6098);
nand U6489 (N_6489,N_6151,N_6003);
xor U6490 (N_6490,N_6123,N_6205);
and U6491 (N_6491,N_6191,N_6097);
or U6492 (N_6492,N_6193,N_6143);
and U6493 (N_6493,N_6014,N_6249);
nand U6494 (N_6494,N_6103,N_6155);
and U6495 (N_6495,N_6084,N_6147);
xnor U6496 (N_6496,N_6118,N_6004);
nand U6497 (N_6497,N_6057,N_6089);
nand U6498 (N_6498,N_6038,N_6018);
xor U6499 (N_6499,N_6090,N_6022);
or U6500 (N_6500,N_6435,N_6446);
and U6501 (N_6501,N_6377,N_6499);
nor U6502 (N_6502,N_6302,N_6402);
and U6503 (N_6503,N_6343,N_6314);
and U6504 (N_6504,N_6409,N_6347);
nand U6505 (N_6505,N_6283,N_6386);
and U6506 (N_6506,N_6296,N_6408);
xor U6507 (N_6507,N_6394,N_6481);
or U6508 (N_6508,N_6256,N_6321);
nand U6509 (N_6509,N_6274,N_6483);
nor U6510 (N_6510,N_6310,N_6259);
or U6511 (N_6511,N_6484,N_6361);
xor U6512 (N_6512,N_6278,N_6497);
or U6513 (N_6513,N_6280,N_6311);
or U6514 (N_6514,N_6488,N_6273);
nor U6515 (N_6515,N_6352,N_6493);
xnor U6516 (N_6516,N_6385,N_6270);
nor U6517 (N_6517,N_6475,N_6458);
or U6518 (N_6518,N_6448,N_6287);
nor U6519 (N_6519,N_6258,N_6348);
nor U6520 (N_6520,N_6353,N_6396);
and U6521 (N_6521,N_6350,N_6495);
nor U6522 (N_6522,N_6308,N_6404);
and U6523 (N_6523,N_6260,N_6468);
xnor U6524 (N_6524,N_6395,N_6432);
and U6525 (N_6525,N_6438,N_6331);
xor U6526 (N_6526,N_6370,N_6410);
xnor U6527 (N_6527,N_6338,N_6285);
xnor U6528 (N_6528,N_6316,N_6471);
and U6529 (N_6529,N_6469,N_6452);
xnor U6530 (N_6530,N_6427,N_6426);
nand U6531 (N_6531,N_6436,N_6450);
nand U6532 (N_6532,N_6263,N_6418);
xor U6533 (N_6533,N_6267,N_6306);
and U6534 (N_6534,N_6362,N_6384);
and U6535 (N_6535,N_6365,N_6463);
nor U6536 (N_6536,N_6332,N_6276);
or U6537 (N_6537,N_6367,N_6466);
xor U6538 (N_6538,N_6369,N_6425);
and U6539 (N_6539,N_6320,N_6455);
or U6540 (N_6540,N_6485,N_6428);
nor U6541 (N_6541,N_6312,N_6376);
nor U6542 (N_6542,N_6407,N_6307);
nor U6543 (N_6543,N_6324,N_6313);
or U6544 (N_6544,N_6295,N_6378);
or U6545 (N_6545,N_6470,N_6303);
and U6546 (N_6546,N_6292,N_6490);
and U6547 (N_6547,N_6337,N_6429);
nand U6548 (N_6548,N_6329,N_6477);
and U6549 (N_6549,N_6380,N_6393);
and U6550 (N_6550,N_6373,N_6299);
xor U6551 (N_6551,N_6264,N_6336);
xor U6552 (N_6552,N_6462,N_6434);
nor U6553 (N_6553,N_6492,N_6479);
xor U6554 (N_6554,N_6326,N_6439);
or U6555 (N_6555,N_6460,N_6279);
nor U6556 (N_6556,N_6251,N_6366);
nand U6557 (N_6557,N_6482,N_6412);
xor U6558 (N_6558,N_6375,N_6415);
xnor U6559 (N_6559,N_6417,N_6431);
nor U6560 (N_6560,N_6391,N_6355);
xnor U6561 (N_6561,N_6345,N_6357);
nand U6562 (N_6562,N_6453,N_6289);
and U6563 (N_6563,N_6486,N_6437);
or U6564 (N_6564,N_6322,N_6489);
nor U6565 (N_6565,N_6464,N_6383);
nand U6566 (N_6566,N_6291,N_6403);
or U6567 (N_6567,N_6317,N_6456);
nand U6568 (N_6568,N_6480,N_6416);
nor U6569 (N_6569,N_6420,N_6271);
nand U6570 (N_6570,N_6398,N_6282);
xor U6571 (N_6571,N_6253,N_6405);
or U6572 (N_6572,N_6359,N_6340);
nor U6573 (N_6573,N_6298,N_6356);
xor U6574 (N_6574,N_6265,N_6284);
and U6575 (N_6575,N_6358,N_6318);
xnor U6576 (N_6576,N_6319,N_6364);
nand U6577 (N_6577,N_6390,N_6309);
nand U6578 (N_6578,N_6371,N_6281);
or U6579 (N_6579,N_6254,N_6323);
nor U6580 (N_6580,N_6419,N_6277);
or U6581 (N_6581,N_6257,N_6443);
nor U6582 (N_6582,N_6328,N_6304);
xnor U6583 (N_6583,N_6440,N_6411);
and U6584 (N_6584,N_6447,N_6368);
and U6585 (N_6585,N_6294,N_6387);
xnor U6586 (N_6586,N_6444,N_6255);
nand U6587 (N_6587,N_6451,N_6334);
xnor U6588 (N_6588,N_6433,N_6413);
xnor U6589 (N_6589,N_6297,N_6467);
nor U6590 (N_6590,N_6250,N_6252);
and U6591 (N_6591,N_6382,N_6293);
nor U6592 (N_6592,N_6454,N_6354);
and U6593 (N_6593,N_6459,N_6478);
xor U6594 (N_6594,N_6339,N_6430);
and U6595 (N_6595,N_6494,N_6423);
nor U6596 (N_6596,N_6275,N_6487);
xor U6597 (N_6597,N_6379,N_6290);
nand U6598 (N_6598,N_6392,N_6341);
or U6599 (N_6599,N_6421,N_6465);
xor U6600 (N_6600,N_6476,N_6330);
or U6601 (N_6601,N_6442,N_6335);
nor U6602 (N_6602,N_6300,N_6288);
nor U6603 (N_6603,N_6406,N_6325);
and U6604 (N_6604,N_6397,N_6388);
nand U6605 (N_6605,N_6445,N_6498);
xnor U6606 (N_6606,N_6400,N_6333);
xor U6607 (N_6607,N_6315,N_6449);
and U6608 (N_6608,N_6363,N_6381);
or U6609 (N_6609,N_6424,N_6457);
nand U6610 (N_6610,N_6344,N_6342);
nand U6611 (N_6611,N_6262,N_6473);
and U6612 (N_6612,N_6269,N_6414);
and U6613 (N_6613,N_6372,N_6360);
or U6614 (N_6614,N_6305,N_6401);
xor U6615 (N_6615,N_6286,N_6374);
or U6616 (N_6616,N_6268,N_6261);
or U6617 (N_6617,N_6327,N_6472);
nand U6618 (N_6618,N_6266,N_6346);
or U6619 (N_6619,N_6441,N_6349);
xnor U6620 (N_6620,N_6301,N_6351);
xor U6621 (N_6621,N_6474,N_6422);
xnor U6622 (N_6622,N_6399,N_6491);
xnor U6623 (N_6623,N_6496,N_6461);
or U6624 (N_6624,N_6389,N_6272);
xnor U6625 (N_6625,N_6437,N_6461);
and U6626 (N_6626,N_6299,N_6489);
and U6627 (N_6627,N_6309,N_6489);
and U6628 (N_6628,N_6434,N_6346);
or U6629 (N_6629,N_6416,N_6352);
nor U6630 (N_6630,N_6455,N_6388);
xor U6631 (N_6631,N_6264,N_6265);
or U6632 (N_6632,N_6409,N_6475);
and U6633 (N_6633,N_6418,N_6354);
nand U6634 (N_6634,N_6394,N_6336);
xnor U6635 (N_6635,N_6468,N_6462);
nor U6636 (N_6636,N_6309,N_6284);
nand U6637 (N_6637,N_6327,N_6335);
xnor U6638 (N_6638,N_6279,N_6482);
nor U6639 (N_6639,N_6272,N_6284);
nand U6640 (N_6640,N_6251,N_6257);
xor U6641 (N_6641,N_6268,N_6338);
or U6642 (N_6642,N_6300,N_6253);
xnor U6643 (N_6643,N_6275,N_6494);
or U6644 (N_6644,N_6289,N_6451);
nor U6645 (N_6645,N_6320,N_6251);
nand U6646 (N_6646,N_6351,N_6417);
or U6647 (N_6647,N_6322,N_6255);
nand U6648 (N_6648,N_6256,N_6472);
and U6649 (N_6649,N_6375,N_6436);
xor U6650 (N_6650,N_6445,N_6424);
xor U6651 (N_6651,N_6272,N_6470);
nand U6652 (N_6652,N_6355,N_6289);
or U6653 (N_6653,N_6466,N_6350);
xnor U6654 (N_6654,N_6376,N_6343);
xor U6655 (N_6655,N_6356,N_6465);
and U6656 (N_6656,N_6304,N_6342);
or U6657 (N_6657,N_6256,N_6376);
nor U6658 (N_6658,N_6370,N_6491);
or U6659 (N_6659,N_6346,N_6413);
and U6660 (N_6660,N_6465,N_6254);
or U6661 (N_6661,N_6366,N_6385);
xnor U6662 (N_6662,N_6478,N_6428);
or U6663 (N_6663,N_6277,N_6337);
nand U6664 (N_6664,N_6404,N_6466);
or U6665 (N_6665,N_6397,N_6477);
and U6666 (N_6666,N_6481,N_6250);
and U6667 (N_6667,N_6368,N_6468);
nand U6668 (N_6668,N_6396,N_6453);
or U6669 (N_6669,N_6398,N_6322);
nor U6670 (N_6670,N_6388,N_6359);
and U6671 (N_6671,N_6313,N_6339);
or U6672 (N_6672,N_6324,N_6303);
and U6673 (N_6673,N_6411,N_6428);
or U6674 (N_6674,N_6377,N_6354);
nor U6675 (N_6675,N_6349,N_6396);
xnor U6676 (N_6676,N_6420,N_6310);
or U6677 (N_6677,N_6375,N_6251);
xnor U6678 (N_6678,N_6477,N_6382);
nor U6679 (N_6679,N_6361,N_6427);
nor U6680 (N_6680,N_6256,N_6455);
nand U6681 (N_6681,N_6469,N_6432);
or U6682 (N_6682,N_6432,N_6325);
or U6683 (N_6683,N_6412,N_6445);
and U6684 (N_6684,N_6290,N_6486);
nand U6685 (N_6685,N_6276,N_6465);
nand U6686 (N_6686,N_6451,N_6312);
and U6687 (N_6687,N_6484,N_6381);
and U6688 (N_6688,N_6303,N_6461);
nand U6689 (N_6689,N_6375,N_6309);
or U6690 (N_6690,N_6343,N_6381);
xnor U6691 (N_6691,N_6342,N_6333);
nand U6692 (N_6692,N_6450,N_6452);
xnor U6693 (N_6693,N_6426,N_6300);
nor U6694 (N_6694,N_6488,N_6461);
and U6695 (N_6695,N_6325,N_6378);
or U6696 (N_6696,N_6383,N_6409);
xor U6697 (N_6697,N_6284,N_6351);
or U6698 (N_6698,N_6464,N_6255);
nand U6699 (N_6699,N_6280,N_6356);
nor U6700 (N_6700,N_6312,N_6484);
and U6701 (N_6701,N_6346,N_6308);
xor U6702 (N_6702,N_6488,N_6294);
nand U6703 (N_6703,N_6336,N_6485);
nor U6704 (N_6704,N_6311,N_6453);
xnor U6705 (N_6705,N_6403,N_6324);
nor U6706 (N_6706,N_6287,N_6301);
xnor U6707 (N_6707,N_6343,N_6334);
nand U6708 (N_6708,N_6416,N_6479);
xnor U6709 (N_6709,N_6449,N_6340);
and U6710 (N_6710,N_6469,N_6349);
or U6711 (N_6711,N_6444,N_6485);
xor U6712 (N_6712,N_6289,N_6398);
nand U6713 (N_6713,N_6456,N_6329);
or U6714 (N_6714,N_6338,N_6434);
nand U6715 (N_6715,N_6417,N_6255);
nand U6716 (N_6716,N_6299,N_6403);
or U6717 (N_6717,N_6326,N_6493);
nand U6718 (N_6718,N_6359,N_6474);
xor U6719 (N_6719,N_6469,N_6279);
xor U6720 (N_6720,N_6272,N_6425);
or U6721 (N_6721,N_6355,N_6276);
xnor U6722 (N_6722,N_6397,N_6350);
nor U6723 (N_6723,N_6394,N_6499);
xor U6724 (N_6724,N_6390,N_6427);
nor U6725 (N_6725,N_6258,N_6455);
nand U6726 (N_6726,N_6252,N_6469);
and U6727 (N_6727,N_6457,N_6306);
nor U6728 (N_6728,N_6471,N_6389);
or U6729 (N_6729,N_6333,N_6336);
and U6730 (N_6730,N_6305,N_6474);
nor U6731 (N_6731,N_6279,N_6480);
xnor U6732 (N_6732,N_6299,N_6273);
nor U6733 (N_6733,N_6278,N_6263);
and U6734 (N_6734,N_6290,N_6436);
or U6735 (N_6735,N_6366,N_6299);
xor U6736 (N_6736,N_6355,N_6419);
or U6737 (N_6737,N_6383,N_6375);
xnor U6738 (N_6738,N_6251,N_6421);
nor U6739 (N_6739,N_6263,N_6463);
or U6740 (N_6740,N_6403,N_6327);
xor U6741 (N_6741,N_6300,N_6287);
and U6742 (N_6742,N_6398,N_6267);
xnor U6743 (N_6743,N_6301,N_6436);
nand U6744 (N_6744,N_6397,N_6411);
xor U6745 (N_6745,N_6410,N_6284);
xor U6746 (N_6746,N_6366,N_6290);
and U6747 (N_6747,N_6445,N_6359);
and U6748 (N_6748,N_6365,N_6319);
and U6749 (N_6749,N_6311,N_6438);
nand U6750 (N_6750,N_6690,N_6558);
nor U6751 (N_6751,N_6706,N_6749);
nor U6752 (N_6752,N_6592,N_6631);
nand U6753 (N_6753,N_6669,N_6704);
nand U6754 (N_6754,N_6716,N_6730);
or U6755 (N_6755,N_6526,N_6542);
xor U6756 (N_6756,N_6667,N_6637);
nand U6757 (N_6757,N_6519,N_6696);
and U6758 (N_6758,N_6737,N_6710);
xor U6759 (N_6759,N_6747,N_6682);
nand U6760 (N_6760,N_6693,N_6717);
or U6761 (N_6761,N_6654,N_6650);
and U6762 (N_6762,N_6613,N_6722);
and U6763 (N_6763,N_6534,N_6676);
and U6764 (N_6764,N_6680,N_6507);
nor U6765 (N_6765,N_6744,N_6570);
nand U6766 (N_6766,N_6614,N_6608);
or U6767 (N_6767,N_6646,N_6617);
nand U6768 (N_6768,N_6713,N_6549);
nand U6769 (N_6769,N_6635,N_6621);
xnor U6770 (N_6770,N_6538,N_6579);
and U6771 (N_6771,N_6514,N_6531);
nand U6772 (N_6772,N_6515,N_6520);
nand U6773 (N_6773,N_6603,N_6639);
nor U6774 (N_6774,N_6628,N_6528);
nand U6775 (N_6775,N_6633,N_6705);
or U6776 (N_6776,N_6670,N_6575);
xnor U6777 (N_6777,N_6529,N_6523);
nand U6778 (N_6778,N_6723,N_6642);
nor U6779 (N_6779,N_6544,N_6552);
and U6780 (N_6780,N_6721,N_6697);
xnor U6781 (N_6781,N_6658,N_6606);
or U6782 (N_6782,N_6521,N_6594);
nand U6783 (N_6783,N_6535,N_6695);
and U6784 (N_6784,N_6708,N_6677);
nand U6785 (N_6785,N_6576,N_6691);
or U6786 (N_6786,N_6591,N_6665);
xor U6787 (N_6787,N_6699,N_6698);
nor U6788 (N_6788,N_6580,N_6601);
nand U6789 (N_6789,N_6636,N_6733);
or U6790 (N_6790,N_6539,N_6609);
nand U6791 (N_6791,N_6584,N_6571);
and U6792 (N_6792,N_6743,N_6746);
nor U6793 (N_6793,N_6707,N_6545);
xor U6794 (N_6794,N_6555,N_6605);
or U6795 (N_6795,N_6562,N_6626);
or U6796 (N_6796,N_6574,N_6648);
and U6797 (N_6797,N_6745,N_6687);
xor U6798 (N_6798,N_6593,N_6551);
xnor U6799 (N_6799,N_6709,N_6662);
nand U6800 (N_6800,N_6663,N_6511);
nor U6801 (N_6801,N_6681,N_6503);
nand U6802 (N_6802,N_6727,N_6632);
xnor U6803 (N_6803,N_6596,N_6627);
or U6804 (N_6804,N_6728,N_6556);
or U6805 (N_6805,N_6530,N_6666);
nand U6806 (N_6806,N_6683,N_6590);
nor U6807 (N_6807,N_6547,N_6563);
and U6808 (N_6808,N_6715,N_6711);
nand U6809 (N_6809,N_6583,N_6600);
or U6810 (N_6810,N_6684,N_6537);
or U6811 (N_6811,N_6572,N_6573);
nand U6812 (N_6812,N_6561,N_6550);
and U6813 (N_6813,N_6527,N_6712);
and U6814 (N_6814,N_6700,N_6504);
nor U6815 (N_6815,N_6647,N_6714);
nor U6816 (N_6816,N_6597,N_6588);
or U6817 (N_6817,N_6578,N_6501);
and U6818 (N_6818,N_6585,N_6599);
and U6819 (N_6819,N_6587,N_6702);
nor U6820 (N_6820,N_6732,N_6565);
nor U6821 (N_6821,N_6622,N_6689);
xnor U6822 (N_6822,N_6739,N_6688);
xor U6823 (N_6823,N_6612,N_6672);
and U6824 (N_6824,N_6736,N_6741);
nor U6825 (N_6825,N_6510,N_6577);
nor U6826 (N_6826,N_6540,N_6657);
xnor U6827 (N_6827,N_6505,N_6671);
nor U6828 (N_6828,N_6624,N_6701);
or U6829 (N_6829,N_6655,N_6607);
or U6830 (N_6830,N_6512,N_6634);
and U6831 (N_6831,N_6649,N_6500);
xor U6832 (N_6832,N_6586,N_6641);
nor U6833 (N_6833,N_6735,N_6566);
xnor U6834 (N_6834,N_6568,N_6543);
nand U6835 (N_6835,N_6652,N_6525);
and U6836 (N_6836,N_6625,N_6731);
nor U6837 (N_6837,N_6725,N_6560);
nand U6838 (N_6838,N_6619,N_6623);
nor U6839 (N_6839,N_6738,N_6589);
and U6840 (N_6840,N_6651,N_6640);
and U6841 (N_6841,N_6615,N_6644);
or U6842 (N_6842,N_6653,N_6679);
nor U6843 (N_6843,N_6581,N_6630);
or U6844 (N_6844,N_6734,N_6719);
and U6845 (N_6845,N_6508,N_6694);
nor U6846 (N_6846,N_6692,N_6569);
xor U6847 (N_6847,N_6610,N_6602);
nand U6848 (N_6848,N_6748,N_6518);
xnor U6849 (N_6849,N_6673,N_6638);
nor U6850 (N_6850,N_6506,N_6598);
nand U6851 (N_6851,N_6685,N_6686);
xnor U6852 (N_6852,N_6536,N_6553);
nand U6853 (N_6853,N_6659,N_6720);
nor U6854 (N_6854,N_6532,N_6645);
nand U6855 (N_6855,N_6516,N_6740);
nand U6856 (N_6856,N_6509,N_6674);
nand U6857 (N_6857,N_6522,N_6554);
nor U6858 (N_6858,N_6567,N_6656);
xor U6859 (N_6859,N_6616,N_6660);
xor U6860 (N_6860,N_6661,N_6502);
xnor U6861 (N_6861,N_6548,N_6724);
xor U6862 (N_6862,N_6629,N_6675);
or U6863 (N_6863,N_6742,N_6557);
or U6864 (N_6864,N_6620,N_6668);
and U6865 (N_6865,N_6524,N_6541);
or U6866 (N_6866,N_6726,N_6513);
or U6867 (N_6867,N_6618,N_6664);
nand U6868 (N_6868,N_6643,N_6718);
and U6869 (N_6869,N_6678,N_6546);
xor U6870 (N_6870,N_6595,N_6517);
and U6871 (N_6871,N_6559,N_6533);
nor U6872 (N_6872,N_6703,N_6582);
nand U6873 (N_6873,N_6604,N_6564);
nor U6874 (N_6874,N_6729,N_6611);
or U6875 (N_6875,N_6588,N_6663);
and U6876 (N_6876,N_6524,N_6706);
or U6877 (N_6877,N_6733,N_6645);
xor U6878 (N_6878,N_6536,N_6674);
or U6879 (N_6879,N_6705,N_6511);
or U6880 (N_6880,N_6707,N_6584);
nand U6881 (N_6881,N_6574,N_6569);
nor U6882 (N_6882,N_6595,N_6576);
nand U6883 (N_6883,N_6624,N_6630);
xor U6884 (N_6884,N_6703,N_6507);
nor U6885 (N_6885,N_6705,N_6502);
xor U6886 (N_6886,N_6575,N_6512);
and U6887 (N_6887,N_6631,N_6550);
and U6888 (N_6888,N_6725,N_6537);
xnor U6889 (N_6889,N_6585,N_6580);
nand U6890 (N_6890,N_6657,N_6527);
and U6891 (N_6891,N_6565,N_6636);
nand U6892 (N_6892,N_6716,N_6617);
or U6893 (N_6893,N_6643,N_6722);
xnor U6894 (N_6894,N_6610,N_6512);
nand U6895 (N_6895,N_6655,N_6618);
or U6896 (N_6896,N_6721,N_6543);
xnor U6897 (N_6897,N_6588,N_6608);
nor U6898 (N_6898,N_6521,N_6629);
and U6899 (N_6899,N_6527,N_6619);
xor U6900 (N_6900,N_6515,N_6626);
nor U6901 (N_6901,N_6679,N_6677);
or U6902 (N_6902,N_6542,N_6569);
or U6903 (N_6903,N_6627,N_6590);
or U6904 (N_6904,N_6583,N_6607);
nand U6905 (N_6905,N_6618,N_6622);
and U6906 (N_6906,N_6632,N_6693);
nand U6907 (N_6907,N_6594,N_6663);
xnor U6908 (N_6908,N_6646,N_6606);
and U6909 (N_6909,N_6635,N_6535);
and U6910 (N_6910,N_6548,N_6582);
or U6911 (N_6911,N_6571,N_6533);
xor U6912 (N_6912,N_6631,N_6722);
and U6913 (N_6913,N_6537,N_6545);
nor U6914 (N_6914,N_6737,N_6607);
or U6915 (N_6915,N_6666,N_6674);
and U6916 (N_6916,N_6699,N_6737);
nand U6917 (N_6917,N_6560,N_6719);
and U6918 (N_6918,N_6701,N_6725);
nor U6919 (N_6919,N_6742,N_6744);
nor U6920 (N_6920,N_6532,N_6742);
nor U6921 (N_6921,N_6596,N_6733);
and U6922 (N_6922,N_6745,N_6593);
and U6923 (N_6923,N_6645,N_6642);
or U6924 (N_6924,N_6563,N_6721);
and U6925 (N_6925,N_6579,N_6673);
or U6926 (N_6926,N_6749,N_6529);
nor U6927 (N_6927,N_6707,N_6506);
nand U6928 (N_6928,N_6572,N_6668);
and U6929 (N_6929,N_6522,N_6561);
nor U6930 (N_6930,N_6543,N_6714);
xnor U6931 (N_6931,N_6676,N_6520);
nand U6932 (N_6932,N_6721,N_6749);
and U6933 (N_6933,N_6700,N_6675);
and U6934 (N_6934,N_6500,N_6665);
or U6935 (N_6935,N_6514,N_6646);
nand U6936 (N_6936,N_6682,N_6555);
nor U6937 (N_6937,N_6532,N_6736);
nand U6938 (N_6938,N_6728,N_6583);
and U6939 (N_6939,N_6712,N_6625);
nor U6940 (N_6940,N_6542,N_6654);
or U6941 (N_6941,N_6661,N_6612);
or U6942 (N_6942,N_6577,N_6737);
nor U6943 (N_6943,N_6654,N_6676);
nor U6944 (N_6944,N_6650,N_6610);
xnor U6945 (N_6945,N_6654,N_6552);
or U6946 (N_6946,N_6680,N_6692);
or U6947 (N_6947,N_6572,N_6519);
and U6948 (N_6948,N_6692,N_6566);
xnor U6949 (N_6949,N_6659,N_6634);
and U6950 (N_6950,N_6586,N_6531);
nand U6951 (N_6951,N_6649,N_6644);
nand U6952 (N_6952,N_6648,N_6703);
xor U6953 (N_6953,N_6710,N_6566);
xor U6954 (N_6954,N_6673,N_6623);
or U6955 (N_6955,N_6699,N_6646);
or U6956 (N_6956,N_6558,N_6651);
and U6957 (N_6957,N_6629,N_6520);
nor U6958 (N_6958,N_6511,N_6658);
and U6959 (N_6959,N_6513,N_6581);
and U6960 (N_6960,N_6593,N_6643);
and U6961 (N_6961,N_6506,N_6565);
and U6962 (N_6962,N_6512,N_6546);
nor U6963 (N_6963,N_6599,N_6520);
xnor U6964 (N_6964,N_6715,N_6652);
nand U6965 (N_6965,N_6607,N_6681);
or U6966 (N_6966,N_6527,N_6609);
and U6967 (N_6967,N_6571,N_6548);
xor U6968 (N_6968,N_6745,N_6657);
and U6969 (N_6969,N_6560,N_6703);
or U6970 (N_6970,N_6679,N_6684);
nor U6971 (N_6971,N_6647,N_6657);
and U6972 (N_6972,N_6540,N_6648);
nand U6973 (N_6973,N_6555,N_6734);
nor U6974 (N_6974,N_6620,N_6672);
or U6975 (N_6975,N_6670,N_6726);
nand U6976 (N_6976,N_6576,N_6607);
nand U6977 (N_6977,N_6737,N_6682);
and U6978 (N_6978,N_6528,N_6525);
and U6979 (N_6979,N_6694,N_6635);
or U6980 (N_6980,N_6629,N_6621);
nand U6981 (N_6981,N_6657,N_6503);
xnor U6982 (N_6982,N_6518,N_6575);
xor U6983 (N_6983,N_6592,N_6601);
and U6984 (N_6984,N_6555,N_6603);
nor U6985 (N_6985,N_6726,N_6611);
or U6986 (N_6986,N_6654,N_6500);
nor U6987 (N_6987,N_6540,N_6709);
nand U6988 (N_6988,N_6561,N_6597);
or U6989 (N_6989,N_6660,N_6658);
nor U6990 (N_6990,N_6512,N_6734);
or U6991 (N_6991,N_6602,N_6743);
or U6992 (N_6992,N_6535,N_6702);
or U6993 (N_6993,N_6728,N_6567);
and U6994 (N_6994,N_6664,N_6627);
or U6995 (N_6995,N_6648,N_6502);
nor U6996 (N_6996,N_6622,N_6537);
nand U6997 (N_6997,N_6543,N_6594);
and U6998 (N_6998,N_6701,N_6722);
or U6999 (N_6999,N_6668,N_6748);
xnor U7000 (N_7000,N_6985,N_6909);
nor U7001 (N_7001,N_6787,N_6993);
or U7002 (N_7002,N_6886,N_6793);
and U7003 (N_7003,N_6913,N_6924);
or U7004 (N_7004,N_6917,N_6914);
xnor U7005 (N_7005,N_6925,N_6973);
and U7006 (N_7006,N_6977,N_6876);
nor U7007 (N_7007,N_6858,N_6939);
nor U7008 (N_7008,N_6838,N_6966);
nor U7009 (N_7009,N_6816,N_6889);
xnor U7010 (N_7010,N_6783,N_6974);
nand U7011 (N_7011,N_6900,N_6954);
nor U7012 (N_7012,N_6775,N_6895);
xor U7013 (N_7013,N_6851,N_6807);
nand U7014 (N_7014,N_6821,N_6841);
nor U7015 (N_7015,N_6879,N_6963);
nand U7016 (N_7016,N_6881,N_6803);
xnor U7017 (N_7017,N_6996,N_6866);
and U7018 (N_7018,N_6877,N_6997);
xor U7019 (N_7019,N_6817,N_6887);
or U7020 (N_7020,N_6782,N_6947);
nor U7021 (N_7021,N_6852,N_6823);
or U7022 (N_7022,N_6897,N_6952);
nor U7023 (N_7023,N_6773,N_6916);
xnor U7024 (N_7024,N_6986,N_6761);
and U7025 (N_7025,N_6830,N_6872);
nor U7026 (N_7026,N_6883,N_6944);
and U7027 (N_7027,N_6848,N_6826);
nor U7028 (N_7028,N_6943,N_6955);
or U7029 (N_7029,N_6829,N_6839);
nand U7030 (N_7030,N_6968,N_6896);
nand U7031 (N_7031,N_6843,N_6970);
or U7032 (N_7032,N_6982,N_6796);
nand U7033 (N_7033,N_6912,N_6983);
or U7034 (N_7034,N_6878,N_6808);
or U7035 (N_7035,N_6804,N_6869);
nor U7036 (N_7036,N_6822,N_6755);
or U7037 (N_7037,N_6950,N_6791);
xor U7038 (N_7038,N_6998,N_6890);
nand U7039 (N_7039,N_6751,N_6921);
or U7040 (N_7040,N_6801,N_6906);
nand U7041 (N_7041,N_6818,N_6922);
or U7042 (N_7042,N_6972,N_6960);
and U7043 (N_7043,N_6784,N_6770);
or U7044 (N_7044,N_6828,N_6846);
nor U7045 (N_7045,N_6893,N_6976);
nor U7046 (N_7046,N_6772,N_6905);
nor U7047 (N_7047,N_6957,N_6932);
nand U7048 (N_7048,N_6812,N_6861);
nand U7049 (N_7049,N_6946,N_6915);
or U7050 (N_7050,N_6929,N_6854);
xor U7051 (N_7051,N_6813,N_6769);
nor U7052 (N_7052,N_6765,N_6989);
nand U7053 (N_7053,N_6999,N_6892);
nand U7054 (N_7054,N_6987,N_6927);
or U7055 (N_7055,N_6837,N_6857);
nand U7056 (N_7056,N_6874,N_6780);
nand U7057 (N_7057,N_6911,N_6918);
or U7058 (N_7058,N_6766,N_6820);
xnor U7059 (N_7059,N_6904,N_6862);
xor U7060 (N_7060,N_6894,N_6980);
and U7061 (N_7061,N_6819,N_6811);
and U7062 (N_7062,N_6781,N_6940);
xnor U7063 (N_7063,N_6867,N_6907);
xor U7064 (N_7064,N_6971,N_6969);
xor U7065 (N_7065,N_6774,N_6964);
or U7066 (N_7066,N_6934,N_6767);
nor U7067 (N_7067,N_6937,N_6790);
xor U7068 (N_7068,N_6938,N_6788);
or U7069 (N_7069,N_6959,N_6880);
and U7070 (N_7070,N_6975,N_6992);
and U7071 (N_7071,N_6832,N_6754);
and U7072 (N_7072,N_6865,N_6825);
nor U7073 (N_7073,N_6951,N_6991);
nor U7074 (N_7074,N_6936,N_6882);
nor U7075 (N_7075,N_6802,N_6844);
xnor U7076 (N_7076,N_6967,N_6794);
nor U7077 (N_7077,N_6923,N_6884);
nand U7078 (N_7078,N_6859,N_6776);
nand U7079 (N_7079,N_6758,N_6849);
xnor U7080 (N_7080,N_6979,N_6930);
xnor U7081 (N_7081,N_6994,N_6785);
xor U7082 (N_7082,N_6910,N_6995);
or U7083 (N_7083,N_6965,N_6863);
or U7084 (N_7084,N_6908,N_6756);
xnor U7085 (N_7085,N_6831,N_6786);
xnor U7086 (N_7086,N_6833,N_6958);
nand U7087 (N_7087,N_6827,N_6805);
nor U7088 (N_7088,N_6888,N_6864);
nand U7089 (N_7089,N_6945,N_6806);
or U7090 (N_7090,N_6856,N_6873);
and U7091 (N_7091,N_6752,N_6764);
and U7092 (N_7092,N_6860,N_6903);
or U7093 (N_7093,N_6953,N_6779);
nor U7094 (N_7094,N_6836,N_6981);
nand U7095 (N_7095,N_6920,N_6926);
nand U7096 (N_7096,N_6797,N_6789);
and U7097 (N_7097,N_6935,N_6902);
nand U7098 (N_7098,N_6948,N_6809);
nor U7099 (N_7099,N_6899,N_6810);
xor U7100 (N_7100,N_6928,N_6753);
nor U7101 (N_7101,N_6799,N_6795);
nor U7102 (N_7102,N_6798,N_6792);
and U7103 (N_7103,N_6949,N_6824);
and U7104 (N_7104,N_6842,N_6763);
or U7105 (N_7105,N_6757,N_6871);
nor U7106 (N_7106,N_6962,N_6778);
xnor U7107 (N_7107,N_6941,N_6875);
xnor U7108 (N_7108,N_6847,N_6850);
or U7109 (N_7109,N_6759,N_6885);
or U7110 (N_7110,N_6870,N_6855);
and U7111 (N_7111,N_6956,N_6933);
nand U7112 (N_7112,N_6834,N_6961);
and U7113 (N_7113,N_6777,N_6800);
nand U7114 (N_7114,N_6760,N_6750);
nand U7115 (N_7115,N_6771,N_6898);
nor U7116 (N_7116,N_6931,N_6901);
xnor U7117 (N_7117,N_6868,N_6919);
or U7118 (N_7118,N_6990,N_6942);
or U7119 (N_7119,N_6815,N_6845);
nand U7120 (N_7120,N_6768,N_6835);
nand U7121 (N_7121,N_6978,N_6853);
xnor U7122 (N_7122,N_6840,N_6984);
nand U7123 (N_7123,N_6814,N_6891);
and U7124 (N_7124,N_6988,N_6762);
nor U7125 (N_7125,N_6998,N_6948);
xnor U7126 (N_7126,N_6926,N_6781);
and U7127 (N_7127,N_6827,N_6911);
nand U7128 (N_7128,N_6778,N_6888);
nor U7129 (N_7129,N_6834,N_6783);
nand U7130 (N_7130,N_6888,N_6769);
xor U7131 (N_7131,N_6878,N_6939);
nand U7132 (N_7132,N_6750,N_6802);
nand U7133 (N_7133,N_6774,N_6905);
and U7134 (N_7134,N_6999,N_6820);
nor U7135 (N_7135,N_6833,N_6775);
nor U7136 (N_7136,N_6991,N_6992);
and U7137 (N_7137,N_6896,N_6914);
and U7138 (N_7138,N_6798,N_6789);
and U7139 (N_7139,N_6921,N_6881);
nor U7140 (N_7140,N_6759,N_6952);
nor U7141 (N_7141,N_6896,N_6811);
or U7142 (N_7142,N_6932,N_6931);
or U7143 (N_7143,N_6972,N_6997);
xor U7144 (N_7144,N_6857,N_6788);
or U7145 (N_7145,N_6827,N_6841);
or U7146 (N_7146,N_6785,N_6828);
and U7147 (N_7147,N_6802,N_6845);
or U7148 (N_7148,N_6788,N_6955);
and U7149 (N_7149,N_6890,N_6820);
nand U7150 (N_7150,N_6968,N_6998);
nand U7151 (N_7151,N_6780,N_6913);
nor U7152 (N_7152,N_6897,N_6875);
or U7153 (N_7153,N_6844,N_6862);
and U7154 (N_7154,N_6898,N_6936);
nor U7155 (N_7155,N_6789,N_6916);
xnor U7156 (N_7156,N_6852,N_6831);
or U7157 (N_7157,N_6810,N_6841);
nor U7158 (N_7158,N_6926,N_6842);
xor U7159 (N_7159,N_6765,N_6900);
nand U7160 (N_7160,N_6854,N_6940);
nand U7161 (N_7161,N_6969,N_6750);
nor U7162 (N_7162,N_6804,N_6772);
xnor U7163 (N_7163,N_6937,N_6767);
nor U7164 (N_7164,N_6980,N_6819);
nand U7165 (N_7165,N_6928,N_6960);
and U7166 (N_7166,N_6908,N_6958);
or U7167 (N_7167,N_6889,N_6762);
nor U7168 (N_7168,N_6799,N_6837);
and U7169 (N_7169,N_6816,N_6918);
or U7170 (N_7170,N_6975,N_6753);
and U7171 (N_7171,N_6890,N_6778);
xor U7172 (N_7172,N_6992,N_6787);
nand U7173 (N_7173,N_6855,N_6781);
nand U7174 (N_7174,N_6865,N_6785);
nand U7175 (N_7175,N_6756,N_6840);
xnor U7176 (N_7176,N_6755,N_6973);
and U7177 (N_7177,N_6984,N_6856);
nor U7178 (N_7178,N_6847,N_6787);
and U7179 (N_7179,N_6911,N_6891);
xor U7180 (N_7180,N_6823,N_6796);
or U7181 (N_7181,N_6785,N_6840);
nand U7182 (N_7182,N_6939,N_6968);
nor U7183 (N_7183,N_6941,N_6764);
nand U7184 (N_7184,N_6842,N_6933);
xnor U7185 (N_7185,N_6995,N_6913);
nand U7186 (N_7186,N_6832,N_6808);
and U7187 (N_7187,N_6885,N_6939);
xnor U7188 (N_7188,N_6999,N_6836);
and U7189 (N_7189,N_6890,N_6856);
xor U7190 (N_7190,N_6949,N_6945);
or U7191 (N_7191,N_6921,N_6809);
nor U7192 (N_7192,N_6793,N_6891);
and U7193 (N_7193,N_6933,N_6954);
xnor U7194 (N_7194,N_6872,N_6843);
xnor U7195 (N_7195,N_6973,N_6963);
nor U7196 (N_7196,N_6996,N_6910);
nor U7197 (N_7197,N_6911,N_6767);
and U7198 (N_7198,N_6833,N_6934);
xor U7199 (N_7199,N_6862,N_6830);
xnor U7200 (N_7200,N_6878,N_6804);
xnor U7201 (N_7201,N_6964,N_6844);
or U7202 (N_7202,N_6767,N_6831);
nand U7203 (N_7203,N_6907,N_6991);
nor U7204 (N_7204,N_6757,N_6886);
nor U7205 (N_7205,N_6808,N_6970);
nand U7206 (N_7206,N_6764,N_6848);
nand U7207 (N_7207,N_6922,N_6869);
and U7208 (N_7208,N_6962,N_6966);
xor U7209 (N_7209,N_6763,N_6899);
nor U7210 (N_7210,N_6750,N_6860);
nor U7211 (N_7211,N_6975,N_6982);
nand U7212 (N_7212,N_6914,N_6817);
nor U7213 (N_7213,N_6799,N_6880);
and U7214 (N_7214,N_6965,N_6927);
and U7215 (N_7215,N_6840,N_6954);
or U7216 (N_7216,N_6778,N_6828);
xor U7217 (N_7217,N_6997,N_6894);
or U7218 (N_7218,N_6779,N_6806);
or U7219 (N_7219,N_6912,N_6754);
or U7220 (N_7220,N_6931,N_6854);
and U7221 (N_7221,N_6965,N_6901);
xnor U7222 (N_7222,N_6923,N_6858);
and U7223 (N_7223,N_6761,N_6966);
and U7224 (N_7224,N_6777,N_6954);
nor U7225 (N_7225,N_6851,N_6894);
nand U7226 (N_7226,N_6954,N_6977);
or U7227 (N_7227,N_6845,N_6902);
and U7228 (N_7228,N_6961,N_6751);
and U7229 (N_7229,N_6850,N_6794);
nor U7230 (N_7230,N_6990,N_6987);
or U7231 (N_7231,N_6926,N_6872);
nor U7232 (N_7232,N_6966,N_6863);
xor U7233 (N_7233,N_6989,N_6919);
xor U7234 (N_7234,N_6966,N_6797);
and U7235 (N_7235,N_6981,N_6928);
and U7236 (N_7236,N_6949,N_6939);
nand U7237 (N_7237,N_6909,N_6842);
xor U7238 (N_7238,N_6960,N_6855);
xor U7239 (N_7239,N_6863,N_6778);
and U7240 (N_7240,N_6877,N_6952);
nand U7241 (N_7241,N_6865,N_6847);
or U7242 (N_7242,N_6815,N_6861);
or U7243 (N_7243,N_6752,N_6854);
and U7244 (N_7244,N_6914,N_6993);
xor U7245 (N_7245,N_6761,N_6840);
and U7246 (N_7246,N_6926,N_6837);
nor U7247 (N_7247,N_6922,N_6945);
xnor U7248 (N_7248,N_6756,N_6811);
nand U7249 (N_7249,N_6906,N_6759);
or U7250 (N_7250,N_7126,N_7191);
nor U7251 (N_7251,N_7090,N_7204);
xnor U7252 (N_7252,N_7249,N_7242);
nand U7253 (N_7253,N_7022,N_7089);
nor U7254 (N_7254,N_7189,N_7247);
nand U7255 (N_7255,N_7026,N_7077);
and U7256 (N_7256,N_7144,N_7131);
xnor U7257 (N_7257,N_7104,N_7074);
xor U7258 (N_7258,N_7045,N_7162);
or U7259 (N_7259,N_7155,N_7093);
nor U7260 (N_7260,N_7017,N_7086);
nor U7261 (N_7261,N_7187,N_7003);
or U7262 (N_7262,N_7206,N_7235);
and U7263 (N_7263,N_7004,N_7071);
or U7264 (N_7264,N_7152,N_7023);
xnor U7265 (N_7265,N_7073,N_7076);
nand U7266 (N_7266,N_7067,N_7112);
and U7267 (N_7267,N_7083,N_7014);
nand U7268 (N_7268,N_7222,N_7215);
and U7269 (N_7269,N_7002,N_7219);
nand U7270 (N_7270,N_7156,N_7012);
nand U7271 (N_7271,N_7185,N_7232);
xnor U7272 (N_7272,N_7122,N_7084);
xor U7273 (N_7273,N_7164,N_7005);
nand U7274 (N_7274,N_7065,N_7016);
and U7275 (N_7275,N_7226,N_7248);
and U7276 (N_7276,N_7107,N_7079);
nand U7277 (N_7277,N_7046,N_7230);
or U7278 (N_7278,N_7054,N_7060);
xor U7279 (N_7279,N_7158,N_7128);
nand U7280 (N_7280,N_7064,N_7244);
nand U7281 (N_7281,N_7062,N_7117);
nand U7282 (N_7282,N_7142,N_7019);
nor U7283 (N_7283,N_7205,N_7186);
and U7284 (N_7284,N_7211,N_7115);
nand U7285 (N_7285,N_7082,N_7029);
nor U7286 (N_7286,N_7195,N_7190);
nand U7287 (N_7287,N_7101,N_7057);
or U7288 (N_7288,N_7140,N_7085);
nand U7289 (N_7289,N_7199,N_7203);
or U7290 (N_7290,N_7143,N_7024);
nor U7291 (N_7291,N_7100,N_7137);
and U7292 (N_7292,N_7224,N_7075);
xnor U7293 (N_7293,N_7007,N_7238);
and U7294 (N_7294,N_7114,N_7092);
xnor U7295 (N_7295,N_7174,N_7037);
xor U7296 (N_7296,N_7116,N_7161);
or U7297 (N_7297,N_7183,N_7125);
nor U7298 (N_7298,N_7154,N_7123);
or U7299 (N_7299,N_7201,N_7139);
nand U7300 (N_7300,N_7127,N_7212);
nand U7301 (N_7301,N_7069,N_7000);
or U7302 (N_7302,N_7106,N_7129);
xnor U7303 (N_7303,N_7148,N_7033);
xnor U7304 (N_7304,N_7109,N_7098);
and U7305 (N_7305,N_7167,N_7216);
xor U7306 (N_7306,N_7111,N_7110);
or U7307 (N_7307,N_7095,N_7207);
or U7308 (N_7308,N_7094,N_7103);
and U7309 (N_7309,N_7170,N_7027);
xnor U7310 (N_7310,N_7202,N_7245);
nand U7311 (N_7311,N_7009,N_7243);
xnor U7312 (N_7312,N_7141,N_7061);
xnor U7313 (N_7313,N_7070,N_7041);
or U7314 (N_7314,N_7231,N_7108);
and U7315 (N_7315,N_7068,N_7192);
and U7316 (N_7316,N_7179,N_7214);
xor U7317 (N_7317,N_7229,N_7198);
and U7318 (N_7318,N_7053,N_7021);
nand U7319 (N_7319,N_7157,N_7239);
xnor U7320 (N_7320,N_7151,N_7138);
nand U7321 (N_7321,N_7088,N_7028);
nor U7322 (N_7322,N_7150,N_7047);
or U7323 (N_7323,N_7039,N_7042);
nand U7324 (N_7324,N_7113,N_7177);
nor U7325 (N_7325,N_7049,N_7124);
and U7326 (N_7326,N_7018,N_7176);
or U7327 (N_7327,N_7063,N_7080);
or U7328 (N_7328,N_7099,N_7237);
nand U7329 (N_7329,N_7119,N_7165);
nand U7330 (N_7330,N_7030,N_7130);
or U7331 (N_7331,N_7097,N_7020);
or U7332 (N_7332,N_7153,N_7163);
and U7333 (N_7333,N_7040,N_7246);
xor U7334 (N_7334,N_7001,N_7178);
xor U7335 (N_7335,N_7105,N_7036);
xor U7336 (N_7336,N_7044,N_7173);
nand U7337 (N_7337,N_7135,N_7210);
or U7338 (N_7338,N_7168,N_7056);
nand U7339 (N_7339,N_7227,N_7134);
and U7340 (N_7340,N_7149,N_7169);
xnor U7341 (N_7341,N_7121,N_7220);
and U7342 (N_7342,N_7200,N_7034);
xnor U7343 (N_7343,N_7171,N_7228);
nand U7344 (N_7344,N_7010,N_7008);
xnor U7345 (N_7345,N_7133,N_7166);
nor U7346 (N_7346,N_7043,N_7172);
nand U7347 (N_7347,N_7035,N_7182);
and U7348 (N_7348,N_7196,N_7221);
or U7349 (N_7349,N_7184,N_7120);
or U7350 (N_7350,N_7055,N_7146);
and U7351 (N_7351,N_7194,N_7132);
or U7352 (N_7352,N_7175,N_7236);
and U7353 (N_7353,N_7051,N_7136);
xor U7354 (N_7354,N_7147,N_7066);
or U7355 (N_7355,N_7096,N_7159);
or U7356 (N_7356,N_7188,N_7193);
or U7357 (N_7357,N_7081,N_7091);
and U7358 (N_7358,N_7209,N_7240);
and U7359 (N_7359,N_7160,N_7015);
xor U7360 (N_7360,N_7208,N_7197);
nor U7361 (N_7361,N_7118,N_7213);
nand U7362 (N_7362,N_7025,N_7223);
and U7363 (N_7363,N_7145,N_7052);
nand U7364 (N_7364,N_7032,N_7218);
nand U7365 (N_7365,N_7059,N_7102);
nor U7366 (N_7366,N_7058,N_7087);
or U7367 (N_7367,N_7013,N_7050);
nand U7368 (N_7368,N_7241,N_7038);
nor U7369 (N_7369,N_7180,N_7233);
or U7370 (N_7370,N_7031,N_7234);
nor U7371 (N_7371,N_7078,N_7006);
xor U7372 (N_7372,N_7011,N_7181);
and U7373 (N_7373,N_7217,N_7048);
nand U7374 (N_7374,N_7072,N_7225);
xnor U7375 (N_7375,N_7166,N_7227);
and U7376 (N_7376,N_7007,N_7235);
and U7377 (N_7377,N_7205,N_7159);
xor U7378 (N_7378,N_7081,N_7100);
nor U7379 (N_7379,N_7160,N_7085);
and U7380 (N_7380,N_7138,N_7100);
or U7381 (N_7381,N_7245,N_7087);
nand U7382 (N_7382,N_7129,N_7138);
or U7383 (N_7383,N_7072,N_7201);
or U7384 (N_7384,N_7219,N_7016);
xnor U7385 (N_7385,N_7156,N_7208);
xor U7386 (N_7386,N_7038,N_7041);
nand U7387 (N_7387,N_7203,N_7236);
and U7388 (N_7388,N_7190,N_7098);
nand U7389 (N_7389,N_7199,N_7117);
nand U7390 (N_7390,N_7033,N_7102);
nor U7391 (N_7391,N_7234,N_7141);
or U7392 (N_7392,N_7127,N_7144);
nand U7393 (N_7393,N_7029,N_7075);
nor U7394 (N_7394,N_7061,N_7045);
or U7395 (N_7395,N_7127,N_7069);
xor U7396 (N_7396,N_7039,N_7113);
xor U7397 (N_7397,N_7105,N_7249);
nand U7398 (N_7398,N_7246,N_7199);
or U7399 (N_7399,N_7235,N_7241);
xnor U7400 (N_7400,N_7166,N_7196);
nand U7401 (N_7401,N_7053,N_7073);
xnor U7402 (N_7402,N_7015,N_7071);
nor U7403 (N_7403,N_7167,N_7227);
nand U7404 (N_7404,N_7244,N_7154);
or U7405 (N_7405,N_7227,N_7073);
and U7406 (N_7406,N_7125,N_7008);
and U7407 (N_7407,N_7080,N_7043);
or U7408 (N_7408,N_7024,N_7177);
xor U7409 (N_7409,N_7173,N_7052);
xnor U7410 (N_7410,N_7139,N_7024);
xnor U7411 (N_7411,N_7001,N_7031);
nand U7412 (N_7412,N_7151,N_7114);
and U7413 (N_7413,N_7129,N_7084);
nor U7414 (N_7414,N_7143,N_7001);
xor U7415 (N_7415,N_7208,N_7086);
or U7416 (N_7416,N_7119,N_7063);
nor U7417 (N_7417,N_7216,N_7029);
nor U7418 (N_7418,N_7185,N_7046);
or U7419 (N_7419,N_7138,N_7148);
nand U7420 (N_7420,N_7046,N_7017);
or U7421 (N_7421,N_7228,N_7185);
or U7422 (N_7422,N_7115,N_7143);
or U7423 (N_7423,N_7125,N_7087);
or U7424 (N_7424,N_7193,N_7123);
nand U7425 (N_7425,N_7201,N_7059);
and U7426 (N_7426,N_7146,N_7028);
or U7427 (N_7427,N_7114,N_7055);
nand U7428 (N_7428,N_7157,N_7219);
or U7429 (N_7429,N_7174,N_7189);
or U7430 (N_7430,N_7073,N_7011);
xor U7431 (N_7431,N_7209,N_7210);
and U7432 (N_7432,N_7182,N_7086);
or U7433 (N_7433,N_7249,N_7057);
nor U7434 (N_7434,N_7147,N_7172);
xnor U7435 (N_7435,N_7224,N_7208);
or U7436 (N_7436,N_7120,N_7103);
nor U7437 (N_7437,N_7009,N_7131);
or U7438 (N_7438,N_7149,N_7233);
xor U7439 (N_7439,N_7239,N_7071);
or U7440 (N_7440,N_7225,N_7202);
or U7441 (N_7441,N_7028,N_7003);
or U7442 (N_7442,N_7207,N_7124);
and U7443 (N_7443,N_7047,N_7015);
or U7444 (N_7444,N_7153,N_7139);
nor U7445 (N_7445,N_7072,N_7157);
and U7446 (N_7446,N_7087,N_7098);
xor U7447 (N_7447,N_7158,N_7211);
nor U7448 (N_7448,N_7085,N_7145);
and U7449 (N_7449,N_7069,N_7066);
and U7450 (N_7450,N_7114,N_7145);
and U7451 (N_7451,N_7135,N_7017);
nand U7452 (N_7452,N_7071,N_7196);
or U7453 (N_7453,N_7094,N_7240);
nor U7454 (N_7454,N_7190,N_7097);
nor U7455 (N_7455,N_7244,N_7047);
nand U7456 (N_7456,N_7068,N_7163);
and U7457 (N_7457,N_7131,N_7041);
xor U7458 (N_7458,N_7246,N_7135);
or U7459 (N_7459,N_7243,N_7064);
nand U7460 (N_7460,N_7248,N_7124);
xor U7461 (N_7461,N_7080,N_7112);
xnor U7462 (N_7462,N_7154,N_7100);
xor U7463 (N_7463,N_7226,N_7234);
nor U7464 (N_7464,N_7182,N_7110);
and U7465 (N_7465,N_7110,N_7128);
xnor U7466 (N_7466,N_7180,N_7113);
or U7467 (N_7467,N_7025,N_7185);
nand U7468 (N_7468,N_7116,N_7024);
or U7469 (N_7469,N_7202,N_7228);
and U7470 (N_7470,N_7090,N_7033);
and U7471 (N_7471,N_7014,N_7113);
or U7472 (N_7472,N_7014,N_7171);
nand U7473 (N_7473,N_7042,N_7091);
nand U7474 (N_7474,N_7066,N_7071);
and U7475 (N_7475,N_7160,N_7037);
and U7476 (N_7476,N_7015,N_7208);
nor U7477 (N_7477,N_7087,N_7079);
nor U7478 (N_7478,N_7136,N_7183);
nor U7479 (N_7479,N_7168,N_7024);
and U7480 (N_7480,N_7239,N_7078);
and U7481 (N_7481,N_7121,N_7080);
nand U7482 (N_7482,N_7114,N_7030);
or U7483 (N_7483,N_7002,N_7205);
nor U7484 (N_7484,N_7101,N_7192);
nand U7485 (N_7485,N_7196,N_7029);
xor U7486 (N_7486,N_7223,N_7222);
nor U7487 (N_7487,N_7095,N_7078);
nor U7488 (N_7488,N_7060,N_7114);
nor U7489 (N_7489,N_7152,N_7119);
xor U7490 (N_7490,N_7099,N_7082);
nand U7491 (N_7491,N_7072,N_7189);
xor U7492 (N_7492,N_7227,N_7223);
xor U7493 (N_7493,N_7141,N_7226);
and U7494 (N_7494,N_7166,N_7216);
or U7495 (N_7495,N_7243,N_7039);
or U7496 (N_7496,N_7029,N_7015);
or U7497 (N_7497,N_7244,N_7102);
or U7498 (N_7498,N_7062,N_7110);
and U7499 (N_7499,N_7142,N_7237);
xor U7500 (N_7500,N_7491,N_7398);
or U7501 (N_7501,N_7262,N_7464);
or U7502 (N_7502,N_7383,N_7352);
and U7503 (N_7503,N_7393,N_7302);
nor U7504 (N_7504,N_7479,N_7328);
and U7505 (N_7505,N_7336,N_7255);
nor U7506 (N_7506,N_7317,N_7439);
nand U7507 (N_7507,N_7420,N_7409);
or U7508 (N_7508,N_7370,N_7469);
or U7509 (N_7509,N_7440,N_7446);
xnor U7510 (N_7510,N_7384,N_7364);
and U7511 (N_7511,N_7273,N_7362);
nor U7512 (N_7512,N_7371,N_7312);
xnor U7513 (N_7513,N_7458,N_7277);
or U7514 (N_7514,N_7397,N_7429);
nor U7515 (N_7515,N_7492,N_7338);
and U7516 (N_7516,N_7496,N_7379);
or U7517 (N_7517,N_7326,N_7381);
xor U7518 (N_7518,N_7291,N_7374);
nand U7519 (N_7519,N_7419,N_7426);
nand U7520 (N_7520,N_7292,N_7299);
nor U7521 (N_7521,N_7257,N_7276);
and U7522 (N_7522,N_7499,N_7319);
xnor U7523 (N_7523,N_7263,N_7261);
and U7524 (N_7524,N_7411,N_7355);
nor U7525 (N_7525,N_7349,N_7265);
or U7526 (N_7526,N_7478,N_7278);
nand U7527 (N_7527,N_7253,N_7380);
xor U7528 (N_7528,N_7417,N_7414);
nor U7529 (N_7529,N_7449,N_7477);
nor U7530 (N_7530,N_7396,N_7366);
or U7531 (N_7531,N_7467,N_7325);
nand U7532 (N_7532,N_7363,N_7268);
and U7533 (N_7533,N_7444,N_7269);
xnor U7534 (N_7534,N_7301,N_7394);
or U7535 (N_7535,N_7311,N_7475);
and U7536 (N_7536,N_7494,N_7422);
nor U7537 (N_7537,N_7388,N_7286);
nand U7538 (N_7538,N_7495,N_7450);
nand U7539 (N_7539,N_7314,N_7421);
xnor U7540 (N_7540,N_7425,N_7353);
xor U7541 (N_7541,N_7303,N_7270);
nand U7542 (N_7542,N_7392,N_7365);
or U7543 (N_7543,N_7448,N_7455);
and U7544 (N_7544,N_7308,N_7315);
nor U7545 (N_7545,N_7424,N_7341);
xnor U7546 (N_7546,N_7264,N_7445);
and U7547 (N_7547,N_7462,N_7285);
nor U7548 (N_7548,N_7368,N_7342);
xor U7549 (N_7549,N_7406,N_7474);
xnor U7550 (N_7550,N_7454,N_7360);
and U7551 (N_7551,N_7346,N_7433);
and U7552 (N_7552,N_7373,N_7386);
nor U7553 (N_7553,N_7348,N_7497);
nor U7554 (N_7554,N_7442,N_7498);
and U7555 (N_7555,N_7487,N_7300);
or U7556 (N_7556,N_7438,N_7481);
nor U7557 (N_7557,N_7361,N_7337);
and U7558 (N_7558,N_7340,N_7405);
nand U7559 (N_7559,N_7436,N_7482);
xor U7560 (N_7560,N_7313,N_7254);
xor U7561 (N_7561,N_7401,N_7320);
xnor U7562 (N_7562,N_7347,N_7281);
or U7563 (N_7563,N_7333,N_7332);
and U7564 (N_7564,N_7287,N_7316);
and U7565 (N_7565,N_7324,N_7274);
xnor U7566 (N_7566,N_7294,N_7375);
nor U7567 (N_7567,N_7290,N_7318);
and U7568 (N_7568,N_7463,N_7327);
nand U7569 (N_7569,N_7430,N_7297);
nand U7570 (N_7570,N_7282,N_7307);
and U7571 (N_7571,N_7385,N_7404);
and U7572 (N_7572,N_7266,N_7283);
or U7573 (N_7573,N_7457,N_7335);
nor U7574 (N_7574,N_7387,N_7447);
and U7575 (N_7575,N_7296,N_7259);
and U7576 (N_7576,N_7305,N_7407);
nand U7577 (N_7577,N_7345,N_7376);
nor U7578 (N_7578,N_7258,N_7460);
and U7579 (N_7579,N_7459,N_7413);
nand U7580 (N_7580,N_7412,N_7382);
xor U7581 (N_7581,N_7339,N_7369);
xor U7582 (N_7582,N_7322,N_7321);
or U7583 (N_7583,N_7289,N_7323);
nand U7584 (N_7584,N_7359,N_7372);
or U7585 (N_7585,N_7434,N_7480);
nor U7586 (N_7586,N_7284,N_7416);
nor U7587 (N_7587,N_7486,N_7476);
or U7588 (N_7588,N_7488,N_7485);
and U7589 (N_7589,N_7367,N_7389);
nor U7590 (N_7590,N_7428,N_7280);
and U7591 (N_7591,N_7295,N_7484);
nand U7592 (N_7592,N_7489,N_7399);
and U7593 (N_7593,N_7441,N_7354);
and U7594 (N_7594,N_7453,N_7343);
nor U7595 (N_7595,N_7395,N_7351);
and U7596 (N_7596,N_7298,N_7250);
nand U7597 (N_7597,N_7408,N_7252);
nor U7598 (N_7598,N_7344,N_7452);
and U7599 (N_7599,N_7260,N_7329);
nand U7600 (N_7600,N_7490,N_7410);
and U7601 (N_7601,N_7466,N_7451);
or U7602 (N_7602,N_7483,N_7279);
nor U7603 (N_7603,N_7304,N_7288);
and U7604 (N_7604,N_7461,N_7468);
and U7605 (N_7605,N_7470,N_7431);
nor U7606 (N_7606,N_7356,N_7391);
nand U7607 (N_7607,N_7437,N_7390);
and U7608 (N_7608,N_7251,N_7256);
and U7609 (N_7609,N_7330,N_7465);
xor U7610 (N_7610,N_7415,N_7402);
or U7611 (N_7611,N_7293,N_7267);
nand U7612 (N_7612,N_7272,N_7275);
xor U7613 (N_7613,N_7427,N_7331);
nand U7614 (N_7614,N_7358,N_7435);
xnor U7615 (N_7615,N_7334,N_7403);
nand U7616 (N_7616,N_7350,N_7309);
nand U7617 (N_7617,N_7472,N_7473);
xor U7618 (N_7618,N_7377,N_7423);
nand U7619 (N_7619,N_7456,N_7418);
and U7620 (N_7620,N_7271,N_7306);
or U7621 (N_7621,N_7310,N_7378);
or U7622 (N_7622,N_7357,N_7493);
and U7623 (N_7623,N_7443,N_7432);
xor U7624 (N_7624,N_7400,N_7471);
and U7625 (N_7625,N_7273,N_7263);
or U7626 (N_7626,N_7447,N_7376);
nand U7627 (N_7627,N_7280,N_7392);
and U7628 (N_7628,N_7417,N_7455);
or U7629 (N_7629,N_7251,N_7387);
xnor U7630 (N_7630,N_7388,N_7346);
xor U7631 (N_7631,N_7430,N_7287);
xor U7632 (N_7632,N_7376,N_7367);
or U7633 (N_7633,N_7456,N_7373);
nor U7634 (N_7634,N_7442,N_7430);
or U7635 (N_7635,N_7350,N_7331);
xor U7636 (N_7636,N_7446,N_7317);
or U7637 (N_7637,N_7344,N_7442);
xnor U7638 (N_7638,N_7299,N_7367);
or U7639 (N_7639,N_7363,N_7301);
xor U7640 (N_7640,N_7365,N_7348);
xnor U7641 (N_7641,N_7337,N_7460);
or U7642 (N_7642,N_7445,N_7325);
or U7643 (N_7643,N_7418,N_7257);
nor U7644 (N_7644,N_7438,N_7416);
xnor U7645 (N_7645,N_7313,N_7299);
or U7646 (N_7646,N_7284,N_7486);
nor U7647 (N_7647,N_7379,N_7335);
and U7648 (N_7648,N_7271,N_7454);
nand U7649 (N_7649,N_7433,N_7382);
nand U7650 (N_7650,N_7352,N_7288);
nor U7651 (N_7651,N_7263,N_7296);
and U7652 (N_7652,N_7462,N_7445);
nor U7653 (N_7653,N_7309,N_7426);
xnor U7654 (N_7654,N_7411,N_7259);
xor U7655 (N_7655,N_7345,N_7421);
nor U7656 (N_7656,N_7441,N_7327);
or U7657 (N_7657,N_7431,N_7316);
or U7658 (N_7658,N_7268,N_7349);
and U7659 (N_7659,N_7445,N_7423);
and U7660 (N_7660,N_7497,N_7401);
or U7661 (N_7661,N_7493,N_7359);
nor U7662 (N_7662,N_7483,N_7347);
or U7663 (N_7663,N_7402,N_7438);
xnor U7664 (N_7664,N_7395,N_7288);
nor U7665 (N_7665,N_7271,N_7408);
nand U7666 (N_7666,N_7367,N_7333);
and U7667 (N_7667,N_7364,N_7414);
and U7668 (N_7668,N_7254,N_7263);
or U7669 (N_7669,N_7464,N_7357);
nand U7670 (N_7670,N_7445,N_7453);
nand U7671 (N_7671,N_7279,N_7418);
and U7672 (N_7672,N_7272,N_7328);
nand U7673 (N_7673,N_7282,N_7455);
nor U7674 (N_7674,N_7385,N_7431);
and U7675 (N_7675,N_7305,N_7314);
xnor U7676 (N_7676,N_7326,N_7445);
nand U7677 (N_7677,N_7331,N_7352);
nor U7678 (N_7678,N_7455,N_7262);
nor U7679 (N_7679,N_7303,N_7413);
or U7680 (N_7680,N_7270,N_7413);
nand U7681 (N_7681,N_7316,N_7343);
nor U7682 (N_7682,N_7324,N_7298);
and U7683 (N_7683,N_7321,N_7332);
xnor U7684 (N_7684,N_7252,N_7388);
xnor U7685 (N_7685,N_7448,N_7381);
nor U7686 (N_7686,N_7488,N_7451);
nor U7687 (N_7687,N_7379,N_7332);
and U7688 (N_7688,N_7268,N_7478);
nand U7689 (N_7689,N_7433,N_7348);
nand U7690 (N_7690,N_7340,N_7478);
and U7691 (N_7691,N_7396,N_7316);
or U7692 (N_7692,N_7461,N_7466);
nand U7693 (N_7693,N_7449,N_7445);
xor U7694 (N_7694,N_7455,N_7405);
or U7695 (N_7695,N_7398,N_7457);
xor U7696 (N_7696,N_7405,N_7288);
xor U7697 (N_7697,N_7322,N_7339);
and U7698 (N_7698,N_7253,N_7300);
or U7699 (N_7699,N_7436,N_7342);
and U7700 (N_7700,N_7300,N_7328);
xnor U7701 (N_7701,N_7411,N_7494);
and U7702 (N_7702,N_7348,N_7292);
and U7703 (N_7703,N_7300,N_7316);
or U7704 (N_7704,N_7449,N_7472);
nand U7705 (N_7705,N_7408,N_7330);
nor U7706 (N_7706,N_7270,N_7421);
and U7707 (N_7707,N_7437,N_7378);
xnor U7708 (N_7708,N_7409,N_7280);
or U7709 (N_7709,N_7416,N_7327);
or U7710 (N_7710,N_7318,N_7426);
nor U7711 (N_7711,N_7477,N_7312);
xnor U7712 (N_7712,N_7303,N_7398);
or U7713 (N_7713,N_7355,N_7306);
or U7714 (N_7714,N_7452,N_7320);
nor U7715 (N_7715,N_7331,N_7346);
nand U7716 (N_7716,N_7261,N_7262);
nand U7717 (N_7717,N_7447,N_7465);
nor U7718 (N_7718,N_7291,N_7495);
xnor U7719 (N_7719,N_7431,N_7390);
and U7720 (N_7720,N_7295,N_7335);
nor U7721 (N_7721,N_7485,N_7373);
xnor U7722 (N_7722,N_7407,N_7257);
or U7723 (N_7723,N_7427,N_7406);
nand U7724 (N_7724,N_7301,N_7356);
and U7725 (N_7725,N_7297,N_7383);
xor U7726 (N_7726,N_7449,N_7282);
or U7727 (N_7727,N_7290,N_7462);
nand U7728 (N_7728,N_7493,N_7497);
xor U7729 (N_7729,N_7258,N_7399);
nor U7730 (N_7730,N_7322,N_7264);
or U7731 (N_7731,N_7480,N_7392);
and U7732 (N_7732,N_7304,N_7290);
nand U7733 (N_7733,N_7419,N_7424);
xor U7734 (N_7734,N_7278,N_7499);
xor U7735 (N_7735,N_7260,N_7384);
nand U7736 (N_7736,N_7470,N_7316);
nand U7737 (N_7737,N_7447,N_7276);
or U7738 (N_7738,N_7360,N_7377);
xnor U7739 (N_7739,N_7375,N_7350);
nor U7740 (N_7740,N_7400,N_7448);
nor U7741 (N_7741,N_7422,N_7493);
and U7742 (N_7742,N_7415,N_7499);
xnor U7743 (N_7743,N_7355,N_7469);
and U7744 (N_7744,N_7383,N_7337);
and U7745 (N_7745,N_7425,N_7452);
xor U7746 (N_7746,N_7346,N_7281);
xnor U7747 (N_7747,N_7275,N_7314);
and U7748 (N_7748,N_7256,N_7476);
or U7749 (N_7749,N_7401,N_7327);
nor U7750 (N_7750,N_7675,N_7684);
xnor U7751 (N_7751,N_7670,N_7571);
nor U7752 (N_7752,N_7551,N_7736);
xor U7753 (N_7753,N_7657,N_7673);
and U7754 (N_7754,N_7696,N_7703);
xnor U7755 (N_7755,N_7734,N_7535);
xor U7756 (N_7756,N_7531,N_7614);
and U7757 (N_7757,N_7648,N_7723);
xnor U7758 (N_7758,N_7682,N_7624);
xor U7759 (N_7759,N_7605,N_7737);
nand U7760 (N_7760,N_7699,N_7610);
and U7761 (N_7761,N_7503,N_7709);
xnor U7762 (N_7762,N_7749,N_7591);
nor U7763 (N_7763,N_7617,N_7658);
and U7764 (N_7764,N_7615,N_7688);
xnor U7765 (N_7765,N_7649,N_7598);
or U7766 (N_7766,N_7621,N_7567);
and U7767 (N_7767,N_7564,N_7548);
nor U7768 (N_7768,N_7597,N_7679);
nand U7769 (N_7769,N_7582,N_7522);
nor U7770 (N_7770,N_7524,N_7630);
or U7771 (N_7771,N_7672,N_7525);
nor U7772 (N_7772,N_7706,N_7747);
nor U7773 (N_7773,N_7659,N_7646);
xnor U7774 (N_7774,N_7619,N_7500);
and U7775 (N_7775,N_7642,N_7546);
xor U7776 (N_7776,N_7550,N_7544);
or U7777 (N_7777,N_7739,N_7586);
or U7778 (N_7778,N_7746,N_7695);
and U7779 (N_7779,N_7729,N_7620);
nor U7780 (N_7780,N_7708,N_7633);
nand U7781 (N_7781,N_7512,N_7575);
nand U7782 (N_7782,N_7622,N_7536);
or U7783 (N_7783,N_7711,N_7725);
xor U7784 (N_7784,N_7574,N_7634);
and U7785 (N_7785,N_7523,N_7680);
nand U7786 (N_7786,N_7521,N_7733);
nand U7787 (N_7787,N_7545,N_7580);
or U7788 (N_7788,N_7678,N_7509);
nor U7789 (N_7789,N_7629,N_7553);
nand U7790 (N_7790,N_7702,N_7539);
nor U7791 (N_7791,N_7537,N_7596);
nand U7792 (N_7792,N_7595,N_7655);
or U7793 (N_7793,N_7645,N_7713);
xnor U7794 (N_7794,N_7669,N_7566);
and U7795 (N_7795,N_7681,N_7508);
nand U7796 (N_7796,N_7583,N_7529);
nand U7797 (N_7797,N_7549,N_7609);
and U7798 (N_7798,N_7743,N_7511);
nor U7799 (N_7799,N_7554,N_7518);
and U7800 (N_7800,N_7611,N_7715);
and U7801 (N_7801,N_7541,N_7560);
nor U7802 (N_7802,N_7540,N_7731);
xnor U7803 (N_7803,N_7676,N_7641);
nor U7804 (N_7804,N_7654,N_7573);
and U7805 (N_7805,N_7744,N_7643);
and U7806 (N_7806,N_7661,N_7674);
nand U7807 (N_7807,N_7712,N_7741);
nor U7808 (N_7808,N_7569,N_7728);
xnor U7809 (N_7809,N_7662,N_7603);
nor U7810 (N_7810,N_7516,N_7602);
nand U7811 (N_7811,N_7552,N_7578);
nor U7812 (N_7812,N_7697,N_7592);
or U7813 (N_7813,N_7640,N_7727);
and U7814 (N_7814,N_7700,N_7730);
xnor U7815 (N_7815,N_7543,N_7519);
or U7816 (N_7816,N_7502,N_7530);
nand U7817 (N_7817,N_7722,N_7636);
xor U7818 (N_7818,N_7718,N_7714);
nor U7819 (N_7819,N_7572,N_7565);
xor U7820 (N_7820,N_7600,N_7726);
nand U7821 (N_7821,N_7720,N_7510);
xnor U7822 (N_7822,N_7542,N_7692);
nand U7823 (N_7823,N_7528,N_7698);
nand U7824 (N_7824,N_7538,N_7637);
or U7825 (N_7825,N_7506,N_7557);
xor U7826 (N_7826,N_7579,N_7590);
xor U7827 (N_7827,N_7685,N_7668);
and U7828 (N_7828,N_7740,N_7660);
nor U7829 (N_7829,N_7589,N_7639);
nand U7830 (N_7830,N_7534,N_7532);
nand U7831 (N_7831,N_7667,N_7513);
xnor U7832 (N_7832,N_7555,N_7587);
and U7833 (N_7833,N_7504,N_7745);
or U7834 (N_7834,N_7748,N_7717);
nor U7835 (N_7835,N_7585,N_7710);
nand U7836 (N_7836,N_7665,N_7563);
or U7837 (N_7837,N_7738,N_7568);
and U7838 (N_7838,N_7704,N_7635);
or U7839 (N_7839,N_7533,N_7570);
nor U7840 (N_7840,N_7687,N_7719);
nor U7841 (N_7841,N_7593,N_7742);
xnor U7842 (N_7842,N_7625,N_7653);
nand U7843 (N_7843,N_7732,N_7705);
xor U7844 (N_7844,N_7647,N_7663);
or U7845 (N_7845,N_7626,N_7693);
nor U7846 (N_7846,N_7716,N_7607);
or U7847 (N_7847,N_7558,N_7721);
nand U7848 (N_7848,N_7683,N_7691);
nor U7849 (N_7849,N_7584,N_7628);
and U7850 (N_7850,N_7724,N_7581);
or U7851 (N_7851,N_7608,N_7686);
xnor U7852 (N_7852,N_7694,N_7547);
xnor U7853 (N_7853,N_7650,N_7652);
and U7854 (N_7854,N_7735,N_7601);
or U7855 (N_7855,N_7599,N_7562);
nor U7856 (N_7856,N_7701,N_7689);
nor U7857 (N_7857,N_7656,N_7559);
and U7858 (N_7858,N_7623,N_7613);
nand U7859 (N_7859,N_7594,N_7690);
or U7860 (N_7860,N_7651,N_7588);
and U7861 (N_7861,N_7612,N_7505);
nor U7862 (N_7862,N_7627,N_7520);
or U7863 (N_7863,N_7664,N_7616);
xnor U7864 (N_7864,N_7576,N_7644);
xor U7865 (N_7865,N_7515,N_7556);
and U7866 (N_7866,N_7561,N_7666);
or U7867 (N_7867,N_7707,N_7631);
nand U7868 (N_7868,N_7514,N_7577);
nor U7869 (N_7869,N_7606,N_7527);
nor U7870 (N_7870,N_7638,N_7501);
xnor U7871 (N_7871,N_7604,N_7618);
and U7872 (N_7872,N_7507,N_7677);
nand U7873 (N_7873,N_7526,N_7632);
nor U7874 (N_7874,N_7671,N_7517);
or U7875 (N_7875,N_7545,N_7574);
nand U7876 (N_7876,N_7687,N_7662);
or U7877 (N_7877,N_7524,N_7552);
nand U7878 (N_7878,N_7560,N_7727);
nor U7879 (N_7879,N_7696,N_7702);
or U7880 (N_7880,N_7619,N_7708);
nand U7881 (N_7881,N_7576,N_7650);
nor U7882 (N_7882,N_7634,N_7655);
xor U7883 (N_7883,N_7626,N_7617);
nand U7884 (N_7884,N_7708,N_7601);
and U7885 (N_7885,N_7715,N_7642);
xnor U7886 (N_7886,N_7546,N_7629);
and U7887 (N_7887,N_7696,N_7523);
nor U7888 (N_7888,N_7597,N_7722);
or U7889 (N_7889,N_7594,N_7592);
and U7890 (N_7890,N_7559,N_7576);
and U7891 (N_7891,N_7577,N_7593);
nand U7892 (N_7892,N_7726,N_7626);
xor U7893 (N_7893,N_7522,N_7588);
or U7894 (N_7894,N_7606,N_7636);
or U7895 (N_7895,N_7654,N_7567);
or U7896 (N_7896,N_7644,N_7616);
nor U7897 (N_7897,N_7681,N_7524);
nor U7898 (N_7898,N_7626,N_7609);
or U7899 (N_7899,N_7652,N_7736);
nand U7900 (N_7900,N_7627,N_7537);
nand U7901 (N_7901,N_7534,N_7681);
nor U7902 (N_7902,N_7695,N_7659);
nor U7903 (N_7903,N_7551,N_7535);
nor U7904 (N_7904,N_7665,N_7654);
xor U7905 (N_7905,N_7693,N_7647);
and U7906 (N_7906,N_7731,N_7503);
nor U7907 (N_7907,N_7619,N_7570);
or U7908 (N_7908,N_7596,N_7674);
xnor U7909 (N_7909,N_7630,N_7522);
xor U7910 (N_7910,N_7549,N_7602);
or U7911 (N_7911,N_7514,N_7673);
xor U7912 (N_7912,N_7743,N_7716);
nand U7913 (N_7913,N_7525,N_7719);
nor U7914 (N_7914,N_7629,N_7568);
or U7915 (N_7915,N_7677,N_7704);
nand U7916 (N_7916,N_7517,N_7717);
and U7917 (N_7917,N_7588,N_7725);
and U7918 (N_7918,N_7554,N_7548);
nor U7919 (N_7919,N_7564,N_7687);
nor U7920 (N_7920,N_7557,N_7564);
nand U7921 (N_7921,N_7571,N_7631);
and U7922 (N_7922,N_7684,N_7600);
xor U7923 (N_7923,N_7649,N_7529);
or U7924 (N_7924,N_7673,N_7617);
and U7925 (N_7925,N_7516,N_7665);
and U7926 (N_7926,N_7520,N_7577);
xor U7927 (N_7927,N_7671,N_7663);
nand U7928 (N_7928,N_7703,N_7701);
and U7929 (N_7929,N_7571,N_7673);
and U7930 (N_7930,N_7717,N_7529);
nor U7931 (N_7931,N_7673,N_7745);
and U7932 (N_7932,N_7686,N_7707);
and U7933 (N_7933,N_7601,N_7548);
xnor U7934 (N_7934,N_7562,N_7577);
nand U7935 (N_7935,N_7681,N_7540);
nor U7936 (N_7936,N_7562,N_7533);
or U7937 (N_7937,N_7507,N_7684);
nor U7938 (N_7938,N_7652,N_7673);
nor U7939 (N_7939,N_7653,N_7524);
nand U7940 (N_7940,N_7544,N_7657);
xor U7941 (N_7941,N_7580,N_7581);
and U7942 (N_7942,N_7532,N_7559);
xnor U7943 (N_7943,N_7747,N_7678);
nor U7944 (N_7944,N_7686,N_7566);
xor U7945 (N_7945,N_7676,N_7629);
or U7946 (N_7946,N_7564,N_7590);
or U7947 (N_7947,N_7623,N_7585);
and U7948 (N_7948,N_7701,N_7574);
or U7949 (N_7949,N_7716,N_7695);
nand U7950 (N_7950,N_7555,N_7631);
nand U7951 (N_7951,N_7677,N_7619);
and U7952 (N_7952,N_7713,N_7647);
and U7953 (N_7953,N_7626,N_7505);
nor U7954 (N_7954,N_7627,N_7572);
nor U7955 (N_7955,N_7656,N_7605);
nor U7956 (N_7956,N_7501,N_7603);
and U7957 (N_7957,N_7736,N_7564);
and U7958 (N_7958,N_7561,N_7651);
nand U7959 (N_7959,N_7573,N_7539);
or U7960 (N_7960,N_7545,N_7589);
or U7961 (N_7961,N_7515,N_7546);
xnor U7962 (N_7962,N_7546,N_7607);
and U7963 (N_7963,N_7534,N_7536);
and U7964 (N_7964,N_7741,N_7631);
xnor U7965 (N_7965,N_7646,N_7585);
and U7966 (N_7966,N_7602,N_7702);
and U7967 (N_7967,N_7693,N_7522);
xnor U7968 (N_7968,N_7695,N_7563);
nand U7969 (N_7969,N_7520,N_7549);
nand U7970 (N_7970,N_7625,N_7631);
nand U7971 (N_7971,N_7568,N_7656);
xnor U7972 (N_7972,N_7517,N_7664);
or U7973 (N_7973,N_7512,N_7613);
or U7974 (N_7974,N_7696,N_7714);
xor U7975 (N_7975,N_7722,N_7606);
nor U7976 (N_7976,N_7521,N_7661);
and U7977 (N_7977,N_7683,N_7636);
nand U7978 (N_7978,N_7721,N_7657);
nor U7979 (N_7979,N_7700,N_7628);
nand U7980 (N_7980,N_7536,N_7717);
or U7981 (N_7981,N_7724,N_7534);
xor U7982 (N_7982,N_7614,N_7703);
xor U7983 (N_7983,N_7626,N_7506);
nor U7984 (N_7984,N_7515,N_7630);
or U7985 (N_7985,N_7608,N_7556);
nand U7986 (N_7986,N_7603,N_7719);
nor U7987 (N_7987,N_7739,N_7547);
nor U7988 (N_7988,N_7620,N_7563);
nand U7989 (N_7989,N_7703,N_7506);
nand U7990 (N_7990,N_7714,N_7508);
nand U7991 (N_7991,N_7535,N_7523);
and U7992 (N_7992,N_7621,N_7530);
xor U7993 (N_7993,N_7686,N_7733);
and U7994 (N_7994,N_7722,N_7617);
or U7995 (N_7995,N_7684,N_7549);
xnor U7996 (N_7996,N_7570,N_7506);
xor U7997 (N_7997,N_7621,N_7519);
nor U7998 (N_7998,N_7501,N_7736);
nor U7999 (N_7999,N_7719,N_7553);
xor U8000 (N_8000,N_7863,N_7962);
xor U8001 (N_8001,N_7778,N_7839);
and U8002 (N_8002,N_7775,N_7837);
nor U8003 (N_8003,N_7953,N_7854);
nor U8004 (N_8004,N_7828,N_7967);
nand U8005 (N_8005,N_7858,N_7860);
nor U8006 (N_8006,N_7920,N_7800);
nor U8007 (N_8007,N_7955,N_7798);
nand U8008 (N_8008,N_7867,N_7905);
nand U8009 (N_8009,N_7842,N_7992);
or U8010 (N_8010,N_7779,N_7898);
nor U8011 (N_8011,N_7978,N_7819);
nand U8012 (N_8012,N_7784,N_7813);
nand U8013 (N_8013,N_7853,N_7838);
or U8014 (N_8014,N_7806,N_7919);
nor U8015 (N_8015,N_7895,N_7763);
nand U8016 (N_8016,N_7830,N_7794);
or U8017 (N_8017,N_7793,N_7768);
or U8018 (N_8018,N_7886,N_7769);
nor U8019 (N_8019,N_7892,N_7818);
or U8020 (N_8020,N_7807,N_7796);
xor U8021 (N_8021,N_7889,N_7900);
and U8022 (N_8022,N_7890,N_7856);
xnor U8023 (N_8023,N_7909,N_7976);
xnor U8024 (N_8024,N_7902,N_7951);
nand U8025 (N_8025,N_7773,N_7761);
nand U8026 (N_8026,N_7971,N_7833);
nand U8027 (N_8027,N_7981,N_7804);
nand U8028 (N_8028,N_7934,N_7991);
xor U8029 (N_8029,N_7824,N_7915);
nand U8030 (N_8030,N_7767,N_7820);
or U8031 (N_8031,N_7937,N_7946);
or U8032 (N_8032,N_7827,N_7811);
or U8033 (N_8033,N_7885,N_7988);
xor U8034 (N_8034,N_7787,N_7947);
nor U8035 (N_8035,N_7985,N_7986);
xor U8036 (N_8036,N_7913,N_7999);
nor U8037 (N_8037,N_7954,N_7871);
nand U8038 (N_8038,N_7810,N_7751);
nand U8039 (N_8039,N_7911,N_7753);
and U8040 (N_8040,N_7914,N_7846);
xor U8041 (N_8041,N_7997,N_7990);
nand U8042 (N_8042,N_7755,N_7869);
and U8043 (N_8043,N_7759,N_7843);
nand U8044 (N_8044,N_7961,N_7850);
or U8045 (N_8045,N_7906,N_7907);
or U8046 (N_8046,N_7994,N_7965);
nand U8047 (N_8047,N_7812,N_7910);
and U8048 (N_8048,N_7896,N_7829);
and U8049 (N_8049,N_7979,N_7832);
xor U8050 (N_8050,N_7912,N_7777);
nand U8051 (N_8051,N_7974,N_7802);
nor U8052 (N_8052,N_7795,N_7814);
nor U8053 (N_8053,N_7958,N_7956);
nand U8054 (N_8054,N_7754,N_7957);
or U8055 (N_8055,N_7866,N_7941);
and U8056 (N_8056,N_7980,N_7792);
nor U8057 (N_8057,N_7805,N_7879);
xor U8058 (N_8058,N_7844,N_7799);
and U8059 (N_8059,N_7916,N_7904);
nor U8060 (N_8060,N_7882,N_7880);
and U8061 (N_8061,N_7816,N_7903);
and U8062 (N_8062,N_7935,N_7780);
xor U8063 (N_8063,N_7940,N_7925);
xnor U8064 (N_8064,N_7931,N_7918);
and U8065 (N_8065,N_7924,N_7801);
nor U8066 (N_8066,N_7848,N_7884);
nand U8067 (N_8067,N_7786,N_7845);
xor U8068 (N_8068,N_7944,N_7982);
nand U8069 (N_8069,N_7772,N_7859);
nor U8070 (N_8070,N_7762,N_7888);
xnor U8071 (N_8071,N_7809,N_7969);
nand U8072 (N_8072,N_7932,N_7826);
nand U8073 (N_8073,N_7891,N_7864);
nor U8074 (N_8074,N_7921,N_7861);
nor U8075 (N_8075,N_7803,N_7949);
or U8076 (N_8076,N_7783,N_7774);
and U8077 (N_8077,N_7901,N_7883);
and U8078 (N_8078,N_7788,N_7899);
nor U8079 (N_8079,N_7760,N_7948);
nand U8080 (N_8080,N_7873,N_7752);
or U8081 (N_8081,N_7757,N_7952);
or U8082 (N_8082,N_7939,N_7834);
nand U8083 (N_8083,N_7943,N_7968);
nand U8084 (N_8084,N_7950,N_7923);
nand U8085 (N_8085,N_7817,N_7849);
or U8086 (N_8086,N_7995,N_7821);
nor U8087 (N_8087,N_7928,N_7836);
nand U8088 (N_8088,N_7942,N_7825);
nor U8089 (N_8089,N_7887,N_7959);
xor U8090 (N_8090,N_7897,N_7789);
and U8091 (N_8091,N_7938,N_7797);
or U8092 (N_8092,N_7835,N_7770);
xor U8093 (N_8093,N_7865,N_7933);
xnor U8094 (N_8094,N_7862,N_7960);
nor U8095 (N_8095,N_7765,N_7973);
and U8096 (N_8096,N_7771,N_7984);
nor U8097 (N_8097,N_7963,N_7808);
nor U8098 (N_8098,N_7847,N_7929);
nor U8099 (N_8099,N_7881,N_7750);
and U8100 (N_8100,N_7851,N_7840);
or U8101 (N_8101,N_7972,N_7975);
or U8102 (N_8102,N_7977,N_7776);
or U8103 (N_8103,N_7790,N_7870);
and U8104 (N_8104,N_7930,N_7781);
and U8105 (N_8105,N_7922,N_7917);
or U8106 (N_8106,N_7758,N_7872);
xnor U8107 (N_8107,N_7831,N_7908);
nand U8108 (N_8108,N_7936,N_7876);
nor U8109 (N_8109,N_7785,N_7766);
xor U8110 (N_8110,N_7782,N_7970);
nor U8111 (N_8111,N_7878,N_7841);
nand U8112 (N_8112,N_7877,N_7987);
xnor U8113 (N_8113,N_7964,N_7989);
nor U8114 (N_8114,N_7855,N_7893);
or U8115 (N_8115,N_7857,N_7926);
and U8116 (N_8116,N_7998,N_7996);
and U8117 (N_8117,N_7822,N_7823);
or U8118 (N_8118,N_7756,N_7791);
nor U8119 (N_8119,N_7894,N_7875);
nand U8120 (N_8120,N_7945,N_7874);
or U8121 (N_8121,N_7927,N_7993);
xnor U8122 (N_8122,N_7852,N_7764);
xnor U8123 (N_8123,N_7983,N_7815);
nor U8124 (N_8124,N_7868,N_7966);
nand U8125 (N_8125,N_7781,N_7790);
nand U8126 (N_8126,N_7933,N_7759);
nand U8127 (N_8127,N_7791,N_7970);
nor U8128 (N_8128,N_7931,N_7912);
and U8129 (N_8129,N_7810,N_7983);
and U8130 (N_8130,N_7925,N_7966);
nor U8131 (N_8131,N_7753,N_7963);
nand U8132 (N_8132,N_7764,N_7865);
or U8133 (N_8133,N_7999,N_7983);
and U8134 (N_8134,N_7889,N_7867);
xnor U8135 (N_8135,N_7995,N_7890);
nand U8136 (N_8136,N_7805,N_7779);
nor U8137 (N_8137,N_7805,N_7797);
or U8138 (N_8138,N_7860,N_7884);
xnor U8139 (N_8139,N_7977,N_7757);
xor U8140 (N_8140,N_7991,N_7883);
xor U8141 (N_8141,N_7763,N_7833);
or U8142 (N_8142,N_7976,N_7989);
and U8143 (N_8143,N_7761,N_7993);
nor U8144 (N_8144,N_7916,N_7915);
xor U8145 (N_8145,N_7827,N_7991);
nor U8146 (N_8146,N_7842,N_7969);
and U8147 (N_8147,N_7844,N_7785);
nand U8148 (N_8148,N_7897,N_7921);
or U8149 (N_8149,N_7979,N_7809);
nor U8150 (N_8150,N_7767,N_7887);
nand U8151 (N_8151,N_7937,N_7998);
xnor U8152 (N_8152,N_7801,N_7851);
xnor U8153 (N_8153,N_7950,N_7910);
nor U8154 (N_8154,N_7884,N_7916);
and U8155 (N_8155,N_7835,N_7841);
or U8156 (N_8156,N_7877,N_7978);
or U8157 (N_8157,N_7795,N_7803);
or U8158 (N_8158,N_7996,N_7814);
nand U8159 (N_8159,N_7765,N_7888);
nor U8160 (N_8160,N_7961,N_7821);
xnor U8161 (N_8161,N_7931,N_7767);
nor U8162 (N_8162,N_7788,N_7882);
nand U8163 (N_8163,N_7756,N_7753);
or U8164 (N_8164,N_7852,N_7834);
or U8165 (N_8165,N_7851,N_7760);
or U8166 (N_8166,N_7784,N_7822);
or U8167 (N_8167,N_7874,N_7791);
and U8168 (N_8168,N_7878,N_7921);
or U8169 (N_8169,N_7806,N_7769);
xor U8170 (N_8170,N_7896,N_7795);
xor U8171 (N_8171,N_7754,N_7804);
xor U8172 (N_8172,N_7911,N_7950);
nand U8173 (N_8173,N_7758,N_7948);
and U8174 (N_8174,N_7976,N_7946);
nand U8175 (N_8175,N_7930,N_7805);
xor U8176 (N_8176,N_7816,N_7841);
nor U8177 (N_8177,N_7879,N_7986);
xnor U8178 (N_8178,N_7883,N_7900);
or U8179 (N_8179,N_7754,N_7808);
nand U8180 (N_8180,N_7929,N_7931);
and U8181 (N_8181,N_7790,N_7995);
and U8182 (N_8182,N_7902,N_7968);
xnor U8183 (N_8183,N_7755,N_7766);
nor U8184 (N_8184,N_7815,N_7934);
or U8185 (N_8185,N_7988,N_7792);
nor U8186 (N_8186,N_7965,N_7750);
nor U8187 (N_8187,N_7964,N_7874);
nor U8188 (N_8188,N_7800,N_7963);
nand U8189 (N_8189,N_7932,N_7766);
or U8190 (N_8190,N_7992,N_7968);
xor U8191 (N_8191,N_7768,N_7816);
nand U8192 (N_8192,N_7773,N_7925);
or U8193 (N_8193,N_7851,N_7809);
and U8194 (N_8194,N_7925,N_7868);
nor U8195 (N_8195,N_7973,N_7848);
or U8196 (N_8196,N_7807,N_7779);
nor U8197 (N_8197,N_7926,N_7757);
and U8198 (N_8198,N_7879,N_7969);
and U8199 (N_8199,N_7946,N_7941);
xnor U8200 (N_8200,N_7758,N_7765);
nor U8201 (N_8201,N_7990,N_7818);
xor U8202 (N_8202,N_7994,N_7800);
or U8203 (N_8203,N_7966,N_7806);
nor U8204 (N_8204,N_7989,N_7765);
or U8205 (N_8205,N_7997,N_7939);
and U8206 (N_8206,N_7859,N_7935);
xor U8207 (N_8207,N_7960,N_7946);
xor U8208 (N_8208,N_7988,N_7852);
nor U8209 (N_8209,N_7817,N_7808);
and U8210 (N_8210,N_7971,N_7912);
xor U8211 (N_8211,N_7833,N_7823);
nand U8212 (N_8212,N_7949,N_7900);
and U8213 (N_8213,N_7775,N_7962);
nand U8214 (N_8214,N_7917,N_7906);
nor U8215 (N_8215,N_7983,N_7882);
nor U8216 (N_8216,N_7973,N_7910);
nand U8217 (N_8217,N_7777,N_7758);
nand U8218 (N_8218,N_7947,N_7779);
nand U8219 (N_8219,N_7977,N_7819);
nand U8220 (N_8220,N_7964,N_7851);
or U8221 (N_8221,N_7768,N_7833);
or U8222 (N_8222,N_7886,N_7905);
and U8223 (N_8223,N_7966,N_7855);
xnor U8224 (N_8224,N_7980,N_7968);
nor U8225 (N_8225,N_7959,N_7937);
nand U8226 (N_8226,N_7774,N_7790);
xnor U8227 (N_8227,N_7775,N_7965);
or U8228 (N_8228,N_7972,N_7940);
xnor U8229 (N_8229,N_7904,N_7779);
nand U8230 (N_8230,N_7900,N_7780);
or U8231 (N_8231,N_7935,N_7976);
xnor U8232 (N_8232,N_7868,N_7852);
or U8233 (N_8233,N_7880,N_7956);
nor U8234 (N_8234,N_7943,N_7900);
xor U8235 (N_8235,N_7796,N_7922);
nand U8236 (N_8236,N_7934,N_7890);
xnor U8237 (N_8237,N_7903,N_7815);
xor U8238 (N_8238,N_7894,N_7810);
nand U8239 (N_8239,N_7791,N_7919);
xor U8240 (N_8240,N_7953,N_7830);
nor U8241 (N_8241,N_7907,N_7865);
nand U8242 (N_8242,N_7935,N_7900);
nand U8243 (N_8243,N_7944,N_7921);
and U8244 (N_8244,N_7798,N_7757);
nand U8245 (N_8245,N_7950,N_7887);
nand U8246 (N_8246,N_7972,N_7755);
or U8247 (N_8247,N_7932,N_7804);
and U8248 (N_8248,N_7761,N_7792);
or U8249 (N_8249,N_7887,N_7829);
and U8250 (N_8250,N_8176,N_8181);
nor U8251 (N_8251,N_8211,N_8059);
or U8252 (N_8252,N_8030,N_8036);
nor U8253 (N_8253,N_8223,N_8183);
or U8254 (N_8254,N_8219,N_8165);
nand U8255 (N_8255,N_8106,N_8168);
nand U8256 (N_8256,N_8009,N_8131);
nor U8257 (N_8257,N_8062,N_8102);
and U8258 (N_8258,N_8020,N_8225);
nor U8259 (N_8259,N_8127,N_8079);
or U8260 (N_8260,N_8205,N_8217);
and U8261 (N_8261,N_8175,N_8031);
xor U8262 (N_8262,N_8004,N_8002);
nand U8263 (N_8263,N_8184,N_8249);
nor U8264 (N_8264,N_8034,N_8063);
and U8265 (N_8265,N_8187,N_8024);
xor U8266 (N_8266,N_8060,N_8015);
xor U8267 (N_8267,N_8143,N_8247);
xor U8268 (N_8268,N_8076,N_8226);
nor U8269 (N_8269,N_8058,N_8144);
or U8270 (N_8270,N_8068,N_8227);
nor U8271 (N_8271,N_8081,N_8235);
nor U8272 (N_8272,N_8220,N_8041);
or U8273 (N_8273,N_8082,N_8019);
nand U8274 (N_8274,N_8180,N_8095);
nor U8275 (N_8275,N_8003,N_8174);
or U8276 (N_8276,N_8051,N_8149);
nand U8277 (N_8277,N_8126,N_8084);
or U8278 (N_8278,N_8115,N_8246);
xnor U8279 (N_8279,N_8201,N_8139);
and U8280 (N_8280,N_8080,N_8173);
xnor U8281 (N_8281,N_8075,N_8240);
nor U8282 (N_8282,N_8212,N_8236);
and U8283 (N_8283,N_8088,N_8186);
nor U8284 (N_8284,N_8132,N_8027);
and U8285 (N_8285,N_8072,N_8204);
nand U8286 (N_8286,N_8229,N_8094);
nor U8287 (N_8287,N_8099,N_8142);
nand U8288 (N_8288,N_8044,N_8233);
and U8289 (N_8289,N_8156,N_8237);
or U8290 (N_8290,N_8158,N_8100);
and U8291 (N_8291,N_8189,N_8023);
nand U8292 (N_8292,N_8207,N_8054);
and U8293 (N_8293,N_8116,N_8045);
nor U8294 (N_8294,N_8029,N_8218);
or U8295 (N_8295,N_8104,N_8089);
nor U8296 (N_8296,N_8097,N_8129);
and U8297 (N_8297,N_8133,N_8206);
xnor U8298 (N_8298,N_8078,N_8118);
nor U8299 (N_8299,N_8043,N_8047);
and U8300 (N_8300,N_8224,N_8141);
xnor U8301 (N_8301,N_8083,N_8052);
nand U8302 (N_8302,N_8198,N_8208);
xnor U8303 (N_8303,N_8248,N_8120);
xor U8304 (N_8304,N_8122,N_8145);
and U8305 (N_8305,N_8007,N_8150);
and U8306 (N_8306,N_8077,N_8101);
or U8307 (N_8307,N_8146,N_8025);
nand U8308 (N_8308,N_8238,N_8182);
nand U8309 (N_8309,N_8163,N_8130);
or U8310 (N_8310,N_8178,N_8221);
and U8311 (N_8311,N_8037,N_8232);
nand U8312 (N_8312,N_8177,N_8245);
nand U8313 (N_8313,N_8162,N_8048);
and U8314 (N_8314,N_8216,N_8055);
nor U8315 (N_8315,N_8006,N_8073);
xnor U8316 (N_8316,N_8065,N_8241);
xor U8317 (N_8317,N_8137,N_8016);
nand U8318 (N_8318,N_8109,N_8140);
or U8319 (N_8319,N_8185,N_8191);
nand U8320 (N_8320,N_8010,N_8056);
xnor U8321 (N_8321,N_8107,N_8157);
or U8322 (N_8322,N_8119,N_8243);
and U8323 (N_8323,N_8155,N_8021);
xor U8324 (N_8324,N_8091,N_8110);
or U8325 (N_8325,N_8042,N_8172);
or U8326 (N_8326,N_8194,N_8199);
or U8327 (N_8327,N_8028,N_8012);
xor U8328 (N_8328,N_8167,N_8053);
or U8329 (N_8329,N_8192,N_8200);
nand U8330 (N_8330,N_8231,N_8135);
or U8331 (N_8331,N_8090,N_8092);
or U8332 (N_8332,N_8169,N_8166);
or U8333 (N_8333,N_8000,N_8013);
and U8334 (N_8334,N_8040,N_8114);
nor U8335 (N_8335,N_8125,N_8136);
or U8336 (N_8336,N_8147,N_8202);
xor U8337 (N_8337,N_8230,N_8179);
nand U8338 (N_8338,N_8134,N_8188);
nor U8339 (N_8339,N_8105,N_8121);
or U8340 (N_8340,N_8113,N_8103);
and U8341 (N_8341,N_8196,N_8160);
nand U8342 (N_8342,N_8171,N_8039);
nor U8343 (N_8343,N_8018,N_8005);
nand U8344 (N_8344,N_8117,N_8203);
or U8345 (N_8345,N_8159,N_8022);
and U8346 (N_8346,N_8087,N_8057);
nand U8347 (N_8347,N_8234,N_8128);
and U8348 (N_8348,N_8112,N_8066);
xor U8349 (N_8349,N_8001,N_8108);
nor U8350 (N_8350,N_8164,N_8242);
or U8351 (N_8351,N_8038,N_8070);
or U8352 (N_8352,N_8035,N_8071);
and U8353 (N_8353,N_8195,N_8170);
xor U8354 (N_8354,N_8161,N_8098);
or U8355 (N_8355,N_8096,N_8244);
or U8356 (N_8356,N_8190,N_8014);
and U8357 (N_8357,N_8049,N_8222);
and U8358 (N_8358,N_8067,N_8111);
nor U8359 (N_8359,N_8032,N_8153);
nor U8360 (N_8360,N_8154,N_8210);
and U8361 (N_8361,N_8011,N_8026);
or U8362 (N_8362,N_8064,N_8093);
nand U8363 (N_8363,N_8152,N_8148);
and U8364 (N_8364,N_8138,N_8124);
and U8365 (N_8365,N_8209,N_8123);
and U8366 (N_8366,N_8193,N_8074);
and U8367 (N_8367,N_8069,N_8008);
nand U8368 (N_8368,N_8228,N_8197);
nand U8369 (N_8369,N_8214,N_8050);
or U8370 (N_8370,N_8033,N_8061);
or U8371 (N_8371,N_8085,N_8151);
or U8372 (N_8372,N_8215,N_8239);
and U8373 (N_8373,N_8086,N_8017);
xnor U8374 (N_8374,N_8046,N_8213);
xnor U8375 (N_8375,N_8112,N_8124);
nand U8376 (N_8376,N_8235,N_8171);
and U8377 (N_8377,N_8215,N_8223);
nand U8378 (N_8378,N_8163,N_8141);
xor U8379 (N_8379,N_8141,N_8159);
or U8380 (N_8380,N_8166,N_8066);
nand U8381 (N_8381,N_8088,N_8082);
and U8382 (N_8382,N_8163,N_8202);
or U8383 (N_8383,N_8217,N_8234);
or U8384 (N_8384,N_8172,N_8187);
or U8385 (N_8385,N_8218,N_8188);
xor U8386 (N_8386,N_8247,N_8033);
xnor U8387 (N_8387,N_8067,N_8227);
and U8388 (N_8388,N_8132,N_8189);
xnor U8389 (N_8389,N_8214,N_8035);
nor U8390 (N_8390,N_8181,N_8183);
nor U8391 (N_8391,N_8190,N_8044);
and U8392 (N_8392,N_8147,N_8086);
nor U8393 (N_8393,N_8071,N_8146);
nand U8394 (N_8394,N_8006,N_8144);
xor U8395 (N_8395,N_8169,N_8245);
xnor U8396 (N_8396,N_8141,N_8185);
or U8397 (N_8397,N_8247,N_8214);
nand U8398 (N_8398,N_8022,N_8063);
and U8399 (N_8399,N_8203,N_8046);
xnor U8400 (N_8400,N_8067,N_8160);
nand U8401 (N_8401,N_8117,N_8027);
xor U8402 (N_8402,N_8124,N_8190);
xor U8403 (N_8403,N_8237,N_8155);
xnor U8404 (N_8404,N_8182,N_8227);
nor U8405 (N_8405,N_8046,N_8163);
nand U8406 (N_8406,N_8249,N_8080);
nand U8407 (N_8407,N_8216,N_8148);
nor U8408 (N_8408,N_8220,N_8077);
nor U8409 (N_8409,N_8124,N_8146);
xor U8410 (N_8410,N_8086,N_8054);
xnor U8411 (N_8411,N_8218,N_8127);
nor U8412 (N_8412,N_8019,N_8223);
nor U8413 (N_8413,N_8177,N_8045);
xnor U8414 (N_8414,N_8229,N_8210);
xor U8415 (N_8415,N_8179,N_8069);
nand U8416 (N_8416,N_8056,N_8107);
nor U8417 (N_8417,N_8203,N_8097);
nand U8418 (N_8418,N_8111,N_8198);
or U8419 (N_8419,N_8236,N_8213);
nand U8420 (N_8420,N_8162,N_8088);
nor U8421 (N_8421,N_8186,N_8245);
xnor U8422 (N_8422,N_8017,N_8020);
or U8423 (N_8423,N_8230,N_8166);
and U8424 (N_8424,N_8153,N_8075);
nor U8425 (N_8425,N_8218,N_8131);
or U8426 (N_8426,N_8026,N_8186);
nor U8427 (N_8427,N_8106,N_8018);
or U8428 (N_8428,N_8045,N_8198);
and U8429 (N_8429,N_8057,N_8090);
nor U8430 (N_8430,N_8205,N_8156);
nand U8431 (N_8431,N_8229,N_8228);
xnor U8432 (N_8432,N_8114,N_8106);
nand U8433 (N_8433,N_8138,N_8230);
or U8434 (N_8434,N_8103,N_8187);
nand U8435 (N_8435,N_8236,N_8017);
or U8436 (N_8436,N_8077,N_8178);
nand U8437 (N_8437,N_8229,N_8216);
and U8438 (N_8438,N_8166,N_8204);
and U8439 (N_8439,N_8197,N_8131);
nor U8440 (N_8440,N_8090,N_8068);
nand U8441 (N_8441,N_8110,N_8106);
xor U8442 (N_8442,N_8238,N_8134);
nor U8443 (N_8443,N_8069,N_8040);
xnor U8444 (N_8444,N_8142,N_8123);
nand U8445 (N_8445,N_8036,N_8022);
xnor U8446 (N_8446,N_8112,N_8053);
nand U8447 (N_8447,N_8227,N_8111);
nor U8448 (N_8448,N_8178,N_8053);
or U8449 (N_8449,N_8125,N_8006);
nand U8450 (N_8450,N_8017,N_8013);
nor U8451 (N_8451,N_8062,N_8084);
xor U8452 (N_8452,N_8020,N_8077);
nor U8453 (N_8453,N_8066,N_8171);
nand U8454 (N_8454,N_8222,N_8032);
xnor U8455 (N_8455,N_8010,N_8027);
xor U8456 (N_8456,N_8117,N_8050);
and U8457 (N_8457,N_8107,N_8239);
nand U8458 (N_8458,N_8089,N_8047);
and U8459 (N_8459,N_8003,N_8091);
xnor U8460 (N_8460,N_8041,N_8091);
nand U8461 (N_8461,N_8151,N_8047);
and U8462 (N_8462,N_8094,N_8044);
xor U8463 (N_8463,N_8152,N_8028);
and U8464 (N_8464,N_8232,N_8102);
or U8465 (N_8465,N_8132,N_8160);
nand U8466 (N_8466,N_8237,N_8053);
nor U8467 (N_8467,N_8162,N_8053);
and U8468 (N_8468,N_8241,N_8077);
and U8469 (N_8469,N_8177,N_8124);
and U8470 (N_8470,N_8091,N_8072);
nor U8471 (N_8471,N_8061,N_8173);
nand U8472 (N_8472,N_8156,N_8074);
and U8473 (N_8473,N_8100,N_8177);
nor U8474 (N_8474,N_8042,N_8140);
or U8475 (N_8475,N_8211,N_8232);
or U8476 (N_8476,N_8230,N_8165);
nor U8477 (N_8477,N_8001,N_8147);
nand U8478 (N_8478,N_8105,N_8091);
xnor U8479 (N_8479,N_8162,N_8174);
or U8480 (N_8480,N_8149,N_8206);
nor U8481 (N_8481,N_8013,N_8150);
nand U8482 (N_8482,N_8209,N_8129);
and U8483 (N_8483,N_8107,N_8173);
nand U8484 (N_8484,N_8235,N_8094);
and U8485 (N_8485,N_8108,N_8039);
nand U8486 (N_8486,N_8238,N_8160);
nor U8487 (N_8487,N_8087,N_8014);
xnor U8488 (N_8488,N_8041,N_8094);
and U8489 (N_8489,N_8243,N_8051);
and U8490 (N_8490,N_8119,N_8222);
and U8491 (N_8491,N_8228,N_8051);
nor U8492 (N_8492,N_8093,N_8020);
xnor U8493 (N_8493,N_8145,N_8100);
nor U8494 (N_8494,N_8120,N_8157);
nor U8495 (N_8495,N_8000,N_8026);
or U8496 (N_8496,N_8024,N_8121);
xor U8497 (N_8497,N_8236,N_8182);
and U8498 (N_8498,N_8221,N_8024);
xor U8499 (N_8499,N_8084,N_8127);
nand U8500 (N_8500,N_8318,N_8480);
or U8501 (N_8501,N_8364,N_8390);
or U8502 (N_8502,N_8389,N_8305);
or U8503 (N_8503,N_8277,N_8320);
nand U8504 (N_8504,N_8419,N_8498);
and U8505 (N_8505,N_8388,N_8291);
xnor U8506 (N_8506,N_8259,N_8307);
and U8507 (N_8507,N_8363,N_8407);
nor U8508 (N_8508,N_8403,N_8470);
or U8509 (N_8509,N_8271,N_8288);
or U8510 (N_8510,N_8386,N_8327);
xnor U8511 (N_8511,N_8460,N_8395);
nor U8512 (N_8512,N_8349,N_8435);
nor U8513 (N_8513,N_8452,N_8340);
and U8514 (N_8514,N_8287,N_8383);
nand U8515 (N_8515,N_8377,N_8267);
and U8516 (N_8516,N_8272,N_8289);
nor U8517 (N_8517,N_8339,N_8309);
or U8518 (N_8518,N_8285,N_8464);
xor U8519 (N_8519,N_8336,N_8469);
nor U8520 (N_8520,N_8302,N_8373);
xnor U8521 (N_8521,N_8448,N_8374);
and U8522 (N_8522,N_8334,N_8379);
xor U8523 (N_8523,N_8496,N_8481);
or U8524 (N_8524,N_8428,N_8476);
nor U8525 (N_8525,N_8445,N_8286);
and U8526 (N_8526,N_8468,N_8495);
and U8527 (N_8527,N_8298,N_8399);
or U8528 (N_8528,N_8250,N_8489);
xor U8529 (N_8529,N_8257,N_8366);
nand U8530 (N_8530,N_8409,N_8438);
and U8531 (N_8531,N_8343,N_8412);
nor U8532 (N_8532,N_8268,N_8442);
nor U8533 (N_8533,N_8465,N_8322);
and U8534 (N_8534,N_8375,N_8492);
nand U8535 (N_8535,N_8304,N_8361);
nand U8536 (N_8536,N_8311,N_8353);
xnor U8537 (N_8537,N_8437,N_8342);
xor U8538 (N_8538,N_8325,N_8385);
nand U8539 (N_8539,N_8433,N_8345);
xor U8540 (N_8540,N_8253,N_8434);
nand U8541 (N_8541,N_8279,N_8341);
and U8542 (N_8542,N_8328,N_8326);
or U8543 (N_8543,N_8485,N_8404);
nand U8544 (N_8544,N_8494,N_8424);
xnor U8545 (N_8545,N_8256,N_8453);
nor U8546 (N_8546,N_8446,N_8406);
and U8547 (N_8547,N_8461,N_8411);
or U8548 (N_8548,N_8357,N_8312);
nor U8549 (N_8549,N_8264,N_8283);
or U8550 (N_8550,N_8432,N_8417);
or U8551 (N_8551,N_8497,N_8332);
nand U8552 (N_8552,N_8344,N_8449);
xnor U8553 (N_8553,N_8423,N_8261);
and U8554 (N_8554,N_8258,N_8387);
or U8555 (N_8555,N_8393,N_8354);
nand U8556 (N_8556,N_8324,N_8441);
or U8557 (N_8557,N_8313,N_8251);
nor U8558 (N_8558,N_8301,N_8472);
nand U8559 (N_8559,N_8352,N_8265);
or U8560 (N_8560,N_8362,N_8463);
or U8561 (N_8561,N_8474,N_8331);
xnor U8562 (N_8562,N_8260,N_8273);
xnor U8563 (N_8563,N_8262,N_8381);
or U8564 (N_8564,N_8457,N_8360);
nand U8565 (N_8565,N_8338,N_8405);
xor U8566 (N_8566,N_8369,N_8276);
or U8567 (N_8567,N_8347,N_8380);
xor U8568 (N_8568,N_8459,N_8430);
nor U8569 (N_8569,N_8348,N_8408);
and U8570 (N_8570,N_8479,N_8436);
nor U8571 (N_8571,N_8490,N_8447);
nand U8572 (N_8572,N_8297,N_8475);
or U8573 (N_8573,N_8416,N_8323);
and U8574 (N_8574,N_8455,N_8482);
nor U8575 (N_8575,N_8367,N_8333);
nand U8576 (N_8576,N_8275,N_8319);
xor U8577 (N_8577,N_8278,N_8358);
or U8578 (N_8578,N_8372,N_8365);
xnor U8579 (N_8579,N_8292,N_8422);
nor U8580 (N_8580,N_8293,N_8402);
nand U8581 (N_8581,N_8414,N_8451);
xor U8582 (N_8582,N_8270,N_8299);
or U8583 (N_8583,N_8290,N_8443);
nand U8584 (N_8584,N_8308,N_8378);
xor U8585 (N_8585,N_8477,N_8281);
and U8586 (N_8586,N_8368,N_8394);
and U8587 (N_8587,N_8426,N_8488);
or U8588 (N_8588,N_8300,N_8382);
nor U8589 (N_8589,N_8493,N_8484);
xnor U8590 (N_8590,N_8266,N_8351);
xor U8591 (N_8591,N_8410,N_8350);
xor U8592 (N_8592,N_8413,N_8486);
nand U8593 (N_8593,N_8254,N_8370);
or U8594 (N_8594,N_8356,N_8487);
and U8595 (N_8595,N_8392,N_8429);
nor U8596 (N_8596,N_8314,N_8294);
nand U8597 (N_8597,N_8391,N_8491);
or U8598 (N_8598,N_8439,N_8315);
or U8599 (N_8599,N_8346,N_8466);
or U8600 (N_8600,N_8483,N_8473);
nor U8601 (N_8601,N_8458,N_8263);
xnor U8602 (N_8602,N_8444,N_8337);
or U8603 (N_8603,N_8316,N_8420);
or U8604 (N_8604,N_8252,N_8282);
nor U8605 (N_8605,N_8371,N_8467);
nand U8606 (N_8606,N_8355,N_8306);
and U8607 (N_8607,N_8303,N_8471);
nor U8608 (N_8608,N_8330,N_8418);
or U8609 (N_8609,N_8269,N_8359);
xor U8610 (N_8610,N_8431,N_8415);
nor U8611 (N_8611,N_8317,N_8321);
xnor U8612 (N_8612,N_8421,N_8295);
nand U8613 (N_8613,N_8425,N_8456);
nor U8614 (N_8614,N_8440,N_8499);
nor U8615 (N_8615,N_8450,N_8478);
or U8616 (N_8616,N_8296,N_8427);
xnor U8617 (N_8617,N_8280,N_8284);
and U8618 (N_8618,N_8255,N_8335);
nand U8619 (N_8619,N_8454,N_8329);
nand U8620 (N_8620,N_8398,N_8376);
nand U8621 (N_8621,N_8274,N_8310);
xor U8622 (N_8622,N_8396,N_8400);
nor U8623 (N_8623,N_8401,N_8384);
nand U8624 (N_8624,N_8462,N_8397);
nor U8625 (N_8625,N_8384,N_8456);
nor U8626 (N_8626,N_8487,N_8471);
and U8627 (N_8627,N_8347,N_8423);
or U8628 (N_8628,N_8373,N_8455);
nor U8629 (N_8629,N_8319,N_8368);
nor U8630 (N_8630,N_8350,N_8401);
nor U8631 (N_8631,N_8491,N_8483);
nand U8632 (N_8632,N_8288,N_8270);
nand U8633 (N_8633,N_8325,N_8456);
xor U8634 (N_8634,N_8355,N_8278);
nor U8635 (N_8635,N_8481,N_8379);
or U8636 (N_8636,N_8494,N_8425);
or U8637 (N_8637,N_8417,N_8265);
or U8638 (N_8638,N_8354,N_8359);
or U8639 (N_8639,N_8290,N_8260);
or U8640 (N_8640,N_8293,N_8429);
xnor U8641 (N_8641,N_8349,N_8396);
xor U8642 (N_8642,N_8358,N_8329);
nor U8643 (N_8643,N_8311,N_8283);
xor U8644 (N_8644,N_8416,N_8415);
and U8645 (N_8645,N_8477,N_8432);
xor U8646 (N_8646,N_8329,N_8403);
or U8647 (N_8647,N_8474,N_8307);
nand U8648 (N_8648,N_8379,N_8422);
nor U8649 (N_8649,N_8363,N_8422);
nand U8650 (N_8650,N_8300,N_8472);
and U8651 (N_8651,N_8441,N_8481);
and U8652 (N_8652,N_8463,N_8385);
nor U8653 (N_8653,N_8496,N_8325);
nand U8654 (N_8654,N_8393,N_8310);
nand U8655 (N_8655,N_8480,N_8256);
or U8656 (N_8656,N_8395,N_8479);
xor U8657 (N_8657,N_8342,N_8415);
and U8658 (N_8658,N_8385,N_8276);
nor U8659 (N_8659,N_8442,N_8383);
nand U8660 (N_8660,N_8299,N_8466);
and U8661 (N_8661,N_8415,N_8344);
and U8662 (N_8662,N_8409,N_8426);
and U8663 (N_8663,N_8393,N_8384);
nor U8664 (N_8664,N_8490,N_8252);
or U8665 (N_8665,N_8474,N_8403);
or U8666 (N_8666,N_8302,N_8266);
xor U8667 (N_8667,N_8493,N_8489);
or U8668 (N_8668,N_8492,N_8417);
or U8669 (N_8669,N_8331,N_8481);
or U8670 (N_8670,N_8260,N_8271);
or U8671 (N_8671,N_8291,N_8477);
or U8672 (N_8672,N_8401,N_8456);
nor U8673 (N_8673,N_8381,N_8324);
and U8674 (N_8674,N_8388,N_8257);
xnor U8675 (N_8675,N_8335,N_8455);
or U8676 (N_8676,N_8442,N_8498);
nand U8677 (N_8677,N_8440,N_8269);
and U8678 (N_8678,N_8347,N_8375);
nor U8679 (N_8679,N_8434,N_8265);
xnor U8680 (N_8680,N_8271,N_8383);
and U8681 (N_8681,N_8491,N_8383);
or U8682 (N_8682,N_8309,N_8436);
nor U8683 (N_8683,N_8308,N_8272);
or U8684 (N_8684,N_8418,N_8487);
nand U8685 (N_8685,N_8392,N_8474);
nand U8686 (N_8686,N_8433,N_8290);
or U8687 (N_8687,N_8406,N_8326);
nand U8688 (N_8688,N_8254,N_8413);
or U8689 (N_8689,N_8498,N_8330);
and U8690 (N_8690,N_8391,N_8446);
nand U8691 (N_8691,N_8441,N_8289);
nor U8692 (N_8692,N_8396,N_8323);
xor U8693 (N_8693,N_8274,N_8426);
xor U8694 (N_8694,N_8401,N_8479);
nor U8695 (N_8695,N_8306,N_8411);
nor U8696 (N_8696,N_8449,N_8315);
and U8697 (N_8697,N_8469,N_8433);
xnor U8698 (N_8698,N_8463,N_8333);
nor U8699 (N_8699,N_8399,N_8368);
nor U8700 (N_8700,N_8262,N_8317);
xor U8701 (N_8701,N_8379,N_8409);
xor U8702 (N_8702,N_8286,N_8298);
xnor U8703 (N_8703,N_8372,N_8445);
xnor U8704 (N_8704,N_8488,N_8409);
nor U8705 (N_8705,N_8408,N_8251);
or U8706 (N_8706,N_8484,N_8302);
xnor U8707 (N_8707,N_8425,N_8356);
or U8708 (N_8708,N_8480,N_8359);
and U8709 (N_8709,N_8309,N_8390);
or U8710 (N_8710,N_8399,N_8483);
nor U8711 (N_8711,N_8370,N_8439);
xor U8712 (N_8712,N_8457,N_8357);
nor U8713 (N_8713,N_8406,N_8464);
nand U8714 (N_8714,N_8361,N_8352);
or U8715 (N_8715,N_8491,N_8424);
and U8716 (N_8716,N_8434,N_8486);
or U8717 (N_8717,N_8322,N_8294);
xnor U8718 (N_8718,N_8336,N_8434);
nand U8719 (N_8719,N_8283,N_8352);
or U8720 (N_8720,N_8309,N_8417);
nor U8721 (N_8721,N_8324,N_8404);
xor U8722 (N_8722,N_8366,N_8499);
and U8723 (N_8723,N_8348,N_8434);
nand U8724 (N_8724,N_8299,N_8298);
and U8725 (N_8725,N_8407,N_8415);
and U8726 (N_8726,N_8267,N_8272);
and U8727 (N_8727,N_8423,N_8497);
xnor U8728 (N_8728,N_8295,N_8348);
xnor U8729 (N_8729,N_8304,N_8472);
nor U8730 (N_8730,N_8429,N_8273);
or U8731 (N_8731,N_8403,N_8251);
xnor U8732 (N_8732,N_8349,N_8416);
and U8733 (N_8733,N_8295,N_8388);
and U8734 (N_8734,N_8291,N_8287);
nor U8735 (N_8735,N_8336,N_8358);
xor U8736 (N_8736,N_8482,N_8444);
and U8737 (N_8737,N_8412,N_8400);
and U8738 (N_8738,N_8421,N_8346);
xor U8739 (N_8739,N_8463,N_8370);
or U8740 (N_8740,N_8479,N_8261);
xnor U8741 (N_8741,N_8258,N_8305);
nand U8742 (N_8742,N_8491,N_8420);
or U8743 (N_8743,N_8310,N_8489);
nand U8744 (N_8744,N_8419,N_8340);
xnor U8745 (N_8745,N_8336,N_8316);
nand U8746 (N_8746,N_8333,N_8338);
nand U8747 (N_8747,N_8485,N_8465);
and U8748 (N_8748,N_8364,N_8257);
or U8749 (N_8749,N_8370,N_8419);
or U8750 (N_8750,N_8505,N_8700);
nand U8751 (N_8751,N_8642,N_8509);
nand U8752 (N_8752,N_8687,N_8574);
xor U8753 (N_8753,N_8726,N_8660);
nand U8754 (N_8754,N_8556,N_8522);
nand U8755 (N_8755,N_8667,N_8537);
xnor U8756 (N_8756,N_8547,N_8518);
nor U8757 (N_8757,N_8592,N_8539);
and U8758 (N_8758,N_8723,N_8521);
or U8759 (N_8759,N_8631,N_8729);
nor U8760 (N_8760,N_8719,N_8678);
and U8761 (N_8761,N_8571,N_8581);
nand U8762 (N_8762,N_8689,N_8637);
and U8763 (N_8763,N_8665,N_8559);
xor U8764 (N_8764,N_8683,N_8705);
or U8765 (N_8765,N_8652,N_8595);
and U8766 (N_8766,N_8638,N_8711);
nand U8767 (N_8767,N_8557,N_8546);
or U8768 (N_8768,N_8603,N_8658);
xor U8769 (N_8769,N_8702,N_8610);
or U8770 (N_8770,N_8746,N_8629);
xor U8771 (N_8771,N_8523,N_8675);
or U8772 (N_8772,N_8730,N_8524);
xor U8773 (N_8773,N_8500,N_8623);
nand U8774 (N_8774,N_8715,N_8601);
or U8775 (N_8775,N_8604,N_8747);
and U8776 (N_8776,N_8618,N_8538);
and U8777 (N_8777,N_8517,N_8591);
and U8778 (N_8778,N_8632,N_8575);
nand U8779 (N_8779,N_8616,N_8553);
and U8780 (N_8780,N_8731,N_8541);
and U8781 (N_8781,N_8703,N_8606);
and U8782 (N_8782,N_8662,N_8691);
or U8783 (N_8783,N_8635,N_8664);
xor U8784 (N_8784,N_8596,N_8572);
or U8785 (N_8785,N_8657,N_8584);
nor U8786 (N_8786,N_8552,N_8578);
or U8787 (N_8787,N_8636,N_8607);
or U8788 (N_8788,N_8513,N_8716);
xor U8789 (N_8789,N_8542,N_8706);
and U8790 (N_8790,N_8699,N_8644);
nand U8791 (N_8791,N_8551,N_8588);
nor U8792 (N_8792,N_8520,N_8564);
nand U8793 (N_8793,N_8554,N_8555);
nand U8794 (N_8794,N_8531,N_8686);
or U8795 (N_8795,N_8568,N_8580);
nand U8796 (N_8796,N_8736,N_8621);
and U8797 (N_8797,N_8530,N_8680);
or U8798 (N_8798,N_8504,N_8684);
nand U8799 (N_8799,N_8708,N_8615);
xor U8800 (N_8800,N_8620,N_8685);
or U8801 (N_8801,N_8676,N_8614);
nor U8802 (N_8802,N_8690,N_8516);
xnor U8803 (N_8803,N_8749,N_8647);
nor U8804 (N_8804,N_8672,N_8712);
or U8805 (N_8805,N_8668,N_8656);
nand U8806 (N_8806,N_8732,N_8694);
and U8807 (N_8807,N_8728,N_8720);
nand U8808 (N_8808,N_8589,N_8501);
nor U8809 (N_8809,N_8585,N_8593);
nand U8810 (N_8810,N_8558,N_8645);
or U8811 (N_8811,N_8677,N_8561);
or U8812 (N_8812,N_8543,N_8602);
or U8813 (N_8813,N_8718,N_8735);
and U8814 (N_8814,N_8506,N_8669);
nor U8815 (N_8815,N_8682,N_8624);
xnor U8816 (N_8816,N_8560,N_8533);
and U8817 (N_8817,N_8740,N_8653);
xor U8818 (N_8818,N_8649,N_8577);
and U8819 (N_8819,N_8650,N_8579);
xnor U8820 (N_8820,N_8654,N_8674);
or U8821 (N_8821,N_8704,N_8625);
xor U8822 (N_8822,N_8655,N_8534);
and U8823 (N_8823,N_8717,N_8576);
xnor U8824 (N_8824,N_8548,N_8748);
nand U8825 (N_8825,N_8527,N_8619);
nor U8826 (N_8826,N_8696,N_8605);
nor U8827 (N_8827,N_8651,N_8611);
and U8828 (N_8828,N_8695,N_8535);
and U8829 (N_8829,N_8598,N_8510);
xnor U8830 (N_8830,N_8525,N_8587);
xnor U8831 (N_8831,N_8663,N_8608);
nand U8832 (N_8832,N_8550,N_8633);
nand U8833 (N_8833,N_8640,N_8565);
or U8834 (N_8834,N_8670,N_8563);
and U8835 (N_8835,N_8528,N_8511);
nor U8836 (N_8836,N_8743,N_8582);
or U8837 (N_8837,N_8627,N_8724);
xor U8838 (N_8838,N_8681,N_8583);
nor U8839 (N_8839,N_8692,N_8661);
nor U8840 (N_8840,N_8721,N_8515);
or U8841 (N_8841,N_8566,N_8609);
xor U8842 (N_8842,N_8512,N_8710);
and U8843 (N_8843,N_8639,N_8722);
nand U8844 (N_8844,N_8714,N_8709);
nand U8845 (N_8845,N_8725,N_8713);
nand U8846 (N_8846,N_8626,N_8697);
and U8847 (N_8847,N_8540,N_8549);
xor U8848 (N_8848,N_8741,N_8529);
or U8849 (N_8849,N_8698,N_8745);
nor U8850 (N_8850,N_8648,N_8679);
nor U8851 (N_8851,N_8742,N_8634);
or U8852 (N_8852,N_8599,N_8536);
nor U8853 (N_8853,N_8600,N_8570);
nand U8854 (N_8854,N_8659,N_8590);
or U8855 (N_8855,N_8594,N_8503);
and U8856 (N_8856,N_8701,N_8507);
or U8857 (N_8857,N_8630,N_8628);
and U8858 (N_8858,N_8744,N_8707);
or U8859 (N_8859,N_8597,N_8622);
xnor U8860 (N_8860,N_8673,N_8567);
xor U8861 (N_8861,N_8526,N_8544);
nor U8862 (N_8862,N_8545,N_8586);
and U8863 (N_8863,N_8643,N_8532);
nor U8864 (N_8864,N_8519,N_8666);
and U8865 (N_8865,N_8502,N_8738);
and U8866 (N_8866,N_8739,N_8573);
and U8867 (N_8867,N_8508,N_8562);
nor U8868 (N_8868,N_8733,N_8569);
nor U8869 (N_8869,N_8734,N_8737);
nand U8870 (N_8870,N_8612,N_8617);
or U8871 (N_8871,N_8671,N_8693);
nor U8872 (N_8872,N_8641,N_8688);
nor U8873 (N_8873,N_8613,N_8646);
xor U8874 (N_8874,N_8514,N_8727);
nand U8875 (N_8875,N_8553,N_8726);
and U8876 (N_8876,N_8538,N_8686);
xnor U8877 (N_8877,N_8584,N_8554);
and U8878 (N_8878,N_8515,N_8550);
xnor U8879 (N_8879,N_8645,N_8698);
and U8880 (N_8880,N_8618,N_8709);
nor U8881 (N_8881,N_8599,N_8573);
and U8882 (N_8882,N_8585,N_8564);
or U8883 (N_8883,N_8741,N_8631);
nand U8884 (N_8884,N_8554,N_8607);
nand U8885 (N_8885,N_8682,N_8652);
and U8886 (N_8886,N_8588,N_8705);
and U8887 (N_8887,N_8500,N_8676);
nor U8888 (N_8888,N_8625,N_8639);
or U8889 (N_8889,N_8673,N_8709);
nor U8890 (N_8890,N_8745,N_8639);
nor U8891 (N_8891,N_8526,N_8580);
or U8892 (N_8892,N_8718,N_8699);
nand U8893 (N_8893,N_8651,N_8587);
nor U8894 (N_8894,N_8602,N_8680);
and U8895 (N_8895,N_8735,N_8566);
nor U8896 (N_8896,N_8620,N_8584);
or U8897 (N_8897,N_8569,N_8576);
xnor U8898 (N_8898,N_8539,N_8657);
nor U8899 (N_8899,N_8699,N_8743);
xor U8900 (N_8900,N_8658,N_8541);
nand U8901 (N_8901,N_8718,N_8509);
and U8902 (N_8902,N_8730,N_8542);
xnor U8903 (N_8903,N_8615,N_8510);
xor U8904 (N_8904,N_8569,N_8564);
nand U8905 (N_8905,N_8541,N_8720);
and U8906 (N_8906,N_8529,N_8618);
xor U8907 (N_8907,N_8639,N_8589);
nor U8908 (N_8908,N_8709,N_8639);
and U8909 (N_8909,N_8637,N_8701);
nand U8910 (N_8910,N_8714,N_8684);
xor U8911 (N_8911,N_8526,N_8730);
or U8912 (N_8912,N_8711,N_8674);
and U8913 (N_8913,N_8511,N_8652);
or U8914 (N_8914,N_8565,N_8635);
or U8915 (N_8915,N_8595,N_8577);
or U8916 (N_8916,N_8698,N_8670);
and U8917 (N_8917,N_8719,N_8706);
or U8918 (N_8918,N_8569,N_8708);
xnor U8919 (N_8919,N_8711,N_8624);
and U8920 (N_8920,N_8577,N_8714);
nand U8921 (N_8921,N_8589,N_8527);
nor U8922 (N_8922,N_8615,N_8743);
or U8923 (N_8923,N_8514,N_8742);
xor U8924 (N_8924,N_8747,N_8530);
nand U8925 (N_8925,N_8507,N_8512);
nand U8926 (N_8926,N_8531,N_8649);
nand U8927 (N_8927,N_8734,N_8572);
and U8928 (N_8928,N_8709,N_8579);
or U8929 (N_8929,N_8641,N_8668);
nand U8930 (N_8930,N_8648,N_8675);
or U8931 (N_8931,N_8693,N_8508);
or U8932 (N_8932,N_8507,N_8553);
and U8933 (N_8933,N_8732,N_8609);
nand U8934 (N_8934,N_8574,N_8536);
nor U8935 (N_8935,N_8703,N_8677);
nand U8936 (N_8936,N_8592,N_8504);
or U8937 (N_8937,N_8522,N_8617);
xor U8938 (N_8938,N_8549,N_8524);
nor U8939 (N_8939,N_8671,N_8634);
or U8940 (N_8940,N_8545,N_8683);
nor U8941 (N_8941,N_8673,N_8514);
and U8942 (N_8942,N_8629,N_8668);
or U8943 (N_8943,N_8526,N_8616);
or U8944 (N_8944,N_8643,N_8522);
xor U8945 (N_8945,N_8702,N_8698);
xnor U8946 (N_8946,N_8512,N_8522);
xnor U8947 (N_8947,N_8700,N_8605);
nor U8948 (N_8948,N_8658,N_8534);
nand U8949 (N_8949,N_8587,N_8674);
or U8950 (N_8950,N_8747,N_8647);
and U8951 (N_8951,N_8511,N_8635);
or U8952 (N_8952,N_8500,N_8713);
xnor U8953 (N_8953,N_8554,N_8559);
or U8954 (N_8954,N_8647,N_8712);
nor U8955 (N_8955,N_8697,N_8678);
nand U8956 (N_8956,N_8588,N_8671);
xor U8957 (N_8957,N_8625,N_8737);
or U8958 (N_8958,N_8519,N_8741);
xor U8959 (N_8959,N_8663,N_8701);
or U8960 (N_8960,N_8688,N_8627);
or U8961 (N_8961,N_8510,N_8578);
or U8962 (N_8962,N_8652,N_8555);
nand U8963 (N_8963,N_8503,N_8653);
and U8964 (N_8964,N_8623,N_8732);
xor U8965 (N_8965,N_8553,N_8724);
nor U8966 (N_8966,N_8529,N_8513);
xnor U8967 (N_8967,N_8715,N_8626);
nor U8968 (N_8968,N_8507,N_8673);
nand U8969 (N_8969,N_8580,N_8745);
or U8970 (N_8970,N_8528,N_8653);
nand U8971 (N_8971,N_8505,N_8678);
nor U8972 (N_8972,N_8568,N_8720);
or U8973 (N_8973,N_8591,N_8638);
nor U8974 (N_8974,N_8555,N_8657);
nor U8975 (N_8975,N_8696,N_8738);
nand U8976 (N_8976,N_8542,N_8552);
xnor U8977 (N_8977,N_8701,N_8600);
nor U8978 (N_8978,N_8739,N_8512);
nand U8979 (N_8979,N_8555,N_8597);
nor U8980 (N_8980,N_8627,N_8653);
or U8981 (N_8981,N_8519,N_8571);
xnor U8982 (N_8982,N_8544,N_8575);
or U8983 (N_8983,N_8544,N_8635);
nor U8984 (N_8984,N_8647,N_8696);
nand U8985 (N_8985,N_8570,N_8598);
or U8986 (N_8986,N_8585,N_8748);
nand U8987 (N_8987,N_8517,N_8544);
and U8988 (N_8988,N_8660,N_8625);
nor U8989 (N_8989,N_8656,N_8623);
or U8990 (N_8990,N_8561,N_8509);
nand U8991 (N_8991,N_8640,N_8501);
and U8992 (N_8992,N_8525,N_8559);
nor U8993 (N_8993,N_8509,N_8503);
nand U8994 (N_8994,N_8658,N_8517);
or U8995 (N_8995,N_8508,N_8573);
xor U8996 (N_8996,N_8605,N_8681);
or U8997 (N_8997,N_8652,N_8627);
nand U8998 (N_8998,N_8734,N_8749);
nand U8999 (N_8999,N_8675,N_8599);
or U9000 (N_9000,N_8909,N_8971);
xnor U9001 (N_9001,N_8860,N_8756);
and U9002 (N_9002,N_8919,N_8799);
nand U9003 (N_9003,N_8849,N_8961);
and U9004 (N_9004,N_8975,N_8892);
xor U9005 (N_9005,N_8783,N_8894);
and U9006 (N_9006,N_8808,N_8788);
xor U9007 (N_9007,N_8811,N_8801);
nand U9008 (N_9008,N_8882,N_8976);
xor U9009 (N_9009,N_8965,N_8809);
xnor U9010 (N_9010,N_8934,N_8914);
nand U9011 (N_9011,N_8873,N_8956);
or U9012 (N_9012,N_8770,N_8985);
or U9013 (N_9013,N_8939,N_8883);
xor U9014 (N_9014,N_8822,N_8853);
nand U9015 (N_9015,N_8871,N_8750);
or U9016 (N_9016,N_8780,N_8893);
or U9017 (N_9017,N_8998,N_8837);
or U9018 (N_9018,N_8765,N_8823);
xor U9019 (N_9019,N_8784,N_8973);
or U9020 (N_9020,N_8833,N_8997);
nor U9021 (N_9021,N_8898,N_8854);
nand U9022 (N_9022,N_8758,N_8754);
nand U9023 (N_9023,N_8847,N_8793);
or U9024 (N_9024,N_8879,N_8974);
nor U9025 (N_9025,N_8922,N_8924);
xnor U9026 (N_9026,N_8995,N_8928);
and U9027 (N_9027,N_8766,N_8941);
nor U9028 (N_9028,N_8960,N_8864);
and U9029 (N_9029,N_8888,N_8778);
nor U9030 (N_9030,N_8927,N_8987);
nor U9031 (N_9031,N_8870,N_8897);
nand U9032 (N_9032,N_8910,N_8918);
or U9033 (N_9033,N_8805,N_8906);
or U9034 (N_9034,N_8986,N_8978);
xnor U9035 (N_9035,N_8787,N_8966);
nand U9036 (N_9036,N_8830,N_8955);
nand U9037 (N_9037,N_8814,N_8962);
or U9038 (N_9038,N_8921,N_8845);
nand U9039 (N_9039,N_8862,N_8948);
xor U9040 (N_9040,N_8872,N_8957);
xnor U9041 (N_9041,N_8877,N_8929);
nand U9042 (N_9042,N_8803,N_8856);
and U9043 (N_9043,N_8861,N_8838);
or U9044 (N_9044,N_8775,N_8869);
or U9045 (N_9045,N_8797,N_8958);
or U9046 (N_9046,N_8984,N_8874);
nor U9047 (N_9047,N_8900,N_8891);
and U9048 (N_9048,N_8990,N_8970);
or U9049 (N_9049,N_8846,N_8887);
or U9050 (N_9050,N_8881,N_8959);
or U9051 (N_9051,N_8800,N_8826);
xor U9052 (N_9052,N_8824,N_8867);
nand U9053 (N_9053,N_8949,N_8968);
nand U9054 (N_9054,N_8991,N_8762);
nand U9055 (N_9055,N_8777,N_8875);
xnor U9056 (N_9056,N_8821,N_8763);
nor U9057 (N_9057,N_8781,N_8753);
or U9058 (N_9058,N_8884,N_8905);
nor U9059 (N_9059,N_8851,N_8908);
nand U9060 (N_9060,N_8930,N_8913);
nand U9061 (N_9061,N_8752,N_8768);
and U9062 (N_9062,N_8802,N_8992);
or U9063 (N_9063,N_8795,N_8946);
and U9064 (N_9064,N_8932,N_8977);
nand U9065 (N_9065,N_8843,N_8996);
or U9066 (N_9066,N_8755,N_8764);
nand U9067 (N_9067,N_8767,N_8865);
and U9068 (N_9068,N_8896,N_8828);
or U9069 (N_9069,N_8967,N_8885);
nor U9070 (N_9070,N_8831,N_8989);
or U9071 (N_9071,N_8839,N_8840);
or U9072 (N_9072,N_8857,N_8848);
nor U9073 (N_9073,N_8776,N_8931);
nor U9074 (N_9074,N_8940,N_8771);
or U9075 (N_9075,N_8911,N_8993);
xnor U9076 (N_9076,N_8850,N_8842);
nor U9077 (N_9077,N_8926,N_8855);
nor U9078 (N_9078,N_8785,N_8816);
nor U9079 (N_9079,N_8827,N_8904);
or U9080 (N_9080,N_8792,N_8912);
or U9081 (N_9081,N_8943,N_8980);
nand U9082 (N_9082,N_8760,N_8901);
nand U9083 (N_9083,N_8773,N_8751);
xor U9084 (N_9084,N_8988,N_8925);
nand U9085 (N_9085,N_8806,N_8804);
and U9086 (N_9086,N_8945,N_8817);
xnor U9087 (N_9087,N_8915,N_8944);
nor U9088 (N_9088,N_8963,N_8972);
nand U9089 (N_9089,N_8994,N_8815);
or U9090 (N_9090,N_8825,N_8829);
xor U9091 (N_9091,N_8789,N_8836);
or U9092 (N_9092,N_8841,N_8886);
or U9093 (N_9093,N_8791,N_8880);
nand U9094 (N_9094,N_8757,N_8933);
nor U9095 (N_9095,N_8923,N_8794);
and U9096 (N_9096,N_8761,N_8798);
xor U9097 (N_9097,N_8951,N_8890);
xor U9098 (N_9098,N_8902,N_8920);
and U9099 (N_9099,N_8935,N_8999);
xnor U9100 (N_9100,N_8868,N_8813);
and U9101 (N_9101,N_8952,N_8863);
or U9102 (N_9102,N_8899,N_8782);
nor U9103 (N_9103,N_8832,N_8796);
and U9104 (N_9104,N_8917,N_8969);
nand U9105 (N_9105,N_8954,N_8866);
nor U9106 (N_9106,N_8947,N_8979);
nand U9107 (N_9107,N_8876,N_8772);
or U9108 (N_9108,N_8895,N_8759);
and U9109 (N_9109,N_8982,N_8953);
nor U9110 (N_9110,N_8818,N_8950);
nor U9111 (N_9111,N_8852,N_8878);
xnor U9112 (N_9112,N_8889,N_8812);
nand U9113 (N_9113,N_8820,N_8819);
nor U9114 (N_9114,N_8810,N_8936);
and U9115 (N_9115,N_8786,N_8835);
nor U9116 (N_9116,N_8938,N_8903);
nand U9117 (N_9117,N_8790,N_8844);
or U9118 (N_9118,N_8858,N_8859);
nand U9119 (N_9119,N_8942,N_8834);
and U9120 (N_9120,N_8807,N_8981);
and U9121 (N_9121,N_8916,N_8964);
and U9122 (N_9122,N_8937,N_8769);
or U9123 (N_9123,N_8774,N_8907);
nand U9124 (N_9124,N_8983,N_8779);
nand U9125 (N_9125,N_8827,N_8862);
xor U9126 (N_9126,N_8962,N_8941);
nand U9127 (N_9127,N_8968,N_8750);
nor U9128 (N_9128,N_8936,N_8813);
nand U9129 (N_9129,N_8878,N_8846);
nor U9130 (N_9130,N_8945,N_8873);
or U9131 (N_9131,N_8791,N_8885);
and U9132 (N_9132,N_8867,N_8924);
and U9133 (N_9133,N_8961,N_8915);
nor U9134 (N_9134,N_8773,N_8796);
or U9135 (N_9135,N_8859,N_8876);
and U9136 (N_9136,N_8920,N_8994);
xnor U9137 (N_9137,N_8964,N_8995);
nor U9138 (N_9138,N_8803,N_8770);
nor U9139 (N_9139,N_8847,N_8805);
nor U9140 (N_9140,N_8886,N_8893);
nor U9141 (N_9141,N_8785,N_8773);
nand U9142 (N_9142,N_8781,N_8876);
nor U9143 (N_9143,N_8958,N_8848);
or U9144 (N_9144,N_8909,N_8861);
xnor U9145 (N_9145,N_8967,N_8827);
nand U9146 (N_9146,N_8974,N_8806);
and U9147 (N_9147,N_8990,N_8789);
and U9148 (N_9148,N_8752,N_8791);
nand U9149 (N_9149,N_8957,N_8991);
or U9150 (N_9150,N_8917,N_8892);
or U9151 (N_9151,N_8971,N_8780);
nor U9152 (N_9152,N_8837,N_8787);
or U9153 (N_9153,N_8908,N_8926);
nand U9154 (N_9154,N_8766,N_8802);
and U9155 (N_9155,N_8893,N_8797);
nand U9156 (N_9156,N_8978,N_8998);
or U9157 (N_9157,N_8923,N_8763);
nor U9158 (N_9158,N_8832,N_8959);
xnor U9159 (N_9159,N_8950,N_8934);
xor U9160 (N_9160,N_8763,N_8978);
nand U9161 (N_9161,N_8980,N_8938);
xnor U9162 (N_9162,N_8753,N_8977);
or U9163 (N_9163,N_8783,N_8901);
xnor U9164 (N_9164,N_8949,N_8759);
nor U9165 (N_9165,N_8890,N_8855);
xnor U9166 (N_9166,N_8954,N_8763);
nor U9167 (N_9167,N_8768,N_8868);
nand U9168 (N_9168,N_8902,N_8976);
nand U9169 (N_9169,N_8803,N_8949);
nand U9170 (N_9170,N_8882,N_8885);
nor U9171 (N_9171,N_8964,N_8825);
or U9172 (N_9172,N_8923,N_8886);
or U9173 (N_9173,N_8801,N_8807);
xor U9174 (N_9174,N_8850,N_8908);
or U9175 (N_9175,N_8872,N_8834);
and U9176 (N_9176,N_8877,N_8892);
xor U9177 (N_9177,N_8923,N_8925);
or U9178 (N_9178,N_8900,N_8983);
nand U9179 (N_9179,N_8991,N_8820);
or U9180 (N_9180,N_8907,N_8891);
and U9181 (N_9181,N_8937,N_8830);
and U9182 (N_9182,N_8778,N_8865);
nand U9183 (N_9183,N_8959,N_8983);
xor U9184 (N_9184,N_8792,N_8854);
nor U9185 (N_9185,N_8997,N_8925);
or U9186 (N_9186,N_8934,N_8750);
nor U9187 (N_9187,N_8944,N_8765);
xnor U9188 (N_9188,N_8817,N_8840);
nand U9189 (N_9189,N_8994,N_8820);
nand U9190 (N_9190,N_8942,N_8763);
or U9191 (N_9191,N_8775,N_8968);
nand U9192 (N_9192,N_8800,N_8892);
or U9193 (N_9193,N_8945,N_8909);
nand U9194 (N_9194,N_8940,N_8881);
xnor U9195 (N_9195,N_8847,N_8777);
nor U9196 (N_9196,N_8792,N_8835);
or U9197 (N_9197,N_8958,N_8758);
nand U9198 (N_9198,N_8993,N_8847);
xor U9199 (N_9199,N_8843,N_8912);
nor U9200 (N_9200,N_8822,N_8793);
xor U9201 (N_9201,N_8851,N_8911);
and U9202 (N_9202,N_8787,N_8891);
nor U9203 (N_9203,N_8998,N_8850);
or U9204 (N_9204,N_8799,N_8867);
xor U9205 (N_9205,N_8900,N_8878);
nand U9206 (N_9206,N_8752,N_8778);
nor U9207 (N_9207,N_8917,N_8769);
or U9208 (N_9208,N_8760,N_8769);
nor U9209 (N_9209,N_8810,N_8771);
xnor U9210 (N_9210,N_8899,N_8948);
nor U9211 (N_9211,N_8922,N_8868);
nand U9212 (N_9212,N_8854,N_8756);
nand U9213 (N_9213,N_8984,N_8811);
nor U9214 (N_9214,N_8936,N_8902);
nor U9215 (N_9215,N_8808,N_8905);
xor U9216 (N_9216,N_8887,N_8882);
nand U9217 (N_9217,N_8836,N_8918);
nand U9218 (N_9218,N_8772,N_8883);
or U9219 (N_9219,N_8852,N_8978);
or U9220 (N_9220,N_8800,N_8942);
nor U9221 (N_9221,N_8919,N_8938);
nor U9222 (N_9222,N_8839,N_8814);
nand U9223 (N_9223,N_8949,N_8795);
nor U9224 (N_9224,N_8771,N_8925);
nor U9225 (N_9225,N_8750,N_8867);
xor U9226 (N_9226,N_8963,N_8806);
nor U9227 (N_9227,N_8860,N_8977);
or U9228 (N_9228,N_8989,N_8894);
and U9229 (N_9229,N_8762,N_8954);
nor U9230 (N_9230,N_8960,N_8879);
and U9231 (N_9231,N_8926,N_8782);
or U9232 (N_9232,N_8911,N_8949);
nor U9233 (N_9233,N_8837,N_8799);
nand U9234 (N_9234,N_8909,N_8821);
or U9235 (N_9235,N_8947,N_8978);
nand U9236 (N_9236,N_8842,N_8835);
or U9237 (N_9237,N_8825,N_8960);
or U9238 (N_9238,N_8890,N_8997);
xnor U9239 (N_9239,N_8892,N_8937);
or U9240 (N_9240,N_8847,N_8998);
nor U9241 (N_9241,N_8766,N_8903);
nand U9242 (N_9242,N_8951,N_8866);
xor U9243 (N_9243,N_8912,N_8752);
nor U9244 (N_9244,N_8895,N_8919);
xor U9245 (N_9245,N_8834,N_8832);
xnor U9246 (N_9246,N_8880,N_8836);
and U9247 (N_9247,N_8958,N_8795);
or U9248 (N_9248,N_8969,N_8977);
or U9249 (N_9249,N_8832,N_8991);
nand U9250 (N_9250,N_9176,N_9031);
xnor U9251 (N_9251,N_9116,N_9226);
or U9252 (N_9252,N_9187,N_9097);
xor U9253 (N_9253,N_9223,N_9208);
nor U9254 (N_9254,N_9067,N_9153);
and U9255 (N_9255,N_9183,N_9142);
xor U9256 (N_9256,N_9147,N_9089);
nor U9257 (N_9257,N_9242,N_9047);
and U9258 (N_9258,N_9109,N_9212);
or U9259 (N_9259,N_9201,N_9000);
or U9260 (N_9260,N_9209,N_9117);
xor U9261 (N_9261,N_9186,N_9100);
nor U9262 (N_9262,N_9001,N_9199);
or U9263 (N_9263,N_9177,N_9085);
xnor U9264 (N_9264,N_9235,N_9055);
and U9265 (N_9265,N_9137,N_9015);
xor U9266 (N_9266,N_9210,N_9146);
and U9267 (N_9267,N_9049,N_9114);
xnor U9268 (N_9268,N_9006,N_9019);
and U9269 (N_9269,N_9119,N_9014);
or U9270 (N_9270,N_9035,N_9038);
and U9271 (N_9271,N_9048,N_9057);
and U9272 (N_9272,N_9036,N_9082);
and U9273 (N_9273,N_9103,N_9196);
nand U9274 (N_9274,N_9012,N_9034);
nor U9275 (N_9275,N_9013,N_9213);
or U9276 (N_9276,N_9245,N_9053);
and U9277 (N_9277,N_9044,N_9219);
or U9278 (N_9278,N_9099,N_9132);
nor U9279 (N_9279,N_9064,N_9078);
nor U9280 (N_9280,N_9069,N_9152);
xor U9281 (N_9281,N_9131,N_9168);
and U9282 (N_9282,N_9096,N_9042);
nand U9283 (N_9283,N_9232,N_9225);
nand U9284 (N_9284,N_9198,N_9102);
nand U9285 (N_9285,N_9181,N_9243);
nand U9286 (N_9286,N_9138,N_9005);
nand U9287 (N_9287,N_9002,N_9238);
nand U9288 (N_9288,N_9237,N_9125);
nor U9289 (N_9289,N_9045,N_9113);
xnor U9290 (N_9290,N_9192,N_9091);
and U9291 (N_9291,N_9222,N_9018);
xnor U9292 (N_9292,N_9039,N_9028);
and U9293 (N_9293,N_9227,N_9108);
xnor U9294 (N_9294,N_9126,N_9093);
and U9295 (N_9295,N_9170,N_9065);
and U9296 (N_9296,N_9189,N_9083);
xor U9297 (N_9297,N_9180,N_9090);
nor U9298 (N_9298,N_9215,N_9094);
xor U9299 (N_9299,N_9111,N_9241);
nor U9300 (N_9300,N_9145,N_9249);
and U9301 (N_9301,N_9063,N_9188);
or U9302 (N_9302,N_9092,N_9071);
xor U9303 (N_9303,N_9139,N_9033);
nand U9304 (N_9304,N_9110,N_9229);
or U9305 (N_9305,N_9072,N_9007);
and U9306 (N_9306,N_9143,N_9204);
and U9307 (N_9307,N_9056,N_9163);
or U9308 (N_9308,N_9095,N_9112);
or U9309 (N_9309,N_9107,N_9160);
nand U9310 (N_9310,N_9123,N_9121);
nand U9311 (N_9311,N_9182,N_9133);
or U9312 (N_9312,N_9203,N_9068);
and U9313 (N_9313,N_9193,N_9076);
nor U9314 (N_9314,N_9003,N_9221);
or U9315 (N_9315,N_9043,N_9134);
nand U9316 (N_9316,N_9118,N_9009);
nand U9317 (N_9317,N_9171,N_9061);
xnor U9318 (N_9318,N_9054,N_9079);
nor U9319 (N_9319,N_9026,N_9140);
nand U9320 (N_9320,N_9244,N_9017);
and U9321 (N_9321,N_9141,N_9008);
xor U9322 (N_9322,N_9220,N_9080);
and U9323 (N_9323,N_9032,N_9173);
or U9324 (N_9324,N_9128,N_9024);
nand U9325 (N_9325,N_9016,N_9155);
and U9326 (N_9326,N_9217,N_9247);
xnor U9327 (N_9327,N_9151,N_9148);
or U9328 (N_9328,N_9185,N_9101);
or U9329 (N_9329,N_9234,N_9029);
nand U9330 (N_9330,N_9023,N_9156);
nand U9331 (N_9331,N_9073,N_9202);
or U9332 (N_9332,N_9154,N_9205);
and U9333 (N_9333,N_9030,N_9224);
nor U9334 (N_9334,N_9074,N_9246);
or U9335 (N_9335,N_9248,N_9240);
xor U9336 (N_9336,N_9086,N_9233);
nor U9337 (N_9337,N_9041,N_9127);
and U9338 (N_9338,N_9158,N_9236);
nor U9339 (N_9339,N_9070,N_9179);
nor U9340 (N_9340,N_9075,N_9051);
and U9341 (N_9341,N_9084,N_9169);
nand U9342 (N_9342,N_9011,N_9060);
nand U9343 (N_9343,N_9159,N_9228);
nor U9344 (N_9344,N_9066,N_9010);
or U9345 (N_9345,N_9120,N_9037);
and U9346 (N_9346,N_9175,N_9115);
xor U9347 (N_9347,N_9178,N_9214);
and U9348 (N_9348,N_9239,N_9122);
nor U9349 (N_9349,N_9194,N_9218);
xnor U9350 (N_9350,N_9129,N_9197);
nor U9351 (N_9351,N_9207,N_9191);
nor U9352 (N_9352,N_9166,N_9020);
or U9353 (N_9353,N_9195,N_9081);
nor U9354 (N_9354,N_9062,N_9136);
xnor U9355 (N_9355,N_9206,N_9150);
nor U9356 (N_9356,N_9230,N_9104);
and U9357 (N_9357,N_9022,N_9164);
and U9358 (N_9358,N_9046,N_9087);
or U9359 (N_9359,N_9124,N_9098);
and U9360 (N_9360,N_9040,N_9021);
nor U9361 (N_9361,N_9050,N_9004);
nand U9362 (N_9362,N_9231,N_9216);
nand U9363 (N_9363,N_9157,N_9174);
nor U9364 (N_9364,N_9135,N_9165);
nand U9365 (N_9365,N_9184,N_9149);
nor U9366 (N_9366,N_9130,N_9162);
nor U9367 (N_9367,N_9144,N_9172);
nand U9368 (N_9368,N_9211,N_9077);
and U9369 (N_9369,N_9200,N_9167);
nor U9370 (N_9370,N_9106,N_9025);
and U9371 (N_9371,N_9105,N_9052);
nand U9372 (N_9372,N_9027,N_9161);
xnor U9373 (N_9373,N_9059,N_9190);
or U9374 (N_9374,N_9058,N_9088);
nand U9375 (N_9375,N_9125,N_9193);
xor U9376 (N_9376,N_9160,N_9053);
nor U9377 (N_9377,N_9096,N_9203);
nand U9378 (N_9378,N_9229,N_9130);
nand U9379 (N_9379,N_9189,N_9208);
and U9380 (N_9380,N_9171,N_9082);
xor U9381 (N_9381,N_9033,N_9246);
or U9382 (N_9382,N_9004,N_9059);
and U9383 (N_9383,N_9021,N_9246);
xor U9384 (N_9384,N_9130,N_9147);
nor U9385 (N_9385,N_9007,N_9193);
nor U9386 (N_9386,N_9095,N_9105);
nor U9387 (N_9387,N_9233,N_9188);
and U9388 (N_9388,N_9009,N_9086);
or U9389 (N_9389,N_9249,N_9191);
xnor U9390 (N_9390,N_9206,N_9107);
and U9391 (N_9391,N_9099,N_9067);
and U9392 (N_9392,N_9020,N_9151);
nand U9393 (N_9393,N_9237,N_9119);
nand U9394 (N_9394,N_9046,N_9086);
and U9395 (N_9395,N_9240,N_9165);
and U9396 (N_9396,N_9144,N_9152);
nor U9397 (N_9397,N_9247,N_9237);
xor U9398 (N_9398,N_9015,N_9234);
or U9399 (N_9399,N_9159,N_9058);
and U9400 (N_9400,N_9156,N_9130);
xor U9401 (N_9401,N_9113,N_9084);
or U9402 (N_9402,N_9002,N_9107);
nor U9403 (N_9403,N_9125,N_9192);
nor U9404 (N_9404,N_9223,N_9109);
and U9405 (N_9405,N_9213,N_9248);
xnor U9406 (N_9406,N_9073,N_9031);
and U9407 (N_9407,N_9247,N_9121);
or U9408 (N_9408,N_9037,N_9096);
nor U9409 (N_9409,N_9236,N_9244);
nor U9410 (N_9410,N_9016,N_9018);
and U9411 (N_9411,N_9004,N_9214);
nand U9412 (N_9412,N_9228,N_9139);
nor U9413 (N_9413,N_9162,N_9122);
and U9414 (N_9414,N_9244,N_9221);
nor U9415 (N_9415,N_9166,N_9207);
xnor U9416 (N_9416,N_9209,N_9119);
nand U9417 (N_9417,N_9034,N_9133);
nor U9418 (N_9418,N_9116,N_9169);
and U9419 (N_9419,N_9079,N_9070);
or U9420 (N_9420,N_9003,N_9049);
nand U9421 (N_9421,N_9182,N_9191);
and U9422 (N_9422,N_9125,N_9011);
and U9423 (N_9423,N_9181,N_9096);
xor U9424 (N_9424,N_9196,N_9040);
xnor U9425 (N_9425,N_9236,N_9091);
nand U9426 (N_9426,N_9243,N_9215);
and U9427 (N_9427,N_9124,N_9182);
or U9428 (N_9428,N_9187,N_9209);
and U9429 (N_9429,N_9243,N_9132);
nor U9430 (N_9430,N_9198,N_9004);
nor U9431 (N_9431,N_9117,N_9242);
nor U9432 (N_9432,N_9217,N_9139);
nor U9433 (N_9433,N_9213,N_9005);
and U9434 (N_9434,N_9011,N_9184);
and U9435 (N_9435,N_9049,N_9181);
and U9436 (N_9436,N_9164,N_9004);
nand U9437 (N_9437,N_9153,N_9147);
nor U9438 (N_9438,N_9084,N_9075);
xnor U9439 (N_9439,N_9009,N_9126);
xnor U9440 (N_9440,N_9037,N_9063);
and U9441 (N_9441,N_9214,N_9204);
and U9442 (N_9442,N_9044,N_9101);
and U9443 (N_9443,N_9236,N_9008);
nor U9444 (N_9444,N_9095,N_9015);
nor U9445 (N_9445,N_9239,N_9201);
nand U9446 (N_9446,N_9006,N_9155);
nor U9447 (N_9447,N_9220,N_9072);
nand U9448 (N_9448,N_9009,N_9236);
nor U9449 (N_9449,N_9129,N_9037);
and U9450 (N_9450,N_9060,N_9067);
nor U9451 (N_9451,N_9049,N_9092);
and U9452 (N_9452,N_9093,N_9105);
nand U9453 (N_9453,N_9216,N_9104);
xor U9454 (N_9454,N_9244,N_9010);
or U9455 (N_9455,N_9124,N_9131);
and U9456 (N_9456,N_9187,N_9170);
xor U9457 (N_9457,N_9126,N_9060);
xor U9458 (N_9458,N_9038,N_9225);
or U9459 (N_9459,N_9174,N_9056);
nor U9460 (N_9460,N_9227,N_9137);
or U9461 (N_9461,N_9072,N_9164);
and U9462 (N_9462,N_9189,N_9146);
or U9463 (N_9463,N_9147,N_9177);
or U9464 (N_9464,N_9031,N_9113);
nand U9465 (N_9465,N_9110,N_9066);
xnor U9466 (N_9466,N_9083,N_9118);
nand U9467 (N_9467,N_9156,N_9057);
and U9468 (N_9468,N_9038,N_9090);
or U9469 (N_9469,N_9096,N_9010);
or U9470 (N_9470,N_9048,N_9197);
xnor U9471 (N_9471,N_9143,N_9232);
or U9472 (N_9472,N_9198,N_9030);
nor U9473 (N_9473,N_9079,N_9113);
and U9474 (N_9474,N_9064,N_9023);
nand U9475 (N_9475,N_9212,N_9169);
nor U9476 (N_9476,N_9245,N_9226);
xor U9477 (N_9477,N_9070,N_9192);
nor U9478 (N_9478,N_9032,N_9086);
nor U9479 (N_9479,N_9050,N_9035);
or U9480 (N_9480,N_9169,N_9030);
or U9481 (N_9481,N_9215,N_9100);
nor U9482 (N_9482,N_9189,N_9216);
or U9483 (N_9483,N_9243,N_9063);
xor U9484 (N_9484,N_9246,N_9096);
nor U9485 (N_9485,N_9009,N_9207);
xor U9486 (N_9486,N_9058,N_9133);
and U9487 (N_9487,N_9094,N_9075);
nor U9488 (N_9488,N_9008,N_9196);
xnor U9489 (N_9489,N_9130,N_9054);
xnor U9490 (N_9490,N_9105,N_9171);
or U9491 (N_9491,N_9180,N_9043);
xnor U9492 (N_9492,N_9070,N_9038);
nor U9493 (N_9493,N_9121,N_9093);
nor U9494 (N_9494,N_9025,N_9131);
or U9495 (N_9495,N_9238,N_9094);
nand U9496 (N_9496,N_9215,N_9027);
nor U9497 (N_9497,N_9187,N_9167);
and U9498 (N_9498,N_9170,N_9004);
and U9499 (N_9499,N_9142,N_9018);
xnor U9500 (N_9500,N_9333,N_9369);
or U9501 (N_9501,N_9496,N_9472);
nand U9502 (N_9502,N_9430,N_9274);
nor U9503 (N_9503,N_9345,N_9417);
xor U9504 (N_9504,N_9438,N_9282);
and U9505 (N_9505,N_9475,N_9416);
and U9506 (N_9506,N_9289,N_9306);
or U9507 (N_9507,N_9436,N_9442);
and U9508 (N_9508,N_9497,N_9311);
nor U9509 (N_9509,N_9488,N_9255);
xor U9510 (N_9510,N_9317,N_9343);
xor U9511 (N_9511,N_9457,N_9395);
xnor U9512 (N_9512,N_9304,N_9371);
xnor U9513 (N_9513,N_9370,N_9490);
nand U9514 (N_9514,N_9277,N_9264);
nand U9515 (N_9515,N_9331,N_9290);
or U9516 (N_9516,N_9480,N_9366);
or U9517 (N_9517,N_9466,N_9335);
nand U9518 (N_9518,N_9251,N_9435);
or U9519 (N_9519,N_9283,N_9387);
xnor U9520 (N_9520,N_9263,N_9315);
nor U9521 (N_9521,N_9257,N_9271);
or U9522 (N_9522,N_9347,N_9461);
nand U9523 (N_9523,N_9307,N_9272);
nor U9524 (N_9524,N_9405,N_9467);
xnor U9525 (N_9525,N_9250,N_9465);
and U9526 (N_9526,N_9486,N_9326);
xor U9527 (N_9527,N_9252,N_9273);
xor U9528 (N_9528,N_9339,N_9278);
nand U9529 (N_9529,N_9493,N_9396);
xnor U9530 (N_9530,N_9449,N_9403);
nor U9531 (N_9531,N_9288,N_9427);
nor U9532 (N_9532,N_9437,N_9477);
xor U9533 (N_9533,N_9494,N_9286);
xnor U9534 (N_9534,N_9441,N_9412);
nand U9535 (N_9535,N_9492,N_9364);
or U9536 (N_9536,N_9470,N_9330);
nand U9537 (N_9537,N_9433,N_9385);
nor U9538 (N_9538,N_9294,N_9381);
or U9539 (N_9539,N_9275,N_9499);
nand U9540 (N_9540,N_9266,N_9359);
nor U9541 (N_9541,N_9404,N_9293);
and U9542 (N_9542,N_9388,N_9365);
or U9543 (N_9543,N_9352,N_9408);
nand U9544 (N_9544,N_9316,N_9353);
xor U9545 (N_9545,N_9386,N_9355);
nand U9546 (N_9546,N_9270,N_9262);
nor U9547 (N_9547,N_9422,N_9479);
xor U9548 (N_9548,N_9414,N_9302);
or U9549 (N_9549,N_9305,N_9367);
or U9550 (N_9550,N_9340,N_9253);
nand U9551 (N_9551,N_9406,N_9428);
xor U9552 (N_9552,N_9469,N_9318);
xnor U9553 (N_9553,N_9308,N_9350);
or U9554 (N_9554,N_9314,N_9322);
nand U9555 (N_9555,N_9292,N_9482);
nor U9556 (N_9556,N_9346,N_9476);
and U9557 (N_9557,N_9267,N_9354);
xor U9558 (N_9558,N_9324,N_9368);
nor U9559 (N_9559,N_9285,N_9407);
nand U9560 (N_9560,N_9393,N_9382);
nand U9561 (N_9561,N_9374,N_9454);
and U9562 (N_9562,N_9372,N_9474);
and U9563 (N_9563,N_9348,N_9390);
and U9564 (N_9564,N_9483,N_9261);
or U9565 (N_9565,N_9327,N_9418);
nor U9566 (N_9566,N_9341,N_9310);
or U9567 (N_9567,N_9455,N_9399);
and U9568 (N_9568,N_9415,N_9409);
or U9569 (N_9569,N_9284,N_9384);
xnor U9570 (N_9570,N_9485,N_9377);
or U9571 (N_9571,N_9321,N_9498);
nor U9572 (N_9572,N_9325,N_9258);
xnor U9573 (N_9573,N_9487,N_9298);
nand U9574 (N_9574,N_9334,N_9401);
nor U9575 (N_9575,N_9313,N_9453);
xnor U9576 (N_9576,N_9478,N_9363);
nand U9577 (N_9577,N_9419,N_9397);
or U9578 (N_9578,N_9376,N_9423);
or U9579 (N_9579,N_9276,N_9447);
xor U9580 (N_9580,N_9464,N_9450);
nor U9581 (N_9581,N_9260,N_9459);
nand U9582 (N_9582,N_9495,N_9434);
or U9583 (N_9583,N_9379,N_9440);
and U9584 (N_9584,N_9380,N_9329);
nor U9585 (N_9585,N_9473,N_9320);
xnor U9586 (N_9586,N_9463,N_9254);
nand U9587 (N_9587,N_9481,N_9458);
or U9588 (N_9588,N_9421,N_9394);
xor U9589 (N_9589,N_9429,N_9426);
and U9590 (N_9590,N_9373,N_9360);
and U9591 (N_9591,N_9448,N_9425);
and U9592 (N_9592,N_9391,N_9484);
or U9593 (N_9593,N_9309,N_9351);
and U9594 (N_9594,N_9256,N_9375);
and U9595 (N_9595,N_9462,N_9468);
nand U9596 (N_9596,N_9491,N_9489);
xnor U9597 (N_9597,N_9319,N_9456);
and U9598 (N_9598,N_9356,N_9268);
and U9599 (N_9599,N_9342,N_9411);
and U9600 (N_9600,N_9420,N_9280);
xor U9601 (N_9601,N_9398,N_9432);
or U9602 (N_9602,N_9392,N_9410);
and U9603 (N_9603,N_9362,N_9349);
and U9604 (N_9604,N_9265,N_9439);
or U9605 (N_9605,N_9338,N_9424);
xnor U9606 (N_9606,N_9336,N_9378);
nor U9607 (N_9607,N_9299,N_9296);
nand U9608 (N_9608,N_9287,N_9443);
xor U9609 (N_9609,N_9361,N_9295);
nor U9610 (N_9610,N_9328,N_9281);
xnor U9611 (N_9611,N_9344,N_9446);
nand U9612 (N_9612,N_9358,N_9300);
or U9613 (N_9613,N_9279,N_9337);
xor U9614 (N_9614,N_9323,N_9445);
nor U9615 (N_9615,N_9297,N_9301);
and U9616 (N_9616,N_9269,N_9402);
nand U9617 (N_9617,N_9303,N_9413);
or U9618 (N_9618,N_9431,N_9452);
and U9619 (N_9619,N_9460,N_9444);
xor U9620 (N_9620,N_9332,N_9400);
or U9621 (N_9621,N_9312,N_9357);
nand U9622 (N_9622,N_9471,N_9383);
nand U9623 (N_9623,N_9451,N_9291);
or U9624 (N_9624,N_9389,N_9259);
or U9625 (N_9625,N_9361,N_9411);
xor U9626 (N_9626,N_9298,N_9371);
nand U9627 (N_9627,N_9312,N_9330);
xnor U9628 (N_9628,N_9432,N_9350);
nor U9629 (N_9629,N_9479,N_9358);
nor U9630 (N_9630,N_9386,N_9358);
or U9631 (N_9631,N_9321,N_9297);
or U9632 (N_9632,N_9405,N_9478);
or U9633 (N_9633,N_9403,N_9480);
or U9634 (N_9634,N_9460,N_9455);
or U9635 (N_9635,N_9477,N_9356);
or U9636 (N_9636,N_9345,N_9430);
or U9637 (N_9637,N_9445,N_9266);
nand U9638 (N_9638,N_9432,N_9374);
nor U9639 (N_9639,N_9401,N_9367);
and U9640 (N_9640,N_9459,N_9386);
or U9641 (N_9641,N_9255,N_9348);
xnor U9642 (N_9642,N_9316,N_9394);
xor U9643 (N_9643,N_9270,N_9408);
and U9644 (N_9644,N_9410,N_9288);
or U9645 (N_9645,N_9367,N_9276);
nor U9646 (N_9646,N_9448,N_9342);
nand U9647 (N_9647,N_9325,N_9266);
xor U9648 (N_9648,N_9259,N_9476);
nor U9649 (N_9649,N_9338,N_9468);
nand U9650 (N_9650,N_9332,N_9308);
nand U9651 (N_9651,N_9367,N_9479);
nor U9652 (N_9652,N_9473,N_9478);
xor U9653 (N_9653,N_9364,N_9313);
xor U9654 (N_9654,N_9374,N_9300);
xor U9655 (N_9655,N_9479,N_9366);
nor U9656 (N_9656,N_9274,N_9465);
and U9657 (N_9657,N_9494,N_9458);
nor U9658 (N_9658,N_9304,N_9494);
nor U9659 (N_9659,N_9462,N_9471);
or U9660 (N_9660,N_9341,N_9405);
or U9661 (N_9661,N_9496,N_9430);
xor U9662 (N_9662,N_9320,N_9345);
or U9663 (N_9663,N_9377,N_9314);
nand U9664 (N_9664,N_9432,N_9456);
and U9665 (N_9665,N_9338,N_9488);
nand U9666 (N_9666,N_9449,N_9364);
nand U9667 (N_9667,N_9383,N_9337);
nand U9668 (N_9668,N_9353,N_9485);
or U9669 (N_9669,N_9341,N_9408);
or U9670 (N_9670,N_9269,N_9480);
and U9671 (N_9671,N_9443,N_9395);
and U9672 (N_9672,N_9319,N_9439);
xor U9673 (N_9673,N_9319,N_9299);
nor U9674 (N_9674,N_9458,N_9409);
and U9675 (N_9675,N_9281,N_9458);
and U9676 (N_9676,N_9380,N_9492);
or U9677 (N_9677,N_9389,N_9289);
nand U9678 (N_9678,N_9267,N_9381);
or U9679 (N_9679,N_9437,N_9445);
nor U9680 (N_9680,N_9477,N_9484);
nand U9681 (N_9681,N_9447,N_9274);
nor U9682 (N_9682,N_9424,N_9335);
xnor U9683 (N_9683,N_9282,N_9325);
or U9684 (N_9684,N_9499,N_9393);
and U9685 (N_9685,N_9417,N_9307);
xnor U9686 (N_9686,N_9384,N_9323);
xnor U9687 (N_9687,N_9469,N_9341);
xnor U9688 (N_9688,N_9408,N_9373);
or U9689 (N_9689,N_9398,N_9464);
nand U9690 (N_9690,N_9325,N_9382);
or U9691 (N_9691,N_9291,N_9490);
nand U9692 (N_9692,N_9476,N_9396);
and U9693 (N_9693,N_9260,N_9352);
and U9694 (N_9694,N_9313,N_9426);
or U9695 (N_9695,N_9339,N_9471);
xnor U9696 (N_9696,N_9258,N_9454);
nor U9697 (N_9697,N_9318,N_9358);
or U9698 (N_9698,N_9434,N_9299);
nand U9699 (N_9699,N_9475,N_9269);
nor U9700 (N_9700,N_9396,N_9333);
xnor U9701 (N_9701,N_9418,N_9448);
and U9702 (N_9702,N_9369,N_9471);
or U9703 (N_9703,N_9312,N_9402);
or U9704 (N_9704,N_9329,N_9253);
and U9705 (N_9705,N_9489,N_9314);
nor U9706 (N_9706,N_9368,N_9337);
xnor U9707 (N_9707,N_9497,N_9424);
and U9708 (N_9708,N_9281,N_9393);
nor U9709 (N_9709,N_9395,N_9308);
nand U9710 (N_9710,N_9494,N_9454);
xnor U9711 (N_9711,N_9272,N_9277);
nand U9712 (N_9712,N_9479,N_9480);
nand U9713 (N_9713,N_9391,N_9430);
and U9714 (N_9714,N_9392,N_9367);
xnor U9715 (N_9715,N_9306,N_9477);
xor U9716 (N_9716,N_9489,N_9315);
and U9717 (N_9717,N_9399,N_9365);
or U9718 (N_9718,N_9261,N_9280);
and U9719 (N_9719,N_9446,N_9416);
or U9720 (N_9720,N_9355,N_9298);
nor U9721 (N_9721,N_9498,N_9269);
or U9722 (N_9722,N_9392,N_9428);
and U9723 (N_9723,N_9357,N_9439);
xnor U9724 (N_9724,N_9344,N_9364);
and U9725 (N_9725,N_9374,N_9275);
xor U9726 (N_9726,N_9408,N_9422);
xnor U9727 (N_9727,N_9270,N_9384);
and U9728 (N_9728,N_9391,N_9342);
and U9729 (N_9729,N_9378,N_9430);
nand U9730 (N_9730,N_9296,N_9341);
nor U9731 (N_9731,N_9452,N_9284);
or U9732 (N_9732,N_9324,N_9466);
or U9733 (N_9733,N_9262,N_9393);
nand U9734 (N_9734,N_9306,N_9452);
xnor U9735 (N_9735,N_9411,N_9372);
nor U9736 (N_9736,N_9357,N_9455);
or U9737 (N_9737,N_9270,N_9481);
xnor U9738 (N_9738,N_9357,N_9255);
xnor U9739 (N_9739,N_9359,N_9317);
xor U9740 (N_9740,N_9278,N_9367);
and U9741 (N_9741,N_9264,N_9430);
or U9742 (N_9742,N_9468,N_9472);
nand U9743 (N_9743,N_9433,N_9494);
nand U9744 (N_9744,N_9435,N_9311);
xor U9745 (N_9745,N_9453,N_9391);
nor U9746 (N_9746,N_9442,N_9372);
xnor U9747 (N_9747,N_9360,N_9492);
xnor U9748 (N_9748,N_9402,N_9375);
xnor U9749 (N_9749,N_9317,N_9442);
nor U9750 (N_9750,N_9701,N_9506);
nand U9751 (N_9751,N_9708,N_9738);
xor U9752 (N_9752,N_9561,N_9525);
and U9753 (N_9753,N_9746,N_9658);
or U9754 (N_9754,N_9505,N_9538);
nand U9755 (N_9755,N_9733,N_9619);
nand U9756 (N_9756,N_9672,N_9673);
and U9757 (N_9757,N_9583,N_9715);
or U9758 (N_9758,N_9594,N_9516);
nand U9759 (N_9759,N_9500,N_9634);
nand U9760 (N_9760,N_9636,N_9573);
nor U9761 (N_9761,N_9557,N_9651);
and U9762 (N_9762,N_9680,N_9534);
and U9763 (N_9763,N_9693,N_9676);
or U9764 (N_9764,N_9705,N_9580);
nand U9765 (N_9765,N_9621,N_9514);
and U9766 (N_9766,N_9623,N_9718);
and U9767 (N_9767,N_9508,N_9523);
xnor U9768 (N_9768,N_9569,N_9574);
xor U9769 (N_9769,N_9663,N_9618);
xnor U9770 (N_9770,N_9625,N_9710);
and U9771 (N_9771,N_9552,N_9731);
nor U9772 (N_9772,N_9616,N_9595);
or U9773 (N_9773,N_9597,N_9732);
and U9774 (N_9774,N_9681,N_9567);
nor U9775 (N_9775,N_9596,N_9665);
and U9776 (N_9776,N_9504,N_9632);
and U9777 (N_9777,N_9515,N_9620);
or U9778 (N_9778,N_9503,N_9686);
xnor U9779 (N_9779,N_9531,N_9622);
nor U9780 (N_9780,N_9586,N_9641);
nor U9781 (N_9781,N_9502,N_9691);
xor U9782 (N_9782,N_9645,N_9602);
and U9783 (N_9783,N_9566,N_9570);
xnor U9784 (N_9784,N_9749,N_9736);
and U9785 (N_9785,N_9614,N_9649);
or U9786 (N_9786,N_9543,N_9565);
xor U9787 (N_9787,N_9741,N_9551);
or U9788 (N_9788,N_9707,N_9541);
nand U9789 (N_9789,N_9593,N_9698);
and U9790 (N_9790,N_9631,N_9706);
or U9791 (N_9791,N_9716,N_9745);
nand U9792 (N_9792,N_9743,N_9739);
xnor U9793 (N_9793,N_9646,N_9656);
or U9794 (N_9794,N_9519,N_9696);
nand U9795 (N_9795,N_9692,N_9657);
nand U9796 (N_9796,N_9722,N_9627);
and U9797 (N_9797,N_9662,N_9650);
nor U9798 (N_9798,N_9725,N_9638);
and U9799 (N_9799,N_9695,N_9664);
nor U9800 (N_9800,N_9737,N_9590);
and U9801 (N_9801,N_9548,N_9603);
or U9802 (N_9802,N_9704,N_9575);
nand U9803 (N_9803,N_9713,N_9568);
and U9804 (N_9804,N_9585,N_9501);
nor U9805 (N_9805,N_9529,N_9702);
or U9806 (N_9806,N_9635,N_9724);
or U9807 (N_9807,N_9532,N_9744);
xnor U9808 (N_9808,N_9678,N_9610);
and U9809 (N_9809,N_9588,N_9688);
nand U9810 (N_9810,N_9675,N_9699);
or U9811 (N_9811,N_9535,N_9671);
nor U9812 (N_9812,N_9611,N_9640);
xnor U9813 (N_9813,N_9729,N_9723);
or U9814 (N_9814,N_9526,N_9512);
or U9815 (N_9815,N_9629,N_9666);
nand U9816 (N_9816,N_9612,N_9518);
xnor U9817 (N_9817,N_9742,N_9556);
xnor U9818 (N_9818,N_9579,N_9539);
xnor U9819 (N_9819,N_9684,N_9558);
or U9820 (N_9820,N_9604,N_9727);
nor U9821 (N_9821,N_9669,N_9547);
and U9822 (N_9822,N_9637,N_9717);
xnor U9823 (N_9823,N_9639,N_9578);
xnor U9824 (N_9824,N_9674,N_9513);
or U9825 (N_9825,N_9572,N_9660);
nor U9826 (N_9826,N_9679,N_9559);
and U9827 (N_9827,N_9682,N_9542);
xnor U9828 (N_9828,N_9517,N_9687);
nand U9829 (N_9829,N_9677,N_9533);
nand U9830 (N_9830,N_9606,N_9601);
xnor U9831 (N_9831,N_9562,N_9700);
nor U9832 (N_9832,N_9554,N_9626);
nand U9833 (N_9833,N_9726,N_9714);
and U9834 (N_9834,N_9652,N_9633);
nand U9835 (N_9835,N_9553,N_9510);
and U9836 (N_9836,N_9520,N_9546);
nor U9837 (N_9837,N_9599,N_9536);
xnor U9838 (N_9838,N_9628,N_9624);
xor U9839 (N_9839,N_9537,N_9697);
nand U9840 (N_9840,N_9540,N_9643);
nor U9841 (N_9841,N_9592,N_9609);
or U9842 (N_9842,N_9549,N_9581);
nor U9843 (N_9843,N_9582,N_9740);
or U9844 (N_9844,N_9527,N_9689);
or U9845 (N_9845,N_9587,N_9670);
xnor U9846 (N_9846,N_9734,N_9591);
nor U9847 (N_9847,N_9735,N_9617);
nor U9848 (N_9848,N_9608,N_9644);
xnor U9849 (N_9849,N_9703,N_9668);
and U9850 (N_9850,N_9550,N_9522);
or U9851 (N_9851,N_9654,N_9659);
or U9852 (N_9852,N_9564,N_9748);
nor U9853 (N_9853,N_9521,N_9613);
nand U9854 (N_9854,N_9642,N_9560);
or U9855 (N_9855,N_9607,N_9728);
nand U9856 (N_9856,N_9528,N_9530);
nor U9857 (N_9857,N_9709,N_9667);
nor U9858 (N_9858,N_9690,N_9511);
and U9859 (N_9859,N_9584,N_9747);
nor U9860 (N_9860,N_9605,N_9563);
xor U9861 (N_9861,N_9655,N_9555);
nor U9862 (N_9862,N_9600,N_9694);
nand U9863 (N_9863,N_9589,N_9524);
nand U9864 (N_9864,N_9648,N_9577);
or U9865 (N_9865,N_9661,N_9544);
nor U9866 (N_9866,N_9545,N_9576);
xnor U9867 (N_9867,N_9711,N_9683);
and U9868 (N_9868,N_9653,N_9730);
xnor U9869 (N_9869,N_9712,N_9647);
nor U9870 (N_9870,N_9721,N_9507);
xnor U9871 (N_9871,N_9685,N_9719);
or U9872 (N_9872,N_9615,N_9720);
and U9873 (N_9873,N_9571,N_9630);
or U9874 (N_9874,N_9509,N_9598);
and U9875 (N_9875,N_9604,N_9523);
and U9876 (N_9876,N_9530,N_9720);
nor U9877 (N_9877,N_9703,N_9727);
or U9878 (N_9878,N_9528,N_9502);
nor U9879 (N_9879,N_9605,N_9722);
or U9880 (N_9880,N_9631,N_9669);
xnor U9881 (N_9881,N_9612,N_9556);
xnor U9882 (N_9882,N_9701,N_9605);
and U9883 (N_9883,N_9665,N_9509);
xnor U9884 (N_9884,N_9737,N_9641);
and U9885 (N_9885,N_9563,N_9649);
nor U9886 (N_9886,N_9622,N_9631);
or U9887 (N_9887,N_9697,N_9648);
nor U9888 (N_9888,N_9712,N_9512);
xor U9889 (N_9889,N_9689,N_9726);
nor U9890 (N_9890,N_9584,N_9666);
and U9891 (N_9891,N_9574,N_9669);
xor U9892 (N_9892,N_9677,N_9538);
or U9893 (N_9893,N_9584,N_9677);
nor U9894 (N_9894,N_9661,N_9675);
nand U9895 (N_9895,N_9632,N_9550);
and U9896 (N_9896,N_9689,N_9568);
nand U9897 (N_9897,N_9652,N_9602);
and U9898 (N_9898,N_9658,N_9514);
nand U9899 (N_9899,N_9533,N_9547);
and U9900 (N_9900,N_9723,N_9627);
and U9901 (N_9901,N_9686,N_9704);
nand U9902 (N_9902,N_9558,N_9698);
and U9903 (N_9903,N_9620,N_9744);
and U9904 (N_9904,N_9573,N_9587);
nand U9905 (N_9905,N_9607,N_9637);
xnor U9906 (N_9906,N_9604,N_9684);
and U9907 (N_9907,N_9676,N_9710);
and U9908 (N_9908,N_9718,N_9682);
and U9909 (N_9909,N_9517,N_9600);
and U9910 (N_9910,N_9526,N_9527);
nor U9911 (N_9911,N_9695,N_9645);
xnor U9912 (N_9912,N_9517,N_9737);
or U9913 (N_9913,N_9564,N_9532);
or U9914 (N_9914,N_9590,N_9633);
nand U9915 (N_9915,N_9603,N_9739);
nor U9916 (N_9916,N_9634,N_9744);
nor U9917 (N_9917,N_9640,N_9691);
nand U9918 (N_9918,N_9537,N_9748);
nand U9919 (N_9919,N_9671,N_9662);
nand U9920 (N_9920,N_9714,N_9584);
nand U9921 (N_9921,N_9674,N_9592);
nor U9922 (N_9922,N_9745,N_9676);
or U9923 (N_9923,N_9723,N_9547);
or U9924 (N_9924,N_9707,N_9504);
nand U9925 (N_9925,N_9661,N_9628);
xor U9926 (N_9926,N_9573,N_9565);
xor U9927 (N_9927,N_9577,N_9673);
xnor U9928 (N_9928,N_9717,N_9574);
and U9929 (N_9929,N_9681,N_9602);
and U9930 (N_9930,N_9555,N_9597);
and U9931 (N_9931,N_9593,N_9581);
xor U9932 (N_9932,N_9622,N_9502);
and U9933 (N_9933,N_9708,N_9555);
nor U9934 (N_9934,N_9595,N_9731);
xor U9935 (N_9935,N_9579,N_9600);
xor U9936 (N_9936,N_9609,N_9703);
or U9937 (N_9937,N_9599,N_9523);
nand U9938 (N_9938,N_9523,N_9665);
or U9939 (N_9939,N_9684,N_9630);
nor U9940 (N_9940,N_9744,N_9736);
xnor U9941 (N_9941,N_9583,N_9559);
nand U9942 (N_9942,N_9652,N_9727);
or U9943 (N_9943,N_9513,N_9694);
nand U9944 (N_9944,N_9685,N_9549);
nor U9945 (N_9945,N_9725,N_9646);
and U9946 (N_9946,N_9502,N_9640);
and U9947 (N_9947,N_9731,N_9541);
nand U9948 (N_9948,N_9662,N_9529);
nor U9949 (N_9949,N_9722,N_9684);
and U9950 (N_9950,N_9551,N_9707);
xor U9951 (N_9951,N_9521,N_9744);
xor U9952 (N_9952,N_9681,N_9698);
and U9953 (N_9953,N_9579,N_9542);
and U9954 (N_9954,N_9702,N_9675);
nor U9955 (N_9955,N_9590,N_9718);
or U9956 (N_9956,N_9725,N_9624);
xor U9957 (N_9957,N_9668,N_9690);
or U9958 (N_9958,N_9704,N_9630);
nor U9959 (N_9959,N_9548,N_9715);
xnor U9960 (N_9960,N_9548,N_9674);
or U9961 (N_9961,N_9713,N_9666);
and U9962 (N_9962,N_9706,N_9621);
or U9963 (N_9963,N_9554,N_9645);
xnor U9964 (N_9964,N_9557,N_9749);
nor U9965 (N_9965,N_9581,N_9543);
or U9966 (N_9966,N_9665,N_9525);
nor U9967 (N_9967,N_9614,N_9695);
nand U9968 (N_9968,N_9609,N_9633);
xor U9969 (N_9969,N_9648,N_9641);
nand U9970 (N_9970,N_9548,N_9528);
nand U9971 (N_9971,N_9653,N_9713);
nand U9972 (N_9972,N_9587,N_9660);
nor U9973 (N_9973,N_9728,N_9644);
nand U9974 (N_9974,N_9661,N_9662);
or U9975 (N_9975,N_9701,N_9527);
xnor U9976 (N_9976,N_9653,N_9654);
or U9977 (N_9977,N_9643,N_9699);
or U9978 (N_9978,N_9706,N_9683);
xnor U9979 (N_9979,N_9670,N_9599);
xnor U9980 (N_9980,N_9548,N_9605);
or U9981 (N_9981,N_9556,N_9741);
xnor U9982 (N_9982,N_9602,N_9664);
nor U9983 (N_9983,N_9657,N_9691);
nor U9984 (N_9984,N_9501,N_9742);
and U9985 (N_9985,N_9632,N_9531);
nand U9986 (N_9986,N_9644,N_9629);
or U9987 (N_9987,N_9524,N_9656);
and U9988 (N_9988,N_9549,N_9564);
or U9989 (N_9989,N_9732,N_9711);
and U9990 (N_9990,N_9728,N_9724);
and U9991 (N_9991,N_9573,N_9550);
or U9992 (N_9992,N_9563,N_9638);
nand U9993 (N_9993,N_9670,N_9543);
nand U9994 (N_9994,N_9700,N_9645);
and U9995 (N_9995,N_9724,N_9647);
nand U9996 (N_9996,N_9641,N_9519);
nand U9997 (N_9997,N_9515,N_9731);
or U9998 (N_9998,N_9504,N_9735);
nor U9999 (N_9999,N_9535,N_9519);
nor U10000 (N_10000,N_9852,N_9936);
and U10001 (N_10001,N_9784,N_9762);
and U10002 (N_10002,N_9870,N_9783);
and U10003 (N_10003,N_9901,N_9974);
xnor U10004 (N_10004,N_9794,N_9860);
xnor U10005 (N_10005,N_9853,N_9805);
and U10006 (N_10006,N_9777,N_9915);
and U10007 (N_10007,N_9996,N_9835);
nor U10008 (N_10008,N_9815,N_9782);
nand U10009 (N_10009,N_9800,N_9897);
nor U10010 (N_10010,N_9920,N_9957);
nand U10011 (N_10011,N_9766,N_9804);
xnor U10012 (N_10012,N_9846,N_9908);
nor U10013 (N_10013,N_9814,N_9898);
or U10014 (N_10014,N_9992,N_9856);
nor U10015 (N_10015,N_9861,N_9880);
xnor U10016 (N_10016,N_9820,N_9891);
and U10017 (N_10017,N_9775,N_9997);
or U10018 (N_10018,N_9801,N_9885);
and U10019 (N_10019,N_9904,N_9943);
and U10020 (N_10020,N_9931,N_9771);
or U10021 (N_10021,N_9914,N_9985);
xor U10022 (N_10022,N_9892,N_9813);
nor U10023 (N_10023,N_9995,N_9905);
xor U10024 (N_10024,N_9790,N_9811);
and U10025 (N_10025,N_9940,N_9906);
and U10026 (N_10026,N_9823,N_9899);
nand U10027 (N_10027,N_9817,N_9765);
nand U10028 (N_10028,N_9888,N_9971);
and U10029 (N_10029,N_9850,N_9955);
xor U10030 (N_10030,N_9930,N_9787);
and U10031 (N_10031,N_9977,N_9865);
and U10032 (N_10032,N_9867,N_9827);
xnor U10033 (N_10033,N_9954,N_9958);
nor U10034 (N_10034,N_9761,N_9960);
nand U10035 (N_10035,N_9951,N_9791);
nor U10036 (N_10036,N_9941,N_9886);
and U10037 (N_10037,N_9963,N_9840);
nor U10038 (N_10038,N_9768,N_9975);
or U10039 (N_10039,N_9987,N_9798);
nor U10040 (N_10040,N_9767,N_9900);
xnor U10041 (N_10041,N_9789,N_9844);
nand U10042 (N_10042,N_9998,N_9809);
and U10043 (N_10043,N_9925,N_9903);
xnor U10044 (N_10044,N_9887,N_9845);
or U10045 (N_10045,N_9822,N_9764);
nor U10046 (N_10046,N_9829,N_9956);
xnor U10047 (N_10047,N_9882,N_9758);
and U10048 (N_10048,N_9834,N_9988);
and U10049 (N_10049,N_9857,N_9873);
and U10050 (N_10050,N_9889,N_9788);
and U10051 (N_10051,N_9763,N_9894);
nand U10052 (N_10052,N_9911,N_9973);
nand U10053 (N_10053,N_9893,N_9948);
and U10054 (N_10054,N_9979,N_9944);
xor U10055 (N_10055,N_9816,N_9916);
or U10056 (N_10056,N_9797,N_9831);
nor U10057 (N_10057,N_9842,N_9890);
or U10058 (N_10058,N_9803,N_9753);
xnor U10059 (N_10059,N_9863,N_9778);
and U10060 (N_10060,N_9808,N_9802);
or U10061 (N_10061,N_9983,N_9825);
or U10062 (N_10062,N_9769,N_9984);
nand U10063 (N_10063,N_9933,N_9843);
xor U10064 (N_10064,N_9770,N_9858);
nand U10065 (N_10065,N_9991,N_9877);
xnor U10066 (N_10066,N_9895,N_9913);
or U10067 (N_10067,N_9839,N_9851);
and U10068 (N_10068,N_9939,N_9907);
and U10069 (N_10069,N_9918,N_9981);
nand U10070 (N_10070,N_9875,N_9962);
nor U10071 (N_10071,N_9772,N_9795);
or U10072 (N_10072,N_9757,N_9912);
or U10073 (N_10073,N_9952,N_9796);
nand U10074 (N_10074,N_9819,N_9755);
nor U10075 (N_10075,N_9935,N_9866);
and U10076 (N_10076,N_9751,N_9937);
nand U10077 (N_10077,N_9953,N_9883);
nor U10078 (N_10078,N_9786,N_9970);
nor U10079 (N_10079,N_9967,N_9964);
and U10080 (N_10080,N_9750,N_9989);
and U10081 (N_10081,N_9869,N_9993);
or U10082 (N_10082,N_9760,N_9965);
nand U10083 (N_10083,N_9968,N_9879);
nand U10084 (N_10084,N_9836,N_9793);
nand U10085 (N_10085,N_9854,N_9756);
and U10086 (N_10086,N_9752,N_9878);
and U10087 (N_10087,N_9929,N_9799);
and U10088 (N_10088,N_9862,N_9947);
and U10089 (N_10089,N_9961,N_9773);
and U10090 (N_10090,N_9976,N_9932);
xor U10091 (N_10091,N_9759,N_9859);
and U10092 (N_10092,N_9806,N_9833);
xor U10093 (N_10093,N_9874,N_9927);
or U10094 (N_10094,N_9871,N_9780);
and U10095 (N_10095,N_9838,N_9824);
nand U10096 (N_10096,N_9959,N_9966);
nand U10097 (N_10097,N_9934,N_9949);
nand U10098 (N_10098,N_9884,N_9978);
xor U10099 (N_10099,N_9849,N_9807);
and U10100 (N_10100,N_9832,N_9922);
nand U10101 (N_10101,N_9902,N_9986);
and U10102 (N_10102,N_9994,N_9792);
nor U10103 (N_10103,N_9855,N_9818);
nor U10104 (N_10104,N_9926,N_9837);
nand U10105 (N_10105,N_9921,N_9923);
nor U10106 (N_10106,N_9950,N_9828);
or U10107 (N_10107,N_9990,N_9779);
nor U10108 (N_10108,N_9781,N_9910);
nor U10109 (N_10109,N_9909,N_9821);
nand U10110 (N_10110,N_9919,N_9928);
nand U10111 (N_10111,N_9982,N_9917);
and U10112 (N_10112,N_9810,N_9785);
xnor U10113 (N_10113,N_9938,N_9924);
nor U10114 (N_10114,N_9872,N_9864);
xor U10115 (N_10115,N_9868,N_9896);
and U10116 (N_10116,N_9942,N_9999);
or U10117 (N_10117,N_9881,N_9972);
nand U10118 (N_10118,N_9776,N_9830);
xnor U10119 (N_10119,N_9980,N_9945);
and U10120 (N_10120,N_9848,N_9826);
nor U10121 (N_10121,N_9847,N_9774);
or U10122 (N_10122,N_9946,N_9969);
xnor U10123 (N_10123,N_9876,N_9841);
xnor U10124 (N_10124,N_9754,N_9812);
and U10125 (N_10125,N_9945,N_9818);
and U10126 (N_10126,N_9750,N_9847);
xnor U10127 (N_10127,N_9961,N_9988);
nand U10128 (N_10128,N_9804,N_9910);
nand U10129 (N_10129,N_9931,N_9895);
or U10130 (N_10130,N_9793,N_9825);
and U10131 (N_10131,N_9793,N_9935);
and U10132 (N_10132,N_9817,N_9908);
and U10133 (N_10133,N_9799,N_9920);
or U10134 (N_10134,N_9948,N_9986);
xor U10135 (N_10135,N_9956,N_9881);
nor U10136 (N_10136,N_9803,N_9893);
nand U10137 (N_10137,N_9877,N_9983);
nor U10138 (N_10138,N_9819,N_9896);
and U10139 (N_10139,N_9975,N_9888);
nor U10140 (N_10140,N_9773,N_9929);
nand U10141 (N_10141,N_9923,N_9869);
nor U10142 (N_10142,N_9858,N_9867);
nand U10143 (N_10143,N_9808,N_9795);
or U10144 (N_10144,N_9768,N_9929);
xor U10145 (N_10145,N_9970,N_9850);
nand U10146 (N_10146,N_9875,N_9840);
or U10147 (N_10147,N_9819,N_9860);
xor U10148 (N_10148,N_9867,N_9869);
and U10149 (N_10149,N_9965,N_9845);
and U10150 (N_10150,N_9903,N_9860);
or U10151 (N_10151,N_9932,N_9846);
nand U10152 (N_10152,N_9902,N_9925);
nor U10153 (N_10153,N_9953,N_9980);
nor U10154 (N_10154,N_9808,N_9995);
xnor U10155 (N_10155,N_9979,N_9880);
and U10156 (N_10156,N_9839,N_9751);
nand U10157 (N_10157,N_9817,N_9968);
or U10158 (N_10158,N_9777,N_9993);
and U10159 (N_10159,N_9808,N_9914);
or U10160 (N_10160,N_9895,N_9769);
xnor U10161 (N_10161,N_9802,N_9992);
xor U10162 (N_10162,N_9930,N_9925);
or U10163 (N_10163,N_9846,N_9775);
xor U10164 (N_10164,N_9929,N_9904);
or U10165 (N_10165,N_9994,N_9975);
nor U10166 (N_10166,N_9995,N_9997);
nand U10167 (N_10167,N_9887,N_9781);
nor U10168 (N_10168,N_9931,N_9965);
nor U10169 (N_10169,N_9914,N_9870);
nand U10170 (N_10170,N_9965,N_9982);
or U10171 (N_10171,N_9826,N_9921);
and U10172 (N_10172,N_9761,N_9964);
nand U10173 (N_10173,N_9753,N_9785);
nand U10174 (N_10174,N_9927,N_9843);
nor U10175 (N_10175,N_9831,N_9883);
or U10176 (N_10176,N_9868,N_9875);
or U10177 (N_10177,N_9838,N_9949);
nand U10178 (N_10178,N_9819,N_9785);
nand U10179 (N_10179,N_9921,N_9867);
and U10180 (N_10180,N_9833,N_9891);
or U10181 (N_10181,N_9811,N_9921);
nand U10182 (N_10182,N_9921,N_9956);
nor U10183 (N_10183,N_9783,N_9972);
xnor U10184 (N_10184,N_9982,N_9756);
and U10185 (N_10185,N_9860,N_9911);
nand U10186 (N_10186,N_9830,N_9975);
nand U10187 (N_10187,N_9901,N_9792);
nand U10188 (N_10188,N_9866,N_9775);
or U10189 (N_10189,N_9911,N_9972);
nor U10190 (N_10190,N_9787,N_9803);
nor U10191 (N_10191,N_9825,N_9853);
nor U10192 (N_10192,N_9924,N_9768);
or U10193 (N_10193,N_9931,N_9982);
nor U10194 (N_10194,N_9896,N_9921);
and U10195 (N_10195,N_9848,N_9953);
or U10196 (N_10196,N_9878,N_9854);
nor U10197 (N_10197,N_9775,N_9804);
xor U10198 (N_10198,N_9962,N_9916);
xor U10199 (N_10199,N_9763,N_9910);
xnor U10200 (N_10200,N_9887,N_9806);
xor U10201 (N_10201,N_9920,N_9917);
nor U10202 (N_10202,N_9980,N_9999);
or U10203 (N_10203,N_9833,N_9768);
xnor U10204 (N_10204,N_9782,N_9938);
nand U10205 (N_10205,N_9828,N_9904);
and U10206 (N_10206,N_9985,N_9852);
and U10207 (N_10207,N_9933,N_9935);
or U10208 (N_10208,N_9834,N_9806);
xor U10209 (N_10209,N_9999,N_9760);
or U10210 (N_10210,N_9919,N_9973);
and U10211 (N_10211,N_9779,N_9941);
xnor U10212 (N_10212,N_9858,N_9997);
xnor U10213 (N_10213,N_9843,N_9856);
nand U10214 (N_10214,N_9865,N_9900);
nor U10215 (N_10215,N_9955,N_9992);
and U10216 (N_10216,N_9929,N_9888);
and U10217 (N_10217,N_9824,N_9895);
or U10218 (N_10218,N_9845,N_9826);
xor U10219 (N_10219,N_9997,N_9792);
nor U10220 (N_10220,N_9857,N_9789);
and U10221 (N_10221,N_9992,N_9932);
nand U10222 (N_10222,N_9933,N_9978);
nor U10223 (N_10223,N_9963,N_9933);
xnor U10224 (N_10224,N_9936,N_9913);
xor U10225 (N_10225,N_9972,N_9929);
and U10226 (N_10226,N_9838,N_9891);
or U10227 (N_10227,N_9905,N_9847);
or U10228 (N_10228,N_9879,N_9885);
xor U10229 (N_10229,N_9924,N_9866);
and U10230 (N_10230,N_9775,N_9772);
or U10231 (N_10231,N_9929,N_9879);
nor U10232 (N_10232,N_9793,N_9937);
nor U10233 (N_10233,N_9800,N_9942);
nand U10234 (N_10234,N_9811,N_9913);
or U10235 (N_10235,N_9917,N_9790);
xnor U10236 (N_10236,N_9869,N_9916);
nand U10237 (N_10237,N_9936,N_9903);
and U10238 (N_10238,N_9840,N_9821);
nor U10239 (N_10239,N_9895,N_9808);
xnor U10240 (N_10240,N_9830,N_9819);
and U10241 (N_10241,N_9887,N_9798);
or U10242 (N_10242,N_9982,N_9807);
and U10243 (N_10243,N_9803,N_9840);
nand U10244 (N_10244,N_9901,N_9778);
or U10245 (N_10245,N_9950,N_9857);
nor U10246 (N_10246,N_9924,N_9758);
or U10247 (N_10247,N_9903,N_9854);
nand U10248 (N_10248,N_9770,N_9906);
or U10249 (N_10249,N_9944,N_9882);
nand U10250 (N_10250,N_10154,N_10094);
xor U10251 (N_10251,N_10041,N_10222);
or U10252 (N_10252,N_10088,N_10069);
xnor U10253 (N_10253,N_10204,N_10238);
nand U10254 (N_10254,N_10208,N_10107);
xor U10255 (N_10255,N_10077,N_10162);
nor U10256 (N_10256,N_10091,N_10037);
or U10257 (N_10257,N_10000,N_10227);
nor U10258 (N_10258,N_10101,N_10123);
nand U10259 (N_10259,N_10167,N_10232);
or U10260 (N_10260,N_10008,N_10130);
nor U10261 (N_10261,N_10070,N_10236);
or U10262 (N_10262,N_10136,N_10104);
nor U10263 (N_10263,N_10151,N_10023);
and U10264 (N_10264,N_10071,N_10131);
or U10265 (N_10265,N_10206,N_10020);
and U10266 (N_10266,N_10244,N_10202);
or U10267 (N_10267,N_10047,N_10110);
and U10268 (N_10268,N_10172,N_10155);
and U10269 (N_10269,N_10097,N_10178);
or U10270 (N_10270,N_10175,N_10144);
xnor U10271 (N_10271,N_10054,N_10239);
xnor U10272 (N_10272,N_10125,N_10160);
xor U10273 (N_10273,N_10109,N_10142);
and U10274 (N_10274,N_10242,N_10192);
or U10275 (N_10275,N_10066,N_10212);
xnor U10276 (N_10276,N_10039,N_10198);
nor U10277 (N_10277,N_10114,N_10011);
xor U10278 (N_10278,N_10146,N_10128);
nand U10279 (N_10279,N_10149,N_10196);
xor U10280 (N_10280,N_10119,N_10159);
nand U10281 (N_10281,N_10213,N_10132);
nand U10282 (N_10282,N_10225,N_10118);
xnor U10283 (N_10283,N_10072,N_10189);
or U10284 (N_10284,N_10171,N_10035);
and U10285 (N_10285,N_10106,N_10089);
nand U10286 (N_10286,N_10191,N_10139);
xnor U10287 (N_10287,N_10223,N_10186);
xor U10288 (N_10288,N_10161,N_10032);
nor U10289 (N_10289,N_10027,N_10217);
or U10290 (N_10290,N_10040,N_10224);
xnor U10291 (N_10291,N_10180,N_10201);
nand U10292 (N_10292,N_10122,N_10061);
and U10293 (N_10293,N_10105,N_10113);
nor U10294 (N_10294,N_10016,N_10219);
nor U10295 (N_10295,N_10177,N_10055);
nor U10296 (N_10296,N_10193,N_10065);
nand U10297 (N_10297,N_10141,N_10190);
or U10298 (N_10298,N_10076,N_10004);
nor U10299 (N_10299,N_10140,N_10169);
nor U10300 (N_10300,N_10233,N_10220);
xnor U10301 (N_10301,N_10166,N_10188);
nor U10302 (N_10302,N_10048,N_10228);
or U10303 (N_10303,N_10246,N_10057);
nand U10304 (N_10304,N_10199,N_10126);
nand U10305 (N_10305,N_10147,N_10045);
nor U10306 (N_10306,N_10095,N_10143);
and U10307 (N_10307,N_10165,N_10093);
nand U10308 (N_10308,N_10099,N_10163);
or U10309 (N_10309,N_10006,N_10015);
nand U10310 (N_10310,N_10215,N_10184);
nand U10311 (N_10311,N_10187,N_10112);
or U10312 (N_10312,N_10083,N_10026);
or U10313 (N_10313,N_10235,N_10134);
xor U10314 (N_10314,N_10025,N_10010);
and U10315 (N_10315,N_10124,N_10121);
and U10316 (N_10316,N_10115,N_10084);
xor U10317 (N_10317,N_10053,N_10231);
xor U10318 (N_10318,N_10195,N_10229);
and U10319 (N_10319,N_10194,N_10150);
nor U10320 (N_10320,N_10174,N_10017);
nor U10321 (N_10321,N_10241,N_10062);
nor U10322 (N_10322,N_10043,N_10207);
nand U10323 (N_10323,N_10030,N_10173);
nand U10324 (N_10324,N_10156,N_10085);
nand U10325 (N_10325,N_10133,N_10100);
or U10326 (N_10326,N_10096,N_10157);
and U10327 (N_10327,N_10137,N_10024);
or U10328 (N_10328,N_10240,N_10226);
nand U10329 (N_10329,N_10018,N_10216);
and U10330 (N_10330,N_10033,N_10209);
and U10331 (N_10331,N_10152,N_10002);
and U10332 (N_10332,N_10056,N_10247);
nand U10333 (N_10333,N_10080,N_10028);
nand U10334 (N_10334,N_10073,N_10249);
and U10335 (N_10335,N_10031,N_10090);
nand U10336 (N_10336,N_10116,N_10185);
nor U10337 (N_10337,N_10098,N_10176);
or U10338 (N_10338,N_10129,N_10183);
and U10339 (N_10339,N_10086,N_10164);
or U10340 (N_10340,N_10036,N_10058);
and U10341 (N_10341,N_10197,N_10009);
and U10342 (N_10342,N_10153,N_10042);
or U10343 (N_10343,N_10203,N_10127);
or U10344 (N_10344,N_10170,N_10158);
nor U10345 (N_10345,N_10179,N_10074);
nand U10346 (N_10346,N_10051,N_10079);
or U10347 (N_10347,N_10230,N_10034);
and U10348 (N_10348,N_10012,N_10078);
nand U10349 (N_10349,N_10029,N_10092);
or U10350 (N_10350,N_10103,N_10117);
and U10351 (N_10351,N_10182,N_10214);
nor U10352 (N_10352,N_10068,N_10049);
nand U10353 (N_10353,N_10138,N_10064);
nand U10354 (N_10354,N_10081,N_10102);
nand U10355 (N_10355,N_10168,N_10237);
nand U10356 (N_10356,N_10145,N_10108);
nand U10357 (N_10357,N_10044,N_10200);
nand U10358 (N_10358,N_10003,N_10221);
or U10359 (N_10359,N_10087,N_10052);
nor U10360 (N_10360,N_10210,N_10205);
nor U10361 (N_10361,N_10014,N_10111);
nand U10362 (N_10362,N_10007,N_10038);
nand U10363 (N_10363,N_10120,N_10001);
xor U10364 (N_10364,N_10022,N_10148);
nor U10365 (N_10365,N_10021,N_10046);
nor U10366 (N_10366,N_10060,N_10218);
xor U10367 (N_10367,N_10181,N_10005);
nor U10368 (N_10368,N_10245,N_10013);
or U10369 (N_10369,N_10211,N_10243);
xor U10370 (N_10370,N_10063,N_10067);
nand U10371 (N_10371,N_10075,N_10059);
xor U10372 (N_10372,N_10019,N_10248);
and U10373 (N_10373,N_10050,N_10135);
or U10374 (N_10374,N_10234,N_10082);
or U10375 (N_10375,N_10220,N_10071);
nor U10376 (N_10376,N_10204,N_10028);
or U10377 (N_10377,N_10216,N_10066);
nor U10378 (N_10378,N_10052,N_10067);
and U10379 (N_10379,N_10177,N_10020);
and U10380 (N_10380,N_10093,N_10074);
and U10381 (N_10381,N_10237,N_10149);
or U10382 (N_10382,N_10035,N_10166);
and U10383 (N_10383,N_10050,N_10159);
xnor U10384 (N_10384,N_10235,N_10014);
nor U10385 (N_10385,N_10168,N_10217);
xnor U10386 (N_10386,N_10244,N_10148);
xor U10387 (N_10387,N_10122,N_10137);
nand U10388 (N_10388,N_10005,N_10033);
nor U10389 (N_10389,N_10229,N_10013);
xnor U10390 (N_10390,N_10059,N_10065);
or U10391 (N_10391,N_10249,N_10187);
nand U10392 (N_10392,N_10058,N_10177);
and U10393 (N_10393,N_10137,N_10041);
and U10394 (N_10394,N_10211,N_10238);
nand U10395 (N_10395,N_10016,N_10058);
nor U10396 (N_10396,N_10032,N_10180);
xor U10397 (N_10397,N_10028,N_10101);
nor U10398 (N_10398,N_10153,N_10046);
and U10399 (N_10399,N_10171,N_10145);
or U10400 (N_10400,N_10194,N_10206);
nor U10401 (N_10401,N_10147,N_10031);
nor U10402 (N_10402,N_10091,N_10085);
and U10403 (N_10403,N_10155,N_10044);
and U10404 (N_10404,N_10005,N_10135);
and U10405 (N_10405,N_10083,N_10207);
xor U10406 (N_10406,N_10070,N_10127);
and U10407 (N_10407,N_10084,N_10074);
xnor U10408 (N_10408,N_10247,N_10185);
xor U10409 (N_10409,N_10055,N_10223);
xor U10410 (N_10410,N_10004,N_10215);
nand U10411 (N_10411,N_10231,N_10111);
xnor U10412 (N_10412,N_10231,N_10132);
and U10413 (N_10413,N_10035,N_10160);
nand U10414 (N_10414,N_10189,N_10099);
xnor U10415 (N_10415,N_10205,N_10072);
nor U10416 (N_10416,N_10116,N_10086);
xor U10417 (N_10417,N_10181,N_10066);
or U10418 (N_10418,N_10228,N_10136);
nor U10419 (N_10419,N_10012,N_10047);
or U10420 (N_10420,N_10178,N_10167);
or U10421 (N_10421,N_10071,N_10059);
nand U10422 (N_10422,N_10186,N_10054);
nand U10423 (N_10423,N_10031,N_10175);
nand U10424 (N_10424,N_10206,N_10153);
xor U10425 (N_10425,N_10034,N_10025);
or U10426 (N_10426,N_10025,N_10089);
xnor U10427 (N_10427,N_10164,N_10156);
or U10428 (N_10428,N_10229,N_10031);
xnor U10429 (N_10429,N_10021,N_10060);
nand U10430 (N_10430,N_10103,N_10024);
and U10431 (N_10431,N_10193,N_10116);
xnor U10432 (N_10432,N_10033,N_10215);
or U10433 (N_10433,N_10132,N_10209);
or U10434 (N_10434,N_10148,N_10238);
and U10435 (N_10435,N_10088,N_10086);
nor U10436 (N_10436,N_10023,N_10184);
or U10437 (N_10437,N_10083,N_10087);
or U10438 (N_10438,N_10007,N_10089);
nor U10439 (N_10439,N_10186,N_10097);
and U10440 (N_10440,N_10072,N_10035);
xor U10441 (N_10441,N_10036,N_10205);
nor U10442 (N_10442,N_10219,N_10207);
or U10443 (N_10443,N_10085,N_10137);
nor U10444 (N_10444,N_10235,N_10216);
nand U10445 (N_10445,N_10136,N_10100);
or U10446 (N_10446,N_10142,N_10217);
nand U10447 (N_10447,N_10025,N_10120);
and U10448 (N_10448,N_10242,N_10141);
xor U10449 (N_10449,N_10122,N_10228);
nand U10450 (N_10450,N_10149,N_10134);
nand U10451 (N_10451,N_10050,N_10190);
and U10452 (N_10452,N_10079,N_10243);
and U10453 (N_10453,N_10034,N_10095);
xor U10454 (N_10454,N_10182,N_10117);
nor U10455 (N_10455,N_10220,N_10100);
and U10456 (N_10456,N_10022,N_10176);
and U10457 (N_10457,N_10242,N_10136);
xnor U10458 (N_10458,N_10150,N_10088);
nand U10459 (N_10459,N_10049,N_10167);
xnor U10460 (N_10460,N_10057,N_10102);
and U10461 (N_10461,N_10243,N_10002);
nand U10462 (N_10462,N_10114,N_10197);
and U10463 (N_10463,N_10028,N_10220);
and U10464 (N_10464,N_10132,N_10183);
nor U10465 (N_10465,N_10166,N_10095);
nand U10466 (N_10466,N_10115,N_10101);
nand U10467 (N_10467,N_10032,N_10081);
xnor U10468 (N_10468,N_10104,N_10001);
nand U10469 (N_10469,N_10181,N_10224);
nand U10470 (N_10470,N_10172,N_10025);
nor U10471 (N_10471,N_10101,N_10048);
nand U10472 (N_10472,N_10059,N_10052);
nand U10473 (N_10473,N_10160,N_10184);
nor U10474 (N_10474,N_10037,N_10027);
or U10475 (N_10475,N_10032,N_10163);
and U10476 (N_10476,N_10146,N_10121);
nand U10477 (N_10477,N_10026,N_10123);
xor U10478 (N_10478,N_10129,N_10011);
xnor U10479 (N_10479,N_10162,N_10160);
xor U10480 (N_10480,N_10215,N_10102);
nand U10481 (N_10481,N_10161,N_10145);
xnor U10482 (N_10482,N_10243,N_10236);
xor U10483 (N_10483,N_10068,N_10154);
or U10484 (N_10484,N_10070,N_10201);
xor U10485 (N_10485,N_10168,N_10193);
nor U10486 (N_10486,N_10035,N_10077);
xnor U10487 (N_10487,N_10067,N_10235);
nand U10488 (N_10488,N_10180,N_10188);
xor U10489 (N_10489,N_10115,N_10141);
xor U10490 (N_10490,N_10139,N_10082);
xnor U10491 (N_10491,N_10203,N_10147);
and U10492 (N_10492,N_10069,N_10035);
or U10493 (N_10493,N_10061,N_10237);
or U10494 (N_10494,N_10088,N_10050);
and U10495 (N_10495,N_10029,N_10233);
nand U10496 (N_10496,N_10018,N_10192);
nand U10497 (N_10497,N_10192,N_10113);
and U10498 (N_10498,N_10149,N_10183);
nor U10499 (N_10499,N_10033,N_10142);
nor U10500 (N_10500,N_10406,N_10274);
nor U10501 (N_10501,N_10391,N_10255);
xor U10502 (N_10502,N_10395,N_10303);
xnor U10503 (N_10503,N_10440,N_10313);
nand U10504 (N_10504,N_10316,N_10467);
or U10505 (N_10505,N_10492,N_10307);
and U10506 (N_10506,N_10481,N_10382);
or U10507 (N_10507,N_10390,N_10432);
nand U10508 (N_10508,N_10396,N_10328);
or U10509 (N_10509,N_10287,N_10374);
or U10510 (N_10510,N_10314,N_10459);
or U10511 (N_10511,N_10368,N_10433);
and U10512 (N_10512,N_10366,N_10372);
and U10513 (N_10513,N_10329,N_10379);
and U10514 (N_10514,N_10480,N_10326);
or U10515 (N_10515,N_10336,N_10405);
or U10516 (N_10516,N_10422,N_10443);
and U10517 (N_10517,N_10387,N_10322);
and U10518 (N_10518,N_10254,N_10334);
or U10519 (N_10519,N_10289,N_10268);
nor U10520 (N_10520,N_10281,N_10337);
and U10521 (N_10521,N_10447,N_10407);
nor U10522 (N_10522,N_10454,N_10449);
or U10523 (N_10523,N_10354,N_10473);
nand U10524 (N_10524,N_10355,N_10394);
and U10525 (N_10525,N_10404,N_10262);
nand U10526 (N_10526,N_10442,N_10305);
or U10527 (N_10527,N_10421,N_10263);
xor U10528 (N_10528,N_10351,N_10450);
nor U10529 (N_10529,N_10439,N_10284);
xnor U10530 (N_10530,N_10403,N_10413);
xor U10531 (N_10531,N_10451,N_10477);
xnor U10532 (N_10532,N_10344,N_10429);
nand U10533 (N_10533,N_10466,N_10294);
nand U10534 (N_10534,N_10410,N_10399);
and U10535 (N_10535,N_10295,N_10359);
xor U10536 (N_10536,N_10258,N_10276);
xnor U10537 (N_10537,N_10486,N_10414);
or U10538 (N_10538,N_10332,N_10409);
nand U10539 (N_10539,N_10487,N_10430);
nor U10540 (N_10540,N_10280,N_10318);
xor U10541 (N_10541,N_10312,N_10308);
or U10542 (N_10542,N_10291,N_10386);
nand U10543 (N_10543,N_10369,N_10371);
nor U10544 (N_10544,N_10455,N_10335);
nor U10545 (N_10545,N_10370,N_10469);
nor U10546 (N_10546,N_10476,N_10438);
nor U10547 (N_10547,N_10488,N_10471);
and U10548 (N_10548,N_10376,N_10427);
xor U10549 (N_10549,N_10426,N_10358);
nor U10550 (N_10550,N_10435,N_10304);
or U10551 (N_10551,N_10350,N_10283);
xnor U10552 (N_10552,N_10299,N_10499);
nand U10553 (N_10553,N_10402,N_10494);
and U10554 (N_10554,N_10261,N_10437);
or U10555 (N_10555,N_10259,N_10356);
nor U10556 (N_10556,N_10484,N_10398);
and U10557 (N_10557,N_10257,N_10453);
and U10558 (N_10558,N_10460,N_10419);
xor U10559 (N_10559,N_10463,N_10448);
or U10560 (N_10560,N_10385,N_10252);
nor U10561 (N_10561,N_10306,N_10320);
nand U10562 (N_10562,N_10286,N_10383);
and U10563 (N_10563,N_10300,N_10345);
or U10564 (N_10564,N_10348,N_10464);
nor U10565 (N_10565,N_10365,N_10397);
or U10566 (N_10566,N_10415,N_10482);
or U10567 (N_10567,N_10330,N_10367);
nor U10568 (N_10568,N_10267,N_10324);
and U10569 (N_10569,N_10290,N_10282);
xnor U10570 (N_10570,N_10485,N_10341);
and U10571 (N_10571,N_10364,N_10317);
nor U10572 (N_10572,N_10444,N_10457);
or U10573 (N_10573,N_10325,N_10462);
or U10574 (N_10574,N_10441,N_10251);
nand U10575 (N_10575,N_10417,N_10333);
or U10576 (N_10576,N_10310,N_10446);
nand U10577 (N_10577,N_10297,N_10293);
nand U10578 (N_10578,N_10434,N_10331);
nand U10579 (N_10579,N_10271,N_10436);
nor U10580 (N_10580,N_10445,N_10381);
or U10581 (N_10581,N_10378,N_10420);
or U10582 (N_10582,N_10264,N_10343);
xnor U10583 (N_10583,N_10408,N_10346);
or U10584 (N_10584,N_10256,N_10270);
nor U10585 (N_10585,N_10323,N_10277);
and U10586 (N_10586,N_10362,N_10357);
and U10587 (N_10587,N_10428,N_10483);
xnor U10588 (N_10588,N_10478,N_10279);
nand U10589 (N_10589,N_10479,N_10465);
xnor U10590 (N_10590,N_10301,N_10302);
xnor U10591 (N_10591,N_10285,N_10470);
or U10592 (N_10592,N_10496,N_10363);
nor U10593 (N_10593,N_10352,N_10400);
nor U10594 (N_10594,N_10377,N_10384);
or U10595 (N_10595,N_10452,N_10265);
nor U10596 (N_10596,N_10416,N_10497);
nand U10597 (N_10597,N_10418,N_10353);
and U10598 (N_10598,N_10423,N_10273);
nor U10599 (N_10599,N_10393,N_10474);
nand U10600 (N_10600,N_10489,N_10361);
nor U10601 (N_10601,N_10425,N_10311);
and U10602 (N_10602,N_10315,N_10389);
xnor U10603 (N_10603,N_10338,N_10269);
nor U10604 (N_10604,N_10342,N_10472);
and U10605 (N_10605,N_10424,N_10412);
nand U10606 (N_10606,N_10347,N_10475);
xnor U10607 (N_10607,N_10349,N_10493);
nand U10608 (N_10608,N_10275,N_10490);
nor U10609 (N_10609,N_10392,N_10288);
xor U10610 (N_10610,N_10491,N_10321);
and U10611 (N_10611,N_10461,N_10375);
or U10612 (N_10612,N_10360,N_10327);
xnor U10613 (N_10613,N_10498,N_10319);
nor U10614 (N_10614,N_10292,N_10339);
or U10615 (N_10615,N_10456,N_10309);
nor U10616 (N_10616,N_10340,N_10495);
nand U10617 (N_10617,N_10401,N_10296);
or U10618 (N_10618,N_10278,N_10250);
nor U10619 (N_10619,N_10431,N_10411);
and U10620 (N_10620,N_10380,N_10388);
and U10621 (N_10621,N_10458,N_10272);
and U10622 (N_10622,N_10468,N_10298);
and U10623 (N_10623,N_10266,N_10373);
xor U10624 (N_10624,N_10260,N_10253);
and U10625 (N_10625,N_10497,N_10407);
nand U10626 (N_10626,N_10484,N_10393);
and U10627 (N_10627,N_10271,N_10267);
nor U10628 (N_10628,N_10329,N_10309);
xnor U10629 (N_10629,N_10383,N_10254);
and U10630 (N_10630,N_10328,N_10417);
nand U10631 (N_10631,N_10322,N_10293);
or U10632 (N_10632,N_10259,N_10256);
xnor U10633 (N_10633,N_10283,N_10275);
nand U10634 (N_10634,N_10295,N_10308);
or U10635 (N_10635,N_10319,N_10460);
and U10636 (N_10636,N_10463,N_10401);
and U10637 (N_10637,N_10254,N_10409);
and U10638 (N_10638,N_10295,N_10378);
nor U10639 (N_10639,N_10346,N_10465);
xor U10640 (N_10640,N_10255,N_10429);
or U10641 (N_10641,N_10311,N_10405);
and U10642 (N_10642,N_10408,N_10445);
and U10643 (N_10643,N_10359,N_10352);
nand U10644 (N_10644,N_10449,N_10465);
and U10645 (N_10645,N_10285,N_10250);
and U10646 (N_10646,N_10385,N_10253);
xnor U10647 (N_10647,N_10306,N_10319);
or U10648 (N_10648,N_10448,N_10271);
nor U10649 (N_10649,N_10306,N_10303);
nor U10650 (N_10650,N_10437,N_10268);
and U10651 (N_10651,N_10434,N_10349);
nor U10652 (N_10652,N_10495,N_10369);
and U10653 (N_10653,N_10447,N_10283);
xor U10654 (N_10654,N_10347,N_10298);
and U10655 (N_10655,N_10488,N_10437);
and U10656 (N_10656,N_10444,N_10422);
xor U10657 (N_10657,N_10326,N_10356);
or U10658 (N_10658,N_10277,N_10465);
nor U10659 (N_10659,N_10305,N_10284);
xnor U10660 (N_10660,N_10261,N_10340);
nand U10661 (N_10661,N_10412,N_10271);
or U10662 (N_10662,N_10303,N_10450);
xnor U10663 (N_10663,N_10304,N_10263);
and U10664 (N_10664,N_10443,N_10322);
or U10665 (N_10665,N_10297,N_10250);
xor U10666 (N_10666,N_10270,N_10306);
nand U10667 (N_10667,N_10271,N_10421);
nor U10668 (N_10668,N_10310,N_10387);
nor U10669 (N_10669,N_10350,N_10260);
or U10670 (N_10670,N_10257,N_10423);
nor U10671 (N_10671,N_10420,N_10377);
or U10672 (N_10672,N_10273,N_10304);
and U10673 (N_10673,N_10267,N_10263);
nand U10674 (N_10674,N_10290,N_10318);
and U10675 (N_10675,N_10325,N_10324);
nor U10676 (N_10676,N_10261,N_10442);
nand U10677 (N_10677,N_10400,N_10320);
nand U10678 (N_10678,N_10320,N_10265);
or U10679 (N_10679,N_10365,N_10403);
xnor U10680 (N_10680,N_10356,N_10367);
nor U10681 (N_10681,N_10424,N_10276);
and U10682 (N_10682,N_10419,N_10328);
and U10683 (N_10683,N_10477,N_10392);
nor U10684 (N_10684,N_10325,N_10315);
xnor U10685 (N_10685,N_10391,N_10344);
or U10686 (N_10686,N_10313,N_10480);
nand U10687 (N_10687,N_10358,N_10270);
and U10688 (N_10688,N_10329,N_10337);
nand U10689 (N_10689,N_10286,N_10330);
nor U10690 (N_10690,N_10310,N_10250);
nor U10691 (N_10691,N_10279,N_10391);
nand U10692 (N_10692,N_10304,N_10325);
and U10693 (N_10693,N_10399,N_10325);
nand U10694 (N_10694,N_10302,N_10417);
nor U10695 (N_10695,N_10371,N_10393);
nand U10696 (N_10696,N_10453,N_10401);
and U10697 (N_10697,N_10450,N_10463);
nand U10698 (N_10698,N_10461,N_10456);
nand U10699 (N_10699,N_10388,N_10288);
or U10700 (N_10700,N_10389,N_10425);
nor U10701 (N_10701,N_10396,N_10461);
or U10702 (N_10702,N_10491,N_10467);
nand U10703 (N_10703,N_10363,N_10325);
xor U10704 (N_10704,N_10251,N_10465);
or U10705 (N_10705,N_10312,N_10373);
nand U10706 (N_10706,N_10491,N_10270);
and U10707 (N_10707,N_10283,N_10411);
nor U10708 (N_10708,N_10304,N_10481);
nor U10709 (N_10709,N_10446,N_10261);
or U10710 (N_10710,N_10304,N_10454);
xnor U10711 (N_10711,N_10269,N_10483);
nor U10712 (N_10712,N_10399,N_10306);
nor U10713 (N_10713,N_10302,N_10351);
nor U10714 (N_10714,N_10438,N_10440);
nor U10715 (N_10715,N_10327,N_10263);
nor U10716 (N_10716,N_10339,N_10476);
or U10717 (N_10717,N_10460,N_10280);
nor U10718 (N_10718,N_10452,N_10496);
nand U10719 (N_10719,N_10288,N_10273);
and U10720 (N_10720,N_10250,N_10332);
or U10721 (N_10721,N_10438,N_10313);
and U10722 (N_10722,N_10477,N_10371);
or U10723 (N_10723,N_10365,N_10421);
xnor U10724 (N_10724,N_10379,N_10468);
nor U10725 (N_10725,N_10435,N_10372);
nor U10726 (N_10726,N_10342,N_10359);
nor U10727 (N_10727,N_10306,N_10333);
or U10728 (N_10728,N_10254,N_10320);
nor U10729 (N_10729,N_10460,N_10281);
xnor U10730 (N_10730,N_10483,N_10434);
nor U10731 (N_10731,N_10456,N_10430);
or U10732 (N_10732,N_10348,N_10305);
or U10733 (N_10733,N_10454,N_10479);
nand U10734 (N_10734,N_10494,N_10399);
and U10735 (N_10735,N_10399,N_10328);
or U10736 (N_10736,N_10360,N_10325);
or U10737 (N_10737,N_10299,N_10447);
xor U10738 (N_10738,N_10496,N_10395);
xnor U10739 (N_10739,N_10384,N_10410);
or U10740 (N_10740,N_10350,N_10378);
or U10741 (N_10741,N_10384,N_10437);
nand U10742 (N_10742,N_10318,N_10321);
or U10743 (N_10743,N_10406,N_10320);
or U10744 (N_10744,N_10423,N_10357);
or U10745 (N_10745,N_10447,N_10313);
nor U10746 (N_10746,N_10345,N_10413);
nor U10747 (N_10747,N_10394,N_10416);
nand U10748 (N_10748,N_10370,N_10273);
or U10749 (N_10749,N_10388,N_10361);
nor U10750 (N_10750,N_10503,N_10567);
nand U10751 (N_10751,N_10511,N_10577);
and U10752 (N_10752,N_10630,N_10593);
or U10753 (N_10753,N_10501,N_10587);
and U10754 (N_10754,N_10608,N_10584);
nand U10755 (N_10755,N_10537,N_10551);
nand U10756 (N_10756,N_10696,N_10609);
xnor U10757 (N_10757,N_10535,N_10582);
or U10758 (N_10758,N_10560,N_10728);
nand U10759 (N_10759,N_10602,N_10627);
nor U10760 (N_10760,N_10644,N_10617);
xor U10761 (N_10761,N_10512,N_10637);
nor U10762 (N_10762,N_10658,N_10685);
nand U10763 (N_10763,N_10682,N_10524);
or U10764 (N_10764,N_10645,N_10723);
or U10765 (N_10765,N_10674,N_10592);
nor U10766 (N_10766,N_10745,N_10739);
and U10767 (N_10767,N_10538,N_10545);
and U10768 (N_10768,N_10746,N_10707);
nand U10769 (N_10769,N_10556,N_10724);
nor U10770 (N_10770,N_10604,N_10588);
nand U10771 (N_10771,N_10607,N_10583);
xnor U10772 (N_10772,N_10736,N_10529);
or U10773 (N_10773,N_10576,N_10650);
nor U10774 (N_10774,N_10549,N_10701);
nand U10775 (N_10775,N_10709,N_10710);
xnor U10776 (N_10776,N_10615,N_10639);
and U10777 (N_10777,N_10695,N_10526);
nand U10778 (N_10778,N_10633,N_10680);
nand U10779 (N_10779,N_10660,N_10548);
xor U10780 (N_10780,N_10613,N_10507);
nand U10781 (N_10781,N_10727,N_10638);
or U10782 (N_10782,N_10666,N_10681);
nor U10783 (N_10783,N_10523,N_10585);
xor U10784 (N_10784,N_10580,N_10743);
or U10785 (N_10785,N_10670,N_10667);
or U10786 (N_10786,N_10561,N_10508);
nor U10787 (N_10787,N_10744,N_10546);
nand U10788 (N_10788,N_10505,N_10568);
and U10789 (N_10789,N_10654,N_10656);
xor U10790 (N_10790,N_10514,N_10694);
nand U10791 (N_10791,N_10601,N_10741);
or U10792 (N_10792,N_10525,N_10502);
nor U10793 (N_10793,N_10732,N_10510);
nand U10794 (N_10794,N_10687,N_10621);
or U10795 (N_10795,N_10530,N_10699);
or U10796 (N_10796,N_10590,N_10622);
and U10797 (N_10797,N_10562,N_10605);
nor U10798 (N_10798,N_10597,N_10726);
and U10799 (N_10799,N_10624,N_10634);
nor U10800 (N_10800,N_10661,N_10737);
xnor U10801 (N_10801,N_10703,N_10669);
nor U10802 (N_10802,N_10657,N_10683);
nor U10803 (N_10803,N_10594,N_10673);
xnor U10804 (N_10804,N_10749,N_10536);
nor U10805 (N_10805,N_10659,N_10702);
xnor U10806 (N_10806,N_10722,N_10611);
xor U10807 (N_10807,N_10714,N_10569);
or U10808 (N_10808,N_10619,N_10572);
nand U10809 (N_10809,N_10693,N_10632);
xor U10810 (N_10810,N_10516,N_10672);
nand U10811 (N_10811,N_10740,N_10653);
nor U10812 (N_10812,N_10628,N_10570);
nor U10813 (N_10813,N_10563,N_10566);
or U10814 (N_10814,N_10500,N_10506);
nor U10815 (N_10815,N_10677,N_10708);
nand U10816 (N_10816,N_10629,N_10547);
and U10817 (N_10817,N_10684,N_10555);
nand U10818 (N_10818,N_10640,N_10618);
nand U10819 (N_10819,N_10649,N_10513);
or U10820 (N_10820,N_10614,N_10571);
or U10821 (N_10821,N_10543,N_10620);
nand U10822 (N_10822,N_10623,N_10747);
or U10823 (N_10823,N_10655,N_10676);
or U10824 (N_10824,N_10531,N_10719);
and U10825 (N_10825,N_10610,N_10733);
and U10826 (N_10826,N_10697,N_10616);
or U10827 (N_10827,N_10641,N_10519);
xor U10828 (N_10828,N_10721,N_10711);
and U10829 (N_10829,N_10731,N_10651);
xnor U10830 (N_10830,N_10573,N_10534);
nand U10831 (N_10831,N_10668,N_10557);
xor U10832 (N_10832,N_10662,N_10678);
or U10833 (N_10833,N_10603,N_10559);
nor U10834 (N_10834,N_10706,N_10663);
or U10835 (N_10835,N_10648,N_10635);
nand U10836 (N_10836,N_10522,N_10586);
nor U10837 (N_10837,N_10717,N_10690);
nand U10838 (N_10838,N_10689,N_10598);
or U10839 (N_10839,N_10518,N_10575);
or U10840 (N_10840,N_10626,N_10558);
and U10841 (N_10841,N_10540,N_10713);
nand U10842 (N_10842,N_10552,N_10544);
nor U10843 (N_10843,N_10675,N_10565);
or U10844 (N_10844,N_10692,N_10679);
xor U10845 (N_10845,N_10718,N_10700);
nor U10846 (N_10846,N_10521,N_10738);
nor U10847 (N_10847,N_10606,N_10730);
and U10848 (N_10848,N_10578,N_10691);
or U10849 (N_10849,N_10642,N_10596);
nor U10850 (N_10850,N_10591,N_10504);
xnor U10851 (N_10851,N_10520,N_10612);
or U10852 (N_10852,N_10665,N_10729);
nor U10853 (N_10853,N_10734,N_10600);
or U10854 (N_10854,N_10712,N_10528);
nor U10855 (N_10855,N_10646,N_10742);
nor U10856 (N_10856,N_10647,N_10595);
or U10857 (N_10857,N_10515,N_10698);
nand U10858 (N_10858,N_10589,N_10564);
nor U10859 (N_10859,N_10625,N_10532);
xnor U10860 (N_10860,N_10509,N_10725);
and U10861 (N_10861,N_10539,N_10704);
and U10862 (N_10862,N_10553,N_10705);
nor U10863 (N_10863,N_10652,N_10735);
nor U10864 (N_10864,N_10542,N_10636);
and U10865 (N_10865,N_10574,N_10631);
nand U10866 (N_10866,N_10748,N_10579);
nand U10867 (N_10867,N_10599,N_10581);
nor U10868 (N_10868,N_10688,N_10550);
and U10869 (N_10869,N_10643,N_10664);
xor U10870 (N_10870,N_10554,N_10541);
nor U10871 (N_10871,N_10533,N_10720);
nor U10872 (N_10872,N_10671,N_10716);
and U10873 (N_10873,N_10715,N_10527);
and U10874 (N_10874,N_10517,N_10686);
xor U10875 (N_10875,N_10652,N_10662);
or U10876 (N_10876,N_10711,N_10553);
and U10877 (N_10877,N_10677,N_10739);
nand U10878 (N_10878,N_10542,N_10626);
xnor U10879 (N_10879,N_10509,N_10674);
nand U10880 (N_10880,N_10545,N_10681);
or U10881 (N_10881,N_10710,N_10731);
or U10882 (N_10882,N_10688,N_10607);
and U10883 (N_10883,N_10566,N_10578);
nand U10884 (N_10884,N_10631,N_10675);
nand U10885 (N_10885,N_10748,N_10594);
nand U10886 (N_10886,N_10503,N_10733);
xnor U10887 (N_10887,N_10554,N_10613);
or U10888 (N_10888,N_10735,N_10658);
and U10889 (N_10889,N_10720,N_10726);
nand U10890 (N_10890,N_10717,N_10708);
nor U10891 (N_10891,N_10549,N_10714);
nand U10892 (N_10892,N_10726,N_10575);
nand U10893 (N_10893,N_10747,N_10545);
and U10894 (N_10894,N_10721,N_10646);
xnor U10895 (N_10895,N_10643,N_10650);
nor U10896 (N_10896,N_10687,N_10563);
xor U10897 (N_10897,N_10586,N_10557);
nand U10898 (N_10898,N_10730,N_10623);
nand U10899 (N_10899,N_10502,N_10655);
and U10900 (N_10900,N_10578,N_10639);
or U10901 (N_10901,N_10610,N_10543);
xnor U10902 (N_10902,N_10527,N_10550);
nand U10903 (N_10903,N_10670,N_10530);
nor U10904 (N_10904,N_10736,N_10724);
and U10905 (N_10905,N_10591,N_10735);
and U10906 (N_10906,N_10694,N_10690);
and U10907 (N_10907,N_10666,N_10673);
nand U10908 (N_10908,N_10612,N_10712);
or U10909 (N_10909,N_10645,N_10548);
xor U10910 (N_10910,N_10500,N_10711);
nor U10911 (N_10911,N_10712,N_10730);
and U10912 (N_10912,N_10673,N_10640);
xor U10913 (N_10913,N_10667,N_10711);
nand U10914 (N_10914,N_10734,N_10507);
and U10915 (N_10915,N_10682,N_10679);
nand U10916 (N_10916,N_10692,N_10706);
xnor U10917 (N_10917,N_10746,N_10749);
xnor U10918 (N_10918,N_10624,N_10567);
nand U10919 (N_10919,N_10523,N_10673);
xor U10920 (N_10920,N_10560,N_10530);
and U10921 (N_10921,N_10523,N_10517);
xnor U10922 (N_10922,N_10616,N_10675);
or U10923 (N_10923,N_10736,N_10718);
or U10924 (N_10924,N_10603,N_10653);
or U10925 (N_10925,N_10552,N_10675);
nor U10926 (N_10926,N_10645,N_10650);
nand U10927 (N_10927,N_10568,N_10694);
or U10928 (N_10928,N_10709,N_10502);
xnor U10929 (N_10929,N_10696,N_10688);
and U10930 (N_10930,N_10693,N_10531);
xor U10931 (N_10931,N_10699,N_10714);
and U10932 (N_10932,N_10617,N_10576);
and U10933 (N_10933,N_10503,N_10532);
and U10934 (N_10934,N_10534,N_10601);
nor U10935 (N_10935,N_10555,N_10614);
and U10936 (N_10936,N_10627,N_10733);
nand U10937 (N_10937,N_10692,N_10510);
or U10938 (N_10938,N_10509,N_10579);
and U10939 (N_10939,N_10716,N_10532);
nor U10940 (N_10940,N_10685,N_10742);
nor U10941 (N_10941,N_10637,N_10604);
xor U10942 (N_10942,N_10594,N_10606);
nor U10943 (N_10943,N_10519,N_10574);
nand U10944 (N_10944,N_10622,N_10648);
and U10945 (N_10945,N_10507,N_10738);
nor U10946 (N_10946,N_10709,N_10591);
and U10947 (N_10947,N_10515,N_10679);
nor U10948 (N_10948,N_10554,N_10638);
xnor U10949 (N_10949,N_10608,N_10684);
xor U10950 (N_10950,N_10671,N_10713);
and U10951 (N_10951,N_10526,N_10589);
and U10952 (N_10952,N_10524,N_10603);
xor U10953 (N_10953,N_10620,N_10622);
or U10954 (N_10954,N_10528,N_10518);
or U10955 (N_10955,N_10637,N_10578);
and U10956 (N_10956,N_10630,N_10505);
nor U10957 (N_10957,N_10535,N_10589);
xnor U10958 (N_10958,N_10673,N_10701);
and U10959 (N_10959,N_10506,N_10537);
nand U10960 (N_10960,N_10549,N_10599);
nor U10961 (N_10961,N_10528,N_10644);
nand U10962 (N_10962,N_10544,N_10688);
and U10963 (N_10963,N_10670,N_10525);
or U10964 (N_10964,N_10537,N_10719);
xnor U10965 (N_10965,N_10635,N_10742);
xnor U10966 (N_10966,N_10531,N_10697);
nand U10967 (N_10967,N_10641,N_10505);
xor U10968 (N_10968,N_10515,N_10526);
nand U10969 (N_10969,N_10744,N_10560);
and U10970 (N_10970,N_10506,N_10731);
nor U10971 (N_10971,N_10506,N_10614);
xor U10972 (N_10972,N_10696,N_10733);
and U10973 (N_10973,N_10575,N_10542);
xor U10974 (N_10974,N_10663,N_10668);
nor U10975 (N_10975,N_10738,N_10656);
xnor U10976 (N_10976,N_10610,N_10629);
nand U10977 (N_10977,N_10563,N_10607);
or U10978 (N_10978,N_10512,N_10722);
xnor U10979 (N_10979,N_10542,N_10624);
or U10980 (N_10980,N_10639,N_10528);
xor U10981 (N_10981,N_10602,N_10641);
or U10982 (N_10982,N_10576,N_10560);
nor U10983 (N_10983,N_10524,N_10730);
or U10984 (N_10984,N_10727,N_10606);
nor U10985 (N_10985,N_10592,N_10583);
or U10986 (N_10986,N_10517,N_10720);
nand U10987 (N_10987,N_10740,N_10726);
or U10988 (N_10988,N_10525,N_10610);
and U10989 (N_10989,N_10697,N_10740);
and U10990 (N_10990,N_10717,N_10608);
nor U10991 (N_10991,N_10721,N_10625);
xnor U10992 (N_10992,N_10739,N_10704);
xor U10993 (N_10993,N_10703,N_10532);
nor U10994 (N_10994,N_10535,N_10532);
nand U10995 (N_10995,N_10743,N_10546);
and U10996 (N_10996,N_10538,N_10521);
nand U10997 (N_10997,N_10588,N_10536);
nor U10998 (N_10998,N_10736,N_10742);
and U10999 (N_10999,N_10742,N_10590);
and U11000 (N_11000,N_10786,N_10763);
nand U11001 (N_11001,N_10964,N_10837);
nor U11002 (N_11002,N_10753,N_10790);
or U11003 (N_11003,N_10810,N_10993);
and U11004 (N_11004,N_10992,N_10808);
and U11005 (N_11005,N_10969,N_10829);
or U11006 (N_11006,N_10978,N_10852);
and U11007 (N_11007,N_10901,N_10777);
xnor U11008 (N_11008,N_10860,N_10856);
or U11009 (N_11009,N_10818,N_10984);
nand U11010 (N_11010,N_10869,N_10922);
or U11011 (N_11011,N_10785,N_10776);
nor U11012 (N_11012,N_10815,N_10890);
and U11013 (N_11013,N_10876,N_10858);
nand U11014 (N_11014,N_10976,N_10887);
nor U11015 (N_11015,N_10755,N_10806);
nand U11016 (N_11016,N_10968,N_10778);
xnor U11017 (N_11017,N_10935,N_10927);
nand U11018 (N_11018,N_10775,N_10816);
nor U11019 (N_11019,N_10881,N_10884);
and U11020 (N_11020,N_10916,N_10904);
nor U11021 (N_11021,N_10934,N_10932);
and U11022 (N_11022,N_10900,N_10991);
xor U11023 (N_11023,N_10765,N_10805);
and U11024 (N_11024,N_10819,N_10854);
or U11025 (N_11025,N_10842,N_10811);
and U11026 (N_11026,N_10908,N_10754);
xnor U11027 (N_11027,N_10960,N_10886);
xor U11028 (N_11028,N_10864,N_10997);
xnor U11029 (N_11029,N_10821,N_10787);
and U11030 (N_11030,N_10871,N_10920);
or U11031 (N_11031,N_10813,N_10836);
or U11032 (N_11032,N_10865,N_10980);
nor U11033 (N_11033,N_10870,N_10803);
nor U11034 (N_11034,N_10918,N_10761);
nor U11035 (N_11035,N_10906,N_10955);
nor U11036 (N_11036,N_10974,N_10767);
and U11037 (N_11037,N_10948,N_10982);
xor U11038 (N_11038,N_10788,N_10781);
nand U11039 (N_11039,N_10970,N_10990);
and U11040 (N_11040,N_10931,N_10863);
xor U11041 (N_11041,N_10894,N_10866);
nand U11042 (N_11042,N_10945,N_10933);
or U11043 (N_11043,N_10757,N_10834);
xor U11044 (N_11044,N_10798,N_10833);
nand U11045 (N_11045,N_10826,N_10942);
nand U11046 (N_11046,N_10999,N_10959);
nor U11047 (N_11047,N_10971,N_10929);
and U11048 (N_11048,N_10950,N_10878);
or U11049 (N_11049,N_10868,N_10921);
xor U11050 (N_11050,N_10953,N_10845);
xor U11051 (N_11051,N_10914,N_10930);
or U11052 (N_11052,N_10941,N_10902);
nor U11053 (N_11053,N_10796,N_10962);
and U11054 (N_11054,N_10897,N_10792);
nor U11055 (N_11055,N_10958,N_10977);
nand U11056 (N_11056,N_10967,N_10907);
or U11057 (N_11057,N_10917,N_10807);
xnor U11058 (N_11058,N_10804,N_10772);
nand U11059 (N_11059,N_10769,N_10831);
nor U11060 (N_11060,N_10812,N_10951);
nand U11061 (N_11061,N_10752,N_10892);
and U11062 (N_11062,N_10986,N_10998);
or U11063 (N_11063,N_10895,N_10764);
or U11064 (N_11064,N_10983,N_10913);
or U11065 (N_11065,N_10972,N_10839);
nor U11066 (N_11066,N_10840,N_10975);
or U11067 (N_11067,N_10928,N_10824);
or U11068 (N_11068,N_10872,N_10938);
xor U11069 (N_11069,N_10989,N_10770);
or U11070 (N_11070,N_10843,N_10957);
nor U11071 (N_11071,N_10943,N_10911);
xor U11072 (N_11072,N_10827,N_10963);
nor U11073 (N_11073,N_10830,N_10793);
or U11074 (N_11074,N_10784,N_10877);
xor U11075 (N_11075,N_10848,N_10924);
nor U11076 (N_11076,N_10995,N_10762);
xnor U11077 (N_11077,N_10853,N_10779);
xnor U11078 (N_11078,N_10954,N_10841);
and U11079 (N_11079,N_10825,N_10783);
xnor U11080 (N_11080,N_10828,N_10800);
xor U11081 (N_11081,N_10956,N_10780);
and U11082 (N_11082,N_10802,N_10889);
xor U11083 (N_11083,N_10799,N_10794);
xor U11084 (N_11084,N_10940,N_10814);
and U11085 (N_11085,N_10979,N_10888);
nand U11086 (N_11086,N_10880,N_10851);
or U11087 (N_11087,N_10883,N_10879);
nor U11088 (N_11088,N_10822,N_10893);
or U11089 (N_11089,N_10909,N_10899);
nand U11090 (N_11090,N_10791,N_10936);
nor U11091 (N_11091,N_10850,N_10905);
or U11092 (N_11092,N_10981,N_10857);
or U11093 (N_11093,N_10823,N_10952);
or U11094 (N_11094,N_10867,N_10875);
and U11095 (N_11095,N_10919,N_10855);
and U11096 (N_11096,N_10771,N_10987);
nor U11097 (N_11097,N_10925,N_10966);
nand U11098 (N_11098,N_10859,N_10861);
xor U11099 (N_11099,N_10797,N_10961);
xnor U11100 (N_11100,N_10944,N_10832);
nor U11101 (N_11101,N_10882,N_10912);
and U11102 (N_11102,N_10846,N_10996);
or U11103 (N_11103,N_10766,N_10873);
xor U11104 (N_11104,N_10891,N_10985);
nor U11105 (N_11105,N_10862,N_10949);
and U11106 (N_11106,N_10903,N_10926);
or U11107 (N_11107,N_10874,N_10896);
xor U11108 (N_11108,N_10835,N_10965);
xor U11109 (N_11109,N_10988,N_10947);
nor U11110 (N_11110,N_10885,N_10939);
and U11111 (N_11111,N_10774,N_10795);
and U11112 (N_11112,N_10915,N_10768);
or U11113 (N_11113,N_10898,N_10751);
nand U11114 (N_11114,N_10809,N_10994);
or U11115 (N_11115,N_10801,N_10844);
xnor U11116 (N_11116,N_10759,N_10789);
xor U11117 (N_11117,N_10817,N_10820);
xor U11118 (N_11118,N_10923,N_10756);
nor U11119 (N_11119,N_10849,N_10782);
or U11120 (N_11120,N_10910,N_10758);
or U11121 (N_11121,N_10773,N_10750);
and U11122 (N_11122,N_10937,N_10847);
or U11123 (N_11123,N_10973,N_10760);
nor U11124 (N_11124,N_10946,N_10838);
xnor U11125 (N_11125,N_10769,N_10972);
xor U11126 (N_11126,N_10886,N_10853);
or U11127 (N_11127,N_10754,N_10770);
nor U11128 (N_11128,N_10760,N_10911);
nor U11129 (N_11129,N_10799,N_10795);
xnor U11130 (N_11130,N_10763,N_10823);
and U11131 (N_11131,N_10881,N_10871);
and U11132 (N_11132,N_10836,N_10762);
and U11133 (N_11133,N_10973,N_10948);
xnor U11134 (N_11134,N_10931,N_10793);
and U11135 (N_11135,N_10941,N_10997);
nor U11136 (N_11136,N_10828,N_10941);
and U11137 (N_11137,N_10873,N_10914);
and U11138 (N_11138,N_10785,N_10830);
xor U11139 (N_11139,N_10963,N_10894);
xnor U11140 (N_11140,N_10894,N_10964);
nand U11141 (N_11141,N_10873,N_10960);
xor U11142 (N_11142,N_10854,N_10993);
and U11143 (N_11143,N_10866,N_10837);
nor U11144 (N_11144,N_10955,N_10823);
and U11145 (N_11145,N_10808,N_10874);
and U11146 (N_11146,N_10830,N_10942);
nand U11147 (N_11147,N_10770,N_10987);
xnor U11148 (N_11148,N_10950,N_10916);
nor U11149 (N_11149,N_10879,N_10928);
nor U11150 (N_11150,N_10981,N_10762);
nand U11151 (N_11151,N_10838,N_10910);
nand U11152 (N_11152,N_10793,N_10846);
or U11153 (N_11153,N_10928,N_10986);
xor U11154 (N_11154,N_10766,N_10966);
or U11155 (N_11155,N_10794,N_10993);
nand U11156 (N_11156,N_10818,N_10956);
and U11157 (N_11157,N_10998,N_10774);
nand U11158 (N_11158,N_10991,N_10904);
xnor U11159 (N_11159,N_10826,N_10903);
xor U11160 (N_11160,N_10950,N_10997);
nand U11161 (N_11161,N_10878,N_10974);
nand U11162 (N_11162,N_10818,N_10969);
xnor U11163 (N_11163,N_10828,N_10970);
nor U11164 (N_11164,N_10917,N_10813);
and U11165 (N_11165,N_10808,N_10954);
nand U11166 (N_11166,N_10831,N_10833);
xor U11167 (N_11167,N_10776,N_10957);
and U11168 (N_11168,N_10918,N_10836);
nand U11169 (N_11169,N_10916,N_10895);
nor U11170 (N_11170,N_10824,N_10971);
or U11171 (N_11171,N_10903,N_10925);
xnor U11172 (N_11172,N_10802,N_10906);
nor U11173 (N_11173,N_10924,N_10854);
and U11174 (N_11174,N_10995,N_10911);
nand U11175 (N_11175,N_10895,N_10921);
and U11176 (N_11176,N_10780,N_10985);
or U11177 (N_11177,N_10948,N_10816);
nor U11178 (N_11178,N_10935,N_10756);
xor U11179 (N_11179,N_10870,N_10999);
or U11180 (N_11180,N_10760,N_10920);
xor U11181 (N_11181,N_10916,N_10933);
xor U11182 (N_11182,N_10941,N_10872);
xor U11183 (N_11183,N_10762,N_10952);
nand U11184 (N_11184,N_10944,N_10767);
nor U11185 (N_11185,N_10997,N_10829);
nor U11186 (N_11186,N_10856,N_10853);
and U11187 (N_11187,N_10960,N_10971);
nor U11188 (N_11188,N_10851,N_10791);
nand U11189 (N_11189,N_10971,N_10886);
nor U11190 (N_11190,N_10800,N_10996);
nor U11191 (N_11191,N_10831,N_10870);
nor U11192 (N_11192,N_10946,N_10990);
nand U11193 (N_11193,N_10944,N_10877);
nand U11194 (N_11194,N_10828,N_10769);
nand U11195 (N_11195,N_10884,N_10990);
nor U11196 (N_11196,N_10871,N_10837);
nand U11197 (N_11197,N_10887,N_10871);
xnor U11198 (N_11198,N_10901,N_10842);
nand U11199 (N_11199,N_10816,N_10820);
nor U11200 (N_11200,N_10785,N_10867);
nand U11201 (N_11201,N_10935,N_10810);
xor U11202 (N_11202,N_10872,N_10811);
xnor U11203 (N_11203,N_10961,N_10791);
xnor U11204 (N_11204,N_10780,N_10879);
xor U11205 (N_11205,N_10910,N_10821);
and U11206 (N_11206,N_10756,N_10830);
nor U11207 (N_11207,N_10941,N_10924);
or U11208 (N_11208,N_10975,N_10920);
nand U11209 (N_11209,N_10911,N_10796);
and U11210 (N_11210,N_10958,N_10801);
and U11211 (N_11211,N_10930,N_10919);
and U11212 (N_11212,N_10757,N_10784);
nand U11213 (N_11213,N_10986,N_10792);
nand U11214 (N_11214,N_10987,N_10784);
xor U11215 (N_11215,N_10862,N_10843);
and U11216 (N_11216,N_10916,N_10934);
nor U11217 (N_11217,N_10834,N_10768);
or U11218 (N_11218,N_10873,N_10915);
nand U11219 (N_11219,N_10978,N_10957);
and U11220 (N_11220,N_10906,N_10932);
and U11221 (N_11221,N_10923,N_10834);
xnor U11222 (N_11222,N_10852,N_10957);
xnor U11223 (N_11223,N_10875,N_10821);
xor U11224 (N_11224,N_10762,N_10887);
and U11225 (N_11225,N_10799,N_10754);
xor U11226 (N_11226,N_10826,N_10787);
xor U11227 (N_11227,N_10837,N_10994);
nor U11228 (N_11228,N_10977,N_10993);
or U11229 (N_11229,N_10804,N_10789);
xor U11230 (N_11230,N_10964,N_10841);
and U11231 (N_11231,N_10785,N_10903);
nand U11232 (N_11232,N_10881,N_10818);
and U11233 (N_11233,N_10991,N_10847);
or U11234 (N_11234,N_10827,N_10750);
or U11235 (N_11235,N_10907,N_10782);
xor U11236 (N_11236,N_10773,N_10908);
nor U11237 (N_11237,N_10987,N_10759);
xor U11238 (N_11238,N_10925,N_10884);
or U11239 (N_11239,N_10882,N_10860);
nor U11240 (N_11240,N_10872,N_10774);
or U11241 (N_11241,N_10994,N_10903);
and U11242 (N_11242,N_10935,N_10892);
or U11243 (N_11243,N_10877,N_10818);
or U11244 (N_11244,N_10849,N_10817);
xor U11245 (N_11245,N_10854,N_10915);
or U11246 (N_11246,N_10809,N_10883);
xnor U11247 (N_11247,N_10969,N_10984);
or U11248 (N_11248,N_10893,N_10966);
nor U11249 (N_11249,N_10893,N_10896);
and U11250 (N_11250,N_11008,N_11146);
nand U11251 (N_11251,N_11129,N_11185);
or U11252 (N_11252,N_11235,N_11144);
and U11253 (N_11253,N_11222,N_11032);
or U11254 (N_11254,N_11111,N_11205);
nand U11255 (N_11255,N_11033,N_11014);
nor U11256 (N_11256,N_11180,N_11124);
nor U11257 (N_11257,N_11175,N_11099);
and U11258 (N_11258,N_11155,N_11041);
xor U11259 (N_11259,N_11031,N_11219);
or U11260 (N_11260,N_11215,N_11081);
or U11261 (N_11261,N_11045,N_11224);
nand U11262 (N_11262,N_11198,N_11104);
xnor U11263 (N_11263,N_11244,N_11236);
nand U11264 (N_11264,N_11165,N_11040);
and U11265 (N_11265,N_11068,N_11039);
or U11266 (N_11266,N_11220,N_11110);
xor U11267 (N_11267,N_11214,N_11054);
and U11268 (N_11268,N_11186,N_11161);
or U11269 (N_11269,N_11107,N_11184);
xor U11270 (N_11270,N_11202,N_11141);
or U11271 (N_11271,N_11140,N_11177);
nand U11272 (N_11272,N_11062,N_11103);
or U11273 (N_11273,N_11150,N_11075);
nand U11274 (N_11274,N_11018,N_11163);
and U11275 (N_11275,N_11006,N_11048);
and U11276 (N_11276,N_11061,N_11022);
nor U11277 (N_11277,N_11097,N_11206);
nand U11278 (N_11278,N_11135,N_11001);
nand U11279 (N_11279,N_11003,N_11195);
or U11280 (N_11280,N_11055,N_11060);
and U11281 (N_11281,N_11194,N_11059);
or U11282 (N_11282,N_11230,N_11171);
nor U11283 (N_11283,N_11197,N_11066);
and U11284 (N_11284,N_11096,N_11020);
nor U11285 (N_11285,N_11080,N_11123);
nand U11286 (N_11286,N_11213,N_11176);
nor U11287 (N_11287,N_11046,N_11094);
xor U11288 (N_11288,N_11083,N_11078);
nand U11289 (N_11289,N_11208,N_11183);
nand U11290 (N_11290,N_11070,N_11173);
nand U11291 (N_11291,N_11145,N_11164);
xnor U11292 (N_11292,N_11121,N_11127);
nor U11293 (N_11293,N_11000,N_11038);
nor U11294 (N_11294,N_11227,N_11226);
nand U11295 (N_11295,N_11034,N_11095);
and U11296 (N_11296,N_11229,N_11026);
and U11297 (N_11297,N_11112,N_11092);
nor U11298 (N_11298,N_11225,N_11168);
nand U11299 (N_11299,N_11147,N_11057);
nor U11300 (N_11300,N_11138,N_11149);
and U11301 (N_11301,N_11241,N_11025);
or U11302 (N_11302,N_11073,N_11212);
and U11303 (N_11303,N_11117,N_11108);
nand U11304 (N_11304,N_11228,N_11119);
nor U11305 (N_11305,N_11148,N_11067);
and U11306 (N_11306,N_11091,N_11203);
nand U11307 (N_11307,N_11114,N_11231);
nand U11308 (N_11308,N_11043,N_11133);
nand U11309 (N_11309,N_11182,N_11063);
xnor U11310 (N_11310,N_11115,N_11088);
nand U11311 (N_11311,N_11120,N_11074);
nor U11312 (N_11312,N_11153,N_11209);
and U11313 (N_11313,N_11101,N_11130);
nand U11314 (N_11314,N_11105,N_11169);
nand U11315 (N_11315,N_11232,N_11102);
nor U11316 (N_11316,N_11207,N_11246);
and U11317 (N_11317,N_11179,N_11056);
and U11318 (N_11318,N_11217,N_11084);
nor U11319 (N_11319,N_11132,N_11223);
nor U11320 (N_11320,N_11024,N_11017);
and U11321 (N_11321,N_11050,N_11089);
xor U11322 (N_11322,N_11154,N_11065);
xor U11323 (N_11323,N_11204,N_11143);
nand U11324 (N_11324,N_11234,N_11052);
nor U11325 (N_11325,N_11239,N_11109);
nand U11326 (N_11326,N_11142,N_11201);
or U11327 (N_11327,N_11100,N_11221);
and U11328 (N_11328,N_11166,N_11023);
nand U11329 (N_11329,N_11245,N_11090);
xnor U11330 (N_11330,N_11192,N_11036);
nor U11331 (N_11331,N_11243,N_11128);
and U11332 (N_11332,N_11113,N_11152);
xnor U11333 (N_11333,N_11072,N_11167);
nand U11334 (N_11334,N_11237,N_11007);
or U11335 (N_11335,N_11016,N_11086);
and U11336 (N_11336,N_11076,N_11122);
xor U11337 (N_11337,N_11051,N_11012);
or U11338 (N_11338,N_11199,N_11210);
nand U11339 (N_11339,N_11188,N_11053);
xor U11340 (N_11340,N_11082,N_11071);
nor U11341 (N_11341,N_11178,N_11170);
nand U11342 (N_11342,N_11189,N_11238);
or U11343 (N_11343,N_11218,N_11044);
or U11344 (N_11344,N_11233,N_11248);
nand U11345 (N_11345,N_11196,N_11042);
xor U11346 (N_11346,N_11029,N_11125);
xor U11347 (N_11347,N_11093,N_11193);
or U11348 (N_11348,N_11240,N_11159);
xnor U11349 (N_11349,N_11191,N_11077);
nor U11350 (N_11350,N_11181,N_11200);
xor U11351 (N_11351,N_11010,N_11158);
nor U11352 (N_11352,N_11162,N_11131);
nor U11353 (N_11353,N_11027,N_11126);
nor U11354 (N_11354,N_11172,N_11058);
nor U11355 (N_11355,N_11009,N_11118);
nor U11356 (N_11356,N_11087,N_11187);
or U11357 (N_11357,N_11019,N_11005);
nor U11358 (N_11358,N_11157,N_11247);
and U11359 (N_11359,N_11211,N_11190);
and U11360 (N_11360,N_11079,N_11002);
nor U11361 (N_11361,N_11030,N_11249);
or U11362 (N_11362,N_11037,N_11151);
or U11363 (N_11363,N_11064,N_11116);
or U11364 (N_11364,N_11098,N_11216);
or U11365 (N_11365,N_11106,N_11174);
nor U11366 (N_11366,N_11013,N_11139);
and U11367 (N_11367,N_11085,N_11160);
or U11368 (N_11368,N_11069,N_11028);
nor U11369 (N_11369,N_11134,N_11047);
or U11370 (N_11370,N_11011,N_11004);
nand U11371 (N_11371,N_11242,N_11015);
and U11372 (N_11372,N_11136,N_11137);
or U11373 (N_11373,N_11035,N_11156);
or U11374 (N_11374,N_11021,N_11049);
and U11375 (N_11375,N_11033,N_11187);
nand U11376 (N_11376,N_11191,N_11203);
xnor U11377 (N_11377,N_11021,N_11186);
nor U11378 (N_11378,N_11058,N_11126);
or U11379 (N_11379,N_11238,N_11010);
nand U11380 (N_11380,N_11237,N_11194);
and U11381 (N_11381,N_11045,N_11056);
and U11382 (N_11382,N_11191,N_11170);
xor U11383 (N_11383,N_11094,N_11164);
xnor U11384 (N_11384,N_11134,N_11077);
nor U11385 (N_11385,N_11051,N_11020);
xor U11386 (N_11386,N_11234,N_11198);
or U11387 (N_11387,N_11076,N_11020);
nand U11388 (N_11388,N_11059,N_11103);
and U11389 (N_11389,N_11083,N_11199);
nor U11390 (N_11390,N_11102,N_11049);
nor U11391 (N_11391,N_11046,N_11127);
nand U11392 (N_11392,N_11112,N_11189);
xor U11393 (N_11393,N_11173,N_11225);
and U11394 (N_11394,N_11163,N_11151);
nand U11395 (N_11395,N_11186,N_11158);
nor U11396 (N_11396,N_11003,N_11172);
xnor U11397 (N_11397,N_11016,N_11200);
nand U11398 (N_11398,N_11034,N_11119);
or U11399 (N_11399,N_11136,N_11008);
xnor U11400 (N_11400,N_11244,N_11083);
xnor U11401 (N_11401,N_11005,N_11211);
xor U11402 (N_11402,N_11185,N_11156);
or U11403 (N_11403,N_11119,N_11127);
xnor U11404 (N_11404,N_11030,N_11108);
nor U11405 (N_11405,N_11072,N_11222);
or U11406 (N_11406,N_11137,N_11112);
nand U11407 (N_11407,N_11159,N_11188);
nor U11408 (N_11408,N_11135,N_11149);
or U11409 (N_11409,N_11230,N_11169);
xor U11410 (N_11410,N_11148,N_11091);
and U11411 (N_11411,N_11073,N_11060);
or U11412 (N_11412,N_11217,N_11150);
or U11413 (N_11413,N_11022,N_11071);
and U11414 (N_11414,N_11186,N_11109);
nand U11415 (N_11415,N_11148,N_11184);
or U11416 (N_11416,N_11224,N_11061);
or U11417 (N_11417,N_11146,N_11129);
xor U11418 (N_11418,N_11061,N_11127);
and U11419 (N_11419,N_11005,N_11070);
nor U11420 (N_11420,N_11174,N_11083);
nor U11421 (N_11421,N_11154,N_11075);
nand U11422 (N_11422,N_11181,N_11053);
and U11423 (N_11423,N_11176,N_11243);
nor U11424 (N_11424,N_11125,N_11087);
nor U11425 (N_11425,N_11018,N_11043);
xor U11426 (N_11426,N_11157,N_11014);
nor U11427 (N_11427,N_11116,N_11170);
nand U11428 (N_11428,N_11003,N_11046);
and U11429 (N_11429,N_11161,N_11059);
nor U11430 (N_11430,N_11192,N_11196);
or U11431 (N_11431,N_11212,N_11247);
or U11432 (N_11432,N_11239,N_11154);
and U11433 (N_11433,N_11091,N_11221);
nor U11434 (N_11434,N_11061,N_11023);
and U11435 (N_11435,N_11024,N_11045);
nand U11436 (N_11436,N_11128,N_11049);
and U11437 (N_11437,N_11191,N_11221);
or U11438 (N_11438,N_11224,N_11155);
xnor U11439 (N_11439,N_11135,N_11228);
and U11440 (N_11440,N_11021,N_11235);
xnor U11441 (N_11441,N_11151,N_11006);
nor U11442 (N_11442,N_11163,N_11027);
nand U11443 (N_11443,N_11249,N_11245);
nand U11444 (N_11444,N_11004,N_11228);
nand U11445 (N_11445,N_11053,N_11195);
nand U11446 (N_11446,N_11095,N_11200);
and U11447 (N_11447,N_11142,N_11023);
or U11448 (N_11448,N_11183,N_11237);
nor U11449 (N_11449,N_11194,N_11179);
nor U11450 (N_11450,N_11063,N_11064);
or U11451 (N_11451,N_11027,N_11244);
nor U11452 (N_11452,N_11194,N_11023);
and U11453 (N_11453,N_11198,N_11173);
nor U11454 (N_11454,N_11068,N_11014);
nor U11455 (N_11455,N_11181,N_11023);
and U11456 (N_11456,N_11236,N_11056);
and U11457 (N_11457,N_11151,N_11023);
nor U11458 (N_11458,N_11130,N_11225);
and U11459 (N_11459,N_11005,N_11022);
nand U11460 (N_11460,N_11205,N_11129);
or U11461 (N_11461,N_11138,N_11115);
or U11462 (N_11462,N_11234,N_11121);
and U11463 (N_11463,N_11199,N_11213);
and U11464 (N_11464,N_11100,N_11159);
and U11465 (N_11465,N_11098,N_11145);
nor U11466 (N_11466,N_11067,N_11194);
or U11467 (N_11467,N_11163,N_11200);
and U11468 (N_11468,N_11247,N_11070);
nor U11469 (N_11469,N_11120,N_11011);
nor U11470 (N_11470,N_11028,N_11188);
nand U11471 (N_11471,N_11086,N_11178);
and U11472 (N_11472,N_11178,N_11186);
xor U11473 (N_11473,N_11237,N_11171);
or U11474 (N_11474,N_11057,N_11046);
xor U11475 (N_11475,N_11224,N_11094);
and U11476 (N_11476,N_11063,N_11009);
nand U11477 (N_11477,N_11097,N_11026);
nand U11478 (N_11478,N_11044,N_11198);
and U11479 (N_11479,N_11039,N_11176);
nand U11480 (N_11480,N_11028,N_11105);
nand U11481 (N_11481,N_11016,N_11133);
or U11482 (N_11482,N_11241,N_11212);
or U11483 (N_11483,N_11156,N_11227);
nor U11484 (N_11484,N_11045,N_11051);
and U11485 (N_11485,N_11237,N_11245);
xor U11486 (N_11486,N_11173,N_11144);
nand U11487 (N_11487,N_11035,N_11139);
nand U11488 (N_11488,N_11125,N_11063);
xor U11489 (N_11489,N_11004,N_11177);
nand U11490 (N_11490,N_11052,N_11235);
nand U11491 (N_11491,N_11023,N_11143);
xor U11492 (N_11492,N_11005,N_11002);
xnor U11493 (N_11493,N_11187,N_11109);
and U11494 (N_11494,N_11217,N_11101);
or U11495 (N_11495,N_11153,N_11086);
nand U11496 (N_11496,N_11118,N_11108);
and U11497 (N_11497,N_11015,N_11110);
xnor U11498 (N_11498,N_11153,N_11136);
and U11499 (N_11499,N_11047,N_11177);
or U11500 (N_11500,N_11407,N_11347);
xnor U11501 (N_11501,N_11382,N_11474);
or U11502 (N_11502,N_11343,N_11399);
and U11503 (N_11503,N_11422,N_11287);
and U11504 (N_11504,N_11278,N_11436);
nor U11505 (N_11505,N_11442,N_11279);
and U11506 (N_11506,N_11440,N_11308);
xor U11507 (N_11507,N_11266,N_11445);
nor U11508 (N_11508,N_11314,N_11448);
and U11509 (N_11509,N_11286,N_11340);
nor U11510 (N_11510,N_11411,N_11482);
nand U11511 (N_11511,N_11403,N_11273);
or U11512 (N_11512,N_11484,N_11318);
nand U11513 (N_11513,N_11370,N_11323);
or U11514 (N_11514,N_11268,N_11424);
nor U11515 (N_11515,N_11470,N_11281);
xnor U11516 (N_11516,N_11313,N_11291);
or U11517 (N_11517,N_11406,N_11401);
nand U11518 (N_11518,N_11414,N_11297);
xor U11519 (N_11519,N_11438,N_11427);
nand U11520 (N_11520,N_11375,N_11489);
or U11521 (N_11521,N_11369,N_11433);
or U11522 (N_11522,N_11439,N_11321);
or U11523 (N_11523,N_11267,N_11367);
xor U11524 (N_11524,N_11296,N_11301);
and U11525 (N_11525,N_11264,N_11376);
xor U11526 (N_11526,N_11263,N_11462);
or U11527 (N_11527,N_11410,N_11345);
and U11528 (N_11528,N_11395,N_11361);
nor U11529 (N_11529,N_11366,N_11451);
nand U11530 (N_11530,N_11430,N_11374);
and U11531 (N_11531,N_11404,N_11255);
xnor U11532 (N_11532,N_11458,N_11312);
nand U11533 (N_11533,N_11260,N_11326);
or U11534 (N_11534,N_11475,N_11276);
and U11535 (N_11535,N_11288,N_11289);
xnor U11536 (N_11536,N_11381,N_11494);
or U11537 (N_11537,N_11311,N_11416);
nand U11538 (N_11538,N_11292,N_11271);
xnor U11539 (N_11539,N_11284,N_11338);
xor U11540 (N_11540,N_11269,N_11394);
nand U11541 (N_11541,N_11274,N_11364);
xor U11542 (N_11542,N_11348,N_11463);
or U11543 (N_11543,N_11473,N_11425);
and U11544 (N_11544,N_11293,N_11490);
xnor U11545 (N_11545,N_11467,N_11342);
xnor U11546 (N_11546,N_11443,N_11402);
nor U11547 (N_11547,N_11421,N_11261);
nand U11548 (N_11548,N_11253,N_11252);
xnor U11549 (N_11549,N_11447,N_11466);
or U11550 (N_11550,N_11455,N_11449);
nor U11551 (N_11551,N_11272,N_11397);
nand U11552 (N_11552,N_11259,N_11275);
nor U11553 (N_11553,N_11486,N_11357);
xor U11554 (N_11554,N_11371,N_11299);
nor U11555 (N_11555,N_11335,N_11251);
or U11556 (N_11556,N_11478,N_11387);
or U11557 (N_11557,N_11302,N_11465);
nand U11558 (N_11558,N_11306,N_11356);
or U11559 (N_11559,N_11454,N_11346);
and U11560 (N_11560,N_11294,N_11295);
nand U11561 (N_11561,N_11457,N_11316);
xor U11562 (N_11562,N_11310,N_11479);
or U11563 (N_11563,N_11483,N_11480);
and U11564 (N_11564,N_11329,N_11488);
xnor U11565 (N_11565,N_11320,N_11354);
nor U11566 (N_11566,N_11363,N_11495);
nand U11567 (N_11567,N_11351,N_11469);
xor U11568 (N_11568,N_11417,N_11352);
and U11569 (N_11569,N_11334,N_11290);
nor U11570 (N_11570,N_11437,N_11336);
nand U11571 (N_11571,N_11464,N_11405);
nor U11572 (N_11572,N_11396,N_11429);
nand U11573 (N_11573,N_11415,N_11420);
nor U11574 (N_11574,N_11383,N_11468);
or U11575 (N_11575,N_11446,N_11377);
or U11576 (N_11576,N_11324,N_11368);
nor U11577 (N_11577,N_11487,N_11280);
nor U11578 (N_11578,N_11325,N_11476);
nand U11579 (N_11579,N_11461,N_11378);
nor U11580 (N_11580,N_11398,N_11389);
and U11581 (N_11581,N_11388,N_11460);
nand U11582 (N_11582,N_11491,N_11331);
nand U11583 (N_11583,N_11258,N_11341);
nand U11584 (N_11584,N_11250,N_11441);
and U11585 (N_11585,N_11477,N_11270);
xnor U11586 (N_11586,N_11315,N_11435);
nor U11587 (N_11587,N_11319,N_11282);
and U11588 (N_11588,N_11283,N_11423);
nand U11589 (N_11589,N_11408,N_11385);
xor U11590 (N_11590,N_11419,N_11365);
nand U11591 (N_11591,N_11358,N_11412);
nand U11592 (N_11592,N_11450,N_11353);
nand U11593 (N_11593,N_11492,N_11328);
xor U11594 (N_11594,N_11392,N_11386);
xnor U11595 (N_11595,N_11355,N_11456);
and U11596 (N_11596,N_11337,N_11426);
nand U11597 (N_11597,N_11307,N_11305);
or U11598 (N_11598,N_11344,N_11384);
and U11599 (N_11599,N_11418,N_11257);
nor U11600 (N_11600,N_11262,N_11360);
nand U11601 (N_11601,N_11327,N_11256);
xor U11602 (N_11602,N_11453,N_11373);
nor U11603 (N_11603,N_11380,N_11409);
and U11604 (N_11604,N_11390,N_11444);
nor U11605 (N_11605,N_11481,N_11330);
xor U11606 (N_11606,N_11304,N_11333);
or U11607 (N_11607,N_11332,N_11362);
xnor U11608 (N_11608,N_11493,N_11413);
xor U11609 (N_11609,N_11372,N_11452);
nand U11610 (N_11610,N_11459,N_11498);
xor U11611 (N_11611,N_11434,N_11391);
xnor U11612 (N_11612,N_11339,N_11285);
and U11613 (N_11613,N_11428,N_11496);
or U11614 (N_11614,N_11298,N_11431);
xor U11615 (N_11615,N_11400,N_11359);
or U11616 (N_11616,N_11471,N_11379);
and U11617 (N_11617,N_11349,N_11254);
or U11618 (N_11618,N_11485,N_11303);
nor U11619 (N_11619,N_11472,N_11499);
nand U11620 (N_11620,N_11432,N_11309);
nand U11621 (N_11621,N_11497,N_11277);
nand U11622 (N_11622,N_11300,N_11393);
xor U11623 (N_11623,N_11322,N_11265);
xnor U11624 (N_11624,N_11317,N_11350);
or U11625 (N_11625,N_11414,N_11301);
and U11626 (N_11626,N_11322,N_11334);
nor U11627 (N_11627,N_11382,N_11292);
and U11628 (N_11628,N_11472,N_11269);
and U11629 (N_11629,N_11276,N_11412);
or U11630 (N_11630,N_11425,N_11397);
nand U11631 (N_11631,N_11354,N_11355);
nor U11632 (N_11632,N_11303,N_11477);
and U11633 (N_11633,N_11267,N_11473);
nor U11634 (N_11634,N_11381,N_11373);
nor U11635 (N_11635,N_11497,N_11387);
or U11636 (N_11636,N_11313,N_11292);
xnor U11637 (N_11637,N_11449,N_11476);
and U11638 (N_11638,N_11373,N_11472);
nand U11639 (N_11639,N_11434,N_11481);
nor U11640 (N_11640,N_11330,N_11479);
or U11641 (N_11641,N_11350,N_11278);
and U11642 (N_11642,N_11403,N_11457);
and U11643 (N_11643,N_11275,N_11398);
or U11644 (N_11644,N_11424,N_11443);
nor U11645 (N_11645,N_11442,N_11381);
nor U11646 (N_11646,N_11496,N_11278);
nor U11647 (N_11647,N_11318,N_11289);
nand U11648 (N_11648,N_11490,N_11382);
or U11649 (N_11649,N_11403,N_11445);
nor U11650 (N_11650,N_11367,N_11394);
nor U11651 (N_11651,N_11466,N_11383);
nor U11652 (N_11652,N_11299,N_11356);
or U11653 (N_11653,N_11485,N_11267);
xor U11654 (N_11654,N_11355,N_11319);
nor U11655 (N_11655,N_11391,N_11492);
or U11656 (N_11656,N_11408,N_11499);
or U11657 (N_11657,N_11330,N_11486);
xor U11658 (N_11658,N_11284,N_11356);
xor U11659 (N_11659,N_11432,N_11379);
xnor U11660 (N_11660,N_11305,N_11383);
nor U11661 (N_11661,N_11499,N_11364);
nor U11662 (N_11662,N_11475,N_11489);
nand U11663 (N_11663,N_11341,N_11433);
nand U11664 (N_11664,N_11262,N_11354);
or U11665 (N_11665,N_11296,N_11434);
and U11666 (N_11666,N_11437,N_11316);
xor U11667 (N_11667,N_11383,N_11460);
nand U11668 (N_11668,N_11423,N_11250);
or U11669 (N_11669,N_11338,N_11458);
and U11670 (N_11670,N_11435,N_11250);
or U11671 (N_11671,N_11276,N_11283);
nor U11672 (N_11672,N_11372,N_11309);
or U11673 (N_11673,N_11356,N_11275);
nand U11674 (N_11674,N_11256,N_11287);
nand U11675 (N_11675,N_11437,N_11284);
nand U11676 (N_11676,N_11255,N_11460);
or U11677 (N_11677,N_11453,N_11271);
nand U11678 (N_11678,N_11316,N_11498);
or U11679 (N_11679,N_11358,N_11319);
xnor U11680 (N_11680,N_11275,N_11413);
or U11681 (N_11681,N_11344,N_11298);
or U11682 (N_11682,N_11388,N_11256);
and U11683 (N_11683,N_11320,N_11381);
xor U11684 (N_11684,N_11489,N_11355);
and U11685 (N_11685,N_11441,N_11432);
and U11686 (N_11686,N_11436,N_11260);
xnor U11687 (N_11687,N_11397,N_11350);
xor U11688 (N_11688,N_11400,N_11431);
nor U11689 (N_11689,N_11254,N_11378);
and U11690 (N_11690,N_11337,N_11480);
and U11691 (N_11691,N_11398,N_11328);
and U11692 (N_11692,N_11257,N_11442);
xnor U11693 (N_11693,N_11380,N_11388);
and U11694 (N_11694,N_11276,N_11368);
nand U11695 (N_11695,N_11490,N_11301);
or U11696 (N_11696,N_11493,N_11444);
or U11697 (N_11697,N_11370,N_11478);
xnor U11698 (N_11698,N_11374,N_11463);
or U11699 (N_11699,N_11381,N_11432);
nor U11700 (N_11700,N_11261,N_11461);
nand U11701 (N_11701,N_11306,N_11256);
nand U11702 (N_11702,N_11286,N_11262);
or U11703 (N_11703,N_11426,N_11343);
or U11704 (N_11704,N_11275,N_11436);
nor U11705 (N_11705,N_11427,N_11406);
and U11706 (N_11706,N_11320,N_11287);
and U11707 (N_11707,N_11388,N_11298);
xnor U11708 (N_11708,N_11446,N_11310);
or U11709 (N_11709,N_11390,N_11257);
nand U11710 (N_11710,N_11285,N_11335);
xor U11711 (N_11711,N_11413,N_11319);
nor U11712 (N_11712,N_11295,N_11438);
nand U11713 (N_11713,N_11349,N_11290);
xnor U11714 (N_11714,N_11457,N_11490);
and U11715 (N_11715,N_11295,N_11465);
or U11716 (N_11716,N_11347,N_11411);
xor U11717 (N_11717,N_11445,N_11417);
nor U11718 (N_11718,N_11411,N_11344);
nor U11719 (N_11719,N_11497,N_11330);
xnor U11720 (N_11720,N_11373,N_11251);
or U11721 (N_11721,N_11329,N_11270);
or U11722 (N_11722,N_11423,N_11340);
xor U11723 (N_11723,N_11377,N_11291);
and U11724 (N_11724,N_11311,N_11398);
and U11725 (N_11725,N_11385,N_11469);
xnor U11726 (N_11726,N_11339,N_11290);
nor U11727 (N_11727,N_11454,N_11401);
nand U11728 (N_11728,N_11274,N_11475);
nor U11729 (N_11729,N_11468,N_11343);
or U11730 (N_11730,N_11470,N_11480);
nor U11731 (N_11731,N_11437,N_11486);
or U11732 (N_11732,N_11255,N_11463);
nand U11733 (N_11733,N_11348,N_11433);
nand U11734 (N_11734,N_11418,N_11492);
nor U11735 (N_11735,N_11403,N_11281);
nor U11736 (N_11736,N_11426,N_11398);
nand U11737 (N_11737,N_11405,N_11369);
nand U11738 (N_11738,N_11467,N_11317);
xor U11739 (N_11739,N_11449,N_11498);
and U11740 (N_11740,N_11252,N_11405);
nor U11741 (N_11741,N_11491,N_11391);
xnor U11742 (N_11742,N_11321,N_11320);
or U11743 (N_11743,N_11361,N_11389);
xnor U11744 (N_11744,N_11334,N_11294);
or U11745 (N_11745,N_11427,N_11268);
nand U11746 (N_11746,N_11337,N_11444);
nor U11747 (N_11747,N_11302,N_11448);
nand U11748 (N_11748,N_11410,N_11486);
nor U11749 (N_11749,N_11333,N_11433);
and U11750 (N_11750,N_11533,N_11726);
nand U11751 (N_11751,N_11746,N_11605);
or U11752 (N_11752,N_11577,N_11601);
nor U11753 (N_11753,N_11509,N_11600);
or U11754 (N_11754,N_11626,N_11570);
and U11755 (N_11755,N_11687,N_11721);
and U11756 (N_11756,N_11650,N_11547);
and U11757 (N_11757,N_11523,N_11546);
nand U11758 (N_11758,N_11707,N_11564);
and U11759 (N_11759,N_11566,N_11619);
nand U11760 (N_11760,N_11514,N_11580);
and U11761 (N_11761,N_11645,N_11696);
and U11762 (N_11762,N_11727,N_11537);
nand U11763 (N_11763,N_11604,N_11544);
or U11764 (N_11764,N_11713,N_11525);
xnor U11765 (N_11765,N_11524,N_11669);
or U11766 (N_11766,N_11730,N_11629);
xnor U11767 (N_11767,N_11723,N_11639);
and U11768 (N_11768,N_11710,N_11584);
and U11769 (N_11769,N_11704,N_11715);
and U11770 (N_11770,N_11505,N_11578);
or U11771 (N_11771,N_11628,N_11586);
or U11772 (N_11772,N_11615,N_11595);
or U11773 (N_11773,N_11722,N_11531);
and U11774 (N_11774,N_11711,N_11582);
xor U11775 (N_11775,N_11656,N_11548);
xor U11776 (N_11776,N_11703,N_11686);
and U11777 (N_11777,N_11611,N_11562);
nor U11778 (N_11778,N_11738,N_11660);
nand U11779 (N_11779,N_11549,N_11596);
and U11780 (N_11780,N_11612,N_11520);
and U11781 (N_11781,N_11624,N_11569);
nor U11782 (N_11782,N_11712,N_11728);
nor U11783 (N_11783,N_11545,N_11672);
and U11784 (N_11784,N_11668,N_11654);
and U11785 (N_11785,N_11517,N_11534);
nor U11786 (N_11786,N_11719,N_11742);
nor U11787 (N_11787,N_11538,N_11695);
and U11788 (N_11788,N_11554,N_11558);
and U11789 (N_11789,N_11732,N_11588);
nand U11790 (N_11790,N_11676,N_11658);
xnor U11791 (N_11791,N_11621,N_11557);
nand U11792 (N_11792,N_11568,N_11593);
xnor U11793 (N_11793,N_11706,N_11617);
nand U11794 (N_11794,N_11653,N_11599);
and U11795 (N_11795,N_11565,N_11683);
nor U11796 (N_11796,N_11607,N_11665);
xor U11797 (N_11797,N_11519,N_11709);
nand U11798 (N_11798,N_11518,N_11510);
or U11799 (N_11799,N_11708,N_11526);
or U11800 (N_11800,N_11512,N_11576);
nor U11801 (N_11801,N_11618,N_11649);
and U11802 (N_11802,N_11583,N_11507);
xnor U11803 (N_11803,N_11684,N_11572);
nand U11804 (N_11804,N_11508,N_11506);
nor U11805 (N_11805,N_11504,N_11725);
nand U11806 (N_11806,N_11671,N_11592);
xor U11807 (N_11807,N_11602,N_11622);
or U11808 (N_11808,N_11674,N_11529);
nor U11809 (N_11809,N_11646,N_11694);
and U11810 (N_11810,N_11530,N_11623);
and U11811 (N_11811,N_11585,N_11736);
nand U11812 (N_11812,N_11643,N_11614);
and U11813 (N_11813,N_11542,N_11731);
nand U11814 (N_11814,N_11527,N_11667);
xnor U11815 (N_11815,N_11535,N_11501);
nor U11816 (N_11816,N_11613,N_11745);
nor U11817 (N_11817,N_11522,N_11589);
or U11818 (N_11818,N_11591,N_11641);
or U11819 (N_11819,N_11692,N_11521);
nor U11820 (N_11820,N_11575,N_11532);
nor U11821 (N_11821,N_11567,N_11636);
xnor U11822 (N_11822,N_11550,N_11733);
or U11823 (N_11823,N_11574,N_11689);
nor U11824 (N_11824,N_11573,N_11740);
xnor U11825 (N_11825,N_11682,N_11563);
nand U11826 (N_11826,N_11515,N_11690);
nor U11827 (N_11827,N_11701,N_11640);
xor U11828 (N_11828,N_11749,N_11632);
xor U11829 (N_11829,N_11555,N_11644);
nand U11830 (N_11830,N_11642,N_11579);
nand U11831 (N_11831,N_11597,N_11729);
and U11832 (N_11832,N_11691,N_11648);
and U11833 (N_11833,N_11541,N_11659);
and U11834 (N_11834,N_11741,N_11747);
nand U11835 (N_11835,N_11528,N_11625);
and U11836 (N_11836,N_11606,N_11657);
or U11837 (N_11837,N_11571,N_11718);
nand U11838 (N_11838,N_11536,N_11551);
xor U11839 (N_11839,N_11697,N_11503);
nand U11840 (N_11840,N_11655,N_11590);
nor U11841 (N_11841,N_11670,N_11699);
or U11842 (N_11842,N_11680,N_11678);
or U11843 (N_11843,N_11664,N_11734);
xnor U11844 (N_11844,N_11502,N_11553);
xor U11845 (N_11845,N_11511,N_11561);
and U11846 (N_11846,N_11717,N_11552);
and U11847 (N_11847,N_11685,N_11610);
nor U11848 (N_11848,N_11702,N_11735);
xnor U11849 (N_11849,N_11603,N_11543);
nor U11850 (N_11850,N_11631,N_11620);
xor U11851 (N_11851,N_11500,N_11705);
xnor U11852 (N_11852,N_11630,N_11673);
xor U11853 (N_11853,N_11666,N_11744);
or U11854 (N_11854,N_11677,N_11587);
or U11855 (N_11855,N_11662,N_11638);
nor U11856 (N_11856,N_11556,N_11516);
nand U11857 (N_11857,N_11609,N_11739);
nand U11858 (N_11858,N_11724,N_11661);
or U11859 (N_11859,N_11616,N_11559);
xor U11860 (N_11860,N_11513,N_11675);
nor U11861 (N_11861,N_11598,N_11647);
or U11862 (N_11862,N_11581,N_11748);
and U11863 (N_11863,N_11540,N_11700);
and U11864 (N_11864,N_11693,N_11743);
or U11865 (N_11865,N_11720,N_11539);
nand U11866 (N_11866,N_11663,N_11637);
nor U11867 (N_11867,N_11633,N_11634);
or U11868 (N_11868,N_11698,N_11681);
or U11869 (N_11869,N_11635,N_11716);
nand U11870 (N_11870,N_11714,N_11679);
and U11871 (N_11871,N_11688,N_11560);
and U11872 (N_11872,N_11737,N_11594);
nand U11873 (N_11873,N_11652,N_11627);
and U11874 (N_11874,N_11651,N_11608);
xnor U11875 (N_11875,N_11681,N_11510);
nand U11876 (N_11876,N_11720,N_11543);
xnor U11877 (N_11877,N_11585,N_11621);
and U11878 (N_11878,N_11611,N_11659);
or U11879 (N_11879,N_11514,N_11550);
and U11880 (N_11880,N_11590,N_11726);
nor U11881 (N_11881,N_11539,N_11629);
and U11882 (N_11882,N_11594,N_11634);
nor U11883 (N_11883,N_11660,N_11596);
nand U11884 (N_11884,N_11589,N_11674);
or U11885 (N_11885,N_11589,N_11664);
xnor U11886 (N_11886,N_11735,N_11502);
or U11887 (N_11887,N_11686,N_11591);
nor U11888 (N_11888,N_11699,N_11661);
nor U11889 (N_11889,N_11734,N_11666);
xnor U11890 (N_11890,N_11555,N_11675);
nand U11891 (N_11891,N_11505,N_11600);
nand U11892 (N_11892,N_11590,N_11503);
and U11893 (N_11893,N_11532,N_11553);
nand U11894 (N_11894,N_11501,N_11738);
xnor U11895 (N_11895,N_11528,N_11507);
xor U11896 (N_11896,N_11506,N_11525);
nand U11897 (N_11897,N_11514,N_11666);
and U11898 (N_11898,N_11655,N_11671);
xor U11899 (N_11899,N_11597,N_11716);
or U11900 (N_11900,N_11553,N_11524);
or U11901 (N_11901,N_11575,N_11656);
or U11902 (N_11902,N_11664,N_11692);
or U11903 (N_11903,N_11648,N_11624);
nand U11904 (N_11904,N_11539,N_11623);
or U11905 (N_11905,N_11587,N_11604);
xnor U11906 (N_11906,N_11733,N_11741);
xor U11907 (N_11907,N_11650,N_11590);
nor U11908 (N_11908,N_11514,N_11604);
xor U11909 (N_11909,N_11530,N_11510);
xnor U11910 (N_11910,N_11694,N_11691);
nand U11911 (N_11911,N_11532,N_11744);
nand U11912 (N_11912,N_11641,N_11539);
xor U11913 (N_11913,N_11611,N_11503);
nand U11914 (N_11914,N_11635,N_11743);
or U11915 (N_11915,N_11576,N_11603);
nor U11916 (N_11916,N_11671,N_11707);
or U11917 (N_11917,N_11741,N_11711);
nand U11918 (N_11918,N_11576,N_11626);
and U11919 (N_11919,N_11596,N_11734);
nand U11920 (N_11920,N_11683,N_11528);
nand U11921 (N_11921,N_11687,N_11739);
nor U11922 (N_11922,N_11603,N_11557);
nor U11923 (N_11923,N_11509,N_11677);
and U11924 (N_11924,N_11743,N_11584);
nand U11925 (N_11925,N_11739,N_11671);
nor U11926 (N_11926,N_11667,N_11661);
or U11927 (N_11927,N_11684,N_11706);
and U11928 (N_11928,N_11617,N_11536);
or U11929 (N_11929,N_11517,N_11732);
nor U11930 (N_11930,N_11520,N_11591);
xor U11931 (N_11931,N_11511,N_11675);
and U11932 (N_11932,N_11602,N_11589);
nand U11933 (N_11933,N_11570,N_11584);
xor U11934 (N_11934,N_11682,N_11621);
or U11935 (N_11935,N_11663,N_11724);
and U11936 (N_11936,N_11635,N_11663);
nor U11937 (N_11937,N_11651,N_11702);
nor U11938 (N_11938,N_11599,N_11594);
or U11939 (N_11939,N_11669,N_11585);
xor U11940 (N_11940,N_11565,N_11702);
and U11941 (N_11941,N_11558,N_11699);
xnor U11942 (N_11942,N_11709,N_11514);
or U11943 (N_11943,N_11680,N_11563);
and U11944 (N_11944,N_11697,N_11685);
nor U11945 (N_11945,N_11728,N_11631);
nand U11946 (N_11946,N_11596,N_11653);
nor U11947 (N_11947,N_11697,N_11742);
xnor U11948 (N_11948,N_11578,N_11687);
or U11949 (N_11949,N_11671,N_11696);
and U11950 (N_11950,N_11608,N_11596);
and U11951 (N_11951,N_11527,N_11676);
xor U11952 (N_11952,N_11679,N_11743);
nand U11953 (N_11953,N_11717,N_11565);
and U11954 (N_11954,N_11646,N_11533);
nor U11955 (N_11955,N_11521,N_11507);
or U11956 (N_11956,N_11520,N_11743);
and U11957 (N_11957,N_11706,N_11570);
xnor U11958 (N_11958,N_11628,N_11504);
or U11959 (N_11959,N_11558,N_11515);
and U11960 (N_11960,N_11637,N_11506);
nand U11961 (N_11961,N_11521,N_11706);
xnor U11962 (N_11962,N_11633,N_11666);
or U11963 (N_11963,N_11709,N_11663);
and U11964 (N_11964,N_11623,N_11629);
nand U11965 (N_11965,N_11610,N_11616);
or U11966 (N_11966,N_11653,N_11518);
xnor U11967 (N_11967,N_11567,N_11701);
xor U11968 (N_11968,N_11705,N_11624);
xnor U11969 (N_11969,N_11729,N_11673);
or U11970 (N_11970,N_11599,N_11749);
and U11971 (N_11971,N_11658,N_11516);
and U11972 (N_11972,N_11652,N_11645);
nor U11973 (N_11973,N_11734,N_11678);
or U11974 (N_11974,N_11654,N_11501);
and U11975 (N_11975,N_11572,N_11542);
nor U11976 (N_11976,N_11503,N_11691);
and U11977 (N_11977,N_11582,N_11573);
and U11978 (N_11978,N_11640,N_11718);
nor U11979 (N_11979,N_11645,N_11708);
and U11980 (N_11980,N_11568,N_11710);
nand U11981 (N_11981,N_11513,N_11554);
nor U11982 (N_11982,N_11739,N_11512);
xor U11983 (N_11983,N_11518,N_11620);
or U11984 (N_11984,N_11679,N_11601);
nor U11985 (N_11985,N_11723,N_11610);
nand U11986 (N_11986,N_11550,N_11743);
and U11987 (N_11987,N_11691,N_11501);
nand U11988 (N_11988,N_11640,N_11630);
nor U11989 (N_11989,N_11686,N_11522);
or U11990 (N_11990,N_11744,N_11509);
or U11991 (N_11991,N_11723,N_11660);
and U11992 (N_11992,N_11574,N_11729);
and U11993 (N_11993,N_11658,N_11683);
xnor U11994 (N_11994,N_11672,N_11729);
xnor U11995 (N_11995,N_11580,N_11737);
and U11996 (N_11996,N_11640,N_11672);
nor U11997 (N_11997,N_11724,N_11727);
xnor U11998 (N_11998,N_11745,N_11719);
xnor U11999 (N_11999,N_11637,N_11666);
nand U12000 (N_12000,N_11847,N_11856);
and U12001 (N_12001,N_11768,N_11939);
nand U12002 (N_12002,N_11761,N_11849);
nand U12003 (N_12003,N_11918,N_11770);
or U12004 (N_12004,N_11931,N_11828);
nand U12005 (N_12005,N_11957,N_11857);
or U12006 (N_12006,N_11899,N_11759);
or U12007 (N_12007,N_11925,N_11995);
nor U12008 (N_12008,N_11907,N_11935);
nand U12009 (N_12009,N_11999,N_11822);
and U12010 (N_12010,N_11982,N_11884);
and U12011 (N_12011,N_11806,N_11959);
and U12012 (N_12012,N_11933,N_11890);
and U12013 (N_12013,N_11989,N_11946);
and U12014 (N_12014,N_11750,N_11795);
nor U12015 (N_12015,N_11930,N_11771);
nor U12016 (N_12016,N_11841,N_11862);
or U12017 (N_12017,N_11868,N_11824);
or U12018 (N_12018,N_11793,N_11814);
and U12019 (N_12019,N_11970,N_11881);
nor U12020 (N_12020,N_11848,N_11823);
or U12021 (N_12021,N_11798,N_11948);
nor U12022 (N_12022,N_11880,N_11858);
nor U12023 (N_12023,N_11764,N_11865);
xnor U12024 (N_12024,N_11943,N_11914);
and U12025 (N_12025,N_11846,N_11830);
or U12026 (N_12026,N_11834,N_11808);
and U12027 (N_12027,N_11753,N_11980);
and U12028 (N_12028,N_11934,N_11983);
xor U12029 (N_12029,N_11818,N_11859);
or U12030 (N_12030,N_11988,N_11920);
xnor U12031 (N_12031,N_11961,N_11962);
nand U12032 (N_12032,N_11754,N_11777);
xor U12033 (N_12033,N_11825,N_11973);
xor U12034 (N_12034,N_11775,N_11885);
nand U12035 (N_12035,N_11792,N_11887);
nor U12036 (N_12036,N_11803,N_11987);
nand U12037 (N_12037,N_11952,N_11840);
nor U12038 (N_12038,N_11984,N_11944);
and U12039 (N_12039,N_11924,N_11904);
and U12040 (N_12040,N_11765,N_11863);
or U12041 (N_12041,N_11917,N_11912);
nor U12042 (N_12042,N_11978,N_11872);
and U12043 (N_12043,N_11758,N_11802);
xnor U12044 (N_12044,N_11928,N_11861);
or U12045 (N_12045,N_11850,N_11902);
xor U12046 (N_12046,N_11981,N_11778);
or U12047 (N_12047,N_11901,N_11871);
nand U12048 (N_12048,N_11938,N_11839);
and U12049 (N_12049,N_11804,N_11760);
nand U12050 (N_12050,N_11896,N_11926);
nand U12051 (N_12051,N_11783,N_11947);
nand U12052 (N_12052,N_11782,N_11854);
xnor U12053 (N_12053,N_11936,N_11786);
and U12054 (N_12054,N_11756,N_11892);
xor U12055 (N_12055,N_11974,N_11893);
xnor U12056 (N_12056,N_11977,N_11831);
nand U12057 (N_12057,N_11968,N_11903);
nand U12058 (N_12058,N_11942,N_11763);
or U12059 (N_12059,N_11811,N_11787);
and U12060 (N_12060,N_11826,N_11784);
nor U12061 (N_12061,N_11867,N_11915);
nor U12062 (N_12062,N_11807,N_11766);
nor U12063 (N_12063,N_11755,N_11801);
or U12064 (N_12064,N_11788,N_11929);
xor U12065 (N_12065,N_11954,N_11975);
nor U12066 (N_12066,N_11965,N_11949);
and U12067 (N_12067,N_11781,N_11866);
xor U12068 (N_12068,N_11972,N_11950);
or U12069 (N_12069,N_11886,N_11853);
or U12070 (N_12070,N_11888,N_11816);
or U12071 (N_12071,N_11875,N_11891);
xor U12072 (N_12072,N_11879,N_11956);
nand U12073 (N_12073,N_11794,N_11911);
xnor U12074 (N_12074,N_11877,N_11955);
or U12075 (N_12075,N_11797,N_11810);
nand U12076 (N_12076,N_11922,N_11927);
and U12077 (N_12077,N_11855,N_11908);
nor U12078 (N_12078,N_11963,N_11773);
xor U12079 (N_12079,N_11769,N_11997);
and U12080 (N_12080,N_11979,N_11843);
and U12081 (N_12081,N_11878,N_11821);
and U12082 (N_12082,N_11895,N_11919);
nor U12083 (N_12083,N_11992,N_11762);
nand U12084 (N_12084,N_11845,N_11860);
nor U12085 (N_12085,N_11998,N_11906);
nor U12086 (N_12086,N_11966,N_11785);
or U12087 (N_12087,N_11945,N_11779);
or U12088 (N_12088,N_11951,N_11772);
or U12089 (N_12089,N_11774,N_11837);
nor U12090 (N_12090,N_11883,N_11960);
nand U12091 (N_12091,N_11905,N_11909);
nor U12092 (N_12092,N_11994,N_11851);
nand U12093 (N_12093,N_11874,N_11889);
nor U12094 (N_12094,N_11876,N_11916);
xnor U12095 (N_12095,N_11991,N_11805);
and U12096 (N_12096,N_11780,N_11913);
nand U12097 (N_12097,N_11910,N_11894);
nand U12098 (N_12098,N_11869,N_11882);
nor U12099 (N_12099,N_11767,N_11967);
nand U12100 (N_12100,N_11835,N_11791);
nor U12101 (N_12101,N_11820,N_11819);
xnor U12102 (N_12102,N_11971,N_11969);
or U12103 (N_12103,N_11799,N_11870);
nor U12104 (N_12104,N_11844,N_11932);
nor U12105 (N_12105,N_11833,N_11897);
nor U12106 (N_12106,N_11752,N_11852);
nor U12107 (N_12107,N_11986,N_11836);
or U12108 (N_12108,N_11990,N_11809);
and U12109 (N_12109,N_11842,N_11940);
nor U12110 (N_12110,N_11898,N_11873);
nor U12111 (N_12111,N_11832,N_11976);
xor U12112 (N_12112,N_11941,N_11838);
and U12113 (N_12113,N_11789,N_11864);
and U12114 (N_12114,N_11815,N_11923);
nand U12115 (N_12115,N_11776,N_11757);
and U12116 (N_12116,N_11993,N_11937);
or U12117 (N_12117,N_11958,N_11827);
nor U12118 (N_12118,N_11921,N_11800);
xnor U12119 (N_12119,N_11790,N_11900);
and U12120 (N_12120,N_11796,N_11817);
and U12121 (N_12121,N_11996,N_11985);
and U12122 (N_12122,N_11751,N_11813);
xnor U12123 (N_12123,N_11812,N_11953);
xor U12124 (N_12124,N_11964,N_11829);
xnor U12125 (N_12125,N_11779,N_11924);
nand U12126 (N_12126,N_11996,N_11872);
nand U12127 (N_12127,N_11904,N_11949);
nand U12128 (N_12128,N_11753,N_11819);
xnor U12129 (N_12129,N_11812,N_11877);
nand U12130 (N_12130,N_11877,N_11759);
nand U12131 (N_12131,N_11859,N_11867);
nor U12132 (N_12132,N_11968,N_11984);
or U12133 (N_12133,N_11955,N_11777);
nor U12134 (N_12134,N_11915,N_11865);
xnor U12135 (N_12135,N_11907,N_11801);
and U12136 (N_12136,N_11846,N_11842);
and U12137 (N_12137,N_11750,N_11769);
xnor U12138 (N_12138,N_11882,N_11785);
and U12139 (N_12139,N_11835,N_11786);
nand U12140 (N_12140,N_11781,N_11832);
or U12141 (N_12141,N_11913,N_11893);
or U12142 (N_12142,N_11808,N_11927);
xor U12143 (N_12143,N_11766,N_11846);
or U12144 (N_12144,N_11803,N_11848);
nor U12145 (N_12145,N_11962,N_11900);
nand U12146 (N_12146,N_11796,N_11775);
xor U12147 (N_12147,N_11959,N_11793);
nor U12148 (N_12148,N_11930,N_11991);
nand U12149 (N_12149,N_11760,N_11772);
and U12150 (N_12150,N_11823,N_11788);
nand U12151 (N_12151,N_11787,N_11786);
nor U12152 (N_12152,N_11807,N_11997);
and U12153 (N_12153,N_11751,N_11952);
or U12154 (N_12154,N_11971,N_11985);
nand U12155 (N_12155,N_11996,N_11892);
nand U12156 (N_12156,N_11846,N_11823);
and U12157 (N_12157,N_11790,N_11907);
xor U12158 (N_12158,N_11808,N_11838);
nor U12159 (N_12159,N_11858,N_11883);
or U12160 (N_12160,N_11950,N_11800);
and U12161 (N_12161,N_11818,N_11930);
or U12162 (N_12162,N_11885,N_11977);
or U12163 (N_12163,N_11867,N_11912);
or U12164 (N_12164,N_11759,N_11892);
and U12165 (N_12165,N_11908,N_11819);
or U12166 (N_12166,N_11765,N_11750);
xnor U12167 (N_12167,N_11987,N_11830);
nor U12168 (N_12168,N_11911,N_11767);
or U12169 (N_12169,N_11796,N_11978);
or U12170 (N_12170,N_11969,N_11991);
xnor U12171 (N_12171,N_11894,N_11794);
nand U12172 (N_12172,N_11973,N_11811);
nand U12173 (N_12173,N_11820,N_11984);
nand U12174 (N_12174,N_11863,N_11886);
xnor U12175 (N_12175,N_11958,N_11873);
or U12176 (N_12176,N_11807,N_11860);
nor U12177 (N_12177,N_11816,N_11894);
nand U12178 (N_12178,N_11898,N_11977);
nor U12179 (N_12179,N_11929,N_11778);
and U12180 (N_12180,N_11835,N_11992);
xor U12181 (N_12181,N_11991,N_11794);
nor U12182 (N_12182,N_11919,N_11902);
nand U12183 (N_12183,N_11946,N_11753);
nand U12184 (N_12184,N_11906,N_11888);
nor U12185 (N_12185,N_11859,N_11757);
nor U12186 (N_12186,N_11763,N_11759);
nand U12187 (N_12187,N_11847,N_11779);
nand U12188 (N_12188,N_11966,N_11937);
or U12189 (N_12189,N_11854,N_11995);
nor U12190 (N_12190,N_11863,N_11760);
nor U12191 (N_12191,N_11765,N_11862);
or U12192 (N_12192,N_11809,N_11858);
nor U12193 (N_12193,N_11821,N_11839);
and U12194 (N_12194,N_11870,N_11867);
nor U12195 (N_12195,N_11838,N_11754);
or U12196 (N_12196,N_11903,N_11878);
and U12197 (N_12197,N_11993,N_11759);
and U12198 (N_12198,N_11924,N_11764);
xnor U12199 (N_12199,N_11935,N_11963);
nor U12200 (N_12200,N_11804,N_11909);
or U12201 (N_12201,N_11849,N_11777);
or U12202 (N_12202,N_11865,N_11982);
nor U12203 (N_12203,N_11799,N_11805);
or U12204 (N_12204,N_11969,N_11968);
nand U12205 (N_12205,N_11800,N_11848);
and U12206 (N_12206,N_11783,N_11893);
nor U12207 (N_12207,N_11781,N_11773);
nor U12208 (N_12208,N_11831,N_11755);
nor U12209 (N_12209,N_11892,N_11991);
or U12210 (N_12210,N_11865,N_11974);
nor U12211 (N_12211,N_11793,N_11822);
xnor U12212 (N_12212,N_11938,N_11942);
nor U12213 (N_12213,N_11907,N_11853);
or U12214 (N_12214,N_11839,N_11793);
nand U12215 (N_12215,N_11977,N_11899);
nor U12216 (N_12216,N_11876,N_11897);
and U12217 (N_12217,N_11902,N_11941);
xor U12218 (N_12218,N_11811,N_11915);
xor U12219 (N_12219,N_11964,N_11767);
xnor U12220 (N_12220,N_11833,N_11930);
nor U12221 (N_12221,N_11965,N_11880);
or U12222 (N_12222,N_11797,N_11892);
nand U12223 (N_12223,N_11766,N_11874);
nand U12224 (N_12224,N_11839,N_11954);
nand U12225 (N_12225,N_11780,N_11974);
and U12226 (N_12226,N_11824,N_11872);
nand U12227 (N_12227,N_11954,N_11991);
xnor U12228 (N_12228,N_11902,N_11930);
and U12229 (N_12229,N_11751,N_11757);
nand U12230 (N_12230,N_11943,N_11816);
and U12231 (N_12231,N_11878,N_11799);
xnor U12232 (N_12232,N_11943,N_11920);
or U12233 (N_12233,N_11926,N_11895);
nor U12234 (N_12234,N_11821,N_11903);
and U12235 (N_12235,N_11783,N_11821);
xnor U12236 (N_12236,N_11968,N_11874);
nor U12237 (N_12237,N_11775,N_11757);
xnor U12238 (N_12238,N_11944,N_11821);
nand U12239 (N_12239,N_11986,N_11844);
nand U12240 (N_12240,N_11863,N_11979);
nand U12241 (N_12241,N_11871,N_11930);
or U12242 (N_12242,N_11829,N_11931);
nor U12243 (N_12243,N_11814,N_11985);
xor U12244 (N_12244,N_11843,N_11760);
xnor U12245 (N_12245,N_11927,N_11755);
or U12246 (N_12246,N_11837,N_11960);
nand U12247 (N_12247,N_11803,N_11938);
or U12248 (N_12248,N_11750,N_11773);
or U12249 (N_12249,N_11877,N_11871);
xor U12250 (N_12250,N_12235,N_12196);
xnor U12251 (N_12251,N_12065,N_12024);
nand U12252 (N_12252,N_12009,N_12231);
or U12253 (N_12253,N_12031,N_12090);
nand U12254 (N_12254,N_12081,N_12193);
nand U12255 (N_12255,N_12216,N_12027);
nor U12256 (N_12256,N_12074,N_12228);
nor U12257 (N_12257,N_12067,N_12079);
and U12258 (N_12258,N_12038,N_12162);
xor U12259 (N_12259,N_12029,N_12134);
nand U12260 (N_12260,N_12171,N_12239);
and U12261 (N_12261,N_12095,N_12033);
xor U12262 (N_12262,N_12108,N_12155);
xor U12263 (N_12263,N_12021,N_12203);
nor U12264 (N_12264,N_12217,N_12148);
nor U12265 (N_12265,N_12016,N_12036);
nor U12266 (N_12266,N_12220,N_12163);
xor U12267 (N_12267,N_12040,N_12156);
xor U12268 (N_12268,N_12169,N_12245);
nand U12269 (N_12269,N_12146,N_12057);
nor U12270 (N_12270,N_12056,N_12145);
nor U12271 (N_12271,N_12041,N_12017);
and U12272 (N_12272,N_12130,N_12136);
or U12273 (N_12273,N_12082,N_12048);
nor U12274 (N_12274,N_12118,N_12075);
or U12275 (N_12275,N_12208,N_12055);
xnor U12276 (N_12276,N_12240,N_12174);
nand U12277 (N_12277,N_12104,N_12100);
xor U12278 (N_12278,N_12177,N_12015);
or U12279 (N_12279,N_12218,N_12018);
nor U12280 (N_12280,N_12210,N_12013);
and U12281 (N_12281,N_12232,N_12141);
nand U12282 (N_12282,N_12023,N_12089);
nor U12283 (N_12283,N_12105,N_12238);
and U12284 (N_12284,N_12010,N_12147);
or U12285 (N_12285,N_12204,N_12135);
nor U12286 (N_12286,N_12049,N_12211);
xnor U12287 (N_12287,N_12236,N_12194);
nand U12288 (N_12288,N_12006,N_12237);
and U12289 (N_12289,N_12022,N_12094);
nor U12290 (N_12290,N_12077,N_12150);
xnor U12291 (N_12291,N_12205,N_12227);
nor U12292 (N_12292,N_12019,N_12172);
nor U12293 (N_12293,N_12122,N_12078);
nor U12294 (N_12294,N_12054,N_12092);
nand U12295 (N_12295,N_12069,N_12059);
xnor U12296 (N_12296,N_12102,N_12087);
nand U12297 (N_12297,N_12061,N_12140);
nand U12298 (N_12298,N_12188,N_12226);
xor U12299 (N_12299,N_12243,N_12192);
xnor U12300 (N_12300,N_12000,N_12215);
or U12301 (N_12301,N_12199,N_12198);
or U12302 (N_12302,N_12225,N_12179);
nand U12303 (N_12303,N_12143,N_12175);
or U12304 (N_12304,N_12173,N_12233);
xor U12305 (N_12305,N_12214,N_12070);
nor U12306 (N_12306,N_12244,N_12088);
and U12307 (N_12307,N_12119,N_12039);
or U12308 (N_12308,N_12044,N_12161);
nor U12309 (N_12309,N_12131,N_12114);
and U12310 (N_12310,N_12042,N_12099);
or U12311 (N_12311,N_12197,N_12116);
and U12312 (N_12312,N_12123,N_12221);
nor U12313 (N_12313,N_12003,N_12124);
nand U12314 (N_12314,N_12160,N_12157);
nor U12315 (N_12315,N_12219,N_12242);
and U12316 (N_12316,N_12012,N_12007);
nand U12317 (N_12317,N_12005,N_12183);
nand U12318 (N_12318,N_12037,N_12170);
xor U12319 (N_12319,N_12206,N_12190);
and U12320 (N_12320,N_12084,N_12248);
xnor U12321 (N_12321,N_12045,N_12052);
xnor U12322 (N_12322,N_12106,N_12154);
xor U12323 (N_12323,N_12066,N_12034);
nor U12324 (N_12324,N_12050,N_12098);
xnor U12325 (N_12325,N_12132,N_12185);
xor U12326 (N_12326,N_12129,N_12230);
nor U12327 (N_12327,N_12166,N_12249);
nand U12328 (N_12328,N_12062,N_12068);
and U12329 (N_12329,N_12229,N_12223);
and U12330 (N_12330,N_12101,N_12241);
nand U12331 (N_12331,N_12153,N_12091);
nand U12332 (N_12332,N_12178,N_12144);
and U12333 (N_12333,N_12085,N_12133);
and U12334 (N_12334,N_12107,N_12246);
and U12335 (N_12335,N_12152,N_12060);
xnor U12336 (N_12336,N_12222,N_12064);
xnor U12337 (N_12337,N_12109,N_12121);
nand U12338 (N_12338,N_12234,N_12182);
xnor U12339 (N_12339,N_12212,N_12167);
and U12340 (N_12340,N_12195,N_12072);
and U12341 (N_12341,N_12247,N_12159);
xor U12342 (N_12342,N_12202,N_12032);
or U12343 (N_12343,N_12014,N_12142);
or U12344 (N_12344,N_12112,N_12011);
and U12345 (N_12345,N_12151,N_12181);
or U12346 (N_12346,N_12149,N_12083);
xor U12347 (N_12347,N_12073,N_12030);
nor U12348 (N_12348,N_12128,N_12168);
or U12349 (N_12349,N_12096,N_12125);
xnor U12350 (N_12350,N_12180,N_12063);
nor U12351 (N_12351,N_12020,N_12127);
and U12352 (N_12352,N_12071,N_12191);
nor U12353 (N_12353,N_12008,N_12086);
or U12354 (N_12354,N_12207,N_12187);
and U12355 (N_12355,N_12184,N_12035);
xnor U12356 (N_12356,N_12103,N_12137);
or U12357 (N_12357,N_12001,N_12164);
nand U12358 (N_12358,N_12126,N_12176);
nand U12359 (N_12359,N_12026,N_12113);
xor U12360 (N_12360,N_12046,N_12201);
and U12361 (N_12361,N_12200,N_12080);
or U12362 (N_12362,N_12058,N_12076);
xnor U12363 (N_12363,N_12004,N_12224);
or U12364 (N_12364,N_12047,N_12028);
nand U12365 (N_12365,N_12139,N_12117);
and U12366 (N_12366,N_12213,N_12158);
and U12367 (N_12367,N_12111,N_12209);
nand U12368 (N_12368,N_12025,N_12120);
and U12369 (N_12369,N_12189,N_12165);
xnor U12370 (N_12370,N_12110,N_12115);
nor U12371 (N_12371,N_12097,N_12051);
or U12372 (N_12372,N_12053,N_12093);
xnor U12373 (N_12373,N_12002,N_12186);
and U12374 (N_12374,N_12138,N_12043);
and U12375 (N_12375,N_12015,N_12007);
and U12376 (N_12376,N_12175,N_12159);
nor U12377 (N_12377,N_12108,N_12240);
nand U12378 (N_12378,N_12129,N_12084);
and U12379 (N_12379,N_12143,N_12156);
xnor U12380 (N_12380,N_12140,N_12180);
nand U12381 (N_12381,N_12232,N_12249);
nand U12382 (N_12382,N_12131,N_12089);
xnor U12383 (N_12383,N_12062,N_12109);
xnor U12384 (N_12384,N_12057,N_12204);
nand U12385 (N_12385,N_12042,N_12181);
or U12386 (N_12386,N_12063,N_12224);
nand U12387 (N_12387,N_12205,N_12073);
nor U12388 (N_12388,N_12235,N_12062);
nand U12389 (N_12389,N_12180,N_12179);
or U12390 (N_12390,N_12045,N_12081);
or U12391 (N_12391,N_12201,N_12008);
and U12392 (N_12392,N_12038,N_12055);
xor U12393 (N_12393,N_12066,N_12221);
nor U12394 (N_12394,N_12011,N_12249);
or U12395 (N_12395,N_12207,N_12006);
nand U12396 (N_12396,N_12220,N_12078);
nor U12397 (N_12397,N_12154,N_12182);
nor U12398 (N_12398,N_12137,N_12246);
nor U12399 (N_12399,N_12221,N_12183);
nor U12400 (N_12400,N_12013,N_12238);
nand U12401 (N_12401,N_12000,N_12126);
and U12402 (N_12402,N_12190,N_12082);
xnor U12403 (N_12403,N_12023,N_12170);
nand U12404 (N_12404,N_12104,N_12054);
or U12405 (N_12405,N_12157,N_12174);
and U12406 (N_12406,N_12047,N_12039);
nor U12407 (N_12407,N_12171,N_12117);
nand U12408 (N_12408,N_12148,N_12143);
nor U12409 (N_12409,N_12236,N_12168);
nand U12410 (N_12410,N_12214,N_12115);
and U12411 (N_12411,N_12143,N_12067);
and U12412 (N_12412,N_12078,N_12051);
nand U12413 (N_12413,N_12074,N_12163);
nand U12414 (N_12414,N_12119,N_12139);
and U12415 (N_12415,N_12240,N_12159);
nand U12416 (N_12416,N_12087,N_12226);
nand U12417 (N_12417,N_12193,N_12198);
nand U12418 (N_12418,N_12082,N_12225);
nor U12419 (N_12419,N_12170,N_12117);
nand U12420 (N_12420,N_12006,N_12135);
nor U12421 (N_12421,N_12117,N_12227);
and U12422 (N_12422,N_12224,N_12156);
or U12423 (N_12423,N_12248,N_12187);
and U12424 (N_12424,N_12107,N_12174);
or U12425 (N_12425,N_12173,N_12134);
nand U12426 (N_12426,N_12156,N_12046);
or U12427 (N_12427,N_12210,N_12127);
and U12428 (N_12428,N_12100,N_12022);
or U12429 (N_12429,N_12064,N_12005);
xor U12430 (N_12430,N_12146,N_12237);
nand U12431 (N_12431,N_12026,N_12185);
and U12432 (N_12432,N_12151,N_12220);
xnor U12433 (N_12433,N_12078,N_12170);
nor U12434 (N_12434,N_12152,N_12131);
xor U12435 (N_12435,N_12112,N_12042);
nand U12436 (N_12436,N_12107,N_12190);
and U12437 (N_12437,N_12217,N_12043);
nand U12438 (N_12438,N_12188,N_12221);
nor U12439 (N_12439,N_12214,N_12029);
xor U12440 (N_12440,N_12079,N_12024);
nor U12441 (N_12441,N_12176,N_12062);
xnor U12442 (N_12442,N_12214,N_12232);
xor U12443 (N_12443,N_12219,N_12129);
xor U12444 (N_12444,N_12204,N_12155);
or U12445 (N_12445,N_12034,N_12014);
nand U12446 (N_12446,N_12123,N_12085);
or U12447 (N_12447,N_12038,N_12093);
nor U12448 (N_12448,N_12229,N_12146);
xor U12449 (N_12449,N_12191,N_12244);
and U12450 (N_12450,N_12118,N_12119);
nand U12451 (N_12451,N_12003,N_12092);
nand U12452 (N_12452,N_12123,N_12139);
or U12453 (N_12453,N_12149,N_12225);
and U12454 (N_12454,N_12003,N_12014);
nor U12455 (N_12455,N_12007,N_12063);
or U12456 (N_12456,N_12173,N_12234);
or U12457 (N_12457,N_12163,N_12028);
or U12458 (N_12458,N_12224,N_12207);
or U12459 (N_12459,N_12192,N_12036);
nand U12460 (N_12460,N_12063,N_12010);
nor U12461 (N_12461,N_12066,N_12026);
and U12462 (N_12462,N_12246,N_12196);
or U12463 (N_12463,N_12190,N_12058);
and U12464 (N_12464,N_12056,N_12043);
nor U12465 (N_12465,N_12048,N_12006);
or U12466 (N_12466,N_12030,N_12096);
xor U12467 (N_12467,N_12170,N_12208);
and U12468 (N_12468,N_12100,N_12079);
or U12469 (N_12469,N_12074,N_12219);
and U12470 (N_12470,N_12198,N_12109);
nand U12471 (N_12471,N_12092,N_12175);
xnor U12472 (N_12472,N_12243,N_12060);
nand U12473 (N_12473,N_12147,N_12210);
xnor U12474 (N_12474,N_12213,N_12070);
or U12475 (N_12475,N_12164,N_12018);
nand U12476 (N_12476,N_12040,N_12101);
nor U12477 (N_12477,N_12183,N_12238);
nand U12478 (N_12478,N_12110,N_12014);
or U12479 (N_12479,N_12178,N_12061);
and U12480 (N_12480,N_12194,N_12047);
and U12481 (N_12481,N_12083,N_12164);
or U12482 (N_12482,N_12006,N_12177);
or U12483 (N_12483,N_12217,N_12121);
nand U12484 (N_12484,N_12214,N_12030);
nand U12485 (N_12485,N_12214,N_12195);
nor U12486 (N_12486,N_12011,N_12184);
and U12487 (N_12487,N_12018,N_12026);
xnor U12488 (N_12488,N_12141,N_12166);
or U12489 (N_12489,N_12040,N_12064);
or U12490 (N_12490,N_12015,N_12208);
and U12491 (N_12491,N_12196,N_12054);
and U12492 (N_12492,N_12212,N_12031);
or U12493 (N_12493,N_12027,N_12191);
nor U12494 (N_12494,N_12106,N_12079);
nand U12495 (N_12495,N_12081,N_12058);
xnor U12496 (N_12496,N_12197,N_12141);
or U12497 (N_12497,N_12153,N_12188);
or U12498 (N_12498,N_12059,N_12165);
and U12499 (N_12499,N_12178,N_12072);
xor U12500 (N_12500,N_12317,N_12292);
nor U12501 (N_12501,N_12495,N_12293);
nand U12502 (N_12502,N_12482,N_12330);
and U12503 (N_12503,N_12463,N_12355);
or U12504 (N_12504,N_12371,N_12256);
nand U12505 (N_12505,N_12489,N_12276);
nand U12506 (N_12506,N_12316,N_12373);
or U12507 (N_12507,N_12344,N_12496);
and U12508 (N_12508,N_12454,N_12382);
xnor U12509 (N_12509,N_12451,N_12265);
nand U12510 (N_12510,N_12263,N_12443);
nor U12511 (N_12511,N_12481,N_12499);
nand U12512 (N_12512,N_12333,N_12427);
and U12513 (N_12513,N_12356,N_12397);
nand U12514 (N_12514,N_12465,N_12250);
nor U12515 (N_12515,N_12322,N_12341);
xnor U12516 (N_12516,N_12484,N_12448);
or U12517 (N_12517,N_12343,N_12415);
nor U12518 (N_12518,N_12264,N_12439);
or U12519 (N_12519,N_12404,N_12392);
nand U12520 (N_12520,N_12393,N_12367);
or U12521 (N_12521,N_12257,N_12444);
or U12522 (N_12522,N_12452,N_12462);
nand U12523 (N_12523,N_12432,N_12424);
or U12524 (N_12524,N_12268,N_12476);
and U12525 (N_12525,N_12417,N_12403);
or U12526 (N_12526,N_12431,N_12251);
nor U12527 (N_12527,N_12430,N_12421);
xnor U12528 (N_12528,N_12376,N_12492);
nor U12529 (N_12529,N_12416,N_12253);
and U12530 (N_12530,N_12347,N_12336);
nor U12531 (N_12531,N_12362,N_12273);
nor U12532 (N_12532,N_12413,N_12487);
nand U12533 (N_12533,N_12386,N_12419);
and U12534 (N_12534,N_12391,N_12426);
nor U12535 (N_12535,N_12304,N_12456);
nor U12536 (N_12536,N_12445,N_12428);
or U12537 (N_12537,N_12475,N_12311);
xnor U12538 (N_12538,N_12387,N_12346);
and U12539 (N_12539,N_12485,N_12446);
xor U12540 (N_12540,N_12457,N_12478);
or U12541 (N_12541,N_12267,N_12433);
and U12542 (N_12542,N_12480,N_12271);
nand U12543 (N_12543,N_12252,N_12472);
nor U12544 (N_12544,N_12493,N_12450);
nand U12545 (N_12545,N_12272,N_12479);
nand U12546 (N_12546,N_12280,N_12477);
nor U12547 (N_12547,N_12339,N_12383);
and U12548 (N_12548,N_12269,N_12498);
and U12549 (N_12549,N_12320,N_12306);
or U12550 (N_12550,N_12464,N_12337);
nor U12551 (N_12551,N_12254,N_12411);
or U12552 (N_12552,N_12281,N_12434);
or U12553 (N_12553,N_12328,N_12258);
nand U12554 (N_12554,N_12379,N_12321);
nor U12555 (N_12555,N_12262,N_12349);
or U12556 (N_12556,N_12318,N_12312);
or U12557 (N_12557,N_12385,N_12301);
nand U12558 (N_12558,N_12358,N_12297);
and U12559 (N_12559,N_12340,N_12368);
or U12560 (N_12560,N_12359,N_12405);
nor U12561 (N_12561,N_12284,N_12327);
and U12562 (N_12562,N_12494,N_12388);
nor U12563 (N_12563,N_12378,N_12410);
and U12564 (N_12564,N_12389,N_12412);
or U12565 (N_12565,N_12422,N_12275);
nand U12566 (N_12566,N_12375,N_12414);
and U12567 (N_12567,N_12338,N_12308);
nand U12568 (N_12568,N_12420,N_12278);
xnor U12569 (N_12569,N_12325,N_12270);
or U12570 (N_12570,N_12300,N_12408);
or U12571 (N_12571,N_12466,N_12396);
and U12572 (N_12572,N_12390,N_12474);
or U12573 (N_12573,N_12294,N_12429);
nand U12574 (N_12574,N_12418,N_12345);
and U12575 (N_12575,N_12365,N_12470);
nor U12576 (N_12576,N_12295,N_12289);
and U12577 (N_12577,N_12319,N_12438);
nor U12578 (N_12578,N_12335,N_12352);
nor U12579 (N_12579,N_12437,N_12395);
nor U12580 (N_12580,N_12360,N_12458);
and U12581 (N_12581,N_12286,N_12324);
or U12582 (N_12582,N_12307,N_12398);
nand U12583 (N_12583,N_12285,N_12302);
nand U12584 (N_12584,N_12473,N_12442);
nor U12585 (N_12585,N_12488,N_12449);
xnor U12586 (N_12586,N_12453,N_12374);
nor U12587 (N_12587,N_12303,N_12313);
xnor U12588 (N_12588,N_12279,N_12423);
nand U12589 (N_12589,N_12288,N_12326);
and U12590 (N_12590,N_12441,N_12334);
xnor U12591 (N_12591,N_12266,N_12353);
and U12592 (N_12592,N_12329,N_12315);
nor U12593 (N_12593,N_12467,N_12361);
nand U12594 (N_12594,N_12497,N_12400);
nor U12595 (N_12595,N_12261,N_12384);
xnor U12596 (N_12596,N_12287,N_12440);
and U12597 (N_12597,N_12461,N_12364);
nand U12598 (N_12598,N_12455,N_12283);
nor U12599 (N_12599,N_12351,N_12259);
or U12600 (N_12600,N_12491,N_12490);
and U12601 (N_12601,N_12486,N_12331);
nand U12602 (N_12602,N_12372,N_12309);
or U12603 (N_12603,N_12291,N_12332);
and U12604 (N_12604,N_12296,N_12277);
or U12605 (N_12605,N_12305,N_12299);
xor U12606 (N_12606,N_12468,N_12402);
or U12607 (N_12607,N_12357,N_12290);
or U12608 (N_12608,N_12435,N_12342);
nor U12609 (N_12609,N_12366,N_12377);
xor U12610 (N_12610,N_12363,N_12436);
and U12611 (N_12611,N_12406,N_12483);
or U12612 (N_12612,N_12310,N_12425);
nor U12613 (N_12613,N_12381,N_12399);
nand U12614 (N_12614,N_12369,N_12447);
xor U12615 (N_12615,N_12471,N_12460);
or U12616 (N_12616,N_12323,N_12298);
or U12617 (N_12617,N_12394,N_12314);
nor U12618 (N_12618,N_12380,N_12401);
and U12619 (N_12619,N_12260,N_12370);
xnor U12620 (N_12620,N_12274,N_12354);
nor U12621 (N_12621,N_12459,N_12282);
and U12622 (N_12622,N_12348,N_12255);
or U12623 (N_12623,N_12407,N_12350);
nand U12624 (N_12624,N_12469,N_12409);
nor U12625 (N_12625,N_12304,N_12268);
or U12626 (N_12626,N_12438,N_12327);
or U12627 (N_12627,N_12365,N_12366);
and U12628 (N_12628,N_12484,N_12305);
nor U12629 (N_12629,N_12276,N_12314);
nand U12630 (N_12630,N_12421,N_12499);
nand U12631 (N_12631,N_12457,N_12276);
xnor U12632 (N_12632,N_12251,N_12493);
or U12633 (N_12633,N_12360,N_12337);
nor U12634 (N_12634,N_12475,N_12466);
or U12635 (N_12635,N_12321,N_12325);
nand U12636 (N_12636,N_12393,N_12466);
xnor U12637 (N_12637,N_12251,N_12328);
nor U12638 (N_12638,N_12320,N_12413);
or U12639 (N_12639,N_12490,N_12308);
nor U12640 (N_12640,N_12477,N_12258);
nand U12641 (N_12641,N_12442,N_12419);
or U12642 (N_12642,N_12301,N_12282);
nand U12643 (N_12643,N_12382,N_12431);
nor U12644 (N_12644,N_12400,N_12448);
nor U12645 (N_12645,N_12349,N_12376);
nand U12646 (N_12646,N_12461,N_12299);
nand U12647 (N_12647,N_12395,N_12270);
xor U12648 (N_12648,N_12296,N_12468);
xnor U12649 (N_12649,N_12303,N_12289);
xor U12650 (N_12650,N_12314,N_12382);
nand U12651 (N_12651,N_12413,N_12319);
xor U12652 (N_12652,N_12420,N_12389);
and U12653 (N_12653,N_12260,N_12407);
or U12654 (N_12654,N_12291,N_12289);
xnor U12655 (N_12655,N_12401,N_12474);
nor U12656 (N_12656,N_12344,N_12340);
or U12657 (N_12657,N_12450,N_12485);
nand U12658 (N_12658,N_12262,N_12400);
and U12659 (N_12659,N_12448,N_12410);
nand U12660 (N_12660,N_12498,N_12496);
nor U12661 (N_12661,N_12409,N_12484);
nor U12662 (N_12662,N_12475,N_12452);
or U12663 (N_12663,N_12404,N_12289);
and U12664 (N_12664,N_12280,N_12387);
nand U12665 (N_12665,N_12302,N_12457);
xnor U12666 (N_12666,N_12267,N_12347);
nand U12667 (N_12667,N_12452,N_12371);
and U12668 (N_12668,N_12341,N_12277);
xor U12669 (N_12669,N_12438,N_12338);
and U12670 (N_12670,N_12337,N_12387);
and U12671 (N_12671,N_12473,N_12399);
nand U12672 (N_12672,N_12362,N_12398);
nor U12673 (N_12673,N_12444,N_12445);
nor U12674 (N_12674,N_12360,N_12397);
nor U12675 (N_12675,N_12284,N_12263);
nand U12676 (N_12676,N_12252,N_12492);
nor U12677 (N_12677,N_12377,N_12487);
or U12678 (N_12678,N_12485,N_12319);
and U12679 (N_12679,N_12327,N_12463);
or U12680 (N_12680,N_12352,N_12331);
nand U12681 (N_12681,N_12464,N_12473);
nand U12682 (N_12682,N_12459,N_12455);
nand U12683 (N_12683,N_12482,N_12265);
and U12684 (N_12684,N_12316,N_12253);
xnor U12685 (N_12685,N_12458,N_12487);
and U12686 (N_12686,N_12453,N_12427);
or U12687 (N_12687,N_12473,N_12314);
nor U12688 (N_12688,N_12371,N_12270);
and U12689 (N_12689,N_12404,N_12268);
nand U12690 (N_12690,N_12436,N_12361);
and U12691 (N_12691,N_12439,N_12481);
nor U12692 (N_12692,N_12283,N_12343);
and U12693 (N_12693,N_12258,N_12476);
xnor U12694 (N_12694,N_12477,N_12291);
xnor U12695 (N_12695,N_12465,N_12370);
nand U12696 (N_12696,N_12383,N_12359);
nor U12697 (N_12697,N_12355,N_12318);
xor U12698 (N_12698,N_12325,N_12474);
nor U12699 (N_12699,N_12380,N_12258);
and U12700 (N_12700,N_12386,N_12344);
or U12701 (N_12701,N_12344,N_12366);
or U12702 (N_12702,N_12315,N_12355);
xnor U12703 (N_12703,N_12442,N_12439);
and U12704 (N_12704,N_12377,N_12337);
and U12705 (N_12705,N_12471,N_12258);
xor U12706 (N_12706,N_12300,N_12314);
nand U12707 (N_12707,N_12318,N_12440);
nor U12708 (N_12708,N_12393,N_12488);
or U12709 (N_12709,N_12488,N_12339);
xnor U12710 (N_12710,N_12250,N_12282);
xor U12711 (N_12711,N_12302,N_12269);
nand U12712 (N_12712,N_12426,N_12250);
nand U12713 (N_12713,N_12280,N_12258);
nand U12714 (N_12714,N_12275,N_12311);
xnor U12715 (N_12715,N_12348,N_12284);
or U12716 (N_12716,N_12347,N_12334);
nor U12717 (N_12717,N_12394,N_12287);
nor U12718 (N_12718,N_12444,N_12301);
nor U12719 (N_12719,N_12395,N_12447);
or U12720 (N_12720,N_12307,N_12470);
nand U12721 (N_12721,N_12308,N_12468);
xor U12722 (N_12722,N_12373,N_12369);
nand U12723 (N_12723,N_12300,N_12499);
and U12724 (N_12724,N_12380,N_12444);
xnor U12725 (N_12725,N_12250,N_12354);
or U12726 (N_12726,N_12355,N_12330);
nand U12727 (N_12727,N_12467,N_12290);
nand U12728 (N_12728,N_12485,N_12407);
and U12729 (N_12729,N_12488,N_12304);
xor U12730 (N_12730,N_12409,N_12274);
nand U12731 (N_12731,N_12481,N_12408);
nor U12732 (N_12732,N_12382,N_12273);
or U12733 (N_12733,N_12367,N_12360);
nor U12734 (N_12734,N_12284,N_12454);
and U12735 (N_12735,N_12484,N_12328);
and U12736 (N_12736,N_12488,N_12272);
or U12737 (N_12737,N_12256,N_12411);
and U12738 (N_12738,N_12264,N_12355);
xnor U12739 (N_12739,N_12278,N_12475);
nand U12740 (N_12740,N_12442,N_12418);
or U12741 (N_12741,N_12344,N_12404);
and U12742 (N_12742,N_12299,N_12451);
nor U12743 (N_12743,N_12303,N_12288);
nand U12744 (N_12744,N_12303,N_12438);
xor U12745 (N_12745,N_12298,N_12292);
nor U12746 (N_12746,N_12399,N_12405);
xnor U12747 (N_12747,N_12449,N_12252);
xnor U12748 (N_12748,N_12404,N_12372);
and U12749 (N_12749,N_12289,N_12388);
and U12750 (N_12750,N_12505,N_12631);
or U12751 (N_12751,N_12602,N_12665);
and U12752 (N_12752,N_12630,N_12674);
nor U12753 (N_12753,N_12620,N_12531);
and U12754 (N_12754,N_12653,N_12571);
xor U12755 (N_12755,N_12676,N_12650);
or U12756 (N_12756,N_12701,N_12550);
nor U12757 (N_12757,N_12512,N_12513);
nand U12758 (N_12758,N_12647,N_12588);
xor U12759 (N_12759,N_12524,N_12523);
xnor U12760 (N_12760,N_12592,N_12641);
xor U12761 (N_12761,N_12656,N_12697);
nand U12762 (N_12762,N_12616,N_12646);
and U12763 (N_12763,N_12560,N_12586);
or U12764 (N_12764,N_12555,N_12577);
or U12765 (N_12765,N_12510,N_12667);
nand U12766 (N_12766,N_12575,N_12734);
and U12767 (N_12767,N_12728,N_12726);
or U12768 (N_12768,N_12596,N_12746);
nand U12769 (N_12769,N_12635,N_12719);
and U12770 (N_12770,N_12669,N_12654);
nand U12771 (N_12771,N_12511,N_12649);
or U12772 (N_12772,N_12670,N_12733);
nor U12773 (N_12773,N_12548,N_12703);
and U12774 (N_12774,N_12578,N_12526);
nor U12775 (N_12775,N_12593,N_12527);
nand U12776 (N_12776,N_12711,N_12668);
or U12777 (N_12777,N_12639,N_12680);
xor U12778 (N_12778,N_12543,N_12706);
and U12779 (N_12779,N_12544,N_12632);
and U12780 (N_12780,N_12606,N_12539);
nand U12781 (N_12781,N_12520,N_12557);
xnor U12782 (N_12782,N_12735,N_12545);
nor U12783 (N_12783,N_12679,N_12612);
nand U12784 (N_12784,N_12643,N_12638);
nor U12785 (N_12785,N_12694,N_12747);
xor U12786 (N_12786,N_12525,N_12690);
nor U12787 (N_12787,N_12625,N_12721);
and U12788 (N_12788,N_12724,N_12615);
and U12789 (N_12789,N_12744,N_12566);
and U12790 (N_12790,N_12698,N_12671);
nand U12791 (N_12791,N_12700,N_12730);
nand U12792 (N_12792,N_12732,N_12637);
xor U12793 (N_12793,N_12619,N_12651);
nor U12794 (N_12794,N_12590,N_12583);
or U12795 (N_12795,N_12572,N_12584);
xnor U12796 (N_12796,N_12514,N_12658);
nor U12797 (N_12797,N_12628,N_12687);
nor U12798 (N_12798,N_12556,N_12562);
and U12799 (N_12799,N_12740,N_12518);
nand U12800 (N_12800,N_12501,N_12585);
or U12801 (N_12801,N_12559,N_12729);
nand U12802 (N_12802,N_12739,N_12691);
xnor U12803 (N_12803,N_12604,N_12558);
nor U12804 (N_12804,N_12693,N_12568);
xnor U12805 (N_12805,N_12538,N_12554);
and U12806 (N_12806,N_12672,N_12516);
xnor U12807 (N_12807,N_12683,N_12608);
xor U12808 (N_12808,N_12540,N_12533);
or U12809 (N_12809,N_12741,N_12657);
nand U12810 (N_12810,N_12574,N_12532);
and U12811 (N_12811,N_12645,N_12552);
nor U12812 (N_12812,N_12599,N_12507);
nand U12813 (N_12813,N_12521,N_12673);
nand U12814 (N_12814,N_12517,N_12573);
or U12815 (N_12815,N_12648,N_12547);
nor U12816 (N_12816,N_12714,N_12537);
xnor U12817 (N_12817,N_12576,N_12666);
xor U12818 (N_12818,N_12522,N_12508);
nand U12819 (N_12819,N_12626,N_12536);
xor U12820 (N_12820,N_12696,N_12553);
nand U12821 (N_12821,N_12662,N_12587);
or U12822 (N_12822,N_12580,N_12504);
and U12823 (N_12823,N_12634,N_12542);
nor U12824 (N_12824,N_12689,N_12709);
or U12825 (N_12825,N_12529,N_12713);
nor U12826 (N_12826,N_12624,N_12660);
xnor U12827 (N_12827,N_12598,N_12715);
and U12828 (N_12828,N_12748,N_12737);
or U12829 (N_12829,N_12551,N_12712);
or U12830 (N_12830,N_12738,N_12717);
xnor U12831 (N_12831,N_12629,N_12609);
nand U12832 (N_12832,N_12500,N_12611);
and U12833 (N_12833,N_12603,N_12582);
nor U12834 (N_12834,N_12565,N_12731);
xor U12835 (N_12835,N_12534,N_12685);
and U12836 (N_12836,N_12564,N_12704);
or U12837 (N_12837,N_12659,N_12675);
and U12838 (N_12838,N_12503,N_12640);
and U12839 (N_12839,N_12636,N_12610);
or U12840 (N_12840,N_12710,N_12614);
and U12841 (N_12841,N_12519,N_12743);
nor U12842 (N_12842,N_12736,N_12607);
nor U12843 (N_12843,N_12699,N_12535);
xnor U12844 (N_12844,N_12718,N_12644);
or U12845 (N_12845,N_12627,N_12589);
and U12846 (N_12846,N_12652,N_12663);
or U12847 (N_12847,N_12681,N_12561);
nor U12848 (N_12848,N_12684,N_12502);
or U12849 (N_12849,N_12506,N_12722);
nor U12850 (N_12850,N_12549,N_12600);
nand U12851 (N_12851,N_12633,N_12581);
or U12852 (N_12852,N_12530,N_12655);
nor U12853 (N_12853,N_12678,N_12528);
or U12854 (N_12854,N_12591,N_12594);
nor U12855 (N_12855,N_12579,N_12707);
xor U12856 (N_12856,N_12563,N_12688);
xor U12857 (N_12857,N_12617,N_12677);
and U12858 (N_12858,N_12570,N_12569);
nor U12859 (N_12859,N_12745,N_12716);
nor U12860 (N_12860,N_12515,N_12686);
xnor U12861 (N_12861,N_12695,N_12567);
nor U12862 (N_12862,N_12702,N_12705);
or U12863 (N_12863,N_12692,N_12597);
and U12864 (N_12864,N_12623,N_12618);
nor U12865 (N_12865,N_12601,N_12708);
nor U12866 (N_12866,N_12661,N_12682);
xnor U12867 (N_12867,N_12613,N_12605);
or U12868 (N_12868,N_12727,N_12749);
and U12869 (N_12869,N_12622,N_12621);
or U12870 (N_12870,N_12725,N_12595);
and U12871 (N_12871,N_12541,N_12720);
nand U12872 (N_12872,N_12509,N_12546);
or U12873 (N_12873,N_12642,N_12742);
nand U12874 (N_12874,N_12664,N_12723);
nand U12875 (N_12875,N_12696,N_12637);
nor U12876 (N_12876,N_12632,N_12709);
nand U12877 (N_12877,N_12654,N_12746);
nand U12878 (N_12878,N_12620,N_12714);
nand U12879 (N_12879,N_12715,N_12588);
nand U12880 (N_12880,N_12642,N_12718);
nand U12881 (N_12881,N_12531,N_12617);
and U12882 (N_12882,N_12682,N_12510);
and U12883 (N_12883,N_12591,N_12678);
nor U12884 (N_12884,N_12577,N_12675);
xor U12885 (N_12885,N_12534,N_12732);
and U12886 (N_12886,N_12572,N_12734);
and U12887 (N_12887,N_12656,N_12731);
nor U12888 (N_12888,N_12658,N_12695);
nor U12889 (N_12889,N_12715,N_12656);
nor U12890 (N_12890,N_12642,N_12581);
and U12891 (N_12891,N_12673,N_12577);
xnor U12892 (N_12892,N_12621,N_12569);
nor U12893 (N_12893,N_12589,N_12551);
nor U12894 (N_12894,N_12504,N_12596);
and U12895 (N_12895,N_12688,N_12647);
xor U12896 (N_12896,N_12662,N_12676);
xor U12897 (N_12897,N_12660,N_12717);
xnor U12898 (N_12898,N_12746,N_12695);
xor U12899 (N_12899,N_12678,N_12699);
nor U12900 (N_12900,N_12502,N_12583);
and U12901 (N_12901,N_12637,N_12734);
or U12902 (N_12902,N_12529,N_12716);
and U12903 (N_12903,N_12587,N_12671);
nor U12904 (N_12904,N_12642,N_12529);
and U12905 (N_12905,N_12660,N_12652);
nor U12906 (N_12906,N_12564,N_12501);
nor U12907 (N_12907,N_12664,N_12670);
nor U12908 (N_12908,N_12637,N_12643);
or U12909 (N_12909,N_12705,N_12657);
nand U12910 (N_12910,N_12518,N_12623);
xor U12911 (N_12911,N_12681,N_12553);
or U12912 (N_12912,N_12503,N_12563);
nand U12913 (N_12913,N_12678,N_12600);
nand U12914 (N_12914,N_12575,N_12646);
or U12915 (N_12915,N_12570,N_12617);
nand U12916 (N_12916,N_12644,N_12587);
or U12917 (N_12917,N_12607,N_12685);
nand U12918 (N_12918,N_12621,N_12670);
nand U12919 (N_12919,N_12539,N_12637);
nor U12920 (N_12920,N_12639,N_12633);
or U12921 (N_12921,N_12545,N_12631);
nand U12922 (N_12922,N_12621,N_12749);
xor U12923 (N_12923,N_12731,N_12748);
and U12924 (N_12924,N_12505,N_12562);
nand U12925 (N_12925,N_12690,N_12726);
and U12926 (N_12926,N_12641,N_12550);
and U12927 (N_12927,N_12503,N_12731);
xnor U12928 (N_12928,N_12711,N_12739);
nor U12929 (N_12929,N_12664,N_12508);
nor U12930 (N_12930,N_12601,N_12513);
xor U12931 (N_12931,N_12739,N_12736);
nor U12932 (N_12932,N_12697,N_12527);
nand U12933 (N_12933,N_12716,N_12601);
and U12934 (N_12934,N_12642,N_12578);
nand U12935 (N_12935,N_12627,N_12569);
or U12936 (N_12936,N_12699,N_12508);
xnor U12937 (N_12937,N_12668,N_12609);
or U12938 (N_12938,N_12584,N_12552);
or U12939 (N_12939,N_12508,N_12510);
and U12940 (N_12940,N_12621,N_12698);
nor U12941 (N_12941,N_12537,N_12526);
nor U12942 (N_12942,N_12623,N_12611);
and U12943 (N_12943,N_12509,N_12588);
xor U12944 (N_12944,N_12697,N_12551);
nor U12945 (N_12945,N_12636,N_12572);
nand U12946 (N_12946,N_12737,N_12665);
nand U12947 (N_12947,N_12642,N_12569);
and U12948 (N_12948,N_12640,N_12615);
or U12949 (N_12949,N_12707,N_12738);
nor U12950 (N_12950,N_12705,N_12531);
xnor U12951 (N_12951,N_12699,N_12658);
and U12952 (N_12952,N_12610,N_12531);
and U12953 (N_12953,N_12522,N_12516);
nand U12954 (N_12954,N_12516,N_12550);
nand U12955 (N_12955,N_12612,N_12663);
and U12956 (N_12956,N_12592,N_12597);
xnor U12957 (N_12957,N_12723,N_12720);
or U12958 (N_12958,N_12708,N_12697);
or U12959 (N_12959,N_12616,N_12683);
or U12960 (N_12960,N_12685,N_12728);
nor U12961 (N_12961,N_12527,N_12630);
or U12962 (N_12962,N_12712,N_12679);
or U12963 (N_12963,N_12610,N_12717);
nor U12964 (N_12964,N_12670,N_12662);
nor U12965 (N_12965,N_12643,N_12576);
nor U12966 (N_12966,N_12628,N_12594);
nand U12967 (N_12967,N_12648,N_12555);
nand U12968 (N_12968,N_12628,N_12559);
and U12969 (N_12969,N_12741,N_12671);
and U12970 (N_12970,N_12522,N_12600);
xnor U12971 (N_12971,N_12654,N_12562);
xnor U12972 (N_12972,N_12531,N_12595);
or U12973 (N_12973,N_12519,N_12539);
xnor U12974 (N_12974,N_12514,N_12622);
nand U12975 (N_12975,N_12724,N_12535);
or U12976 (N_12976,N_12700,N_12537);
xor U12977 (N_12977,N_12662,N_12627);
xor U12978 (N_12978,N_12657,N_12748);
and U12979 (N_12979,N_12704,N_12707);
or U12980 (N_12980,N_12638,N_12581);
or U12981 (N_12981,N_12703,N_12625);
or U12982 (N_12982,N_12634,N_12670);
nand U12983 (N_12983,N_12626,N_12722);
nor U12984 (N_12984,N_12670,N_12526);
xor U12985 (N_12985,N_12661,N_12579);
or U12986 (N_12986,N_12560,N_12585);
and U12987 (N_12987,N_12693,N_12711);
nand U12988 (N_12988,N_12739,N_12648);
or U12989 (N_12989,N_12587,N_12549);
nor U12990 (N_12990,N_12542,N_12627);
nand U12991 (N_12991,N_12644,N_12570);
nor U12992 (N_12992,N_12636,N_12686);
or U12993 (N_12993,N_12660,N_12627);
nand U12994 (N_12994,N_12611,N_12676);
nand U12995 (N_12995,N_12591,N_12588);
nor U12996 (N_12996,N_12708,N_12607);
nand U12997 (N_12997,N_12739,N_12684);
nor U12998 (N_12998,N_12664,N_12661);
nand U12999 (N_12999,N_12702,N_12577);
and U13000 (N_13000,N_12977,N_12955);
and U13001 (N_13001,N_12906,N_12900);
and U13002 (N_13002,N_12831,N_12953);
nand U13003 (N_13003,N_12808,N_12932);
nor U13004 (N_13004,N_12878,N_12875);
and U13005 (N_13005,N_12752,N_12979);
nor U13006 (N_13006,N_12832,N_12936);
nor U13007 (N_13007,N_12861,N_12973);
or U13008 (N_13008,N_12828,N_12902);
and U13009 (N_13009,N_12893,N_12931);
or U13010 (N_13010,N_12886,N_12938);
nor U13011 (N_13011,N_12794,N_12796);
xnor U13012 (N_13012,N_12857,N_12865);
nor U13013 (N_13013,N_12803,N_12918);
nand U13014 (N_13014,N_12759,N_12869);
or U13015 (N_13015,N_12892,N_12856);
nand U13016 (N_13016,N_12905,N_12975);
or U13017 (N_13017,N_12763,N_12756);
nor U13018 (N_13018,N_12835,N_12995);
xor U13019 (N_13019,N_12921,N_12990);
xnor U13020 (N_13020,N_12840,N_12987);
xor U13021 (N_13021,N_12858,N_12937);
nand U13022 (N_13022,N_12915,N_12964);
and U13023 (N_13023,N_12960,N_12791);
nor U13024 (N_13024,N_12996,N_12778);
nor U13025 (N_13025,N_12765,N_12811);
and U13026 (N_13026,N_12952,N_12820);
or U13027 (N_13027,N_12911,N_12750);
nor U13028 (N_13028,N_12883,N_12967);
nor U13029 (N_13029,N_12926,N_12916);
and U13030 (N_13030,N_12919,N_12786);
and U13031 (N_13031,N_12844,N_12945);
and U13032 (N_13032,N_12942,N_12879);
nand U13033 (N_13033,N_12972,N_12813);
nand U13034 (N_13034,N_12805,N_12806);
nor U13035 (N_13035,N_12874,N_12772);
xnor U13036 (N_13036,N_12885,N_12933);
nor U13037 (N_13037,N_12827,N_12837);
or U13038 (N_13038,N_12862,N_12958);
or U13039 (N_13039,N_12845,N_12941);
xnor U13040 (N_13040,N_12962,N_12764);
nor U13041 (N_13041,N_12826,N_12930);
xnor U13042 (N_13042,N_12887,N_12993);
nor U13043 (N_13043,N_12838,N_12961);
nor U13044 (N_13044,N_12779,N_12771);
nand U13045 (N_13045,N_12984,N_12998);
nand U13046 (N_13046,N_12894,N_12947);
and U13047 (N_13047,N_12818,N_12978);
nor U13048 (N_13048,N_12836,N_12850);
and U13049 (N_13049,N_12903,N_12795);
and U13050 (N_13050,N_12966,N_12888);
xor U13051 (N_13051,N_12971,N_12913);
or U13052 (N_13052,N_12788,N_12959);
and U13053 (N_13053,N_12989,N_12766);
or U13054 (N_13054,N_12957,N_12992);
or U13055 (N_13055,N_12775,N_12991);
nor U13056 (N_13056,N_12822,N_12762);
and U13057 (N_13057,N_12760,N_12800);
and U13058 (N_13058,N_12774,N_12935);
or U13059 (N_13059,N_12924,N_12928);
or U13060 (N_13060,N_12849,N_12792);
nand U13061 (N_13061,N_12914,N_12940);
nand U13062 (N_13062,N_12948,N_12970);
or U13063 (N_13063,N_12753,N_12985);
xnor U13064 (N_13064,N_12876,N_12809);
xnor U13065 (N_13065,N_12891,N_12790);
nand U13066 (N_13066,N_12983,N_12859);
nand U13067 (N_13067,N_12854,N_12882);
xor U13068 (N_13068,N_12758,N_12807);
nand U13069 (N_13069,N_12864,N_12872);
nor U13070 (N_13070,N_12798,N_12890);
xor U13071 (N_13071,N_12954,N_12842);
and U13072 (N_13072,N_12949,N_12968);
nand U13073 (N_13073,N_12870,N_12881);
xnor U13074 (N_13074,N_12823,N_12814);
nand U13075 (N_13075,N_12867,N_12793);
nand U13076 (N_13076,N_12839,N_12929);
or U13077 (N_13077,N_12877,N_12787);
nand U13078 (N_13078,N_12855,N_12899);
nand U13079 (N_13079,N_12785,N_12999);
and U13080 (N_13080,N_12841,N_12920);
or U13081 (N_13081,N_12830,N_12815);
and U13082 (N_13082,N_12851,N_12976);
or U13083 (N_13083,N_12801,N_12767);
and U13084 (N_13084,N_12852,N_12819);
nor U13085 (N_13085,N_12768,N_12755);
or U13086 (N_13086,N_12956,N_12904);
xnor U13087 (N_13087,N_12825,N_12843);
xnor U13088 (N_13088,N_12901,N_12910);
nor U13089 (N_13089,N_12868,N_12799);
nor U13090 (N_13090,N_12950,N_12946);
or U13091 (N_13091,N_12751,N_12997);
and U13092 (N_13092,N_12782,N_12897);
or U13093 (N_13093,N_12980,N_12866);
nand U13094 (N_13094,N_12797,N_12969);
or U13095 (N_13095,N_12777,N_12784);
nand U13096 (N_13096,N_12757,N_12817);
xor U13097 (N_13097,N_12884,N_12847);
or U13098 (N_13098,N_12816,N_12982);
or U13099 (N_13099,N_12812,N_12925);
or U13100 (N_13100,N_12895,N_12922);
nand U13101 (N_13101,N_12908,N_12939);
and U13102 (N_13102,N_12907,N_12802);
xnor U13103 (N_13103,N_12934,N_12853);
or U13104 (N_13104,N_12917,N_12804);
nand U13105 (N_13105,N_12923,N_12986);
and U13106 (N_13106,N_12994,N_12821);
nand U13107 (N_13107,N_12776,N_12829);
or U13108 (N_13108,N_12780,N_12889);
and U13109 (N_13109,N_12773,N_12880);
nand U13110 (N_13110,N_12988,N_12846);
xor U13111 (N_13111,N_12770,N_12896);
nand U13112 (N_13112,N_12944,N_12927);
or U13113 (N_13113,N_12871,N_12963);
nand U13114 (N_13114,N_12943,N_12754);
nand U13115 (N_13115,N_12981,N_12974);
or U13116 (N_13116,N_12912,N_12834);
nand U13117 (N_13117,N_12833,N_12783);
and U13118 (N_13118,N_12789,N_12810);
nor U13119 (N_13119,N_12860,N_12965);
and U13120 (N_13120,N_12863,N_12909);
xnor U13121 (N_13121,N_12824,N_12898);
or U13122 (N_13122,N_12781,N_12873);
nand U13123 (N_13123,N_12761,N_12769);
nor U13124 (N_13124,N_12951,N_12848);
and U13125 (N_13125,N_12981,N_12903);
nor U13126 (N_13126,N_12793,N_12978);
nand U13127 (N_13127,N_12763,N_12884);
nand U13128 (N_13128,N_12772,N_12933);
xnor U13129 (N_13129,N_12988,N_12835);
and U13130 (N_13130,N_12913,N_12881);
and U13131 (N_13131,N_12952,N_12757);
nand U13132 (N_13132,N_12899,N_12782);
nand U13133 (N_13133,N_12873,N_12895);
or U13134 (N_13134,N_12789,N_12845);
xor U13135 (N_13135,N_12766,N_12903);
and U13136 (N_13136,N_12927,N_12788);
nor U13137 (N_13137,N_12773,N_12852);
and U13138 (N_13138,N_12841,N_12930);
xor U13139 (N_13139,N_12761,N_12826);
or U13140 (N_13140,N_12895,N_12991);
nand U13141 (N_13141,N_12815,N_12901);
and U13142 (N_13142,N_12891,N_12830);
nand U13143 (N_13143,N_12926,N_12784);
xor U13144 (N_13144,N_12771,N_12833);
and U13145 (N_13145,N_12863,N_12771);
xor U13146 (N_13146,N_12869,N_12794);
or U13147 (N_13147,N_12982,N_12861);
nand U13148 (N_13148,N_12912,N_12769);
or U13149 (N_13149,N_12979,N_12866);
nor U13150 (N_13150,N_12901,N_12919);
and U13151 (N_13151,N_12847,N_12885);
nand U13152 (N_13152,N_12994,N_12759);
nor U13153 (N_13153,N_12884,N_12906);
or U13154 (N_13154,N_12948,N_12814);
and U13155 (N_13155,N_12876,N_12842);
nor U13156 (N_13156,N_12999,N_12903);
nor U13157 (N_13157,N_12973,N_12899);
or U13158 (N_13158,N_12779,N_12892);
xor U13159 (N_13159,N_12813,N_12850);
nor U13160 (N_13160,N_12837,N_12820);
xnor U13161 (N_13161,N_12831,N_12764);
nand U13162 (N_13162,N_12918,N_12940);
nand U13163 (N_13163,N_12820,N_12769);
or U13164 (N_13164,N_12919,N_12956);
nand U13165 (N_13165,N_12832,N_12829);
or U13166 (N_13166,N_12854,N_12887);
or U13167 (N_13167,N_12866,N_12840);
or U13168 (N_13168,N_12880,N_12943);
nor U13169 (N_13169,N_12980,N_12981);
or U13170 (N_13170,N_12878,N_12827);
or U13171 (N_13171,N_12996,N_12763);
xnor U13172 (N_13172,N_12996,N_12973);
nand U13173 (N_13173,N_12990,N_12836);
nor U13174 (N_13174,N_12888,N_12825);
or U13175 (N_13175,N_12918,N_12956);
nand U13176 (N_13176,N_12855,N_12954);
or U13177 (N_13177,N_12995,N_12794);
or U13178 (N_13178,N_12840,N_12986);
nor U13179 (N_13179,N_12879,N_12895);
nand U13180 (N_13180,N_12902,N_12819);
xnor U13181 (N_13181,N_12824,N_12922);
nand U13182 (N_13182,N_12961,N_12992);
nand U13183 (N_13183,N_12792,N_12911);
xor U13184 (N_13184,N_12936,N_12879);
nand U13185 (N_13185,N_12755,N_12841);
nand U13186 (N_13186,N_12970,N_12872);
nor U13187 (N_13187,N_12771,N_12987);
or U13188 (N_13188,N_12915,N_12956);
nor U13189 (N_13189,N_12907,N_12926);
xnor U13190 (N_13190,N_12954,N_12967);
xnor U13191 (N_13191,N_12980,N_12760);
and U13192 (N_13192,N_12850,N_12881);
or U13193 (N_13193,N_12929,N_12935);
and U13194 (N_13194,N_12788,N_12939);
or U13195 (N_13195,N_12858,N_12807);
nor U13196 (N_13196,N_12778,N_12886);
nor U13197 (N_13197,N_12885,N_12794);
and U13198 (N_13198,N_12886,N_12900);
xnor U13199 (N_13199,N_12994,N_12888);
and U13200 (N_13200,N_12920,N_12940);
nand U13201 (N_13201,N_12880,N_12751);
nor U13202 (N_13202,N_12901,N_12761);
or U13203 (N_13203,N_12992,N_12952);
and U13204 (N_13204,N_12944,N_12903);
or U13205 (N_13205,N_12904,N_12756);
nand U13206 (N_13206,N_12968,N_12770);
xnor U13207 (N_13207,N_12827,N_12925);
and U13208 (N_13208,N_12764,N_12872);
and U13209 (N_13209,N_12770,N_12808);
or U13210 (N_13210,N_12937,N_12876);
nor U13211 (N_13211,N_12928,N_12771);
nand U13212 (N_13212,N_12907,N_12793);
nor U13213 (N_13213,N_12753,N_12920);
or U13214 (N_13214,N_12775,N_12857);
or U13215 (N_13215,N_12896,N_12945);
nand U13216 (N_13216,N_12996,N_12881);
nor U13217 (N_13217,N_12843,N_12972);
and U13218 (N_13218,N_12982,N_12905);
and U13219 (N_13219,N_12813,N_12943);
or U13220 (N_13220,N_12766,N_12809);
nor U13221 (N_13221,N_12855,N_12988);
and U13222 (N_13222,N_12916,N_12973);
nor U13223 (N_13223,N_12783,N_12921);
xnor U13224 (N_13224,N_12881,N_12805);
nand U13225 (N_13225,N_12850,N_12880);
nand U13226 (N_13226,N_12815,N_12982);
and U13227 (N_13227,N_12904,N_12844);
or U13228 (N_13228,N_12847,N_12934);
or U13229 (N_13229,N_12975,N_12860);
nor U13230 (N_13230,N_12892,N_12900);
or U13231 (N_13231,N_12854,N_12960);
and U13232 (N_13232,N_12831,N_12888);
and U13233 (N_13233,N_12780,N_12812);
or U13234 (N_13234,N_12924,N_12992);
and U13235 (N_13235,N_12913,N_12798);
xnor U13236 (N_13236,N_12907,N_12807);
nand U13237 (N_13237,N_12931,N_12836);
and U13238 (N_13238,N_12915,N_12924);
nand U13239 (N_13239,N_12963,N_12903);
or U13240 (N_13240,N_12762,N_12849);
nand U13241 (N_13241,N_12957,N_12904);
nor U13242 (N_13242,N_12989,N_12880);
nand U13243 (N_13243,N_12777,N_12988);
nand U13244 (N_13244,N_12770,N_12997);
xnor U13245 (N_13245,N_12825,N_12893);
xnor U13246 (N_13246,N_12862,N_12807);
nor U13247 (N_13247,N_12937,N_12949);
and U13248 (N_13248,N_12940,N_12887);
xnor U13249 (N_13249,N_12880,N_12817);
or U13250 (N_13250,N_13238,N_13185);
nand U13251 (N_13251,N_13015,N_13133);
xnor U13252 (N_13252,N_13011,N_13059);
or U13253 (N_13253,N_13196,N_13160);
nor U13254 (N_13254,N_13028,N_13131);
and U13255 (N_13255,N_13000,N_13064);
and U13256 (N_13256,N_13169,N_13178);
or U13257 (N_13257,N_13051,N_13018);
or U13258 (N_13258,N_13082,N_13054);
or U13259 (N_13259,N_13013,N_13071);
or U13260 (N_13260,N_13139,N_13219);
nand U13261 (N_13261,N_13075,N_13207);
or U13262 (N_13262,N_13126,N_13033);
and U13263 (N_13263,N_13188,N_13100);
xor U13264 (N_13264,N_13201,N_13080);
nand U13265 (N_13265,N_13199,N_13086);
or U13266 (N_13266,N_13066,N_13005);
and U13267 (N_13267,N_13241,N_13115);
or U13268 (N_13268,N_13122,N_13097);
nand U13269 (N_13269,N_13101,N_13065);
or U13270 (N_13270,N_13008,N_13058);
or U13271 (N_13271,N_13129,N_13110);
and U13272 (N_13272,N_13210,N_13150);
nor U13273 (N_13273,N_13056,N_13077);
nor U13274 (N_13274,N_13229,N_13079);
nand U13275 (N_13275,N_13234,N_13181);
nor U13276 (N_13276,N_13104,N_13175);
xnor U13277 (N_13277,N_13039,N_13026);
nor U13278 (N_13278,N_13147,N_13137);
and U13279 (N_13279,N_13030,N_13046);
xor U13280 (N_13280,N_13180,N_13204);
or U13281 (N_13281,N_13246,N_13085);
and U13282 (N_13282,N_13007,N_13083);
and U13283 (N_13283,N_13235,N_13078);
and U13284 (N_13284,N_13105,N_13057);
xnor U13285 (N_13285,N_13248,N_13195);
and U13286 (N_13286,N_13052,N_13036);
nor U13287 (N_13287,N_13116,N_13109);
xnor U13288 (N_13288,N_13192,N_13061);
and U13289 (N_13289,N_13037,N_13024);
and U13290 (N_13290,N_13038,N_13114);
or U13291 (N_13291,N_13073,N_13132);
nand U13292 (N_13292,N_13184,N_13032);
xnor U13293 (N_13293,N_13161,N_13168);
and U13294 (N_13294,N_13165,N_13130);
nor U13295 (N_13295,N_13228,N_13063);
nor U13296 (N_13296,N_13088,N_13009);
or U13297 (N_13297,N_13006,N_13103);
nand U13298 (N_13298,N_13031,N_13021);
or U13299 (N_13299,N_13102,N_13099);
and U13300 (N_13300,N_13186,N_13070);
or U13301 (N_13301,N_13220,N_13060);
nor U13302 (N_13302,N_13243,N_13224);
xnor U13303 (N_13303,N_13156,N_13134);
nor U13304 (N_13304,N_13230,N_13050);
xor U13305 (N_13305,N_13019,N_13242);
nor U13306 (N_13306,N_13172,N_13174);
or U13307 (N_13307,N_13027,N_13208);
or U13308 (N_13308,N_13041,N_13124);
nand U13309 (N_13309,N_13023,N_13245);
and U13310 (N_13310,N_13118,N_13107);
nand U13311 (N_13311,N_13153,N_13183);
and U13312 (N_13312,N_13112,N_13067);
xnor U13313 (N_13313,N_13140,N_13239);
nand U13314 (N_13314,N_13048,N_13221);
xor U13315 (N_13315,N_13092,N_13040);
or U13316 (N_13316,N_13162,N_13249);
and U13317 (N_13317,N_13043,N_13146);
and U13318 (N_13318,N_13232,N_13091);
nor U13319 (N_13319,N_13125,N_13227);
or U13320 (N_13320,N_13187,N_13062);
and U13321 (N_13321,N_13144,N_13016);
and U13322 (N_13322,N_13003,N_13142);
nor U13323 (N_13323,N_13177,N_13136);
nor U13324 (N_13324,N_13081,N_13143);
or U13325 (N_13325,N_13128,N_13226);
and U13326 (N_13326,N_13094,N_13098);
or U13327 (N_13327,N_13049,N_13022);
nor U13328 (N_13328,N_13096,N_13209);
nand U13329 (N_13329,N_13194,N_13069);
nand U13330 (N_13330,N_13089,N_13068);
or U13331 (N_13331,N_13198,N_13108);
nor U13332 (N_13332,N_13035,N_13240);
xor U13333 (N_13333,N_13029,N_13215);
or U13334 (N_13334,N_13123,N_13191);
or U13335 (N_13335,N_13182,N_13166);
or U13336 (N_13336,N_13202,N_13074);
nand U13337 (N_13337,N_13157,N_13211);
xnor U13338 (N_13338,N_13218,N_13151);
nor U13339 (N_13339,N_13145,N_13159);
xnor U13340 (N_13340,N_13164,N_13173);
xor U13341 (N_13341,N_13247,N_13045);
or U13342 (N_13342,N_13152,N_13084);
nor U13343 (N_13343,N_13055,N_13141);
nand U13344 (N_13344,N_13044,N_13190);
nor U13345 (N_13345,N_13206,N_13216);
nor U13346 (N_13346,N_13213,N_13214);
xnor U13347 (N_13347,N_13095,N_13205);
or U13348 (N_13348,N_13217,N_13017);
or U13349 (N_13349,N_13121,N_13117);
nand U13350 (N_13350,N_13179,N_13113);
xor U13351 (N_13351,N_13076,N_13072);
xor U13352 (N_13352,N_13233,N_13197);
or U13353 (N_13353,N_13222,N_13010);
xor U13354 (N_13354,N_13001,N_13193);
and U13355 (N_13355,N_13087,N_13119);
xnor U13356 (N_13356,N_13236,N_13203);
and U13357 (N_13357,N_13154,N_13093);
nand U13358 (N_13358,N_13090,N_13014);
nor U13359 (N_13359,N_13002,N_13025);
nand U13360 (N_13360,N_13111,N_13127);
and U13361 (N_13361,N_13176,N_13200);
and U13362 (N_13362,N_13170,N_13171);
nand U13363 (N_13363,N_13053,N_13120);
xor U13364 (N_13364,N_13212,N_13158);
and U13365 (N_13365,N_13167,N_13148);
and U13366 (N_13366,N_13135,N_13106);
xnor U13367 (N_13367,N_13138,N_13223);
xor U13368 (N_13368,N_13189,N_13163);
or U13369 (N_13369,N_13149,N_13155);
and U13370 (N_13370,N_13020,N_13012);
xor U13371 (N_13371,N_13225,N_13004);
or U13372 (N_13372,N_13047,N_13231);
nor U13373 (N_13373,N_13034,N_13244);
nor U13374 (N_13374,N_13042,N_13237);
xor U13375 (N_13375,N_13190,N_13004);
or U13376 (N_13376,N_13105,N_13120);
and U13377 (N_13377,N_13247,N_13171);
xnor U13378 (N_13378,N_13131,N_13135);
nor U13379 (N_13379,N_13061,N_13155);
nand U13380 (N_13380,N_13008,N_13025);
and U13381 (N_13381,N_13013,N_13190);
xnor U13382 (N_13382,N_13193,N_13026);
nand U13383 (N_13383,N_13232,N_13176);
or U13384 (N_13384,N_13209,N_13086);
nor U13385 (N_13385,N_13119,N_13012);
xor U13386 (N_13386,N_13130,N_13226);
nor U13387 (N_13387,N_13102,N_13173);
and U13388 (N_13388,N_13085,N_13110);
or U13389 (N_13389,N_13003,N_13095);
or U13390 (N_13390,N_13247,N_13038);
nor U13391 (N_13391,N_13127,N_13023);
or U13392 (N_13392,N_13085,N_13122);
xor U13393 (N_13393,N_13124,N_13234);
xor U13394 (N_13394,N_13040,N_13111);
xor U13395 (N_13395,N_13161,N_13085);
and U13396 (N_13396,N_13053,N_13228);
xnor U13397 (N_13397,N_13159,N_13021);
xnor U13398 (N_13398,N_13127,N_13030);
and U13399 (N_13399,N_13100,N_13038);
nor U13400 (N_13400,N_13056,N_13092);
and U13401 (N_13401,N_13010,N_13233);
nor U13402 (N_13402,N_13063,N_13031);
xnor U13403 (N_13403,N_13191,N_13190);
or U13404 (N_13404,N_13230,N_13214);
nor U13405 (N_13405,N_13015,N_13165);
and U13406 (N_13406,N_13245,N_13146);
nand U13407 (N_13407,N_13228,N_13192);
nor U13408 (N_13408,N_13172,N_13202);
nor U13409 (N_13409,N_13134,N_13225);
and U13410 (N_13410,N_13167,N_13200);
or U13411 (N_13411,N_13067,N_13084);
and U13412 (N_13412,N_13137,N_13025);
or U13413 (N_13413,N_13166,N_13054);
and U13414 (N_13414,N_13068,N_13006);
or U13415 (N_13415,N_13102,N_13001);
and U13416 (N_13416,N_13082,N_13095);
nand U13417 (N_13417,N_13087,N_13240);
nor U13418 (N_13418,N_13207,N_13177);
nor U13419 (N_13419,N_13128,N_13038);
and U13420 (N_13420,N_13022,N_13141);
or U13421 (N_13421,N_13046,N_13245);
xor U13422 (N_13422,N_13123,N_13059);
xnor U13423 (N_13423,N_13004,N_13215);
xor U13424 (N_13424,N_13230,N_13115);
nor U13425 (N_13425,N_13068,N_13209);
nor U13426 (N_13426,N_13006,N_13135);
or U13427 (N_13427,N_13230,N_13133);
nand U13428 (N_13428,N_13062,N_13157);
nor U13429 (N_13429,N_13187,N_13019);
nand U13430 (N_13430,N_13234,N_13076);
xor U13431 (N_13431,N_13053,N_13011);
or U13432 (N_13432,N_13146,N_13120);
nand U13433 (N_13433,N_13093,N_13107);
or U13434 (N_13434,N_13137,N_13077);
nor U13435 (N_13435,N_13009,N_13045);
and U13436 (N_13436,N_13095,N_13091);
xor U13437 (N_13437,N_13189,N_13052);
nand U13438 (N_13438,N_13209,N_13036);
nand U13439 (N_13439,N_13058,N_13164);
nor U13440 (N_13440,N_13062,N_13069);
nand U13441 (N_13441,N_13120,N_13022);
xnor U13442 (N_13442,N_13027,N_13037);
nor U13443 (N_13443,N_13176,N_13165);
and U13444 (N_13444,N_13050,N_13105);
and U13445 (N_13445,N_13203,N_13207);
or U13446 (N_13446,N_13130,N_13038);
or U13447 (N_13447,N_13242,N_13247);
and U13448 (N_13448,N_13089,N_13030);
nand U13449 (N_13449,N_13229,N_13247);
nor U13450 (N_13450,N_13182,N_13194);
nand U13451 (N_13451,N_13091,N_13150);
nor U13452 (N_13452,N_13228,N_13090);
or U13453 (N_13453,N_13231,N_13025);
and U13454 (N_13454,N_13202,N_13096);
nand U13455 (N_13455,N_13195,N_13117);
nor U13456 (N_13456,N_13139,N_13160);
nand U13457 (N_13457,N_13004,N_13103);
and U13458 (N_13458,N_13057,N_13084);
and U13459 (N_13459,N_13006,N_13101);
or U13460 (N_13460,N_13222,N_13230);
or U13461 (N_13461,N_13150,N_13119);
nor U13462 (N_13462,N_13016,N_13158);
and U13463 (N_13463,N_13085,N_13069);
or U13464 (N_13464,N_13136,N_13175);
and U13465 (N_13465,N_13042,N_13167);
nand U13466 (N_13466,N_13110,N_13071);
or U13467 (N_13467,N_13229,N_13022);
and U13468 (N_13468,N_13246,N_13029);
nand U13469 (N_13469,N_13235,N_13088);
xnor U13470 (N_13470,N_13056,N_13131);
xor U13471 (N_13471,N_13019,N_13023);
nor U13472 (N_13472,N_13154,N_13102);
nor U13473 (N_13473,N_13198,N_13117);
or U13474 (N_13474,N_13026,N_13156);
and U13475 (N_13475,N_13202,N_13021);
nor U13476 (N_13476,N_13143,N_13117);
or U13477 (N_13477,N_13065,N_13090);
or U13478 (N_13478,N_13161,N_13071);
nor U13479 (N_13479,N_13102,N_13212);
or U13480 (N_13480,N_13078,N_13242);
nor U13481 (N_13481,N_13028,N_13014);
nor U13482 (N_13482,N_13109,N_13125);
or U13483 (N_13483,N_13134,N_13140);
or U13484 (N_13484,N_13007,N_13174);
nand U13485 (N_13485,N_13004,N_13198);
nor U13486 (N_13486,N_13002,N_13028);
nor U13487 (N_13487,N_13176,N_13017);
and U13488 (N_13488,N_13062,N_13104);
nand U13489 (N_13489,N_13247,N_13101);
and U13490 (N_13490,N_13166,N_13171);
or U13491 (N_13491,N_13244,N_13016);
and U13492 (N_13492,N_13232,N_13080);
and U13493 (N_13493,N_13229,N_13139);
xor U13494 (N_13494,N_13045,N_13200);
nor U13495 (N_13495,N_13229,N_13018);
nand U13496 (N_13496,N_13058,N_13160);
xor U13497 (N_13497,N_13072,N_13081);
or U13498 (N_13498,N_13121,N_13153);
nand U13499 (N_13499,N_13177,N_13031);
nor U13500 (N_13500,N_13475,N_13463);
and U13501 (N_13501,N_13396,N_13451);
or U13502 (N_13502,N_13281,N_13390);
and U13503 (N_13503,N_13361,N_13452);
nor U13504 (N_13504,N_13478,N_13370);
nor U13505 (N_13505,N_13365,N_13375);
xor U13506 (N_13506,N_13333,N_13344);
nand U13507 (N_13507,N_13393,N_13360);
nand U13508 (N_13508,N_13261,N_13320);
nor U13509 (N_13509,N_13372,N_13308);
and U13510 (N_13510,N_13420,N_13250);
or U13511 (N_13511,N_13289,N_13258);
nand U13512 (N_13512,N_13432,N_13351);
nor U13513 (N_13513,N_13348,N_13427);
and U13514 (N_13514,N_13262,N_13304);
nand U13515 (N_13515,N_13418,N_13416);
or U13516 (N_13516,N_13378,N_13283);
or U13517 (N_13517,N_13408,N_13411);
nor U13518 (N_13518,N_13291,N_13421);
nand U13519 (N_13519,N_13367,N_13442);
nor U13520 (N_13520,N_13492,N_13286);
xor U13521 (N_13521,N_13434,N_13376);
and U13522 (N_13522,N_13414,N_13430);
xnor U13523 (N_13523,N_13271,N_13465);
nor U13524 (N_13524,N_13406,N_13357);
or U13525 (N_13525,N_13447,N_13340);
xor U13526 (N_13526,N_13288,N_13256);
nand U13527 (N_13527,N_13326,N_13267);
and U13528 (N_13528,N_13436,N_13343);
nand U13529 (N_13529,N_13362,N_13314);
or U13530 (N_13530,N_13356,N_13251);
and U13531 (N_13531,N_13491,N_13377);
nor U13532 (N_13532,N_13481,N_13495);
nor U13533 (N_13533,N_13383,N_13270);
and U13534 (N_13534,N_13309,N_13419);
xnor U13535 (N_13535,N_13327,N_13268);
xnor U13536 (N_13536,N_13473,N_13303);
xnor U13537 (N_13537,N_13347,N_13363);
nand U13538 (N_13538,N_13449,N_13255);
and U13539 (N_13539,N_13282,N_13339);
and U13540 (N_13540,N_13382,N_13423);
or U13541 (N_13541,N_13254,N_13443);
nand U13542 (N_13542,N_13444,N_13269);
nor U13543 (N_13543,N_13457,N_13290);
xnor U13544 (N_13544,N_13470,N_13477);
xnor U13545 (N_13545,N_13467,N_13471);
nor U13546 (N_13546,N_13295,N_13368);
xor U13547 (N_13547,N_13341,N_13428);
or U13548 (N_13548,N_13294,N_13342);
or U13549 (N_13549,N_13431,N_13394);
and U13550 (N_13550,N_13331,N_13300);
nor U13551 (N_13551,N_13392,N_13409);
and U13552 (N_13552,N_13364,N_13305);
xnor U13553 (N_13553,N_13438,N_13429);
nand U13554 (N_13554,N_13276,N_13285);
or U13555 (N_13555,N_13490,N_13358);
nor U13556 (N_13556,N_13301,N_13319);
nand U13557 (N_13557,N_13252,N_13293);
nor U13558 (N_13558,N_13422,N_13260);
nand U13559 (N_13559,N_13337,N_13315);
and U13560 (N_13560,N_13389,N_13456);
xor U13561 (N_13561,N_13381,N_13454);
xnor U13562 (N_13562,N_13401,N_13296);
and U13563 (N_13563,N_13259,N_13455);
nand U13564 (N_13564,N_13403,N_13445);
nand U13565 (N_13565,N_13488,N_13391);
or U13566 (N_13566,N_13410,N_13387);
or U13567 (N_13567,N_13346,N_13323);
or U13568 (N_13568,N_13266,N_13474);
nor U13569 (N_13569,N_13460,N_13379);
nand U13570 (N_13570,N_13277,N_13322);
xnor U13571 (N_13571,N_13352,N_13412);
or U13572 (N_13572,N_13257,N_13446);
and U13573 (N_13573,N_13468,N_13469);
nand U13574 (N_13574,N_13388,N_13310);
nand U13575 (N_13575,N_13426,N_13280);
nand U13576 (N_13576,N_13311,N_13334);
nor U13577 (N_13577,N_13321,N_13279);
xnor U13578 (N_13578,N_13292,N_13329);
nor U13579 (N_13579,N_13253,N_13395);
nor U13580 (N_13580,N_13479,N_13278);
or U13581 (N_13581,N_13464,N_13384);
and U13582 (N_13582,N_13302,N_13450);
nand U13583 (N_13583,N_13458,N_13287);
or U13584 (N_13584,N_13275,N_13398);
xor U13585 (N_13585,N_13484,N_13459);
or U13586 (N_13586,N_13399,N_13359);
and U13587 (N_13587,N_13386,N_13489);
or U13588 (N_13588,N_13273,N_13307);
and U13589 (N_13589,N_13298,N_13274);
nor U13590 (N_13590,N_13485,N_13462);
and U13591 (N_13591,N_13472,N_13264);
and U13592 (N_13592,N_13466,N_13497);
xnor U13593 (N_13593,N_13439,N_13369);
and U13594 (N_13594,N_13480,N_13297);
xnor U13595 (N_13595,N_13366,N_13345);
nand U13596 (N_13596,N_13441,N_13338);
xor U13597 (N_13597,N_13374,N_13415);
or U13598 (N_13598,N_13496,N_13330);
and U13599 (N_13599,N_13325,N_13385);
or U13600 (N_13600,N_13284,N_13413);
xor U13601 (N_13601,N_13354,N_13380);
nand U13602 (N_13602,N_13355,N_13435);
xnor U13603 (N_13603,N_13448,N_13318);
or U13604 (N_13604,N_13350,N_13400);
xor U13605 (N_13605,N_13335,N_13407);
nand U13606 (N_13606,N_13328,N_13316);
or U13607 (N_13607,N_13476,N_13487);
nor U13608 (N_13608,N_13306,N_13317);
xor U13609 (N_13609,N_13265,N_13272);
and U13610 (N_13610,N_13263,N_13397);
and U13611 (N_13611,N_13324,N_13498);
xor U13612 (N_13612,N_13313,N_13373);
or U13613 (N_13613,N_13433,N_13453);
or U13614 (N_13614,N_13482,N_13371);
or U13615 (N_13615,N_13493,N_13349);
nand U13616 (N_13616,N_13299,N_13486);
and U13617 (N_13617,N_13461,N_13494);
or U13618 (N_13618,N_13336,N_13402);
and U13619 (N_13619,N_13437,N_13425);
nand U13620 (N_13620,N_13404,N_13424);
or U13621 (N_13621,N_13499,N_13405);
xor U13622 (N_13622,N_13440,N_13353);
or U13623 (N_13623,N_13332,N_13312);
nand U13624 (N_13624,N_13417,N_13483);
nor U13625 (N_13625,N_13361,N_13308);
xnor U13626 (N_13626,N_13479,N_13487);
and U13627 (N_13627,N_13464,N_13320);
xnor U13628 (N_13628,N_13319,N_13367);
and U13629 (N_13629,N_13271,N_13463);
nand U13630 (N_13630,N_13300,N_13456);
xnor U13631 (N_13631,N_13352,N_13407);
nor U13632 (N_13632,N_13374,N_13488);
nor U13633 (N_13633,N_13423,N_13273);
nor U13634 (N_13634,N_13427,N_13398);
nand U13635 (N_13635,N_13412,N_13278);
or U13636 (N_13636,N_13387,N_13429);
xnor U13637 (N_13637,N_13265,N_13436);
and U13638 (N_13638,N_13431,N_13251);
xnor U13639 (N_13639,N_13468,N_13493);
nand U13640 (N_13640,N_13392,N_13444);
and U13641 (N_13641,N_13494,N_13300);
and U13642 (N_13642,N_13447,N_13344);
nor U13643 (N_13643,N_13472,N_13362);
and U13644 (N_13644,N_13333,N_13413);
and U13645 (N_13645,N_13342,N_13347);
and U13646 (N_13646,N_13398,N_13412);
and U13647 (N_13647,N_13392,N_13332);
and U13648 (N_13648,N_13458,N_13277);
nor U13649 (N_13649,N_13365,N_13411);
nand U13650 (N_13650,N_13382,N_13309);
nand U13651 (N_13651,N_13282,N_13294);
nand U13652 (N_13652,N_13447,N_13342);
or U13653 (N_13653,N_13351,N_13474);
nor U13654 (N_13654,N_13293,N_13417);
nor U13655 (N_13655,N_13466,N_13406);
or U13656 (N_13656,N_13260,N_13348);
xor U13657 (N_13657,N_13485,N_13465);
xnor U13658 (N_13658,N_13483,N_13292);
nor U13659 (N_13659,N_13468,N_13385);
xnor U13660 (N_13660,N_13498,N_13312);
and U13661 (N_13661,N_13316,N_13427);
nand U13662 (N_13662,N_13278,N_13267);
or U13663 (N_13663,N_13336,N_13397);
or U13664 (N_13664,N_13447,N_13359);
and U13665 (N_13665,N_13361,N_13316);
xor U13666 (N_13666,N_13401,N_13322);
or U13667 (N_13667,N_13450,N_13458);
nand U13668 (N_13668,N_13341,N_13432);
nand U13669 (N_13669,N_13380,N_13287);
xor U13670 (N_13670,N_13392,N_13292);
and U13671 (N_13671,N_13418,N_13296);
xor U13672 (N_13672,N_13460,N_13486);
and U13673 (N_13673,N_13495,N_13350);
or U13674 (N_13674,N_13333,N_13308);
or U13675 (N_13675,N_13465,N_13409);
or U13676 (N_13676,N_13380,N_13284);
and U13677 (N_13677,N_13484,N_13269);
or U13678 (N_13678,N_13318,N_13404);
xnor U13679 (N_13679,N_13411,N_13482);
xnor U13680 (N_13680,N_13359,N_13443);
or U13681 (N_13681,N_13345,N_13429);
and U13682 (N_13682,N_13472,N_13320);
nor U13683 (N_13683,N_13250,N_13415);
or U13684 (N_13684,N_13492,N_13476);
nand U13685 (N_13685,N_13488,N_13301);
and U13686 (N_13686,N_13410,N_13386);
or U13687 (N_13687,N_13421,N_13444);
xnor U13688 (N_13688,N_13441,N_13284);
nand U13689 (N_13689,N_13307,N_13301);
or U13690 (N_13690,N_13448,N_13431);
nor U13691 (N_13691,N_13368,N_13408);
nand U13692 (N_13692,N_13437,N_13349);
or U13693 (N_13693,N_13301,N_13462);
nor U13694 (N_13694,N_13368,N_13420);
and U13695 (N_13695,N_13317,N_13458);
nor U13696 (N_13696,N_13280,N_13486);
and U13697 (N_13697,N_13404,N_13433);
xnor U13698 (N_13698,N_13459,N_13483);
and U13699 (N_13699,N_13292,N_13348);
nand U13700 (N_13700,N_13391,N_13336);
and U13701 (N_13701,N_13463,N_13311);
or U13702 (N_13702,N_13324,N_13480);
nand U13703 (N_13703,N_13259,N_13287);
and U13704 (N_13704,N_13392,N_13280);
or U13705 (N_13705,N_13362,N_13490);
or U13706 (N_13706,N_13367,N_13423);
xnor U13707 (N_13707,N_13342,N_13363);
or U13708 (N_13708,N_13335,N_13314);
and U13709 (N_13709,N_13270,N_13280);
xnor U13710 (N_13710,N_13364,N_13311);
nand U13711 (N_13711,N_13400,N_13335);
nand U13712 (N_13712,N_13322,N_13421);
or U13713 (N_13713,N_13406,N_13381);
or U13714 (N_13714,N_13495,N_13439);
nor U13715 (N_13715,N_13329,N_13340);
and U13716 (N_13716,N_13409,N_13424);
and U13717 (N_13717,N_13278,N_13443);
or U13718 (N_13718,N_13458,N_13250);
nand U13719 (N_13719,N_13453,N_13464);
nor U13720 (N_13720,N_13477,N_13485);
nor U13721 (N_13721,N_13288,N_13480);
and U13722 (N_13722,N_13420,N_13307);
and U13723 (N_13723,N_13296,N_13436);
nor U13724 (N_13724,N_13497,N_13311);
or U13725 (N_13725,N_13303,N_13280);
nand U13726 (N_13726,N_13433,N_13375);
and U13727 (N_13727,N_13344,N_13292);
nor U13728 (N_13728,N_13328,N_13307);
xnor U13729 (N_13729,N_13408,N_13427);
nand U13730 (N_13730,N_13481,N_13266);
nand U13731 (N_13731,N_13309,N_13266);
xor U13732 (N_13732,N_13403,N_13423);
nor U13733 (N_13733,N_13317,N_13417);
nand U13734 (N_13734,N_13310,N_13291);
nand U13735 (N_13735,N_13281,N_13267);
xnor U13736 (N_13736,N_13481,N_13462);
xor U13737 (N_13737,N_13480,N_13387);
nor U13738 (N_13738,N_13382,N_13338);
or U13739 (N_13739,N_13337,N_13344);
nand U13740 (N_13740,N_13337,N_13447);
xnor U13741 (N_13741,N_13345,N_13326);
and U13742 (N_13742,N_13321,N_13324);
and U13743 (N_13743,N_13315,N_13332);
nand U13744 (N_13744,N_13256,N_13492);
nor U13745 (N_13745,N_13257,N_13362);
and U13746 (N_13746,N_13489,N_13353);
xor U13747 (N_13747,N_13285,N_13383);
or U13748 (N_13748,N_13254,N_13289);
or U13749 (N_13749,N_13472,N_13437);
nor U13750 (N_13750,N_13727,N_13709);
xor U13751 (N_13751,N_13572,N_13713);
and U13752 (N_13752,N_13603,N_13620);
and U13753 (N_13753,N_13721,N_13519);
xor U13754 (N_13754,N_13518,N_13517);
or U13755 (N_13755,N_13719,N_13502);
nor U13756 (N_13756,N_13629,N_13725);
xnor U13757 (N_13757,N_13748,N_13522);
xnor U13758 (N_13758,N_13500,N_13588);
nor U13759 (N_13759,N_13536,N_13612);
nand U13760 (N_13760,N_13616,N_13574);
nand U13761 (N_13761,N_13706,N_13509);
and U13762 (N_13762,N_13726,N_13557);
xor U13763 (N_13763,N_13635,N_13613);
or U13764 (N_13764,N_13652,N_13569);
and U13765 (N_13765,N_13530,N_13722);
nor U13766 (N_13766,N_13614,N_13567);
nand U13767 (N_13767,N_13589,N_13570);
and U13768 (N_13768,N_13649,N_13657);
nor U13769 (N_13769,N_13523,N_13711);
nor U13770 (N_13770,N_13724,N_13674);
nand U13771 (N_13771,N_13683,N_13609);
and U13772 (N_13772,N_13605,N_13633);
nand U13773 (N_13773,N_13561,N_13704);
or U13774 (N_13774,N_13602,N_13507);
and U13775 (N_13775,N_13545,N_13624);
and U13776 (N_13776,N_13601,N_13640);
xnor U13777 (N_13777,N_13626,N_13556);
and U13778 (N_13778,N_13729,N_13539);
and U13779 (N_13779,N_13648,N_13672);
nand U13780 (N_13780,N_13741,N_13533);
xor U13781 (N_13781,N_13696,N_13693);
and U13782 (N_13782,N_13668,N_13643);
nand U13783 (N_13783,N_13520,N_13645);
xor U13784 (N_13784,N_13511,N_13695);
or U13785 (N_13785,N_13663,N_13506);
nor U13786 (N_13786,N_13733,N_13577);
nand U13787 (N_13787,N_13513,N_13598);
xnor U13788 (N_13788,N_13694,N_13503);
xnor U13789 (N_13789,N_13636,N_13595);
nor U13790 (N_13790,N_13548,N_13720);
or U13791 (N_13791,N_13611,N_13699);
xnor U13792 (N_13792,N_13534,N_13700);
nor U13793 (N_13793,N_13673,N_13591);
nand U13794 (N_13794,N_13714,N_13562);
and U13795 (N_13795,N_13617,N_13580);
nor U13796 (N_13796,N_13527,N_13565);
nand U13797 (N_13797,N_13630,N_13691);
or U13798 (N_13798,N_13615,N_13687);
nor U13799 (N_13799,N_13676,N_13578);
nand U13800 (N_13800,N_13563,N_13701);
nor U13801 (N_13801,N_13553,N_13689);
or U13802 (N_13802,N_13621,N_13690);
nor U13803 (N_13803,N_13610,N_13682);
nor U13804 (N_13804,N_13627,N_13607);
nand U13805 (N_13805,N_13568,N_13708);
nor U13806 (N_13806,N_13728,N_13526);
nor U13807 (N_13807,N_13579,N_13739);
or U13808 (N_13808,N_13505,N_13543);
nand U13809 (N_13809,N_13516,N_13596);
and U13810 (N_13810,N_13535,N_13638);
nor U13811 (N_13811,N_13515,N_13675);
xor U13812 (N_13812,N_13745,N_13504);
xor U13813 (N_13813,N_13524,N_13718);
xnor U13814 (N_13814,N_13743,N_13646);
xor U13815 (N_13815,N_13734,N_13666);
nor U13816 (N_13816,N_13600,N_13552);
nor U13817 (N_13817,N_13512,N_13658);
or U13818 (N_13818,N_13592,N_13514);
or U13819 (N_13819,N_13542,N_13670);
nand U13820 (N_13820,N_13593,N_13537);
or U13821 (N_13821,N_13740,N_13662);
nand U13822 (N_13822,N_13599,N_13508);
nand U13823 (N_13823,N_13597,N_13692);
and U13824 (N_13824,N_13573,N_13684);
nand U13825 (N_13825,N_13678,N_13586);
or U13826 (N_13826,N_13584,N_13650);
nand U13827 (N_13827,N_13501,N_13571);
xor U13828 (N_13828,N_13546,N_13525);
or U13829 (N_13829,N_13558,N_13651);
nor U13830 (N_13830,N_13628,N_13717);
or U13831 (N_13831,N_13744,N_13661);
and U13832 (N_13832,N_13671,N_13698);
nand U13833 (N_13833,N_13669,N_13590);
and U13834 (N_13834,N_13622,N_13712);
and U13835 (N_13835,N_13554,N_13705);
nor U13836 (N_13836,N_13639,N_13685);
xor U13837 (N_13837,N_13654,N_13679);
nor U13838 (N_13838,N_13664,N_13547);
nor U13839 (N_13839,N_13560,N_13581);
nor U13840 (N_13840,N_13555,N_13587);
or U13841 (N_13841,N_13566,N_13715);
nand U13842 (N_13842,N_13528,N_13541);
nand U13843 (N_13843,N_13510,N_13697);
nor U13844 (N_13844,N_13731,N_13551);
and U13845 (N_13845,N_13631,N_13686);
and U13846 (N_13846,N_13608,N_13655);
or U13847 (N_13847,N_13585,N_13730);
nand U13848 (N_13848,N_13642,N_13659);
xor U13849 (N_13849,N_13641,N_13531);
nand U13850 (N_13850,N_13653,N_13688);
nand U13851 (N_13851,N_13660,N_13619);
and U13852 (N_13852,N_13582,N_13576);
or U13853 (N_13853,N_13583,N_13637);
xor U13854 (N_13854,N_13656,N_13550);
nand U13855 (N_13855,N_13737,N_13749);
and U13856 (N_13856,N_13604,N_13742);
nor U13857 (N_13857,N_13540,N_13736);
xor U13858 (N_13858,N_13594,N_13677);
nand U13859 (N_13859,N_13665,N_13564);
and U13860 (N_13860,N_13747,N_13746);
or U13861 (N_13861,N_13707,N_13521);
nor U13862 (N_13862,N_13681,N_13680);
nand U13863 (N_13863,N_13538,N_13716);
xor U13864 (N_13864,N_13606,N_13644);
nand U13865 (N_13865,N_13575,N_13632);
and U13866 (N_13866,N_13703,N_13549);
and U13867 (N_13867,N_13529,N_13623);
or U13868 (N_13868,N_13532,N_13702);
and U13869 (N_13869,N_13710,N_13732);
nor U13870 (N_13870,N_13738,N_13667);
nor U13871 (N_13871,N_13559,N_13544);
xnor U13872 (N_13872,N_13618,N_13634);
or U13873 (N_13873,N_13735,N_13625);
nor U13874 (N_13874,N_13647,N_13723);
xnor U13875 (N_13875,N_13530,N_13695);
xor U13876 (N_13876,N_13694,N_13651);
and U13877 (N_13877,N_13554,N_13565);
nor U13878 (N_13878,N_13523,N_13578);
nand U13879 (N_13879,N_13741,N_13549);
nor U13880 (N_13880,N_13641,N_13562);
nand U13881 (N_13881,N_13702,N_13578);
nand U13882 (N_13882,N_13514,N_13523);
and U13883 (N_13883,N_13641,N_13691);
nor U13884 (N_13884,N_13638,N_13625);
and U13885 (N_13885,N_13510,N_13613);
or U13886 (N_13886,N_13698,N_13661);
xnor U13887 (N_13887,N_13574,N_13533);
and U13888 (N_13888,N_13562,N_13529);
and U13889 (N_13889,N_13662,N_13695);
and U13890 (N_13890,N_13689,N_13635);
xnor U13891 (N_13891,N_13644,N_13601);
or U13892 (N_13892,N_13613,N_13575);
nand U13893 (N_13893,N_13679,N_13599);
or U13894 (N_13894,N_13505,N_13624);
nand U13895 (N_13895,N_13545,N_13661);
nand U13896 (N_13896,N_13514,N_13633);
nor U13897 (N_13897,N_13693,N_13746);
or U13898 (N_13898,N_13618,N_13633);
and U13899 (N_13899,N_13732,N_13529);
and U13900 (N_13900,N_13620,N_13512);
and U13901 (N_13901,N_13629,N_13608);
or U13902 (N_13902,N_13519,N_13549);
xnor U13903 (N_13903,N_13690,N_13640);
nand U13904 (N_13904,N_13588,N_13530);
nand U13905 (N_13905,N_13629,N_13633);
nand U13906 (N_13906,N_13722,N_13640);
or U13907 (N_13907,N_13616,N_13641);
or U13908 (N_13908,N_13536,N_13500);
xor U13909 (N_13909,N_13676,N_13739);
and U13910 (N_13910,N_13698,N_13575);
or U13911 (N_13911,N_13528,N_13709);
nand U13912 (N_13912,N_13656,N_13553);
xnor U13913 (N_13913,N_13717,N_13651);
nand U13914 (N_13914,N_13638,N_13749);
nand U13915 (N_13915,N_13627,N_13642);
xnor U13916 (N_13916,N_13702,N_13607);
nand U13917 (N_13917,N_13733,N_13568);
and U13918 (N_13918,N_13699,N_13674);
nor U13919 (N_13919,N_13668,N_13500);
nand U13920 (N_13920,N_13561,N_13632);
xor U13921 (N_13921,N_13545,N_13532);
nand U13922 (N_13922,N_13546,N_13539);
nor U13923 (N_13923,N_13544,N_13729);
xor U13924 (N_13924,N_13503,N_13709);
xor U13925 (N_13925,N_13632,N_13677);
xnor U13926 (N_13926,N_13616,N_13580);
nand U13927 (N_13927,N_13541,N_13688);
xor U13928 (N_13928,N_13588,N_13722);
xor U13929 (N_13929,N_13506,N_13539);
nand U13930 (N_13930,N_13571,N_13578);
and U13931 (N_13931,N_13550,N_13693);
nand U13932 (N_13932,N_13513,N_13611);
nand U13933 (N_13933,N_13681,N_13661);
or U13934 (N_13934,N_13683,N_13576);
nand U13935 (N_13935,N_13557,N_13533);
nand U13936 (N_13936,N_13610,N_13618);
xnor U13937 (N_13937,N_13648,N_13526);
or U13938 (N_13938,N_13531,N_13629);
xor U13939 (N_13939,N_13719,N_13622);
nand U13940 (N_13940,N_13614,N_13609);
or U13941 (N_13941,N_13607,N_13728);
or U13942 (N_13942,N_13576,N_13714);
and U13943 (N_13943,N_13530,N_13690);
nor U13944 (N_13944,N_13531,N_13737);
xor U13945 (N_13945,N_13545,N_13561);
nor U13946 (N_13946,N_13589,N_13749);
or U13947 (N_13947,N_13510,N_13745);
or U13948 (N_13948,N_13735,N_13546);
and U13949 (N_13949,N_13667,N_13633);
nor U13950 (N_13950,N_13664,N_13616);
and U13951 (N_13951,N_13698,N_13632);
xnor U13952 (N_13952,N_13563,N_13541);
nor U13953 (N_13953,N_13515,N_13560);
nor U13954 (N_13954,N_13549,N_13516);
xor U13955 (N_13955,N_13709,N_13546);
and U13956 (N_13956,N_13514,N_13627);
or U13957 (N_13957,N_13651,N_13551);
and U13958 (N_13958,N_13500,N_13621);
xor U13959 (N_13959,N_13537,N_13578);
xor U13960 (N_13960,N_13527,N_13593);
or U13961 (N_13961,N_13649,N_13608);
and U13962 (N_13962,N_13698,N_13597);
or U13963 (N_13963,N_13615,N_13649);
and U13964 (N_13964,N_13507,N_13541);
or U13965 (N_13965,N_13670,N_13552);
nor U13966 (N_13966,N_13561,N_13723);
nand U13967 (N_13967,N_13614,N_13699);
nor U13968 (N_13968,N_13726,N_13610);
or U13969 (N_13969,N_13715,N_13640);
xor U13970 (N_13970,N_13663,N_13597);
nor U13971 (N_13971,N_13738,N_13505);
or U13972 (N_13972,N_13569,N_13568);
and U13973 (N_13973,N_13698,N_13543);
nor U13974 (N_13974,N_13502,N_13590);
nor U13975 (N_13975,N_13614,N_13521);
and U13976 (N_13976,N_13725,N_13682);
xor U13977 (N_13977,N_13657,N_13530);
or U13978 (N_13978,N_13632,N_13700);
nor U13979 (N_13979,N_13627,N_13502);
nor U13980 (N_13980,N_13627,N_13508);
or U13981 (N_13981,N_13526,N_13698);
or U13982 (N_13982,N_13650,N_13738);
and U13983 (N_13983,N_13634,N_13515);
xor U13984 (N_13984,N_13548,N_13613);
nor U13985 (N_13985,N_13606,N_13744);
and U13986 (N_13986,N_13605,N_13738);
xnor U13987 (N_13987,N_13647,N_13640);
or U13988 (N_13988,N_13513,N_13655);
and U13989 (N_13989,N_13745,N_13700);
nor U13990 (N_13990,N_13525,N_13678);
nor U13991 (N_13991,N_13672,N_13560);
or U13992 (N_13992,N_13590,N_13727);
or U13993 (N_13993,N_13572,N_13554);
nand U13994 (N_13994,N_13648,N_13651);
nand U13995 (N_13995,N_13533,N_13519);
nor U13996 (N_13996,N_13526,N_13675);
and U13997 (N_13997,N_13693,N_13645);
and U13998 (N_13998,N_13545,N_13596);
xnor U13999 (N_13999,N_13722,N_13579);
nor U14000 (N_14000,N_13943,N_13953);
or U14001 (N_14001,N_13913,N_13989);
and U14002 (N_14002,N_13821,N_13757);
nand U14003 (N_14003,N_13944,N_13759);
nor U14004 (N_14004,N_13853,N_13831);
nand U14005 (N_14005,N_13787,N_13959);
and U14006 (N_14006,N_13833,N_13771);
xor U14007 (N_14007,N_13937,N_13889);
nand U14008 (N_14008,N_13870,N_13996);
or U14009 (N_14009,N_13985,N_13804);
nand U14010 (N_14010,N_13849,N_13916);
and U14011 (N_14011,N_13762,N_13756);
or U14012 (N_14012,N_13767,N_13963);
nand U14013 (N_14013,N_13920,N_13835);
nor U14014 (N_14014,N_13842,N_13906);
xnor U14015 (N_14015,N_13967,N_13978);
and U14016 (N_14016,N_13918,N_13784);
or U14017 (N_14017,N_13981,N_13778);
xor U14018 (N_14018,N_13895,N_13919);
nand U14019 (N_14019,N_13817,N_13911);
or U14020 (N_14020,N_13903,N_13823);
xnor U14021 (N_14021,N_13826,N_13798);
or U14022 (N_14022,N_13803,N_13800);
and U14023 (N_14023,N_13936,N_13818);
nand U14024 (N_14024,N_13838,N_13830);
xor U14025 (N_14025,N_13880,N_13984);
nand U14026 (N_14026,N_13884,N_13761);
nor U14027 (N_14027,N_13801,N_13837);
and U14028 (N_14028,N_13930,N_13914);
nor U14029 (N_14029,N_13766,N_13986);
and U14030 (N_14030,N_13777,N_13898);
nor U14031 (N_14031,N_13928,N_13965);
and U14032 (N_14032,N_13949,N_13763);
nor U14033 (N_14033,N_13808,N_13990);
and U14034 (N_14034,N_13956,N_13786);
and U14035 (N_14035,N_13931,N_13793);
nor U14036 (N_14036,N_13910,N_13827);
xnor U14037 (N_14037,N_13902,N_13899);
nand U14038 (N_14038,N_13946,N_13909);
nand U14039 (N_14039,N_13850,N_13754);
or U14040 (N_14040,N_13790,N_13825);
and U14041 (N_14041,N_13845,N_13776);
nor U14042 (N_14042,N_13795,N_13810);
nand U14043 (N_14043,N_13925,N_13952);
and U14044 (N_14044,N_13885,N_13815);
xor U14045 (N_14045,N_13819,N_13950);
nor U14046 (N_14046,N_13980,N_13994);
nand U14047 (N_14047,N_13905,N_13955);
or U14048 (N_14048,N_13875,N_13922);
nor U14049 (N_14049,N_13832,N_13843);
xnor U14050 (N_14050,N_13792,N_13768);
nor U14051 (N_14051,N_13864,N_13901);
nor U14052 (N_14052,N_13893,N_13934);
nand U14053 (N_14053,N_13995,N_13858);
nand U14054 (N_14054,N_13834,N_13775);
or U14055 (N_14055,N_13969,N_13882);
nand U14056 (N_14056,N_13966,N_13781);
and U14057 (N_14057,N_13948,N_13829);
xnor U14058 (N_14058,N_13890,N_13836);
and U14059 (N_14059,N_13824,N_13774);
nand U14060 (N_14060,N_13789,N_13794);
xor U14061 (N_14061,N_13881,N_13957);
nand U14062 (N_14062,N_13813,N_13888);
xor U14063 (N_14063,N_13779,N_13960);
nor U14064 (N_14064,N_13887,N_13961);
nor U14065 (N_14065,N_13846,N_13852);
xor U14066 (N_14066,N_13861,N_13841);
nand U14067 (N_14067,N_13979,N_13924);
nand U14068 (N_14068,N_13886,N_13970);
and U14069 (N_14069,N_13863,N_13942);
nand U14070 (N_14070,N_13806,N_13951);
nor U14071 (N_14071,N_13878,N_13805);
or U14072 (N_14072,N_13879,N_13983);
nor U14073 (N_14073,N_13987,N_13855);
or U14074 (N_14074,N_13788,N_13892);
and U14075 (N_14075,N_13954,N_13859);
nor U14076 (N_14076,N_13972,N_13940);
nand U14077 (N_14077,N_13868,N_13915);
nor U14078 (N_14078,N_13816,N_13927);
nor U14079 (N_14079,N_13993,N_13854);
or U14080 (N_14080,N_13904,N_13783);
or U14081 (N_14081,N_13785,N_13973);
and U14082 (N_14082,N_13932,N_13857);
and U14083 (N_14083,N_13758,N_13769);
xnor U14084 (N_14084,N_13844,N_13753);
xor U14085 (N_14085,N_13802,N_13839);
nor U14086 (N_14086,N_13974,N_13872);
or U14087 (N_14087,N_13917,N_13865);
xor U14088 (N_14088,N_13820,N_13998);
or U14089 (N_14089,N_13772,N_13883);
nor U14090 (N_14090,N_13867,N_13782);
and U14091 (N_14091,N_13938,N_13807);
nor U14092 (N_14092,N_13999,N_13945);
or U14093 (N_14093,N_13897,N_13929);
and U14094 (N_14094,N_13921,N_13939);
xnor U14095 (N_14095,N_13791,N_13991);
nor U14096 (N_14096,N_13780,N_13765);
or U14097 (N_14097,N_13997,N_13796);
xnor U14098 (N_14098,N_13814,N_13866);
and U14099 (N_14099,N_13873,N_13828);
nor U14100 (N_14100,N_13988,N_13962);
nand U14101 (N_14101,N_13975,N_13811);
nor U14102 (N_14102,N_13923,N_13840);
nand U14103 (N_14103,N_13926,N_13812);
nor U14104 (N_14104,N_13822,N_13752);
and U14105 (N_14105,N_13773,N_13977);
nand U14106 (N_14106,N_13847,N_13935);
nand U14107 (N_14107,N_13751,N_13877);
or U14108 (N_14108,N_13976,N_13958);
or U14109 (N_14109,N_13876,N_13851);
and U14110 (N_14110,N_13809,N_13755);
and U14111 (N_14111,N_13860,N_13907);
nor U14112 (N_14112,N_13750,N_13894);
nor U14113 (N_14113,N_13770,N_13900);
or U14114 (N_14114,N_13941,N_13971);
nand U14115 (N_14115,N_13874,N_13871);
nor U14116 (N_14116,N_13760,N_13764);
and U14117 (N_14117,N_13799,N_13896);
or U14118 (N_14118,N_13862,N_13982);
and U14119 (N_14119,N_13908,N_13856);
nand U14120 (N_14120,N_13968,N_13947);
nand U14121 (N_14121,N_13912,N_13964);
nor U14122 (N_14122,N_13891,N_13992);
or U14123 (N_14123,N_13848,N_13869);
or U14124 (N_14124,N_13933,N_13797);
nor U14125 (N_14125,N_13987,N_13872);
and U14126 (N_14126,N_13832,N_13949);
and U14127 (N_14127,N_13794,N_13785);
nor U14128 (N_14128,N_13884,N_13753);
nand U14129 (N_14129,N_13926,N_13854);
xnor U14130 (N_14130,N_13751,N_13942);
nor U14131 (N_14131,N_13890,N_13752);
nor U14132 (N_14132,N_13784,N_13892);
nand U14133 (N_14133,N_13819,N_13947);
or U14134 (N_14134,N_13971,N_13816);
nor U14135 (N_14135,N_13784,N_13951);
or U14136 (N_14136,N_13964,N_13816);
or U14137 (N_14137,N_13880,N_13797);
xnor U14138 (N_14138,N_13880,N_13837);
and U14139 (N_14139,N_13957,N_13771);
or U14140 (N_14140,N_13933,N_13902);
and U14141 (N_14141,N_13917,N_13827);
or U14142 (N_14142,N_13773,N_13973);
xor U14143 (N_14143,N_13807,N_13976);
and U14144 (N_14144,N_13770,N_13792);
xnor U14145 (N_14145,N_13763,N_13956);
and U14146 (N_14146,N_13799,N_13918);
xor U14147 (N_14147,N_13888,N_13864);
nor U14148 (N_14148,N_13828,N_13930);
xnor U14149 (N_14149,N_13946,N_13919);
or U14150 (N_14150,N_13923,N_13864);
nand U14151 (N_14151,N_13996,N_13752);
and U14152 (N_14152,N_13790,N_13817);
nand U14153 (N_14153,N_13985,N_13769);
and U14154 (N_14154,N_13922,N_13928);
xor U14155 (N_14155,N_13881,N_13891);
nor U14156 (N_14156,N_13926,N_13862);
xnor U14157 (N_14157,N_13967,N_13837);
or U14158 (N_14158,N_13765,N_13953);
and U14159 (N_14159,N_13788,N_13841);
xnor U14160 (N_14160,N_13925,N_13915);
and U14161 (N_14161,N_13968,N_13941);
xor U14162 (N_14162,N_13805,N_13981);
nand U14163 (N_14163,N_13789,N_13835);
nand U14164 (N_14164,N_13998,N_13762);
and U14165 (N_14165,N_13826,N_13836);
nor U14166 (N_14166,N_13867,N_13798);
nor U14167 (N_14167,N_13900,N_13854);
nor U14168 (N_14168,N_13863,N_13838);
and U14169 (N_14169,N_13868,N_13877);
nand U14170 (N_14170,N_13803,N_13768);
nand U14171 (N_14171,N_13794,N_13827);
nor U14172 (N_14172,N_13876,N_13795);
nor U14173 (N_14173,N_13777,N_13807);
or U14174 (N_14174,N_13944,N_13812);
or U14175 (N_14175,N_13927,N_13837);
or U14176 (N_14176,N_13881,N_13829);
nor U14177 (N_14177,N_13874,N_13877);
nand U14178 (N_14178,N_13879,N_13909);
nand U14179 (N_14179,N_13975,N_13764);
nor U14180 (N_14180,N_13986,N_13846);
nor U14181 (N_14181,N_13978,N_13761);
or U14182 (N_14182,N_13817,N_13915);
xor U14183 (N_14183,N_13984,N_13977);
nor U14184 (N_14184,N_13977,N_13997);
nor U14185 (N_14185,N_13949,N_13827);
nand U14186 (N_14186,N_13958,N_13908);
nor U14187 (N_14187,N_13800,N_13852);
and U14188 (N_14188,N_13836,N_13916);
or U14189 (N_14189,N_13874,N_13996);
nor U14190 (N_14190,N_13766,N_13997);
xnor U14191 (N_14191,N_13959,N_13889);
and U14192 (N_14192,N_13808,N_13818);
xnor U14193 (N_14193,N_13962,N_13778);
nor U14194 (N_14194,N_13838,N_13869);
nand U14195 (N_14195,N_13793,N_13917);
nor U14196 (N_14196,N_13927,N_13771);
nand U14197 (N_14197,N_13993,N_13957);
or U14198 (N_14198,N_13771,N_13969);
nor U14199 (N_14199,N_13973,N_13881);
nand U14200 (N_14200,N_13906,N_13956);
nand U14201 (N_14201,N_13992,N_13872);
nor U14202 (N_14202,N_13768,N_13964);
nand U14203 (N_14203,N_13980,N_13978);
nor U14204 (N_14204,N_13967,N_13788);
xnor U14205 (N_14205,N_13843,N_13801);
xnor U14206 (N_14206,N_13759,N_13987);
or U14207 (N_14207,N_13774,N_13962);
xor U14208 (N_14208,N_13848,N_13792);
nor U14209 (N_14209,N_13949,N_13966);
nand U14210 (N_14210,N_13907,N_13757);
nor U14211 (N_14211,N_13754,N_13910);
nand U14212 (N_14212,N_13791,N_13940);
nand U14213 (N_14213,N_13927,N_13795);
or U14214 (N_14214,N_13929,N_13885);
nand U14215 (N_14215,N_13872,N_13789);
and U14216 (N_14216,N_13862,N_13997);
and U14217 (N_14217,N_13941,N_13917);
xor U14218 (N_14218,N_13886,N_13792);
and U14219 (N_14219,N_13802,N_13940);
or U14220 (N_14220,N_13832,N_13937);
nand U14221 (N_14221,N_13827,N_13923);
xnor U14222 (N_14222,N_13858,N_13754);
nand U14223 (N_14223,N_13919,N_13768);
nor U14224 (N_14224,N_13835,N_13761);
and U14225 (N_14225,N_13833,N_13809);
nor U14226 (N_14226,N_13779,N_13987);
xor U14227 (N_14227,N_13980,N_13856);
or U14228 (N_14228,N_13860,N_13941);
nor U14229 (N_14229,N_13989,N_13834);
nand U14230 (N_14230,N_13943,N_13777);
and U14231 (N_14231,N_13885,N_13989);
or U14232 (N_14232,N_13964,N_13955);
xor U14233 (N_14233,N_13940,N_13862);
xor U14234 (N_14234,N_13984,N_13949);
and U14235 (N_14235,N_13984,N_13922);
nor U14236 (N_14236,N_13996,N_13810);
and U14237 (N_14237,N_13756,N_13978);
nand U14238 (N_14238,N_13789,N_13881);
nand U14239 (N_14239,N_13922,N_13782);
nand U14240 (N_14240,N_13756,N_13899);
nand U14241 (N_14241,N_13883,N_13895);
or U14242 (N_14242,N_13810,N_13822);
nor U14243 (N_14243,N_13778,N_13800);
or U14244 (N_14244,N_13940,N_13861);
nor U14245 (N_14245,N_13897,N_13957);
and U14246 (N_14246,N_13985,N_13842);
and U14247 (N_14247,N_13934,N_13776);
and U14248 (N_14248,N_13800,N_13938);
and U14249 (N_14249,N_13856,N_13915);
xnor U14250 (N_14250,N_14078,N_14200);
nor U14251 (N_14251,N_14069,N_14008);
xnor U14252 (N_14252,N_14033,N_14100);
nor U14253 (N_14253,N_14026,N_14139);
and U14254 (N_14254,N_14249,N_14160);
nor U14255 (N_14255,N_14117,N_14175);
xor U14256 (N_14256,N_14103,N_14131);
nand U14257 (N_14257,N_14225,N_14212);
xnor U14258 (N_14258,N_14245,N_14232);
nor U14259 (N_14259,N_14099,N_14222);
nor U14260 (N_14260,N_14165,N_14238);
and U14261 (N_14261,N_14063,N_14097);
or U14262 (N_14262,N_14211,N_14068);
or U14263 (N_14263,N_14236,N_14207);
and U14264 (N_14264,N_14040,N_14189);
xnor U14265 (N_14265,N_14151,N_14121);
nor U14266 (N_14266,N_14203,N_14176);
nor U14267 (N_14267,N_14155,N_14054);
nand U14268 (N_14268,N_14029,N_14147);
xnor U14269 (N_14269,N_14055,N_14183);
nor U14270 (N_14270,N_14142,N_14208);
or U14271 (N_14271,N_14169,N_14077);
and U14272 (N_14272,N_14116,N_14037);
nand U14273 (N_14273,N_14237,N_14000);
nand U14274 (N_14274,N_14193,N_14092);
nor U14275 (N_14275,N_14168,N_14070);
and U14276 (N_14276,N_14048,N_14133);
or U14277 (N_14277,N_14135,N_14216);
nand U14278 (N_14278,N_14170,N_14214);
xor U14279 (N_14279,N_14079,N_14132);
and U14280 (N_14280,N_14071,N_14105);
nand U14281 (N_14281,N_14039,N_14177);
xnor U14282 (N_14282,N_14095,N_14109);
nand U14283 (N_14283,N_14228,N_14190);
nand U14284 (N_14284,N_14209,N_14112);
nand U14285 (N_14285,N_14003,N_14060);
nor U14286 (N_14286,N_14015,N_14052);
nand U14287 (N_14287,N_14080,N_14223);
nand U14288 (N_14288,N_14047,N_14224);
nand U14289 (N_14289,N_14085,N_14087);
nand U14290 (N_14290,N_14102,N_14053);
and U14291 (N_14291,N_14219,N_14210);
xor U14292 (N_14292,N_14178,N_14186);
xor U14293 (N_14293,N_14127,N_14025);
and U14294 (N_14294,N_14152,N_14233);
nand U14295 (N_14295,N_14042,N_14050);
and U14296 (N_14296,N_14202,N_14199);
and U14297 (N_14297,N_14163,N_14019);
or U14298 (N_14298,N_14018,N_14240);
nor U14299 (N_14299,N_14179,N_14197);
xnor U14300 (N_14300,N_14130,N_14090);
nor U14301 (N_14301,N_14011,N_14017);
nor U14302 (N_14302,N_14234,N_14196);
nor U14303 (N_14303,N_14122,N_14198);
and U14304 (N_14304,N_14049,N_14098);
or U14305 (N_14305,N_14062,N_14158);
and U14306 (N_14306,N_14192,N_14072);
nand U14307 (N_14307,N_14156,N_14213);
or U14308 (N_14308,N_14244,N_14243);
xor U14309 (N_14309,N_14084,N_14154);
nor U14310 (N_14310,N_14144,N_14138);
nor U14311 (N_14311,N_14114,N_14164);
xor U14312 (N_14312,N_14174,N_14067);
or U14313 (N_14313,N_14239,N_14023);
xnor U14314 (N_14314,N_14153,N_14137);
nand U14315 (N_14315,N_14009,N_14065);
nand U14316 (N_14316,N_14016,N_14043);
nand U14317 (N_14317,N_14013,N_14076);
xnor U14318 (N_14318,N_14027,N_14088);
or U14319 (N_14319,N_14229,N_14094);
xnor U14320 (N_14320,N_14188,N_14045);
or U14321 (N_14321,N_14075,N_14184);
nand U14322 (N_14322,N_14024,N_14226);
nand U14323 (N_14323,N_14206,N_14231);
nand U14324 (N_14324,N_14036,N_14205);
xor U14325 (N_14325,N_14056,N_14248);
nand U14326 (N_14326,N_14140,N_14118);
nor U14327 (N_14327,N_14246,N_14126);
and U14328 (N_14328,N_14031,N_14157);
nor U14329 (N_14329,N_14012,N_14066);
nand U14330 (N_14330,N_14217,N_14150);
or U14331 (N_14331,N_14161,N_14180);
or U14332 (N_14332,N_14030,N_14107);
nor U14333 (N_14333,N_14093,N_14082);
nand U14334 (N_14334,N_14104,N_14001);
or U14335 (N_14335,N_14218,N_14032);
or U14336 (N_14336,N_14145,N_14086);
nand U14337 (N_14337,N_14124,N_14064);
nor U14338 (N_14338,N_14091,N_14148);
nor U14339 (N_14339,N_14215,N_14021);
or U14340 (N_14340,N_14046,N_14081);
nand U14341 (N_14341,N_14007,N_14096);
and U14342 (N_14342,N_14204,N_14182);
nand U14343 (N_14343,N_14172,N_14187);
nand U14344 (N_14344,N_14166,N_14073);
and U14345 (N_14345,N_14028,N_14120);
nor U14346 (N_14346,N_14167,N_14235);
or U14347 (N_14347,N_14241,N_14201);
or U14348 (N_14348,N_14162,N_14128);
and U14349 (N_14349,N_14220,N_14041);
or U14350 (N_14350,N_14185,N_14113);
or U14351 (N_14351,N_14242,N_14221);
xor U14352 (N_14352,N_14141,N_14195);
and U14353 (N_14353,N_14074,N_14171);
or U14354 (N_14354,N_14181,N_14110);
nor U14355 (N_14355,N_14010,N_14006);
xor U14356 (N_14356,N_14038,N_14134);
nor U14357 (N_14357,N_14111,N_14125);
nand U14358 (N_14358,N_14020,N_14083);
nor U14359 (N_14359,N_14159,N_14101);
xor U14360 (N_14360,N_14227,N_14146);
xor U14361 (N_14361,N_14035,N_14143);
nand U14362 (N_14362,N_14014,N_14058);
and U14363 (N_14363,N_14061,N_14005);
or U14364 (N_14364,N_14089,N_14059);
nand U14365 (N_14365,N_14191,N_14051);
and U14366 (N_14366,N_14106,N_14123);
nor U14367 (N_14367,N_14108,N_14136);
xor U14368 (N_14368,N_14194,N_14004);
or U14369 (N_14369,N_14119,N_14129);
or U14370 (N_14370,N_14247,N_14057);
nor U14371 (N_14371,N_14034,N_14044);
and U14372 (N_14372,N_14022,N_14002);
xor U14373 (N_14373,N_14173,N_14230);
nor U14374 (N_14374,N_14149,N_14115);
nand U14375 (N_14375,N_14194,N_14201);
xnor U14376 (N_14376,N_14074,N_14172);
and U14377 (N_14377,N_14220,N_14016);
nor U14378 (N_14378,N_14175,N_14249);
or U14379 (N_14379,N_14044,N_14075);
xnor U14380 (N_14380,N_14194,N_14203);
nand U14381 (N_14381,N_14035,N_14174);
or U14382 (N_14382,N_14194,N_14164);
or U14383 (N_14383,N_14133,N_14049);
and U14384 (N_14384,N_14165,N_14030);
xor U14385 (N_14385,N_14110,N_14204);
xor U14386 (N_14386,N_14204,N_14146);
xor U14387 (N_14387,N_14228,N_14050);
and U14388 (N_14388,N_14106,N_14034);
or U14389 (N_14389,N_14055,N_14152);
nor U14390 (N_14390,N_14039,N_14063);
nor U14391 (N_14391,N_14203,N_14216);
nor U14392 (N_14392,N_14043,N_14081);
xnor U14393 (N_14393,N_14035,N_14214);
nand U14394 (N_14394,N_14211,N_14223);
and U14395 (N_14395,N_14033,N_14193);
and U14396 (N_14396,N_14148,N_14009);
and U14397 (N_14397,N_14034,N_14012);
xnor U14398 (N_14398,N_14029,N_14007);
nor U14399 (N_14399,N_14063,N_14157);
or U14400 (N_14400,N_14031,N_14124);
or U14401 (N_14401,N_14049,N_14190);
nand U14402 (N_14402,N_14133,N_14038);
nand U14403 (N_14403,N_14043,N_14222);
and U14404 (N_14404,N_14091,N_14016);
xnor U14405 (N_14405,N_14239,N_14177);
and U14406 (N_14406,N_14005,N_14101);
or U14407 (N_14407,N_14151,N_14170);
xnor U14408 (N_14408,N_14116,N_14170);
nor U14409 (N_14409,N_14116,N_14006);
nand U14410 (N_14410,N_14094,N_14091);
or U14411 (N_14411,N_14007,N_14210);
xor U14412 (N_14412,N_14131,N_14140);
and U14413 (N_14413,N_14048,N_14064);
and U14414 (N_14414,N_14053,N_14233);
or U14415 (N_14415,N_14194,N_14086);
and U14416 (N_14416,N_14034,N_14023);
nand U14417 (N_14417,N_14232,N_14001);
and U14418 (N_14418,N_14166,N_14181);
xor U14419 (N_14419,N_14009,N_14167);
nor U14420 (N_14420,N_14036,N_14022);
nand U14421 (N_14421,N_14185,N_14053);
and U14422 (N_14422,N_14112,N_14171);
nor U14423 (N_14423,N_14231,N_14112);
and U14424 (N_14424,N_14061,N_14112);
nand U14425 (N_14425,N_14104,N_14118);
or U14426 (N_14426,N_14128,N_14218);
and U14427 (N_14427,N_14176,N_14093);
xor U14428 (N_14428,N_14115,N_14130);
nor U14429 (N_14429,N_14082,N_14142);
and U14430 (N_14430,N_14141,N_14139);
xor U14431 (N_14431,N_14045,N_14174);
nor U14432 (N_14432,N_14244,N_14221);
or U14433 (N_14433,N_14081,N_14102);
and U14434 (N_14434,N_14008,N_14180);
xor U14435 (N_14435,N_14210,N_14224);
and U14436 (N_14436,N_14117,N_14156);
xor U14437 (N_14437,N_14175,N_14204);
nor U14438 (N_14438,N_14003,N_14151);
nand U14439 (N_14439,N_14006,N_14076);
xor U14440 (N_14440,N_14015,N_14070);
and U14441 (N_14441,N_14022,N_14228);
or U14442 (N_14442,N_14138,N_14133);
nand U14443 (N_14443,N_14051,N_14211);
and U14444 (N_14444,N_14049,N_14079);
and U14445 (N_14445,N_14070,N_14114);
and U14446 (N_14446,N_14139,N_14150);
or U14447 (N_14447,N_14054,N_14154);
and U14448 (N_14448,N_14094,N_14112);
or U14449 (N_14449,N_14136,N_14021);
or U14450 (N_14450,N_14201,N_14246);
and U14451 (N_14451,N_14139,N_14014);
nand U14452 (N_14452,N_14248,N_14110);
nor U14453 (N_14453,N_14096,N_14197);
nand U14454 (N_14454,N_14084,N_14249);
nand U14455 (N_14455,N_14058,N_14070);
xnor U14456 (N_14456,N_14119,N_14120);
xnor U14457 (N_14457,N_14071,N_14070);
or U14458 (N_14458,N_14238,N_14176);
nand U14459 (N_14459,N_14142,N_14027);
xor U14460 (N_14460,N_14056,N_14117);
xnor U14461 (N_14461,N_14128,N_14013);
nor U14462 (N_14462,N_14142,N_14103);
xnor U14463 (N_14463,N_14149,N_14215);
nor U14464 (N_14464,N_14200,N_14129);
nand U14465 (N_14465,N_14071,N_14205);
nand U14466 (N_14466,N_14058,N_14101);
xnor U14467 (N_14467,N_14032,N_14182);
nand U14468 (N_14468,N_14232,N_14010);
nand U14469 (N_14469,N_14164,N_14206);
or U14470 (N_14470,N_14113,N_14131);
and U14471 (N_14471,N_14193,N_14211);
or U14472 (N_14472,N_14099,N_14162);
nor U14473 (N_14473,N_14043,N_14205);
or U14474 (N_14474,N_14219,N_14186);
xor U14475 (N_14475,N_14185,N_14196);
nand U14476 (N_14476,N_14126,N_14152);
nor U14477 (N_14477,N_14235,N_14059);
xnor U14478 (N_14478,N_14088,N_14170);
nand U14479 (N_14479,N_14181,N_14119);
xor U14480 (N_14480,N_14031,N_14029);
and U14481 (N_14481,N_14241,N_14062);
xor U14482 (N_14482,N_14216,N_14166);
xnor U14483 (N_14483,N_14214,N_14024);
nand U14484 (N_14484,N_14175,N_14074);
nor U14485 (N_14485,N_14033,N_14141);
nand U14486 (N_14486,N_14243,N_14053);
nor U14487 (N_14487,N_14172,N_14246);
nor U14488 (N_14488,N_14180,N_14115);
nor U14489 (N_14489,N_14240,N_14097);
and U14490 (N_14490,N_14145,N_14166);
xnor U14491 (N_14491,N_14223,N_14096);
nor U14492 (N_14492,N_14158,N_14247);
or U14493 (N_14493,N_14229,N_14080);
or U14494 (N_14494,N_14140,N_14066);
nand U14495 (N_14495,N_14225,N_14067);
and U14496 (N_14496,N_14058,N_14025);
xnor U14497 (N_14497,N_14038,N_14186);
nand U14498 (N_14498,N_14169,N_14196);
and U14499 (N_14499,N_14103,N_14106);
xnor U14500 (N_14500,N_14359,N_14374);
and U14501 (N_14501,N_14390,N_14490);
or U14502 (N_14502,N_14260,N_14413);
and U14503 (N_14503,N_14325,N_14278);
nand U14504 (N_14504,N_14453,N_14371);
and U14505 (N_14505,N_14481,N_14259);
nand U14506 (N_14506,N_14311,N_14312);
or U14507 (N_14507,N_14298,N_14488);
nor U14508 (N_14508,N_14435,N_14433);
or U14509 (N_14509,N_14286,N_14428);
and U14510 (N_14510,N_14302,N_14262);
nor U14511 (N_14511,N_14405,N_14256);
nor U14512 (N_14512,N_14354,N_14279);
or U14513 (N_14513,N_14448,N_14295);
nand U14514 (N_14514,N_14261,N_14389);
nand U14515 (N_14515,N_14330,N_14436);
nor U14516 (N_14516,N_14459,N_14446);
and U14517 (N_14517,N_14494,N_14255);
xnor U14518 (N_14518,N_14417,N_14482);
nor U14519 (N_14519,N_14420,N_14414);
nor U14520 (N_14520,N_14331,N_14437);
and U14521 (N_14521,N_14299,N_14444);
or U14522 (N_14522,N_14442,N_14336);
nor U14523 (N_14523,N_14333,N_14409);
and U14524 (N_14524,N_14328,N_14427);
and U14525 (N_14525,N_14268,N_14475);
and U14526 (N_14526,N_14408,N_14407);
and U14527 (N_14527,N_14350,N_14252);
and U14528 (N_14528,N_14308,N_14347);
nor U14529 (N_14529,N_14309,N_14339);
xnor U14530 (N_14530,N_14478,N_14426);
and U14531 (N_14531,N_14382,N_14440);
nor U14532 (N_14532,N_14445,N_14467);
nand U14533 (N_14533,N_14460,N_14289);
and U14534 (N_14534,N_14280,N_14424);
xor U14535 (N_14535,N_14285,N_14380);
or U14536 (N_14536,N_14469,N_14304);
or U14537 (N_14537,N_14434,N_14348);
or U14538 (N_14538,N_14265,N_14411);
nand U14539 (N_14539,N_14361,N_14263);
xnor U14540 (N_14540,N_14257,N_14485);
nand U14541 (N_14541,N_14476,N_14355);
nand U14542 (N_14542,N_14270,N_14332);
nor U14543 (N_14543,N_14345,N_14383);
nand U14544 (N_14544,N_14254,N_14432);
nand U14545 (N_14545,N_14277,N_14313);
xnor U14546 (N_14546,N_14296,N_14416);
nor U14547 (N_14547,N_14441,N_14321);
nor U14548 (N_14548,N_14492,N_14470);
nor U14549 (N_14549,N_14378,N_14474);
or U14550 (N_14550,N_14461,N_14439);
nand U14551 (N_14551,N_14370,N_14293);
nand U14552 (N_14552,N_14497,N_14449);
nor U14553 (N_14553,N_14307,N_14375);
and U14554 (N_14554,N_14366,N_14360);
and U14555 (N_14555,N_14362,N_14396);
and U14556 (N_14556,N_14251,N_14399);
nor U14557 (N_14557,N_14406,N_14334);
or U14558 (N_14558,N_14338,N_14337);
or U14559 (N_14559,N_14275,N_14273);
xnor U14560 (N_14560,N_14479,N_14466);
nand U14561 (N_14561,N_14316,N_14326);
nand U14562 (N_14562,N_14281,N_14342);
nor U14563 (N_14563,N_14391,N_14465);
xnor U14564 (N_14564,N_14372,N_14463);
or U14565 (N_14565,N_14305,N_14471);
or U14566 (N_14566,N_14423,N_14294);
xnor U14567 (N_14567,N_14450,N_14357);
or U14568 (N_14568,N_14454,N_14292);
xor U14569 (N_14569,N_14329,N_14341);
nor U14570 (N_14570,N_14272,N_14468);
xor U14571 (N_14571,N_14395,N_14483);
and U14572 (N_14572,N_14319,N_14384);
or U14573 (N_14573,N_14353,N_14335);
and U14574 (N_14574,N_14421,N_14376);
nor U14575 (N_14575,N_14373,N_14431);
and U14576 (N_14576,N_14499,N_14397);
nor U14577 (N_14577,N_14303,N_14356);
nand U14578 (N_14578,N_14266,N_14317);
xor U14579 (N_14579,N_14318,N_14379);
xnor U14580 (N_14580,N_14377,N_14425);
nor U14581 (N_14581,N_14352,N_14264);
and U14582 (N_14582,N_14402,N_14394);
nor U14583 (N_14583,N_14415,N_14443);
and U14584 (N_14584,N_14323,N_14287);
nor U14585 (N_14585,N_14472,N_14403);
and U14586 (N_14586,N_14346,N_14457);
nor U14587 (N_14587,N_14487,N_14498);
nand U14588 (N_14588,N_14267,N_14269);
nor U14589 (N_14589,N_14343,N_14340);
and U14590 (N_14590,N_14363,N_14327);
or U14591 (N_14591,N_14400,N_14282);
and U14592 (N_14592,N_14284,N_14410);
and U14593 (N_14593,N_14388,N_14392);
xor U14594 (N_14594,N_14489,N_14430);
nor U14595 (N_14595,N_14412,N_14314);
nand U14596 (N_14596,N_14451,N_14419);
nor U14597 (N_14597,N_14271,N_14456);
or U14598 (N_14598,N_14480,N_14386);
nor U14599 (N_14599,N_14253,N_14306);
and U14600 (N_14600,N_14493,N_14297);
nor U14601 (N_14601,N_14369,N_14365);
and U14602 (N_14602,N_14300,N_14250);
nor U14603 (N_14603,N_14322,N_14422);
nor U14604 (N_14604,N_14447,N_14404);
nand U14605 (N_14605,N_14452,N_14368);
or U14606 (N_14606,N_14315,N_14484);
or U14607 (N_14607,N_14344,N_14393);
nand U14608 (N_14608,N_14349,N_14418);
nand U14609 (N_14609,N_14486,N_14274);
nor U14610 (N_14610,N_14320,N_14367);
nand U14611 (N_14611,N_14496,N_14301);
xnor U14612 (N_14612,N_14491,N_14495);
or U14613 (N_14613,N_14429,N_14438);
and U14614 (N_14614,N_14398,N_14455);
nand U14615 (N_14615,N_14381,N_14276);
nor U14616 (N_14616,N_14258,N_14464);
and U14617 (N_14617,N_14351,N_14462);
or U14618 (N_14618,N_14364,N_14473);
or U14619 (N_14619,N_14385,N_14401);
nor U14620 (N_14620,N_14458,N_14283);
xor U14621 (N_14621,N_14310,N_14291);
xnor U14622 (N_14622,N_14288,N_14324);
and U14623 (N_14623,N_14477,N_14358);
or U14624 (N_14624,N_14290,N_14387);
xor U14625 (N_14625,N_14456,N_14489);
or U14626 (N_14626,N_14439,N_14301);
or U14627 (N_14627,N_14410,N_14287);
or U14628 (N_14628,N_14453,N_14256);
nand U14629 (N_14629,N_14340,N_14327);
xor U14630 (N_14630,N_14358,N_14401);
and U14631 (N_14631,N_14486,N_14260);
nor U14632 (N_14632,N_14455,N_14349);
or U14633 (N_14633,N_14300,N_14461);
nor U14634 (N_14634,N_14439,N_14397);
and U14635 (N_14635,N_14475,N_14330);
or U14636 (N_14636,N_14267,N_14268);
or U14637 (N_14637,N_14471,N_14333);
nor U14638 (N_14638,N_14428,N_14257);
nor U14639 (N_14639,N_14346,N_14400);
or U14640 (N_14640,N_14478,N_14334);
xor U14641 (N_14641,N_14479,N_14302);
and U14642 (N_14642,N_14439,N_14295);
or U14643 (N_14643,N_14299,N_14426);
or U14644 (N_14644,N_14460,N_14454);
and U14645 (N_14645,N_14479,N_14433);
xor U14646 (N_14646,N_14398,N_14286);
and U14647 (N_14647,N_14301,N_14279);
xnor U14648 (N_14648,N_14336,N_14355);
or U14649 (N_14649,N_14488,N_14494);
xnor U14650 (N_14650,N_14484,N_14455);
or U14651 (N_14651,N_14430,N_14296);
nand U14652 (N_14652,N_14492,N_14308);
nor U14653 (N_14653,N_14294,N_14372);
nand U14654 (N_14654,N_14438,N_14497);
or U14655 (N_14655,N_14348,N_14445);
and U14656 (N_14656,N_14296,N_14441);
and U14657 (N_14657,N_14263,N_14446);
xnor U14658 (N_14658,N_14477,N_14289);
xnor U14659 (N_14659,N_14293,N_14269);
and U14660 (N_14660,N_14419,N_14349);
nand U14661 (N_14661,N_14353,N_14424);
xor U14662 (N_14662,N_14380,N_14386);
and U14663 (N_14663,N_14320,N_14281);
and U14664 (N_14664,N_14405,N_14444);
xor U14665 (N_14665,N_14317,N_14429);
nand U14666 (N_14666,N_14284,N_14260);
and U14667 (N_14667,N_14389,N_14412);
nor U14668 (N_14668,N_14257,N_14315);
or U14669 (N_14669,N_14446,N_14429);
xor U14670 (N_14670,N_14475,N_14276);
nor U14671 (N_14671,N_14254,N_14469);
nand U14672 (N_14672,N_14369,N_14292);
nor U14673 (N_14673,N_14488,N_14457);
nand U14674 (N_14674,N_14359,N_14344);
and U14675 (N_14675,N_14316,N_14364);
and U14676 (N_14676,N_14303,N_14256);
nand U14677 (N_14677,N_14348,N_14275);
nor U14678 (N_14678,N_14334,N_14397);
nor U14679 (N_14679,N_14286,N_14314);
xnor U14680 (N_14680,N_14327,N_14430);
and U14681 (N_14681,N_14447,N_14268);
nor U14682 (N_14682,N_14429,N_14282);
or U14683 (N_14683,N_14267,N_14332);
or U14684 (N_14684,N_14479,N_14312);
or U14685 (N_14685,N_14493,N_14358);
nor U14686 (N_14686,N_14317,N_14334);
nor U14687 (N_14687,N_14266,N_14479);
nand U14688 (N_14688,N_14295,N_14387);
and U14689 (N_14689,N_14438,N_14347);
nand U14690 (N_14690,N_14460,N_14438);
nor U14691 (N_14691,N_14290,N_14498);
nor U14692 (N_14692,N_14319,N_14418);
and U14693 (N_14693,N_14282,N_14369);
nor U14694 (N_14694,N_14322,N_14400);
xnor U14695 (N_14695,N_14401,N_14303);
nor U14696 (N_14696,N_14406,N_14299);
or U14697 (N_14697,N_14415,N_14282);
nor U14698 (N_14698,N_14402,N_14457);
xnor U14699 (N_14699,N_14322,N_14390);
xnor U14700 (N_14700,N_14346,N_14402);
and U14701 (N_14701,N_14462,N_14334);
nand U14702 (N_14702,N_14433,N_14281);
xor U14703 (N_14703,N_14462,N_14449);
nor U14704 (N_14704,N_14449,N_14379);
nand U14705 (N_14705,N_14458,N_14367);
and U14706 (N_14706,N_14384,N_14270);
xor U14707 (N_14707,N_14450,N_14256);
and U14708 (N_14708,N_14470,N_14474);
nand U14709 (N_14709,N_14250,N_14262);
nor U14710 (N_14710,N_14255,N_14316);
xnor U14711 (N_14711,N_14381,N_14261);
or U14712 (N_14712,N_14351,N_14412);
and U14713 (N_14713,N_14372,N_14279);
and U14714 (N_14714,N_14418,N_14366);
nand U14715 (N_14715,N_14458,N_14400);
and U14716 (N_14716,N_14279,N_14429);
nor U14717 (N_14717,N_14418,N_14423);
xnor U14718 (N_14718,N_14410,N_14440);
xnor U14719 (N_14719,N_14274,N_14367);
xnor U14720 (N_14720,N_14476,N_14389);
nor U14721 (N_14721,N_14295,N_14265);
or U14722 (N_14722,N_14406,N_14257);
or U14723 (N_14723,N_14300,N_14377);
and U14724 (N_14724,N_14494,N_14309);
nor U14725 (N_14725,N_14275,N_14332);
or U14726 (N_14726,N_14344,N_14278);
nand U14727 (N_14727,N_14307,N_14406);
nand U14728 (N_14728,N_14313,N_14407);
xnor U14729 (N_14729,N_14412,N_14305);
or U14730 (N_14730,N_14499,N_14447);
xor U14731 (N_14731,N_14447,N_14350);
and U14732 (N_14732,N_14251,N_14453);
nor U14733 (N_14733,N_14268,N_14303);
or U14734 (N_14734,N_14304,N_14445);
xnor U14735 (N_14735,N_14486,N_14424);
and U14736 (N_14736,N_14269,N_14396);
or U14737 (N_14737,N_14284,N_14328);
xnor U14738 (N_14738,N_14279,N_14472);
nor U14739 (N_14739,N_14444,N_14439);
nand U14740 (N_14740,N_14469,N_14313);
nor U14741 (N_14741,N_14417,N_14345);
and U14742 (N_14742,N_14301,N_14265);
and U14743 (N_14743,N_14286,N_14328);
xnor U14744 (N_14744,N_14410,N_14274);
or U14745 (N_14745,N_14442,N_14292);
or U14746 (N_14746,N_14436,N_14403);
and U14747 (N_14747,N_14390,N_14398);
xor U14748 (N_14748,N_14369,N_14389);
xor U14749 (N_14749,N_14399,N_14425);
nand U14750 (N_14750,N_14624,N_14721);
nand U14751 (N_14751,N_14530,N_14699);
nand U14752 (N_14752,N_14563,N_14610);
nor U14753 (N_14753,N_14550,N_14510);
nor U14754 (N_14754,N_14564,N_14640);
nand U14755 (N_14755,N_14566,N_14526);
xor U14756 (N_14756,N_14677,N_14691);
or U14757 (N_14757,N_14647,N_14690);
nor U14758 (N_14758,N_14710,N_14614);
nand U14759 (N_14759,N_14725,N_14688);
xor U14760 (N_14760,N_14709,N_14592);
or U14761 (N_14761,N_14649,N_14637);
and U14762 (N_14762,N_14500,N_14621);
nor U14763 (N_14763,N_14532,N_14558);
and U14764 (N_14764,N_14515,N_14533);
xor U14765 (N_14765,N_14713,N_14626);
xor U14766 (N_14766,N_14574,N_14598);
or U14767 (N_14767,N_14737,N_14731);
nand U14768 (N_14768,N_14569,N_14527);
nor U14769 (N_14769,N_14738,N_14539);
nor U14770 (N_14770,N_14501,N_14745);
nor U14771 (N_14771,N_14589,N_14584);
or U14772 (N_14772,N_14580,N_14565);
nand U14773 (N_14773,N_14702,N_14664);
and U14774 (N_14774,N_14572,N_14720);
or U14775 (N_14775,N_14541,N_14612);
nor U14776 (N_14776,N_14605,N_14680);
nand U14777 (N_14777,N_14726,N_14601);
xor U14778 (N_14778,N_14519,N_14682);
xnor U14779 (N_14779,N_14512,N_14553);
nor U14780 (N_14780,N_14525,N_14537);
nand U14781 (N_14781,N_14613,N_14559);
and U14782 (N_14782,N_14562,N_14704);
nor U14783 (N_14783,N_14585,N_14668);
or U14784 (N_14784,N_14618,N_14590);
nand U14785 (N_14785,N_14687,N_14703);
nand U14786 (N_14786,N_14607,N_14744);
or U14787 (N_14787,N_14623,N_14528);
xnor U14788 (N_14788,N_14746,N_14718);
or U14789 (N_14789,N_14735,N_14535);
xor U14790 (N_14790,N_14659,N_14648);
nor U14791 (N_14791,N_14676,N_14685);
xnor U14792 (N_14792,N_14520,N_14638);
and U14793 (N_14793,N_14663,N_14657);
xor U14794 (N_14794,N_14599,N_14724);
nand U14795 (N_14795,N_14579,N_14554);
and U14796 (N_14796,N_14741,N_14630);
nor U14797 (N_14797,N_14555,N_14705);
xnor U14798 (N_14798,N_14567,N_14634);
and U14799 (N_14799,N_14595,N_14549);
and U14800 (N_14800,N_14672,N_14739);
nor U14801 (N_14801,N_14723,N_14669);
and U14802 (N_14802,N_14692,N_14608);
or U14803 (N_14803,N_14671,N_14665);
or U14804 (N_14804,N_14701,N_14653);
or U14805 (N_14805,N_14674,N_14708);
nor U14806 (N_14806,N_14543,N_14587);
xor U14807 (N_14807,N_14611,N_14700);
nand U14808 (N_14808,N_14606,N_14749);
and U14809 (N_14809,N_14732,N_14716);
nor U14810 (N_14810,N_14728,N_14670);
xnor U14811 (N_14811,N_14593,N_14586);
or U14812 (N_14812,N_14531,N_14714);
nand U14813 (N_14813,N_14652,N_14570);
xnor U14814 (N_14814,N_14523,N_14517);
or U14815 (N_14815,N_14508,N_14568);
nor U14816 (N_14816,N_14748,N_14667);
or U14817 (N_14817,N_14609,N_14678);
and U14818 (N_14818,N_14552,N_14706);
nand U14819 (N_14819,N_14662,N_14518);
nand U14820 (N_14820,N_14645,N_14521);
or U14821 (N_14821,N_14711,N_14506);
xnor U14822 (N_14822,N_14502,N_14628);
nand U14823 (N_14823,N_14529,N_14734);
nand U14824 (N_14824,N_14597,N_14602);
nor U14825 (N_14825,N_14505,N_14542);
nand U14826 (N_14826,N_14636,N_14620);
nand U14827 (N_14827,N_14666,N_14696);
nand U14828 (N_14828,N_14644,N_14646);
nand U14829 (N_14829,N_14684,N_14615);
nand U14830 (N_14830,N_14722,N_14536);
xor U14831 (N_14831,N_14582,N_14681);
nand U14832 (N_14832,N_14576,N_14651);
nor U14833 (N_14833,N_14715,N_14573);
nor U14834 (N_14834,N_14504,N_14600);
nor U14835 (N_14835,N_14633,N_14643);
xnor U14836 (N_14836,N_14509,N_14740);
nor U14837 (N_14837,N_14547,N_14544);
xor U14838 (N_14838,N_14712,N_14571);
nand U14839 (N_14839,N_14503,N_14560);
and U14840 (N_14840,N_14743,N_14660);
nand U14841 (N_14841,N_14603,N_14689);
nand U14842 (N_14842,N_14551,N_14686);
and U14843 (N_14843,N_14742,N_14727);
xor U14844 (N_14844,N_14673,N_14516);
nand U14845 (N_14845,N_14588,N_14694);
nand U14846 (N_14846,N_14654,N_14575);
or U14847 (N_14847,N_14683,N_14733);
xor U14848 (N_14848,N_14545,N_14635);
or U14849 (N_14849,N_14534,N_14629);
and U14850 (N_14850,N_14578,N_14679);
or U14851 (N_14851,N_14707,N_14658);
nand U14852 (N_14852,N_14507,N_14693);
or U14853 (N_14853,N_14619,N_14729);
nand U14854 (N_14854,N_14675,N_14594);
and U14855 (N_14855,N_14538,N_14514);
and U14856 (N_14856,N_14522,N_14540);
xor U14857 (N_14857,N_14511,N_14730);
or U14858 (N_14858,N_14639,N_14632);
or U14859 (N_14859,N_14697,N_14561);
nor U14860 (N_14860,N_14642,N_14524);
and U14861 (N_14861,N_14546,N_14581);
nand U14862 (N_14862,N_14604,N_14577);
xor U14863 (N_14863,N_14596,N_14641);
xor U14864 (N_14864,N_14661,N_14513);
or U14865 (N_14865,N_14719,N_14698);
nand U14866 (N_14866,N_14622,N_14695);
nor U14867 (N_14867,N_14616,N_14548);
nor U14868 (N_14868,N_14650,N_14583);
xnor U14869 (N_14869,N_14617,N_14557);
nand U14870 (N_14870,N_14736,N_14655);
nor U14871 (N_14871,N_14627,N_14556);
and U14872 (N_14872,N_14747,N_14717);
nor U14873 (N_14873,N_14631,N_14591);
or U14874 (N_14874,N_14625,N_14656);
xor U14875 (N_14875,N_14726,N_14524);
xnor U14876 (N_14876,N_14510,N_14606);
and U14877 (N_14877,N_14725,N_14691);
and U14878 (N_14878,N_14651,N_14584);
and U14879 (N_14879,N_14679,N_14632);
or U14880 (N_14880,N_14616,N_14679);
and U14881 (N_14881,N_14572,N_14739);
and U14882 (N_14882,N_14549,N_14527);
xor U14883 (N_14883,N_14573,N_14724);
xnor U14884 (N_14884,N_14654,N_14557);
and U14885 (N_14885,N_14692,N_14587);
or U14886 (N_14886,N_14675,N_14530);
nor U14887 (N_14887,N_14733,N_14628);
and U14888 (N_14888,N_14702,N_14563);
and U14889 (N_14889,N_14730,N_14634);
or U14890 (N_14890,N_14530,N_14736);
or U14891 (N_14891,N_14688,N_14591);
xor U14892 (N_14892,N_14674,N_14614);
or U14893 (N_14893,N_14536,N_14743);
and U14894 (N_14894,N_14615,N_14591);
and U14895 (N_14895,N_14554,N_14589);
xor U14896 (N_14896,N_14741,N_14602);
or U14897 (N_14897,N_14721,N_14574);
or U14898 (N_14898,N_14665,N_14560);
nand U14899 (N_14899,N_14640,N_14567);
or U14900 (N_14900,N_14688,N_14716);
xnor U14901 (N_14901,N_14679,N_14696);
or U14902 (N_14902,N_14743,N_14692);
xnor U14903 (N_14903,N_14504,N_14598);
xnor U14904 (N_14904,N_14551,N_14652);
nor U14905 (N_14905,N_14709,N_14726);
nor U14906 (N_14906,N_14651,N_14600);
nor U14907 (N_14907,N_14600,N_14560);
and U14908 (N_14908,N_14596,N_14734);
or U14909 (N_14909,N_14733,N_14651);
nand U14910 (N_14910,N_14580,N_14518);
nand U14911 (N_14911,N_14515,N_14615);
nand U14912 (N_14912,N_14628,N_14708);
or U14913 (N_14913,N_14632,N_14671);
nand U14914 (N_14914,N_14601,N_14725);
xnor U14915 (N_14915,N_14639,N_14502);
and U14916 (N_14916,N_14719,N_14713);
and U14917 (N_14917,N_14649,N_14616);
or U14918 (N_14918,N_14741,N_14582);
or U14919 (N_14919,N_14602,N_14533);
xnor U14920 (N_14920,N_14737,N_14614);
and U14921 (N_14921,N_14553,N_14526);
or U14922 (N_14922,N_14644,N_14563);
and U14923 (N_14923,N_14612,N_14672);
or U14924 (N_14924,N_14517,N_14616);
and U14925 (N_14925,N_14585,N_14638);
nand U14926 (N_14926,N_14512,N_14745);
nor U14927 (N_14927,N_14544,N_14643);
or U14928 (N_14928,N_14681,N_14562);
xnor U14929 (N_14929,N_14613,N_14652);
xnor U14930 (N_14930,N_14526,N_14503);
and U14931 (N_14931,N_14738,N_14658);
nand U14932 (N_14932,N_14608,N_14520);
or U14933 (N_14933,N_14749,N_14615);
xnor U14934 (N_14934,N_14613,N_14636);
or U14935 (N_14935,N_14716,N_14655);
nand U14936 (N_14936,N_14732,N_14518);
nand U14937 (N_14937,N_14735,N_14624);
nor U14938 (N_14938,N_14637,N_14690);
nor U14939 (N_14939,N_14512,N_14714);
and U14940 (N_14940,N_14707,N_14536);
or U14941 (N_14941,N_14681,N_14609);
nor U14942 (N_14942,N_14633,N_14551);
or U14943 (N_14943,N_14589,N_14527);
and U14944 (N_14944,N_14662,N_14729);
nand U14945 (N_14945,N_14542,N_14504);
nor U14946 (N_14946,N_14637,N_14568);
and U14947 (N_14947,N_14599,N_14637);
xnor U14948 (N_14948,N_14731,N_14722);
nand U14949 (N_14949,N_14723,N_14570);
and U14950 (N_14950,N_14714,N_14653);
nor U14951 (N_14951,N_14587,N_14524);
and U14952 (N_14952,N_14627,N_14670);
xnor U14953 (N_14953,N_14550,N_14531);
xnor U14954 (N_14954,N_14591,N_14502);
xor U14955 (N_14955,N_14589,N_14722);
and U14956 (N_14956,N_14561,N_14622);
xnor U14957 (N_14957,N_14588,N_14681);
or U14958 (N_14958,N_14616,N_14614);
or U14959 (N_14959,N_14722,N_14696);
nand U14960 (N_14960,N_14594,N_14735);
and U14961 (N_14961,N_14564,N_14740);
xor U14962 (N_14962,N_14677,N_14505);
xnor U14963 (N_14963,N_14665,N_14568);
nand U14964 (N_14964,N_14594,N_14526);
nand U14965 (N_14965,N_14509,N_14520);
and U14966 (N_14966,N_14529,N_14660);
nor U14967 (N_14967,N_14635,N_14597);
nor U14968 (N_14968,N_14668,N_14747);
xor U14969 (N_14969,N_14529,N_14512);
nand U14970 (N_14970,N_14733,N_14684);
nand U14971 (N_14971,N_14541,N_14589);
or U14972 (N_14972,N_14733,N_14719);
and U14973 (N_14973,N_14551,N_14562);
and U14974 (N_14974,N_14503,N_14580);
or U14975 (N_14975,N_14691,N_14545);
and U14976 (N_14976,N_14569,N_14506);
nand U14977 (N_14977,N_14689,N_14525);
nor U14978 (N_14978,N_14700,N_14506);
nor U14979 (N_14979,N_14586,N_14670);
or U14980 (N_14980,N_14749,N_14578);
nand U14981 (N_14981,N_14702,N_14745);
and U14982 (N_14982,N_14525,N_14663);
nor U14983 (N_14983,N_14616,N_14589);
and U14984 (N_14984,N_14609,N_14697);
or U14985 (N_14985,N_14600,N_14674);
nor U14986 (N_14986,N_14647,N_14702);
or U14987 (N_14987,N_14565,N_14670);
nand U14988 (N_14988,N_14566,N_14620);
nor U14989 (N_14989,N_14534,N_14671);
nand U14990 (N_14990,N_14608,N_14524);
or U14991 (N_14991,N_14746,N_14712);
xor U14992 (N_14992,N_14604,N_14521);
nor U14993 (N_14993,N_14558,N_14509);
and U14994 (N_14994,N_14539,N_14584);
xnor U14995 (N_14995,N_14733,N_14696);
or U14996 (N_14996,N_14747,N_14718);
nor U14997 (N_14997,N_14748,N_14665);
xor U14998 (N_14998,N_14613,N_14572);
or U14999 (N_14999,N_14699,N_14723);
nor U15000 (N_15000,N_14912,N_14976);
and U15001 (N_15001,N_14785,N_14881);
or U15002 (N_15002,N_14887,N_14791);
nand U15003 (N_15003,N_14868,N_14802);
nor U15004 (N_15004,N_14842,N_14797);
or U15005 (N_15005,N_14776,N_14767);
xnor U15006 (N_15006,N_14788,N_14898);
nor U15007 (N_15007,N_14962,N_14917);
or U15008 (N_15008,N_14759,N_14985);
xnor U15009 (N_15009,N_14941,N_14799);
and U15010 (N_15010,N_14831,N_14938);
and U15011 (N_15011,N_14943,N_14801);
xor U15012 (N_15012,N_14808,N_14890);
and U15013 (N_15013,N_14891,N_14953);
or U15014 (N_15014,N_14798,N_14841);
xor U15015 (N_15015,N_14913,N_14993);
xor U15016 (N_15016,N_14853,N_14936);
xnor U15017 (N_15017,N_14770,N_14835);
and U15018 (N_15018,N_14927,N_14821);
xor U15019 (N_15019,N_14816,N_14907);
xor U15020 (N_15020,N_14786,N_14875);
nand U15021 (N_15021,N_14889,N_14815);
xnor U15022 (N_15022,N_14870,N_14848);
nor U15023 (N_15023,N_14974,N_14935);
nor U15024 (N_15024,N_14768,N_14787);
or U15025 (N_15025,N_14897,N_14980);
xnor U15026 (N_15026,N_14924,N_14782);
and U15027 (N_15027,N_14920,N_14800);
or U15028 (N_15028,N_14990,N_14998);
nand U15029 (N_15029,N_14964,N_14901);
or U15030 (N_15030,N_14939,N_14855);
and U15031 (N_15031,N_14774,N_14928);
and U15032 (N_15032,N_14915,N_14940);
nand U15033 (N_15033,N_14858,N_14756);
and U15034 (N_15034,N_14885,N_14983);
nor U15035 (N_15035,N_14862,N_14949);
nor U15036 (N_15036,N_14869,N_14896);
nand U15037 (N_15037,N_14957,N_14878);
and U15038 (N_15038,N_14967,N_14754);
nand U15039 (N_15039,N_14804,N_14908);
xnor U15040 (N_15040,N_14981,N_14761);
nand U15041 (N_15041,N_14921,N_14773);
or U15042 (N_15042,N_14987,N_14775);
nor U15043 (N_15043,N_14795,N_14832);
or U15044 (N_15044,N_14945,N_14857);
nand U15045 (N_15045,N_14757,N_14956);
xor U15046 (N_15046,N_14966,N_14950);
nor U15047 (N_15047,N_14963,N_14982);
and U15048 (N_15048,N_14784,N_14884);
and U15049 (N_15049,N_14902,N_14766);
xnor U15050 (N_15050,N_14984,N_14805);
or U15051 (N_15051,N_14867,N_14865);
xnor U15052 (N_15052,N_14806,N_14910);
xnor U15053 (N_15053,N_14876,N_14872);
and U15054 (N_15054,N_14873,N_14899);
nor U15055 (N_15055,N_14856,N_14854);
nand U15056 (N_15056,N_14790,N_14781);
xor U15057 (N_15057,N_14929,N_14918);
and U15058 (N_15058,N_14793,N_14847);
nor U15059 (N_15059,N_14961,N_14909);
or U15060 (N_15060,N_14914,N_14783);
nand U15061 (N_15061,N_14836,N_14824);
or U15062 (N_15062,N_14792,N_14851);
xor U15063 (N_15063,N_14833,N_14978);
nand U15064 (N_15064,N_14958,N_14819);
nand U15065 (N_15065,N_14861,N_14839);
nand U15066 (N_15066,N_14871,N_14843);
xnor U15067 (N_15067,N_14944,N_14999);
nand U15068 (N_15068,N_14794,N_14825);
nand U15069 (N_15069,N_14951,N_14863);
or U15070 (N_15070,N_14762,N_14880);
xnor U15071 (N_15071,N_14903,N_14970);
and U15072 (N_15072,N_14765,N_14827);
or U15073 (N_15073,N_14779,N_14866);
nand U15074 (N_15074,N_14849,N_14769);
xnor U15075 (N_15075,N_14823,N_14763);
nand U15076 (N_15076,N_14960,N_14977);
nor U15077 (N_15077,N_14965,N_14886);
and U15078 (N_15078,N_14975,N_14826);
nor U15079 (N_15079,N_14905,N_14973);
xnor U15080 (N_15080,N_14859,N_14852);
or U15081 (N_15081,N_14932,N_14758);
xnor U15082 (N_15082,N_14994,N_14916);
and U15083 (N_15083,N_14995,N_14764);
nor U15084 (N_15084,N_14883,N_14772);
nor U15085 (N_15085,N_14971,N_14992);
or U15086 (N_15086,N_14934,N_14860);
nand U15087 (N_15087,N_14930,N_14844);
xnor U15088 (N_15088,N_14750,N_14882);
nand U15089 (N_15089,N_14879,N_14955);
or U15090 (N_15090,N_14926,N_14894);
nand U15091 (N_15091,N_14919,N_14751);
and U15092 (N_15092,N_14893,N_14755);
and U15093 (N_15093,N_14829,N_14923);
and U15094 (N_15094,N_14959,N_14947);
or U15095 (N_15095,N_14809,N_14752);
or U15096 (N_15096,N_14874,N_14771);
and U15097 (N_15097,N_14996,N_14778);
nor U15098 (N_15098,N_14972,N_14892);
xnor U15099 (N_15099,N_14952,N_14840);
or U15100 (N_15100,N_14933,N_14989);
nor U15101 (N_15101,N_14979,N_14968);
nand U15102 (N_15102,N_14906,N_14948);
xnor U15103 (N_15103,N_14997,N_14822);
xor U15104 (N_15104,N_14810,N_14937);
and U15105 (N_15105,N_14850,N_14760);
xnor U15106 (N_15106,N_14925,N_14807);
nor U15107 (N_15107,N_14900,N_14845);
xnor U15108 (N_15108,N_14812,N_14922);
nor U15109 (N_15109,N_14820,N_14814);
or U15110 (N_15110,N_14991,N_14830);
or U15111 (N_15111,N_14942,N_14818);
nand U15112 (N_15112,N_14817,N_14777);
and U15113 (N_15113,N_14904,N_14803);
nor U15114 (N_15114,N_14834,N_14837);
nand U15115 (N_15115,N_14931,N_14877);
nand U15116 (N_15116,N_14838,N_14946);
and U15117 (N_15117,N_14864,N_14811);
nor U15118 (N_15118,N_14986,N_14954);
and U15119 (N_15119,N_14828,N_14895);
xnor U15120 (N_15120,N_14888,N_14969);
nor U15121 (N_15121,N_14789,N_14813);
or U15122 (N_15122,N_14911,N_14753);
or U15123 (N_15123,N_14846,N_14796);
or U15124 (N_15124,N_14780,N_14988);
and U15125 (N_15125,N_14920,N_14949);
and U15126 (N_15126,N_14882,N_14868);
or U15127 (N_15127,N_14974,N_14878);
and U15128 (N_15128,N_14949,N_14771);
xor U15129 (N_15129,N_14969,N_14809);
nor U15130 (N_15130,N_14796,N_14857);
and U15131 (N_15131,N_14981,N_14952);
and U15132 (N_15132,N_14922,N_14896);
xor U15133 (N_15133,N_14834,N_14823);
xor U15134 (N_15134,N_14830,N_14775);
xor U15135 (N_15135,N_14871,N_14879);
xor U15136 (N_15136,N_14971,N_14940);
or U15137 (N_15137,N_14862,N_14910);
nand U15138 (N_15138,N_14766,N_14908);
nor U15139 (N_15139,N_14929,N_14864);
nand U15140 (N_15140,N_14926,N_14965);
nand U15141 (N_15141,N_14894,N_14972);
nand U15142 (N_15142,N_14916,N_14897);
or U15143 (N_15143,N_14824,N_14760);
nand U15144 (N_15144,N_14991,N_14901);
or U15145 (N_15145,N_14868,N_14937);
nand U15146 (N_15146,N_14841,N_14936);
nor U15147 (N_15147,N_14802,N_14926);
xnor U15148 (N_15148,N_14769,N_14750);
nand U15149 (N_15149,N_14875,N_14874);
and U15150 (N_15150,N_14925,N_14839);
and U15151 (N_15151,N_14835,N_14935);
or U15152 (N_15152,N_14876,N_14878);
nand U15153 (N_15153,N_14798,N_14846);
nand U15154 (N_15154,N_14999,N_14750);
xor U15155 (N_15155,N_14800,N_14998);
xnor U15156 (N_15156,N_14859,N_14991);
xnor U15157 (N_15157,N_14865,N_14881);
and U15158 (N_15158,N_14935,N_14791);
or U15159 (N_15159,N_14884,N_14775);
or U15160 (N_15160,N_14750,N_14953);
nor U15161 (N_15161,N_14954,N_14969);
and U15162 (N_15162,N_14820,N_14975);
nand U15163 (N_15163,N_14780,N_14859);
xnor U15164 (N_15164,N_14993,N_14793);
xnor U15165 (N_15165,N_14935,N_14977);
xnor U15166 (N_15166,N_14844,N_14799);
xor U15167 (N_15167,N_14897,N_14772);
or U15168 (N_15168,N_14885,N_14767);
and U15169 (N_15169,N_14894,N_14762);
or U15170 (N_15170,N_14945,N_14908);
xnor U15171 (N_15171,N_14831,N_14891);
or U15172 (N_15172,N_14900,N_14926);
nand U15173 (N_15173,N_14821,N_14912);
xnor U15174 (N_15174,N_14801,N_14818);
nand U15175 (N_15175,N_14863,N_14999);
nand U15176 (N_15176,N_14904,N_14891);
nand U15177 (N_15177,N_14934,N_14944);
xnor U15178 (N_15178,N_14794,N_14982);
nor U15179 (N_15179,N_14861,N_14901);
and U15180 (N_15180,N_14981,N_14921);
nor U15181 (N_15181,N_14756,N_14823);
and U15182 (N_15182,N_14792,N_14971);
or U15183 (N_15183,N_14962,N_14836);
nand U15184 (N_15184,N_14760,N_14770);
nor U15185 (N_15185,N_14897,N_14767);
and U15186 (N_15186,N_14954,N_14916);
xnor U15187 (N_15187,N_14767,N_14789);
nand U15188 (N_15188,N_14893,N_14889);
nand U15189 (N_15189,N_14873,N_14875);
or U15190 (N_15190,N_14771,N_14859);
xor U15191 (N_15191,N_14997,N_14952);
xor U15192 (N_15192,N_14753,N_14967);
xnor U15193 (N_15193,N_14939,N_14997);
xor U15194 (N_15194,N_14834,N_14963);
nor U15195 (N_15195,N_14923,N_14773);
nand U15196 (N_15196,N_14751,N_14777);
and U15197 (N_15197,N_14813,N_14912);
xor U15198 (N_15198,N_14801,N_14770);
nand U15199 (N_15199,N_14909,N_14875);
nand U15200 (N_15200,N_14787,N_14985);
nor U15201 (N_15201,N_14945,N_14860);
xor U15202 (N_15202,N_14814,N_14856);
nand U15203 (N_15203,N_14943,N_14937);
nor U15204 (N_15204,N_14931,N_14883);
xor U15205 (N_15205,N_14844,N_14813);
xor U15206 (N_15206,N_14849,N_14789);
or U15207 (N_15207,N_14986,N_14756);
nand U15208 (N_15208,N_14877,N_14881);
nor U15209 (N_15209,N_14937,N_14908);
or U15210 (N_15210,N_14793,N_14889);
and U15211 (N_15211,N_14905,N_14763);
nand U15212 (N_15212,N_14925,N_14763);
or U15213 (N_15213,N_14970,N_14869);
nand U15214 (N_15214,N_14859,N_14860);
nor U15215 (N_15215,N_14803,N_14823);
nand U15216 (N_15216,N_14942,N_14816);
xnor U15217 (N_15217,N_14891,N_14870);
or U15218 (N_15218,N_14921,N_14879);
or U15219 (N_15219,N_14906,N_14893);
and U15220 (N_15220,N_14915,N_14758);
nand U15221 (N_15221,N_14958,N_14955);
nor U15222 (N_15222,N_14959,N_14929);
and U15223 (N_15223,N_14805,N_14995);
or U15224 (N_15224,N_14904,N_14870);
nand U15225 (N_15225,N_14921,N_14976);
xnor U15226 (N_15226,N_14857,N_14913);
and U15227 (N_15227,N_14783,N_14879);
or U15228 (N_15228,N_14824,N_14993);
nand U15229 (N_15229,N_14860,N_14813);
nand U15230 (N_15230,N_14783,N_14837);
nand U15231 (N_15231,N_14819,N_14995);
xnor U15232 (N_15232,N_14947,N_14797);
xor U15233 (N_15233,N_14971,N_14966);
or U15234 (N_15234,N_14973,N_14953);
or U15235 (N_15235,N_14971,N_14910);
and U15236 (N_15236,N_14791,N_14842);
or U15237 (N_15237,N_14989,N_14930);
nand U15238 (N_15238,N_14825,N_14954);
nor U15239 (N_15239,N_14815,N_14931);
and U15240 (N_15240,N_14754,N_14787);
and U15241 (N_15241,N_14950,N_14972);
nand U15242 (N_15242,N_14935,N_14938);
and U15243 (N_15243,N_14817,N_14995);
xnor U15244 (N_15244,N_14953,N_14963);
xor U15245 (N_15245,N_14768,N_14751);
or U15246 (N_15246,N_14951,N_14969);
and U15247 (N_15247,N_14901,N_14916);
xnor U15248 (N_15248,N_14754,N_14912);
or U15249 (N_15249,N_14945,N_14977);
xnor U15250 (N_15250,N_15237,N_15188);
or U15251 (N_15251,N_15194,N_15078);
or U15252 (N_15252,N_15123,N_15089);
and U15253 (N_15253,N_15247,N_15139);
and U15254 (N_15254,N_15091,N_15057);
or U15255 (N_15255,N_15217,N_15054);
nand U15256 (N_15256,N_15114,N_15079);
xnor U15257 (N_15257,N_15015,N_15164);
or U15258 (N_15258,N_15056,N_15022);
nor U15259 (N_15259,N_15165,N_15147);
or U15260 (N_15260,N_15037,N_15026);
nor U15261 (N_15261,N_15021,N_15019);
nor U15262 (N_15262,N_15199,N_15209);
nor U15263 (N_15263,N_15187,N_15169);
or U15264 (N_15264,N_15096,N_15127);
or U15265 (N_15265,N_15152,N_15025);
and U15266 (N_15266,N_15016,N_15003);
nand U15267 (N_15267,N_15075,N_15062);
xnor U15268 (N_15268,N_15197,N_15102);
and U15269 (N_15269,N_15059,N_15119);
nand U15270 (N_15270,N_15125,N_15048);
nand U15271 (N_15271,N_15043,N_15185);
nand U15272 (N_15272,N_15018,N_15085);
nand U15273 (N_15273,N_15134,N_15160);
and U15274 (N_15274,N_15163,N_15131);
and U15275 (N_15275,N_15146,N_15190);
nand U15276 (N_15276,N_15007,N_15156);
nor U15277 (N_15277,N_15066,N_15176);
or U15278 (N_15278,N_15044,N_15069);
nand U15279 (N_15279,N_15162,N_15116);
and U15280 (N_15280,N_15234,N_15155);
and U15281 (N_15281,N_15099,N_15235);
nor U15282 (N_15282,N_15118,N_15236);
nand U15283 (N_15283,N_15124,N_15072);
nand U15284 (N_15284,N_15074,N_15213);
and U15285 (N_15285,N_15248,N_15142);
xor U15286 (N_15286,N_15005,N_15071);
and U15287 (N_15287,N_15231,N_15201);
and U15288 (N_15288,N_15111,N_15210);
and U15289 (N_15289,N_15204,N_15211);
nor U15290 (N_15290,N_15106,N_15101);
nor U15291 (N_15291,N_15029,N_15112);
xor U15292 (N_15292,N_15017,N_15060);
nand U15293 (N_15293,N_15203,N_15189);
nor U15294 (N_15294,N_15130,N_15088);
or U15295 (N_15295,N_15177,N_15182);
and U15296 (N_15296,N_15168,N_15157);
nand U15297 (N_15297,N_15208,N_15238);
nor U15298 (N_15298,N_15172,N_15195);
or U15299 (N_15299,N_15034,N_15100);
nand U15300 (N_15300,N_15000,N_15171);
xnor U15301 (N_15301,N_15068,N_15076);
xnor U15302 (N_15302,N_15092,N_15198);
xor U15303 (N_15303,N_15122,N_15230);
or U15304 (N_15304,N_15039,N_15178);
nand U15305 (N_15305,N_15002,N_15148);
nor U15306 (N_15306,N_15028,N_15181);
and U15307 (N_15307,N_15227,N_15240);
xor U15308 (N_15308,N_15242,N_15120);
nor U15309 (N_15309,N_15049,N_15140);
nand U15310 (N_15310,N_15086,N_15090);
or U15311 (N_15311,N_15229,N_15024);
and U15312 (N_15312,N_15035,N_15245);
nand U15313 (N_15313,N_15137,N_15202);
or U15314 (N_15314,N_15221,N_15184);
and U15315 (N_15315,N_15061,N_15226);
nand U15316 (N_15316,N_15080,N_15128);
nand U15317 (N_15317,N_15067,N_15047);
and U15318 (N_15318,N_15161,N_15232);
and U15319 (N_15319,N_15097,N_15083);
or U15320 (N_15320,N_15065,N_15023);
or U15321 (N_15321,N_15150,N_15121);
xor U15322 (N_15322,N_15225,N_15233);
nor U15323 (N_15323,N_15173,N_15045);
nor U15324 (N_15324,N_15175,N_15243);
nor U15325 (N_15325,N_15144,N_15215);
xor U15326 (N_15326,N_15108,N_15095);
nand U15327 (N_15327,N_15058,N_15212);
nand U15328 (N_15328,N_15105,N_15115);
and U15329 (N_15329,N_15192,N_15004);
nand U15330 (N_15330,N_15241,N_15170);
nor U15331 (N_15331,N_15104,N_15219);
xnor U15332 (N_15332,N_15126,N_15149);
and U15333 (N_15333,N_15031,N_15153);
and U15334 (N_15334,N_15098,N_15220);
and U15335 (N_15335,N_15081,N_15012);
nand U15336 (N_15336,N_15133,N_15216);
and U15337 (N_15337,N_15082,N_15246);
nor U15338 (N_15338,N_15143,N_15244);
nor U15339 (N_15339,N_15036,N_15214);
xnor U15340 (N_15340,N_15093,N_15151);
xnor U15341 (N_15341,N_15113,N_15135);
or U15342 (N_15342,N_15196,N_15154);
nand U15343 (N_15343,N_15046,N_15027);
nor U15344 (N_15344,N_15009,N_15013);
and U15345 (N_15345,N_15040,N_15129);
or U15346 (N_15346,N_15141,N_15200);
nor U15347 (N_15347,N_15159,N_15055);
nand U15348 (N_15348,N_15239,N_15006);
xor U15349 (N_15349,N_15052,N_15180);
nand U15350 (N_15350,N_15107,N_15020);
and U15351 (N_15351,N_15207,N_15041);
or U15352 (N_15352,N_15205,N_15145);
nand U15353 (N_15353,N_15191,N_15077);
and U15354 (N_15354,N_15064,N_15228);
xor U15355 (N_15355,N_15174,N_15073);
nor U15356 (N_15356,N_15032,N_15167);
nor U15357 (N_15357,N_15103,N_15053);
nand U15358 (N_15358,N_15038,N_15110);
or U15359 (N_15359,N_15030,N_15179);
or U15360 (N_15360,N_15050,N_15117);
nor U15361 (N_15361,N_15222,N_15087);
and U15362 (N_15362,N_15010,N_15011);
nand U15363 (N_15363,N_15132,N_15224);
and U15364 (N_15364,N_15042,N_15166);
xor U15365 (N_15365,N_15063,N_15138);
nand U15366 (N_15366,N_15218,N_15223);
or U15367 (N_15367,N_15183,N_15084);
and U15368 (N_15368,N_15008,N_15158);
nor U15369 (N_15369,N_15206,N_15001);
or U15370 (N_15370,N_15109,N_15186);
nor U15371 (N_15371,N_15136,N_15051);
or U15372 (N_15372,N_15249,N_15193);
xor U15373 (N_15373,N_15094,N_15070);
or U15374 (N_15374,N_15033,N_15014);
or U15375 (N_15375,N_15215,N_15020);
nor U15376 (N_15376,N_15064,N_15024);
nand U15377 (N_15377,N_15161,N_15123);
xnor U15378 (N_15378,N_15016,N_15095);
nand U15379 (N_15379,N_15175,N_15073);
or U15380 (N_15380,N_15096,N_15053);
xnor U15381 (N_15381,N_15168,N_15107);
xnor U15382 (N_15382,N_15177,N_15131);
or U15383 (N_15383,N_15188,N_15133);
or U15384 (N_15384,N_15140,N_15208);
and U15385 (N_15385,N_15063,N_15245);
and U15386 (N_15386,N_15032,N_15021);
nor U15387 (N_15387,N_15223,N_15190);
and U15388 (N_15388,N_15119,N_15240);
and U15389 (N_15389,N_15116,N_15221);
nand U15390 (N_15390,N_15211,N_15234);
nor U15391 (N_15391,N_15096,N_15025);
and U15392 (N_15392,N_15108,N_15116);
xnor U15393 (N_15393,N_15063,N_15057);
and U15394 (N_15394,N_15079,N_15016);
or U15395 (N_15395,N_15089,N_15025);
nor U15396 (N_15396,N_15143,N_15079);
or U15397 (N_15397,N_15207,N_15068);
nor U15398 (N_15398,N_15000,N_15110);
nand U15399 (N_15399,N_15137,N_15224);
nor U15400 (N_15400,N_15062,N_15202);
xnor U15401 (N_15401,N_15150,N_15065);
or U15402 (N_15402,N_15091,N_15150);
nand U15403 (N_15403,N_15192,N_15229);
or U15404 (N_15404,N_15037,N_15219);
or U15405 (N_15405,N_15230,N_15054);
nor U15406 (N_15406,N_15043,N_15153);
and U15407 (N_15407,N_15228,N_15128);
and U15408 (N_15408,N_15187,N_15075);
nand U15409 (N_15409,N_15015,N_15066);
or U15410 (N_15410,N_15136,N_15240);
or U15411 (N_15411,N_15058,N_15061);
nor U15412 (N_15412,N_15018,N_15130);
nor U15413 (N_15413,N_15039,N_15060);
nand U15414 (N_15414,N_15234,N_15145);
nor U15415 (N_15415,N_15023,N_15204);
and U15416 (N_15416,N_15190,N_15064);
nand U15417 (N_15417,N_15195,N_15167);
nand U15418 (N_15418,N_15244,N_15173);
nand U15419 (N_15419,N_15193,N_15001);
nand U15420 (N_15420,N_15056,N_15013);
xnor U15421 (N_15421,N_15041,N_15170);
nor U15422 (N_15422,N_15074,N_15160);
or U15423 (N_15423,N_15055,N_15244);
or U15424 (N_15424,N_15212,N_15068);
xor U15425 (N_15425,N_15103,N_15000);
and U15426 (N_15426,N_15113,N_15151);
or U15427 (N_15427,N_15221,N_15035);
nor U15428 (N_15428,N_15180,N_15201);
xor U15429 (N_15429,N_15019,N_15209);
or U15430 (N_15430,N_15024,N_15105);
xnor U15431 (N_15431,N_15139,N_15113);
nor U15432 (N_15432,N_15137,N_15059);
or U15433 (N_15433,N_15114,N_15039);
and U15434 (N_15434,N_15150,N_15141);
and U15435 (N_15435,N_15174,N_15099);
nor U15436 (N_15436,N_15241,N_15145);
nor U15437 (N_15437,N_15146,N_15157);
and U15438 (N_15438,N_15231,N_15140);
nor U15439 (N_15439,N_15176,N_15179);
and U15440 (N_15440,N_15069,N_15180);
nand U15441 (N_15441,N_15223,N_15136);
xnor U15442 (N_15442,N_15101,N_15190);
xor U15443 (N_15443,N_15004,N_15047);
xor U15444 (N_15444,N_15164,N_15222);
nand U15445 (N_15445,N_15155,N_15244);
and U15446 (N_15446,N_15119,N_15185);
and U15447 (N_15447,N_15063,N_15176);
nand U15448 (N_15448,N_15201,N_15057);
nand U15449 (N_15449,N_15151,N_15174);
and U15450 (N_15450,N_15017,N_15062);
or U15451 (N_15451,N_15008,N_15115);
nand U15452 (N_15452,N_15107,N_15016);
xor U15453 (N_15453,N_15043,N_15208);
or U15454 (N_15454,N_15147,N_15034);
or U15455 (N_15455,N_15202,N_15160);
nor U15456 (N_15456,N_15158,N_15099);
nor U15457 (N_15457,N_15104,N_15195);
and U15458 (N_15458,N_15198,N_15094);
xor U15459 (N_15459,N_15023,N_15042);
or U15460 (N_15460,N_15096,N_15026);
and U15461 (N_15461,N_15152,N_15211);
nand U15462 (N_15462,N_15037,N_15202);
xor U15463 (N_15463,N_15008,N_15098);
or U15464 (N_15464,N_15247,N_15206);
nand U15465 (N_15465,N_15232,N_15162);
nand U15466 (N_15466,N_15177,N_15039);
or U15467 (N_15467,N_15158,N_15046);
xnor U15468 (N_15468,N_15229,N_15148);
or U15469 (N_15469,N_15121,N_15102);
xnor U15470 (N_15470,N_15062,N_15107);
and U15471 (N_15471,N_15005,N_15209);
nor U15472 (N_15472,N_15142,N_15021);
nand U15473 (N_15473,N_15212,N_15172);
nand U15474 (N_15474,N_15016,N_15056);
or U15475 (N_15475,N_15020,N_15244);
nand U15476 (N_15476,N_15209,N_15196);
nor U15477 (N_15477,N_15227,N_15232);
and U15478 (N_15478,N_15159,N_15198);
nor U15479 (N_15479,N_15230,N_15026);
or U15480 (N_15480,N_15111,N_15144);
xnor U15481 (N_15481,N_15039,N_15138);
nand U15482 (N_15482,N_15038,N_15124);
or U15483 (N_15483,N_15123,N_15204);
nand U15484 (N_15484,N_15042,N_15062);
nor U15485 (N_15485,N_15004,N_15082);
nor U15486 (N_15486,N_15115,N_15011);
or U15487 (N_15487,N_15172,N_15186);
nand U15488 (N_15488,N_15167,N_15221);
nor U15489 (N_15489,N_15170,N_15001);
or U15490 (N_15490,N_15226,N_15075);
or U15491 (N_15491,N_15204,N_15075);
nor U15492 (N_15492,N_15188,N_15000);
nand U15493 (N_15493,N_15173,N_15098);
nand U15494 (N_15494,N_15048,N_15145);
nand U15495 (N_15495,N_15125,N_15244);
and U15496 (N_15496,N_15138,N_15199);
or U15497 (N_15497,N_15084,N_15247);
nand U15498 (N_15498,N_15235,N_15112);
nand U15499 (N_15499,N_15112,N_15135);
nand U15500 (N_15500,N_15482,N_15299);
or U15501 (N_15501,N_15328,N_15330);
xor U15502 (N_15502,N_15317,N_15404);
and U15503 (N_15503,N_15284,N_15322);
nor U15504 (N_15504,N_15374,N_15457);
or U15505 (N_15505,N_15495,N_15341);
nor U15506 (N_15506,N_15382,N_15309);
nand U15507 (N_15507,N_15289,N_15453);
nor U15508 (N_15508,N_15366,N_15301);
and U15509 (N_15509,N_15426,N_15261);
and U15510 (N_15510,N_15358,N_15492);
nand U15511 (N_15511,N_15427,N_15402);
xnor U15512 (N_15512,N_15323,N_15263);
nand U15513 (N_15513,N_15367,N_15296);
xor U15514 (N_15514,N_15395,N_15265);
xor U15515 (N_15515,N_15447,N_15262);
and U15516 (N_15516,N_15450,N_15472);
nor U15517 (N_15517,N_15438,N_15313);
nand U15518 (N_15518,N_15415,N_15485);
xnor U15519 (N_15519,N_15336,N_15251);
nand U15520 (N_15520,N_15459,N_15310);
nor U15521 (N_15521,N_15394,N_15344);
and U15522 (N_15522,N_15455,N_15281);
and U15523 (N_15523,N_15412,N_15362);
or U15524 (N_15524,N_15320,N_15392);
and U15525 (N_15525,N_15439,N_15399);
nand U15526 (N_15526,N_15335,N_15490);
or U15527 (N_15527,N_15274,N_15266);
or U15528 (N_15528,N_15391,N_15282);
xnor U15529 (N_15529,N_15488,N_15425);
xnor U15530 (N_15530,N_15290,N_15440);
or U15531 (N_15531,N_15496,N_15338);
nor U15532 (N_15532,N_15435,N_15396);
nor U15533 (N_15533,N_15332,N_15355);
and U15534 (N_15534,N_15304,N_15252);
xnor U15535 (N_15535,N_15291,N_15470);
and U15536 (N_15536,N_15469,N_15286);
nand U15537 (N_15537,N_15258,N_15428);
or U15538 (N_15538,N_15302,N_15321);
nor U15539 (N_15539,N_15257,N_15357);
nor U15540 (N_15540,N_15416,N_15307);
or U15541 (N_15541,N_15387,N_15297);
and U15542 (N_15542,N_15349,N_15350);
xor U15543 (N_15543,N_15292,N_15410);
nor U15544 (N_15544,N_15413,N_15390);
nor U15545 (N_15545,N_15479,N_15294);
or U15546 (N_15546,N_15456,N_15364);
or U15547 (N_15547,N_15377,N_15345);
and U15548 (N_15548,N_15471,N_15461);
nor U15549 (N_15549,N_15465,N_15444);
xor U15550 (N_15550,N_15466,N_15462);
or U15551 (N_15551,N_15422,N_15441);
and U15552 (N_15552,N_15478,N_15371);
xnor U15553 (N_15553,N_15473,N_15268);
xnor U15554 (N_15554,N_15333,N_15311);
nor U15555 (N_15555,N_15445,N_15386);
and U15556 (N_15556,N_15408,N_15474);
xnor U15557 (N_15557,N_15499,N_15365);
or U15558 (N_15558,N_15451,N_15378);
xor U15559 (N_15559,N_15475,N_15295);
xor U15560 (N_15560,N_15418,N_15405);
and U15561 (N_15561,N_15411,N_15318);
nor U15562 (N_15562,N_15273,N_15400);
and U15563 (N_15563,N_15326,N_15433);
nand U15564 (N_15564,N_15437,N_15476);
xnor U15565 (N_15565,N_15430,N_15486);
xor U15566 (N_15566,N_15305,N_15373);
xnor U15567 (N_15567,N_15385,N_15255);
and U15568 (N_15568,N_15409,N_15256);
or U15569 (N_15569,N_15325,N_15259);
or U15570 (N_15570,N_15359,N_15319);
or U15571 (N_15571,N_15340,N_15329);
or U15572 (N_15572,N_15269,N_15351);
nor U15573 (N_15573,N_15487,N_15389);
nand U15574 (N_15574,N_15327,N_15312);
nor U15575 (N_15575,N_15449,N_15452);
xor U15576 (N_15576,N_15460,N_15454);
xor U15577 (N_15577,N_15484,N_15414);
nand U15578 (N_15578,N_15431,N_15393);
nand U15579 (N_15579,N_15316,N_15489);
and U15580 (N_15580,N_15420,N_15354);
xnor U15581 (N_15581,N_15491,N_15346);
xor U15582 (N_15582,N_15343,N_15380);
nor U15583 (N_15583,N_15442,N_15370);
nor U15584 (N_15584,N_15306,N_15375);
and U15585 (N_15585,N_15353,N_15381);
and U15586 (N_15586,N_15397,N_15464);
and U15587 (N_15587,N_15436,N_15363);
and U15588 (N_15588,N_15468,N_15406);
nand U15589 (N_15589,N_15272,N_15324);
nand U15590 (N_15590,N_15264,N_15314);
nand U15591 (N_15591,N_15288,N_15497);
nand U15592 (N_15592,N_15369,N_15270);
and U15593 (N_15593,N_15432,N_15458);
and U15594 (N_15594,N_15443,N_15276);
or U15595 (N_15595,N_15379,N_15398);
xor U15596 (N_15596,N_15342,N_15275);
or U15597 (N_15597,N_15481,N_15483);
xnor U15598 (N_15598,N_15278,N_15407);
xor U15599 (N_15599,N_15494,N_15285);
nand U15600 (N_15600,N_15368,N_15421);
or U15601 (N_15601,N_15372,N_15279);
xor U15602 (N_15602,N_15348,N_15308);
or U15603 (N_15603,N_15448,N_15280);
xnor U15604 (N_15604,N_15250,N_15303);
and U15605 (N_15605,N_15352,N_15388);
xnor U15606 (N_15606,N_15477,N_15271);
or U15607 (N_15607,N_15434,N_15424);
nand U15608 (N_15608,N_15401,N_15298);
xnor U15609 (N_15609,N_15417,N_15446);
nor U15610 (N_15610,N_15498,N_15254);
or U15611 (N_15611,N_15347,N_15384);
and U15612 (N_15612,N_15361,N_15334);
xnor U15613 (N_15613,N_15376,N_15423);
xnor U15614 (N_15614,N_15293,N_15463);
or U15615 (N_15615,N_15331,N_15260);
nor U15616 (N_15616,N_15287,N_15429);
and U15617 (N_15617,N_15493,N_15356);
or U15618 (N_15618,N_15419,N_15300);
xor U15619 (N_15619,N_15360,N_15403);
nor U15620 (N_15620,N_15315,N_15339);
xnor U15621 (N_15621,N_15337,N_15253);
xnor U15622 (N_15622,N_15283,N_15277);
nor U15623 (N_15623,N_15383,N_15267);
xnor U15624 (N_15624,N_15467,N_15480);
and U15625 (N_15625,N_15442,N_15443);
nand U15626 (N_15626,N_15456,N_15266);
nor U15627 (N_15627,N_15432,N_15339);
xor U15628 (N_15628,N_15419,N_15403);
or U15629 (N_15629,N_15315,N_15384);
or U15630 (N_15630,N_15454,N_15273);
nor U15631 (N_15631,N_15443,N_15422);
xor U15632 (N_15632,N_15316,N_15458);
nor U15633 (N_15633,N_15256,N_15285);
nor U15634 (N_15634,N_15265,N_15497);
or U15635 (N_15635,N_15374,N_15268);
or U15636 (N_15636,N_15269,N_15478);
and U15637 (N_15637,N_15400,N_15478);
xor U15638 (N_15638,N_15487,N_15404);
or U15639 (N_15639,N_15301,N_15435);
xor U15640 (N_15640,N_15375,N_15451);
nor U15641 (N_15641,N_15483,N_15425);
nor U15642 (N_15642,N_15451,N_15349);
or U15643 (N_15643,N_15491,N_15362);
or U15644 (N_15644,N_15337,N_15280);
nand U15645 (N_15645,N_15344,N_15459);
and U15646 (N_15646,N_15448,N_15287);
and U15647 (N_15647,N_15388,N_15496);
xor U15648 (N_15648,N_15452,N_15263);
nor U15649 (N_15649,N_15355,N_15422);
xor U15650 (N_15650,N_15456,N_15268);
or U15651 (N_15651,N_15413,N_15416);
nand U15652 (N_15652,N_15252,N_15311);
or U15653 (N_15653,N_15492,N_15475);
nor U15654 (N_15654,N_15486,N_15326);
and U15655 (N_15655,N_15450,N_15378);
or U15656 (N_15656,N_15471,N_15333);
xor U15657 (N_15657,N_15404,N_15276);
nand U15658 (N_15658,N_15469,N_15320);
xnor U15659 (N_15659,N_15401,N_15310);
nand U15660 (N_15660,N_15357,N_15380);
nand U15661 (N_15661,N_15359,N_15310);
xor U15662 (N_15662,N_15341,N_15305);
nand U15663 (N_15663,N_15318,N_15461);
and U15664 (N_15664,N_15466,N_15315);
nor U15665 (N_15665,N_15393,N_15461);
xnor U15666 (N_15666,N_15310,N_15408);
xnor U15667 (N_15667,N_15464,N_15304);
nor U15668 (N_15668,N_15399,N_15421);
nor U15669 (N_15669,N_15455,N_15420);
nand U15670 (N_15670,N_15337,N_15250);
xnor U15671 (N_15671,N_15404,N_15285);
xnor U15672 (N_15672,N_15464,N_15396);
or U15673 (N_15673,N_15274,N_15392);
nand U15674 (N_15674,N_15471,N_15485);
xnor U15675 (N_15675,N_15354,N_15398);
nand U15676 (N_15676,N_15338,N_15498);
and U15677 (N_15677,N_15498,N_15482);
or U15678 (N_15678,N_15417,N_15442);
xor U15679 (N_15679,N_15403,N_15426);
or U15680 (N_15680,N_15282,N_15337);
or U15681 (N_15681,N_15321,N_15488);
or U15682 (N_15682,N_15322,N_15343);
nand U15683 (N_15683,N_15388,N_15367);
xnor U15684 (N_15684,N_15447,N_15389);
or U15685 (N_15685,N_15382,N_15367);
and U15686 (N_15686,N_15339,N_15430);
and U15687 (N_15687,N_15395,N_15458);
and U15688 (N_15688,N_15304,N_15317);
nand U15689 (N_15689,N_15419,N_15331);
and U15690 (N_15690,N_15445,N_15440);
or U15691 (N_15691,N_15440,N_15416);
nand U15692 (N_15692,N_15447,N_15416);
xnor U15693 (N_15693,N_15369,N_15382);
nand U15694 (N_15694,N_15256,N_15411);
and U15695 (N_15695,N_15405,N_15465);
and U15696 (N_15696,N_15252,N_15444);
nand U15697 (N_15697,N_15318,N_15297);
nor U15698 (N_15698,N_15471,N_15483);
nand U15699 (N_15699,N_15269,N_15284);
or U15700 (N_15700,N_15373,N_15387);
and U15701 (N_15701,N_15336,N_15332);
xnor U15702 (N_15702,N_15257,N_15496);
and U15703 (N_15703,N_15478,N_15341);
xnor U15704 (N_15704,N_15313,N_15317);
and U15705 (N_15705,N_15485,N_15306);
or U15706 (N_15706,N_15271,N_15423);
xor U15707 (N_15707,N_15355,N_15373);
nor U15708 (N_15708,N_15454,N_15353);
nand U15709 (N_15709,N_15333,N_15305);
xnor U15710 (N_15710,N_15473,N_15269);
xnor U15711 (N_15711,N_15485,N_15399);
or U15712 (N_15712,N_15446,N_15464);
or U15713 (N_15713,N_15416,N_15344);
and U15714 (N_15714,N_15331,N_15329);
or U15715 (N_15715,N_15456,N_15420);
xor U15716 (N_15716,N_15315,N_15430);
or U15717 (N_15717,N_15342,N_15451);
nor U15718 (N_15718,N_15385,N_15479);
nor U15719 (N_15719,N_15485,N_15433);
xor U15720 (N_15720,N_15346,N_15484);
and U15721 (N_15721,N_15431,N_15290);
nand U15722 (N_15722,N_15305,N_15298);
nand U15723 (N_15723,N_15423,N_15391);
nand U15724 (N_15724,N_15465,N_15470);
or U15725 (N_15725,N_15420,N_15372);
nor U15726 (N_15726,N_15342,N_15497);
or U15727 (N_15727,N_15356,N_15288);
nand U15728 (N_15728,N_15470,N_15460);
and U15729 (N_15729,N_15498,N_15331);
nor U15730 (N_15730,N_15358,N_15471);
or U15731 (N_15731,N_15499,N_15308);
and U15732 (N_15732,N_15437,N_15267);
or U15733 (N_15733,N_15358,N_15348);
xor U15734 (N_15734,N_15489,N_15285);
and U15735 (N_15735,N_15393,N_15410);
nor U15736 (N_15736,N_15275,N_15276);
nand U15737 (N_15737,N_15335,N_15454);
nor U15738 (N_15738,N_15431,N_15262);
or U15739 (N_15739,N_15470,N_15413);
nand U15740 (N_15740,N_15355,N_15330);
and U15741 (N_15741,N_15482,N_15378);
nand U15742 (N_15742,N_15312,N_15409);
and U15743 (N_15743,N_15380,N_15324);
or U15744 (N_15744,N_15487,N_15317);
nand U15745 (N_15745,N_15430,N_15324);
xnor U15746 (N_15746,N_15251,N_15494);
xnor U15747 (N_15747,N_15333,N_15494);
nand U15748 (N_15748,N_15274,N_15288);
or U15749 (N_15749,N_15305,N_15457);
nand U15750 (N_15750,N_15509,N_15633);
and U15751 (N_15751,N_15734,N_15507);
or U15752 (N_15752,N_15699,N_15697);
xnor U15753 (N_15753,N_15652,N_15578);
and U15754 (N_15754,N_15531,N_15516);
nor U15755 (N_15755,N_15610,N_15606);
xor U15756 (N_15756,N_15635,N_15558);
or U15757 (N_15757,N_15536,N_15736);
and U15758 (N_15758,N_15692,N_15743);
and U15759 (N_15759,N_15549,N_15664);
xor U15760 (N_15760,N_15530,N_15571);
xor U15761 (N_15761,N_15691,N_15573);
xor U15762 (N_15762,N_15534,N_15739);
nand U15763 (N_15763,N_15695,N_15658);
xor U15764 (N_15764,N_15568,N_15630);
nor U15765 (N_15765,N_15569,N_15708);
and U15766 (N_15766,N_15645,N_15532);
nor U15767 (N_15767,N_15559,N_15749);
or U15768 (N_15768,N_15628,N_15577);
nand U15769 (N_15769,N_15538,N_15727);
nand U15770 (N_15770,N_15525,N_15522);
and U15771 (N_15771,N_15563,N_15575);
nand U15772 (N_15772,N_15501,N_15683);
xor U15773 (N_15773,N_15637,N_15738);
nor U15774 (N_15774,N_15730,N_15665);
nand U15775 (N_15775,N_15662,N_15524);
nor U15776 (N_15776,N_15639,N_15580);
and U15777 (N_15777,N_15512,N_15729);
or U15778 (N_15778,N_15554,N_15718);
or U15779 (N_15779,N_15682,N_15547);
nand U15780 (N_15780,N_15616,N_15545);
nor U15781 (N_15781,N_15519,N_15688);
xnor U15782 (N_15782,N_15675,N_15701);
or U15783 (N_15783,N_15612,N_15744);
or U15784 (N_15784,N_15506,N_15614);
xor U15785 (N_15785,N_15550,N_15719);
nand U15786 (N_15786,N_15649,N_15667);
nand U15787 (N_15787,N_15587,N_15626);
and U15788 (N_15788,N_15565,N_15654);
and U15789 (N_15789,N_15712,N_15661);
nand U15790 (N_15790,N_15704,N_15663);
nor U15791 (N_15791,N_15741,N_15625);
and U15792 (N_15792,N_15540,N_15690);
nand U15793 (N_15793,N_15604,N_15732);
xor U15794 (N_15794,N_15511,N_15651);
nand U15795 (N_15795,N_15523,N_15517);
or U15796 (N_15796,N_15723,N_15609);
or U15797 (N_15797,N_15582,N_15513);
or U15798 (N_15798,N_15657,N_15647);
and U15799 (N_15799,N_15613,N_15636);
xor U15800 (N_15800,N_15684,N_15602);
nor U15801 (N_15801,N_15584,N_15505);
nand U15802 (N_15802,N_15685,N_15542);
and U15803 (N_15803,N_15728,N_15705);
or U15804 (N_15804,N_15527,N_15556);
nor U15805 (N_15805,N_15648,N_15611);
or U15806 (N_15806,N_15627,N_15555);
and U15807 (N_15807,N_15615,N_15742);
and U15808 (N_15808,N_15595,N_15557);
nand U15809 (N_15809,N_15737,N_15567);
and U15810 (N_15810,N_15521,N_15715);
nor U15811 (N_15811,N_15724,N_15735);
nand U15812 (N_15812,N_15539,N_15607);
xor U15813 (N_15813,N_15677,N_15671);
nor U15814 (N_15814,N_15552,N_15564);
and U15815 (N_15815,N_15535,N_15673);
xnor U15816 (N_15816,N_15641,N_15643);
nor U15817 (N_15817,N_15515,N_15581);
xor U15818 (N_15818,N_15709,N_15589);
and U15819 (N_15819,N_15504,N_15660);
xor U15820 (N_15820,N_15672,N_15726);
nor U15821 (N_15821,N_15676,N_15594);
and U15822 (N_15822,N_15679,N_15631);
nand U15823 (N_15823,N_15680,N_15601);
and U15824 (N_15824,N_15745,N_15674);
nor U15825 (N_15825,N_15621,N_15640);
nor U15826 (N_15826,N_15721,N_15716);
and U15827 (N_15827,N_15711,N_15710);
nand U15828 (N_15828,N_15537,N_15731);
and U15829 (N_15829,N_15543,N_15508);
nor U15830 (N_15830,N_15608,N_15518);
xor U15831 (N_15831,N_15590,N_15574);
nand U15832 (N_15832,N_15510,N_15548);
nor U15833 (N_15833,N_15689,N_15722);
xnor U15834 (N_15834,N_15503,N_15659);
and U15835 (N_15835,N_15605,N_15686);
or U15836 (N_15836,N_15707,N_15703);
nor U15837 (N_15837,N_15603,N_15544);
or U15838 (N_15838,N_15583,N_15666);
nand U15839 (N_15839,N_15551,N_15570);
and U15840 (N_15840,N_15562,N_15579);
nand U15841 (N_15841,N_15632,N_15588);
or U15842 (N_15842,N_15713,N_15678);
nand U15843 (N_15843,N_15546,N_15747);
nand U15844 (N_15844,N_15642,N_15529);
nand U15845 (N_15845,N_15592,N_15696);
and U15846 (N_15846,N_15650,N_15706);
or U15847 (N_15847,N_15681,N_15597);
or U15848 (N_15848,N_15599,N_15528);
xnor U15849 (N_15849,N_15600,N_15655);
nor U15850 (N_15850,N_15622,N_15598);
or U15851 (N_15851,N_15669,N_15717);
or U15852 (N_15852,N_15668,N_15617);
xor U15853 (N_15853,N_15725,N_15638);
nor U15854 (N_15854,N_15698,N_15646);
or U15855 (N_15855,N_15624,N_15629);
xnor U15856 (N_15856,N_15514,N_15572);
or U15857 (N_15857,N_15566,N_15591);
nand U15858 (N_15858,N_15502,N_15586);
nand U15859 (N_15859,N_15733,N_15553);
nand U15860 (N_15860,N_15670,N_15634);
nand U15861 (N_15861,N_15693,N_15656);
nand U15862 (N_15862,N_15746,N_15702);
and U15863 (N_15863,N_15520,N_15561);
and U15864 (N_15864,N_15618,N_15576);
nand U15865 (N_15865,N_15500,N_15700);
nand U15866 (N_15866,N_15687,N_15748);
or U15867 (N_15867,N_15653,N_15620);
nand U15868 (N_15868,N_15541,N_15619);
and U15869 (N_15869,N_15585,N_15644);
nand U15870 (N_15870,N_15694,N_15526);
xor U15871 (N_15871,N_15560,N_15593);
nand U15872 (N_15872,N_15740,N_15596);
xor U15873 (N_15873,N_15623,N_15720);
or U15874 (N_15874,N_15714,N_15533);
xor U15875 (N_15875,N_15685,N_15529);
and U15876 (N_15876,N_15554,N_15509);
or U15877 (N_15877,N_15679,N_15577);
xor U15878 (N_15878,N_15608,N_15537);
and U15879 (N_15879,N_15685,N_15709);
or U15880 (N_15880,N_15559,N_15589);
nand U15881 (N_15881,N_15740,N_15561);
xor U15882 (N_15882,N_15610,N_15569);
xor U15883 (N_15883,N_15733,N_15628);
nand U15884 (N_15884,N_15645,N_15671);
nor U15885 (N_15885,N_15548,N_15672);
xnor U15886 (N_15886,N_15577,N_15651);
nor U15887 (N_15887,N_15508,N_15740);
xnor U15888 (N_15888,N_15651,N_15693);
xnor U15889 (N_15889,N_15748,N_15604);
nand U15890 (N_15890,N_15516,N_15616);
nor U15891 (N_15891,N_15655,N_15608);
nand U15892 (N_15892,N_15556,N_15584);
and U15893 (N_15893,N_15730,N_15504);
and U15894 (N_15894,N_15646,N_15749);
or U15895 (N_15895,N_15742,N_15578);
nand U15896 (N_15896,N_15572,N_15748);
and U15897 (N_15897,N_15548,N_15629);
xor U15898 (N_15898,N_15534,N_15724);
and U15899 (N_15899,N_15520,N_15544);
nor U15900 (N_15900,N_15608,N_15672);
nor U15901 (N_15901,N_15555,N_15628);
and U15902 (N_15902,N_15615,N_15550);
nand U15903 (N_15903,N_15747,N_15576);
and U15904 (N_15904,N_15733,N_15605);
or U15905 (N_15905,N_15644,N_15537);
nand U15906 (N_15906,N_15634,N_15702);
nor U15907 (N_15907,N_15598,N_15654);
nand U15908 (N_15908,N_15589,N_15635);
xor U15909 (N_15909,N_15545,N_15550);
nor U15910 (N_15910,N_15610,N_15587);
nor U15911 (N_15911,N_15643,N_15684);
or U15912 (N_15912,N_15523,N_15656);
nor U15913 (N_15913,N_15674,N_15609);
xor U15914 (N_15914,N_15540,N_15514);
nand U15915 (N_15915,N_15722,N_15720);
nand U15916 (N_15916,N_15609,N_15533);
nand U15917 (N_15917,N_15736,N_15676);
xor U15918 (N_15918,N_15588,N_15626);
xnor U15919 (N_15919,N_15631,N_15692);
nand U15920 (N_15920,N_15644,N_15566);
or U15921 (N_15921,N_15711,N_15550);
xnor U15922 (N_15922,N_15586,N_15587);
and U15923 (N_15923,N_15520,N_15650);
and U15924 (N_15924,N_15691,N_15648);
nand U15925 (N_15925,N_15643,N_15567);
nor U15926 (N_15926,N_15711,N_15632);
nor U15927 (N_15927,N_15506,N_15530);
and U15928 (N_15928,N_15648,N_15692);
or U15929 (N_15929,N_15507,N_15686);
nor U15930 (N_15930,N_15576,N_15653);
xnor U15931 (N_15931,N_15718,N_15547);
xor U15932 (N_15932,N_15699,N_15522);
and U15933 (N_15933,N_15744,N_15746);
nand U15934 (N_15934,N_15626,N_15622);
or U15935 (N_15935,N_15665,N_15502);
nand U15936 (N_15936,N_15736,N_15666);
or U15937 (N_15937,N_15616,N_15627);
xor U15938 (N_15938,N_15638,N_15730);
or U15939 (N_15939,N_15701,N_15515);
nor U15940 (N_15940,N_15685,N_15691);
xnor U15941 (N_15941,N_15564,N_15651);
or U15942 (N_15942,N_15724,N_15574);
xor U15943 (N_15943,N_15700,N_15502);
nand U15944 (N_15944,N_15734,N_15509);
and U15945 (N_15945,N_15569,N_15554);
nor U15946 (N_15946,N_15559,N_15674);
or U15947 (N_15947,N_15710,N_15538);
nand U15948 (N_15948,N_15586,N_15527);
nand U15949 (N_15949,N_15736,N_15530);
or U15950 (N_15950,N_15522,N_15543);
and U15951 (N_15951,N_15568,N_15733);
nand U15952 (N_15952,N_15675,N_15615);
or U15953 (N_15953,N_15640,N_15538);
and U15954 (N_15954,N_15683,N_15545);
xnor U15955 (N_15955,N_15691,N_15528);
nand U15956 (N_15956,N_15606,N_15703);
xnor U15957 (N_15957,N_15526,N_15688);
nor U15958 (N_15958,N_15729,N_15690);
and U15959 (N_15959,N_15729,N_15533);
and U15960 (N_15960,N_15650,N_15579);
and U15961 (N_15961,N_15656,N_15550);
or U15962 (N_15962,N_15560,N_15626);
xnor U15963 (N_15963,N_15723,N_15604);
nor U15964 (N_15964,N_15536,N_15687);
xnor U15965 (N_15965,N_15651,N_15707);
and U15966 (N_15966,N_15566,N_15587);
xor U15967 (N_15967,N_15515,N_15520);
nand U15968 (N_15968,N_15738,N_15510);
and U15969 (N_15969,N_15516,N_15528);
nor U15970 (N_15970,N_15525,N_15573);
nor U15971 (N_15971,N_15526,N_15685);
nand U15972 (N_15972,N_15713,N_15669);
and U15973 (N_15973,N_15681,N_15556);
nand U15974 (N_15974,N_15604,N_15678);
nand U15975 (N_15975,N_15714,N_15574);
or U15976 (N_15976,N_15663,N_15697);
and U15977 (N_15977,N_15702,N_15655);
nor U15978 (N_15978,N_15502,N_15720);
xnor U15979 (N_15979,N_15519,N_15708);
nor U15980 (N_15980,N_15577,N_15509);
nor U15981 (N_15981,N_15693,N_15560);
nor U15982 (N_15982,N_15583,N_15729);
nor U15983 (N_15983,N_15587,N_15697);
nand U15984 (N_15984,N_15708,N_15625);
nand U15985 (N_15985,N_15702,N_15542);
and U15986 (N_15986,N_15557,N_15601);
xor U15987 (N_15987,N_15650,N_15743);
or U15988 (N_15988,N_15680,N_15589);
xnor U15989 (N_15989,N_15581,N_15599);
and U15990 (N_15990,N_15728,N_15528);
or U15991 (N_15991,N_15669,N_15747);
nand U15992 (N_15992,N_15643,N_15735);
xnor U15993 (N_15993,N_15507,N_15665);
nor U15994 (N_15994,N_15607,N_15623);
nand U15995 (N_15995,N_15533,N_15659);
and U15996 (N_15996,N_15652,N_15573);
nand U15997 (N_15997,N_15694,N_15506);
nor U15998 (N_15998,N_15562,N_15561);
or U15999 (N_15999,N_15687,N_15699);
and U16000 (N_16000,N_15889,N_15963);
and U16001 (N_16001,N_15919,N_15949);
nor U16002 (N_16002,N_15796,N_15883);
nor U16003 (N_16003,N_15942,N_15755);
or U16004 (N_16004,N_15774,N_15763);
or U16005 (N_16005,N_15891,N_15819);
xnor U16006 (N_16006,N_15757,N_15927);
or U16007 (N_16007,N_15772,N_15909);
or U16008 (N_16008,N_15779,N_15935);
or U16009 (N_16009,N_15943,N_15920);
nand U16010 (N_16010,N_15952,N_15947);
xnor U16011 (N_16011,N_15954,N_15880);
nor U16012 (N_16012,N_15857,N_15856);
xor U16013 (N_16013,N_15969,N_15967);
or U16014 (N_16014,N_15869,N_15841);
nand U16015 (N_16015,N_15838,N_15959);
and U16016 (N_16016,N_15785,N_15837);
or U16017 (N_16017,N_15921,N_15836);
and U16018 (N_16018,N_15798,N_15769);
xor U16019 (N_16019,N_15764,N_15976);
or U16020 (N_16020,N_15761,N_15953);
xnor U16021 (N_16021,N_15842,N_15860);
nor U16022 (N_16022,N_15813,N_15892);
xnor U16023 (N_16023,N_15923,N_15955);
nand U16024 (N_16024,N_15766,N_15828);
and U16025 (N_16025,N_15876,N_15974);
nor U16026 (N_16026,N_15911,N_15998);
xor U16027 (N_16027,N_15847,N_15815);
nand U16028 (N_16028,N_15936,N_15989);
nor U16029 (N_16029,N_15770,N_15859);
and U16030 (N_16030,N_15972,N_15840);
or U16031 (N_16031,N_15938,N_15754);
or U16032 (N_16032,N_15928,N_15994);
or U16033 (N_16033,N_15906,N_15981);
nor U16034 (N_16034,N_15922,N_15867);
and U16035 (N_16035,N_15956,N_15934);
and U16036 (N_16036,N_15932,N_15853);
xor U16037 (N_16037,N_15870,N_15908);
nor U16038 (N_16038,N_15964,N_15905);
nand U16039 (N_16039,N_15915,N_15816);
xor U16040 (N_16040,N_15799,N_15788);
nand U16041 (N_16041,N_15991,N_15806);
or U16042 (N_16042,N_15780,N_15913);
or U16043 (N_16043,N_15979,N_15961);
or U16044 (N_16044,N_15765,N_15834);
nand U16045 (N_16045,N_15802,N_15965);
and U16046 (N_16046,N_15824,N_15758);
nand U16047 (N_16047,N_15830,N_15917);
nor U16048 (N_16048,N_15821,N_15873);
nor U16049 (N_16049,N_15809,N_15884);
nand U16050 (N_16050,N_15996,N_15924);
and U16051 (N_16051,N_15901,N_15948);
or U16052 (N_16052,N_15878,N_15902);
nor U16053 (N_16053,N_15983,N_15795);
nand U16054 (N_16054,N_15805,N_15791);
or U16055 (N_16055,N_15893,N_15792);
and U16056 (N_16056,N_15845,N_15768);
xnor U16057 (N_16057,N_15897,N_15962);
and U16058 (N_16058,N_15773,N_15812);
xor U16059 (N_16059,N_15817,N_15826);
xor U16060 (N_16060,N_15822,N_15832);
nand U16061 (N_16061,N_15874,N_15868);
and U16062 (N_16062,N_15861,N_15966);
xnor U16063 (N_16063,N_15794,N_15751);
nor U16064 (N_16064,N_15823,N_15930);
or U16065 (N_16065,N_15835,N_15829);
or U16066 (N_16066,N_15848,N_15756);
and U16067 (N_16067,N_15825,N_15851);
nand U16068 (N_16068,N_15960,N_15879);
nor U16069 (N_16069,N_15910,N_15916);
and U16070 (N_16070,N_15980,N_15865);
nor U16071 (N_16071,N_15753,N_15982);
nor U16072 (N_16072,N_15850,N_15877);
or U16073 (N_16073,N_15811,N_15945);
nor U16074 (N_16074,N_15939,N_15925);
nand U16075 (N_16075,N_15904,N_15797);
xnor U16076 (N_16076,N_15767,N_15760);
or U16077 (N_16077,N_15852,N_15975);
nor U16078 (N_16078,N_15790,N_15929);
and U16079 (N_16079,N_15946,N_15807);
nand U16080 (N_16080,N_15885,N_15786);
xor U16081 (N_16081,N_15759,N_15957);
and U16082 (N_16082,N_15970,N_15886);
nand U16083 (N_16083,N_15933,N_15864);
xor U16084 (N_16084,N_15854,N_15793);
and U16085 (N_16085,N_15778,N_15771);
xnor U16086 (N_16086,N_15950,N_15995);
nor U16087 (N_16087,N_15971,N_15752);
or U16088 (N_16088,N_15862,N_15872);
or U16089 (N_16089,N_15931,N_15782);
nor U16090 (N_16090,N_15863,N_15968);
xnor U16091 (N_16091,N_15818,N_15914);
xnor U16092 (N_16092,N_15985,N_15887);
and U16093 (N_16093,N_15762,N_15781);
or U16094 (N_16094,N_15973,N_15750);
xnor U16095 (N_16095,N_15984,N_15881);
xor U16096 (N_16096,N_15803,N_15992);
xor U16097 (N_16097,N_15898,N_15918);
nand U16098 (N_16098,N_15941,N_15987);
nand U16099 (N_16099,N_15871,N_15951);
and U16100 (N_16100,N_15875,N_15958);
xnor U16101 (N_16101,N_15827,N_15843);
or U16102 (N_16102,N_15907,N_15944);
nor U16103 (N_16103,N_15775,N_15844);
or U16104 (N_16104,N_15783,N_15895);
nor U16105 (N_16105,N_15977,N_15784);
and U16106 (N_16106,N_15940,N_15800);
nor U16107 (N_16107,N_15776,N_15997);
xnor U16108 (N_16108,N_15858,N_15839);
and U16109 (N_16109,N_15777,N_15866);
nand U16110 (N_16110,N_15801,N_15988);
nand U16111 (N_16111,N_15896,N_15849);
xnor U16112 (N_16112,N_15926,N_15882);
or U16113 (N_16113,N_15990,N_15903);
and U16114 (N_16114,N_15978,N_15855);
nor U16115 (N_16115,N_15900,N_15814);
and U16116 (N_16116,N_15810,N_15804);
and U16117 (N_16117,N_15808,N_15986);
nor U16118 (N_16118,N_15831,N_15820);
and U16119 (N_16119,N_15894,N_15789);
xnor U16120 (N_16120,N_15999,N_15787);
nand U16121 (N_16121,N_15937,N_15890);
nor U16122 (N_16122,N_15888,N_15833);
and U16123 (N_16123,N_15912,N_15899);
nand U16124 (N_16124,N_15846,N_15993);
and U16125 (N_16125,N_15864,N_15907);
and U16126 (N_16126,N_15787,N_15996);
and U16127 (N_16127,N_15894,N_15840);
nand U16128 (N_16128,N_15839,N_15935);
or U16129 (N_16129,N_15815,N_15800);
or U16130 (N_16130,N_15776,N_15845);
xor U16131 (N_16131,N_15964,N_15875);
or U16132 (N_16132,N_15920,N_15807);
nor U16133 (N_16133,N_15833,N_15857);
nor U16134 (N_16134,N_15966,N_15828);
or U16135 (N_16135,N_15829,N_15795);
and U16136 (N_16136,N_15898,N_15949);
xnor U16137 (N_16137,N_15871,N_15864);
and U16138 (N_16138,N_15823,N_15988);
and U16139 (N_16139,N_15883,N_15941);
nor U16140 (N_16140,N_15776,N_15902);
nor U16141 (N_16141,N_15954,N_15871);
nor U16142 (N_16142,N_15938,N_15775);
nand U16143 (N_16143,N_15843,N_15822);
nor U16144 (N_16144,N_15942,N_15937);
nor U16145 (N_16145,N_15856,N_15891);
nor U16146 (N_16146,N_15811,N_15893);
or U16147 (N_16147,N_15785,N_15911);
and U16148 (N_16148,N_15993,N_15997);
and U16149 (N_16149,N_15918,N_15758);
or U16150 (N_16150,N_15971,N_15821);
or U16151 (N_16151,N_15841,N_15802);
nor U16152 (N_16152,N_15937,N_15769);
and U16153 (N_16153,N_15804,N_15840);
and U16154 (N_16154,N_15931,N_15826);
nand U16155 (N_16155,N_15882,N_15765);
nand U16156 (N_16156,N_15778,N_15777);
xor U16157 (N_16157,N_15918,N_15808);
nand U16158 (N_16158,N_15951,N_15866);
nor U16159 (N_16159,N_15823,N_15893);
nor U16160 (N_16160,N_15818,N_15979);
or U16161 (N_16161,N_15759,N_15889);
or U16162 (N_16162,N_15758,N_15893);
nand U16163 (N_16163,N_15931,N_15895);
or U16164 (N_16164,N_15852,N_15824);
or U16165 (N_16165,N_15753,N_15944);
and U16166 (N_16166,N_15764,N_15909);
nor U16167 (N_16167,N_15764,N_15848);
and U16168 (N_16168,N_15914,N_15877);
xnor U16169 (N_16169,N_15828,N_15878);
nand U16170 (N_16170,N_15805,N_15778);
and U16171 (N_16171,N_15976,N_15784);
and U16172 (N_16172,N_15845,N_15866);
nand U16173 (N_16173,N_15891,N_15826);
nand U16174 (N_16174,N_15960,N_15762);
and U16175 (N_16175,N_15845,N_15815);
and U16176 (N_16176,N_15932,N_15936);
and U16177 (N_16177,N_15787,N_15897);
xor U16178 (N_16178,N_15777,N_15831);
nor U16179 (N_16179,N_15988,N_15783);
nor U16180 (N_16180,N_15838,N_15936);
or U16181 (N_16181,N_15956,N_15981);
nor U16182 (N_16182,N_15968,N_15828);
nand U16183 (N_16183,N_15952,N_15883);
and U16184 (N_16184,N_15784,N_15895);
nor U16185 (N_16185,N_15770,N_15925);
nor U16186 (N_16186,N_15775,N_15847);
nor U16187 (N_16187,N_15996,N_15816);
and U16188 (N_16188,N_15766,N_15829);
nand U16189 (N_16189,N_15773,N_15935);
nand U16190 (N_16190,N_15856,N_15951);
or U16191 (N_16191,N_15992,N_15765);
nor U16192 (N_16192,N_15943,N_15881);
xnor U16193 (N_16193,N_15972,N_15855);
or U16194 (N_16194,N_15754,N_15796);
or U16195 (N_16195,N_15969,N_15890);
or U16196 (N_16196,N_15930,N_15895);
nand U16197 (N_16197,N_15986,N_15766);
xnor U16198 (N_16198,N_15971,N_15988);
nor U16199 (N_16199,N_15802,N_15809);
nor U16200 (N_16200,N_15991,N_15963);
nand U16201 (N_16201,N_15949,N_15937);
and U16202 (N_16202,N_15898,N_15915);
nand U16203 (N_16203,N_15926,N_15788);
nand U16204 (N_16204,N_15776,N_15806);
or U16205 (N_16205,N_15851,N_15827);
xor U16206 (N_16206,N_15781,N_15884);
xor U16207 (N_16207,N_15779,N_15778);
xor U16208 (N_16208,N_15865,N_15838);
nand U16209 (N_16209,N_15898,N_15998);
nor U16210 (N_16210,N_15813,N_15886);
nor U16211 (N_16211,N_15940,N_15978);
nand U16212 (N_16212,N_15790,N_15910);
nand U16213 (N_16213,N_15912,N_15943);
or U16214 (N_16214,N_15940,N_15850);
or U16215 (N_16215,N_15954,N_15920);
xor U16216 (N_16216,N_15785,N_15910);
xor U16217 (N_16217,N_15937,N_15806);
or U16218 (N_16218,N_15964,N_15853);
nand U16219 (N_16219,N_15906,N_15862);
nor U16220 (N_16220,N_15855,N_15854);
nand U16221 (N_16221,N_15901,N_15807);
nand U16222 (N_16222,N_15897,N_15900);
nor U16223 (N_16223,N_15789,N_15774);
or U16224 (N_16224,N_15870,N_15990);
or U16225 (N_16225,N_15950,N_15836);
nor U16226 (N_16226,N_15901,N_15985);
nand U16227 (N_16227,N_15956,N_15908);
nor U16228 (N_16228,N_15901,N_15959);
and U16229 (N_16229,N_15920,N_15882);
xor U16230 (N_16230,N_15930,N_15933);
or U16231 (N_16231,N_15856,N_15936);
nand U16232 (N_16232,N_15765,N_15830);
or U16233 (N_16233,N_15767,N_15960);
nor U16234 (N_16234,N_15791,N_15895);
nand U16235 (N_16235,N_15998,N_15895);
and U16236 (N_16236,N_15977,N_15990);
and U16237 (N_16237,N_15993,N_15877);
and U16238 (N_16238,N_15862,N_15767);
xor U16239 (N_16239,N_15850,N_15975);
xnor U16240 (N_16240,N_15950,N_15952);
nand U16241 (N_16241,N_15990,N_15750);
nor U16242 (N_16242,N_15790,N_15869);
xnor U16243 (N_16243,N_15886,N_15800);
xor U16244 (N_16244,N_15786,N_15997);
nand U16245 (N_16245,N_15956,N_15815);
nand U16246 (N_16246,N_15880,N_15918);
and U16247 (N_16247,N_15850,N_15780);
and U16248 (N_16248,N_15867,N_15905);
nand U16249 (N_16249,N_15825,N_15751);
nand U16250 (N_16250,N_16083,N_16200);
and U16251 (N_16251,N_16212,N_16051);
nand U16252 (N_16252,N_16201,N_16236);
xnor U16253 (N_16253,N_16171,N_16085);
or U16254 (N_16254,N_16165,N_16075);
and U16255 (N_16255,N_16166,N_16109);
nand U16256 (N_16256,N_16007,N_16010);
nand U16257 (N_16257,N_16242,N_16037);
xnor U16258 (N_16258,N_16193,N_16145);
nor U16259 (N_16259,N_16240,N_16057);
and U16260 (N_16260,N_16207,N_16078);
or U16261 (N_16261,N_16024,N_16219);
nor U16262 (N_16262,N_16068,N_16152);
nand U16263 (N_16263,N_16062,N_16061);
or U16264 (N_16264,N_16033,N_16064);
nor U16265 (N_16265,N_16170,N_16004);
and U16266 (N_16266,N_16153,N_16117);
nor U16267 (N_16267,N_16139,N_16183);
nor U16268 (N_16268,N_16189,N_16054);
nand U16269 (N_16269,N_16150,N_16012);
or U16270 (N_16270,N_16087,N_16103);
and U16271 (N_16271,N_16040,N_16175);
nor U16272 (N_16272,N_16048,N_16003);
and U16273 (N_16273,N_16009,N_16228);
xor U16274 (N_16274,N_16106,N_16072);
xor U16275 (N_16275,N_16158,N_16137);
or U16276 (N_16276,N_16135,N_16247);
xnor U16277 (N_16277,N_16186,N_16126);
and U16278 (N_16278,N_16167,N_16076);
and U16279 (N_16279,N_16202,N_16190);
and U16280 (N_16280,N_16063,N_16128);
xor U16281 (N_16281,N_16029,N_16047);
or U16282 (N_16282,N_16177,N_16125);
and U16283 (N_16283,N_16000,N_16235);
or U16284 (N_16284,N_16133,N_16074);
or U16285 (N_16285,N_16208,N_16131);
nand U16286 (N_16286,N_16232,N_16173);
nor U16287 (N_16287,N_16237,N_16213);
and U16288 (N_16288,N_16222,N_16089);
and U16289 (N_16289,N_16215,N_16161);
nand U16290 (N_16290,N_16226,N_16136);
and U16291 (N_16291,N_16116,N_16034);
nor U16292 (N_16292,N_16070,N_16112);
nor U16293 (N_16293,N_16230,N_16084);
xnor U16294 (N_16294,N_16097,N_16023);
and U16295 (N_16295,N_16082,N_16229);
or U16296 (N_16296,N_16108,N_16221);
xor U16297 (N_16297,N_16060,N_16055);
nand U16298 (N_16298,N_16043,N_16144);
nand U16299 (N_16299,N_16102,N_16141);
xor U16300 (N_16300,N_16099,N_16111);
and U16301 (N_16301,N_16036,N_16067);
or U16302 (N_16302,N_16233,N_16017);
and U16303 (N_16303,N_16239,N_16231);
nand U16304 (N_16304,N_16011,N_16143);
nor U16305 (N_16305,N_16008,N_16073);
nand U16306 (N_16306,N_16032,N_16022);
nand U16307 (N_16307,N_16042,N_16025);
nor U16308 (N_16308,N_16091,N_16154);
nor U16309 (N_16309,N_16142,N_16049);
and U16310 (N_16310,N_16196,N_16249);
and U16311 (N_16311,N_16002,N_16113);
or U16312 (N_16312,N_16129,N_16058);
and U16313 (N_16313,N_16206,N_16174);
and U16314 (N_16314,N_16019,N_16238);
xor U16315 (N_16315,N_16122,N_16188);
nor U16316 (N_16316,N_16118,N_16163);
nand U16317 (N_16317,N_16005,N_16077);
nand U16318 (N_16318,N_16181,N_16162);
xnor U16319 (N_16319,N_16050,N_16092);
nor U16320 (N_16320,N_16147,N_16114);
or U16321 (N_16321,N_16046,N_16093);
nor U16322 (N_16322,N_16096,N_16182);
and U16323 (N_16323,N_16115,N_16066);
nor U16324 (N_16324,N_16194,N_16041);
nand U16325 (N_16325,N_16119,N_16148);
nor U16326 (N_16326,N_16098,N_16100);
or U16327 (N_16327,N_16071,N_16026);
nand U16328 (N_16328,N_16027,N_16243);
and U16329 (N_16329,N_16107,N_16218);
nor U16330 (N_16330,N_16020,N_16168);
nand U16331 (N_16331,N_16105,N_16156);
and U16332 (N_16332,N_16014,N_16045);
nor U16333 (N_16333,N_16246,N_16138);
nand U16334 (N_16334,N_16191,N_16104);
xnor U16335 (N_16335,N_16210,N_16248);
or U16336 (N_16336,N_16223,N_16245);
and U16337 (N_16337,N_16069,N_16080);
or U16338 (N_16338,N_16184,N_16101);
nor U16339 (N_16339,N_16094,N_16185);
and U16340 (N_16340,N_16127,N_16079);
nand U16341 (N_16341,N_16164,N_16110);
xor U16342 (N_16342,N_16124,N_16180);
xor U16343 (N_16343,N_16001,N_16160);
or U16344 (N_16344,N_16176,N_16157);
nand U16345 (N_16345,N_16123,N_16224);
nor U16346 (N_16346,N_16028,N_16130);
xor U16347 (N_16347,N_16081,N_16021);
or U16348 (N_16348,N_16220,N_16044);
xnor U16349 (N_16349,N_16018,N_16178);
and U16350 (N_16350,N_16149,N_16155);
or U16351 (N_16351,N_16216,N_16169);
xnor U16352 (N_16352,N_16203,N_16016);
nor U16353 (N_16353,N_16086,N_16192);
or U16354 (N_16354,N_16187,N_16244);
xor U16355 (N_16355,N_16065,N_16134);
or U16356 (N_16356,N_16056,N_16204);
nor U16357 (N_16357,N_16197,N_16013);
nand U16358 (N_16358,N_16038,N_16088);
xnor U16359 (N_16359,N_16172,N_16211);
and U16360 (N_16360,N_16030,N_16132);
nand U16361 (N_16361,N_16205,N_16031);
or U16362 (N_16362,N_16179,N_16006);
or U16363 (N_16363,N_16209,N_16214);
nor U16364 (N_16364,N_16053,N_16059);
or U16365 (N_16365,N_16095,N_16052);
xnor U16366 (N_16366,N_16217,N_16121);
nor U16367 (N_16367,N_16035,N_16140);
or U16368 (N_16368,N_16195,N_16198);
and U16369 (N_16369,N_16234,N_16159);
xnor U16370 (N_16370,N_16225,N_16227);
or U16371 (N_16371,N_16146,N_16120);
and U16372 (N_16372,N_16199,N_16151);
or U16373 (N_16373,N_16241,N_16090);
and U16374 (N_16374,N_16015,N_16039);
nand U16375 (N_16375,N_16104,N_16160);
or U16376 (N_16376,N_16096,N_16128);
and U16377 (N_16377,N_16042,N_16227);
and U16378 (N_16378,N_16230,N_16141);
xor U16379 (N_16379,N_16207,N_16126);
or U16380 (N_16380,N_16027,N_16130);
or U16381 (N_16381,N_16152,N_16139);
nand U16382 (N_16382,N_16123,N_16182);
xor U16383 (N_16383,N_16057,N_16065);
or U16384 (N_16384,N_16135,N_16131);
and U16385 (N_16385,N_16062,N_16193);
nand U16386 (N_16386,N_16150,N_16198);
or U16387 (N_16387,N_16155,N_16043);
and U16388 (N_16388,N_16193,N_16000);
xnor U16389 (N_16389,N_16157,N_16135);
nand U16390 (N_16390,N_16022,N_16175);
or U16391 (N_16391,N_16079,N_16057);
nor U16392 (N_16392,N_16169,N_16144);
xnor U16393 (N_16393,N_16085,N_16094);
nor U16394 (N_16394,N_16170,N_16202);
nand U16395 (N_16395,N_16034,N_16182);
or U16396 (N_16396,N_16086,N_16150);
xor U16397 (N_16397,N_16208,N_16241);
nor U16398 (N_16398,N_16120,N_16106);
or U16399 (N_16399,N_16043,N_16026);
or U16400 (N_16400,N_16170,N_16005);
nand U16401 (N_16401,N_16119,N_16212);
or U16402 (N_16402,N_16094,N_16059);
or U16403 (N_16403,N_16143,N_16066);
or U16404 (N_16404,N_16060,N_16172);
nor U16405 (N_16405,N_16100,N_16109);
or U16406 (N_16406,N_16087,N_16105);
xnor U16407 (N_16407,N_16011,N_16036);
xnor U16408 (N_16408,N_16088,N_16160);
or U16409 (N_16409,N_16079,N_16046);
or U16410 (N_16410,N_16058,N_16014);
nor U16411 (N_16411,N_16127,N_16080);
nor U16412 (N_16412,N_16030,N_16019);
nor U16413 (N_16413,N_16180,N_16141);
and U16414 (N_16414,N_16196,N_16142);
nand U16415 (N_16415,N_16049,N_16036);
or U16416 (N_16416,N_16020,N_16098);
nor U16417 (N_16417,N_16118,N_16016);
and U16418 (N_16418,N_16193,N_16190);
nor U16419 (N_16419,N_16178,N_16231);
nand U16420 (N_16420,N_16079,N_16092);
or U16421 (N_16421,N_16204,N_16111);
xnor U16422 (N_16422,N_16117,N_16067);
nand U16423 (N_16423,N_16088,N_16112);
nand U16424 (N_16424,N_16224,N_16247);
nor U16425 (N_16425,N_16245,N_16128);
or U16426 (N_16426,N_16084,N_16017);
nor U16427 (N_16427,N_16188,N_16098);
xnor U16428 (N_16428,N_16121,N_16184);
xor U16429 (N_16429,N_16157,N_16137);
nand U16430 (N_16430,N_16136,N_16174);
nand U16431 (N_16431,N_16174,N_16144);
nand U16432 (N_16432,N_16042,N_16075);
nor U16433 (N_16433,N_16011,N_16173);
and U16434 (N_16434,N_16181,N_16051);
nor U16435 (N_16435,N_16236,N_16131);
nor U16436 (N_16436,N_16237,N_16036);
xor U16437 (N_16437,N_16008,N_16069);
nand U16438 (N_16438,N_16168,N_16030);
nor U16439 (N_16439,N_16130,N_16037);
nor U16440 (N_16440,N_16118,N_16028);
nor U16441 (N_16441,N_16137,N_16069);
nand U16442 (N_16442,N_16023,N_16056);
nor U16443 (N_16443,N_16173,N_16126);
xor U16444 (N_16444,N_16139,N_16023);
xor U16445 (N_16445,N_16199,N_16138);
and U16446 (N_16446,N_16024,N_16136);
xor U16447 (N_16447,N_16054,N_16174);
or U16448 (N_16448,N_16130,N_16014);
or U16449 (N_16449,N_16181,N_16099);
xnor U16450 (N_16450,N_16221,N_16058);
or U16451 (N_16451,N_16208,N_16085);
nand U16452 (N_16452,N_16040,N_16063);
xnor U16453 (N_16453,N_16173,N_16024);
and U16454 (N_16454,N_16061,N_16127);
and U16455 (N_16455,N_16162,N_16152);
nor U16456 (N_16456,N_16160,N_16091);
nor U16457 (N_16457,N_16050,N_16244);
nand U16458 (N_16458,N_16244,N_16142);
nand U16459 (N_16459,N_16163,N_16200);
nor U16460 (N_16460,N_16087,N_16076);
nor U16461 (N_16461,N_16219,N_16236);
nor U16462 (N_16462,N_16218,N_16207);
xnor U16463 (N_16463,N_16236,N_16067);
nor U16464 (N_16464,N_16023,N_16242);
and U16465 (N_16465,N_16038,N_16110);
nand U16466 (N_16466,N_16193,N_16040);
or U16467 (N_16467,N_16169,N_16193);
or U16468 (N_16468,N_16219,N_16137);
nand U16469 (N_16469,N_16049,N_16092);
or U16470 (N_16470,N_16242,N_16216);
nor U16471 (N_16471,N_16048,N_16019);
and U16472 (N_16472,N_16217,N_16171);
nor U16473 (N_16473,N_16070,N_16233);
or U16474 (N_16474,N_16066,N_16202);
nor U16475 (N_16475,N_16042,N_16185);
xnor U16476 (N_16476,N_16091,N_16094);
nor U16477 (N_16477,N_16163,N_16007);
nand U16478 (N_16478,N_16028,N_16014);
nor U16479 (N_16479,N_16077,N_16040);
or U16480 (N_16480,N_16204,N_16219);
and U16481 (N_16481,N_16168,N_16133);
nor U16482 (N_16482,N_16134,N_16112);
nand U16483 (N_16483,N_16021,N_16232);
xnor U16484 (N_16484,N_16136,N_16148);
nor U16485 (N_16485,N_16015,N_16107);
nand U16486 (N_16486,N_16055,N_16023);
xnor U16487 (N_16487,N_16127,N_16118);
nand U16488 (N_16488,N_16215,N_16186);
nor U16489 (N_16489,N_16221,N_16193);
xor U16490 (N_16490,N_16120,N_16115);
nand U16491 (N_16491,N_16135,N_16089);
and U16492 (N_16492,N_16223,N_16019);
and U16493 (N_16493,N_16027,N_16081);
nand U16494 (N_16494,N_16237,N_16120);
nand U16495 (N_16495,N_16189,N_16137);
and U16496 (N_16496,N_16164,N_16163);
or U16497 (N_16497,N_16034,N_16002);
nor U16498 (N_16498,N_16006,N_16013);
nand U16499 (N_16499,N_16120,N_16179);
nor U16500 (N_16500,N_16420,N_16465);
nand U16501 (N_16501,N_16377,N_16393);
or U16502 (N_16502,N_16471,N_16392);
nor U16503 (N_16503,N_16331,N_16328);
and U16504 (N_16504,N_16404,N_16468);
xnor U16505 (N_16505,N_16326,N_16397);
nor U16506 (N_16506,N_16297,N_16269);
xnor U16507 (N_16507,N_16321,N_16348);
and U16508 (N_16508,N_16286,N_16351);
nand U16509 (N_16509,N_16312,N_16256);
nor U16510 (N_16510,N_16479,N_16371);
nand U16511 (N_16511,N_16433,N_16448);
and U16512 (N_16512,N_16439,N_16462);
nor U16513 (N_16513,N_16411,N_16385);
and U16514 (N_16514,N_16254,N_16271);
or U16515 (N_16515,N_16273,N_16325);
nand U16516 (N_16516,N_16492,N_16442);
and U16517 (N_16517,N_16444,N_16352);
and U16518 (N_16518,N_16381,N_16401);
and U16519 (N_16519,N_16414,N_16417);
nor U16520 (N_16520,N_16270,N_16403);
and U16521 (N_16521,N_16282,N_16423);
or U16522 (N_16522,N_16283,N_16274);
and U16523 (N_16523,N_16339,N_16315);
xor U16524 (N_16524,N_16376,N_16380);
xor U16525 (N_16525,N_16470,N_16298);
nor U16526 (N_16526,N_16494,N_16412);
nand U16527 (N_16527,N_16388,N_16374);
and U16528 (N_16528,N_16285,N_16426);
or U16529 (N_16529,N_16344,N_16322);
nor U16530 (N_16530,N_16364,N_16338);
xor U16531 (N_16531,N_16261,N_16280);
nor U16532 (N_16532,N_16354,N_16264);
or U16533 (N_16533,N_16436,N_16478);
or U16534 (N_16534,N_16424,N_16309);
and U16535 (N_16535,N_16455,N_16487);
nor U16536 (N_16536,N_16382,N_16451);
nand U16537 (N_16537,N_16265,N_16292);
and U16538 (N_16538,N_16258,N_16260);
xnor U16539 (N_16539,N_16454,N_16373);
xnor U16540 (N_16540,N_16337,N_16394);
nor U16541 (N_16541,N_16317,N_16358);
or U16542 (N_16542,N_16275,N_16350);
and U16543 (N_16543,N_16294,N_16257);
nand U16544 (N_16544,N_16342,N_16303);
or U16545 (N_16545,N_16480,N_16482);
nor U16546 (N_16546,N_16356,N_16333);
xnor U16547 (N_16547,N_16489,N_16266);
xor U16548 (N_16548,N_16262,N_16277);
nor U16549 (N_16549,N_16304,N_16418);
nor U16550 (N_16550,N_16390,N_16483);
or U16551 (N_16551,N_16367,N_16476);
or U16552 (N_16552,N_16413,N_16316);
nand U16553 (N_16553,N_16449,N_16360);
nand U16554 (N_16554,N_16250,N_16375);
xor U16555 (N_16555,N_16293,N_16495);
xnor U16556 (N_16556,N_16437,N_16335);
xnor U16557 (N_16557,N_16332,N_16450);
nor U16558 (N_16558,N_16384,N_16314);
xor U16559 (N_16559,N_16432,N_16281);
nand U16560 (N_16560,N_16343,N_16425);
and U16561 (N_16561,N_16363,N_16368);
and U16562 (N_16562,N_16389,N_16369);
nor U16563 (N_16563,N_16399,N_16308);
xnor U16564 (N_16564,N_16340,N_16336);
xor U16565 (N_16565,N_16284,N_16313);
xor U16566 (N_16566,N_16330,N_16301);
or U16567 (N_16567,N_16365,N_16459);
nor U16568 (N_16568,N_16435,N_16290);
nand U16569 (N_16569,N_16383,N_16327);
and U16570 (N_16570,N_16463,N_16410);
nand U16571 (N_16571,N_16355,N_16405);
nor U16572 (N_16572,N_16460,N_16430);
nor U16573 (N_16573,N_16268,N_16473);
nor U16574 (N_16574,N_16452,N_16319);
and U16575 (N_16575,N_16440,N_16307);
xor U16576 (N_16576,N_16251,N_16310);
and U16577 (N_16577,N_16457,N_16406);
and U16578 (N_16578,N_16395,N_16387);
or U16579 (N_16579,N_16300,N_16461);
and U16580 (N_16580,N_16311,N_16474);
nor U16581 (N_16581,N_16386,N_16396);
nand U16582 (N_16582,N_16259,N_16429);
nor U16583 (N_16583,N_16359,N_16408);
xor U16584 (N_16584,N_16378,N_16353);
xor U16585 (N_16585,N_16347,N_16469);
and U16586 (N_16586,N_16324,N_16296);
nor U16587 (N_16587,N_16434,N_16415);
nand U16588 (N_16588,N_16295,N_16464);
nand U16589 (N_16589,N_16402,N_16446);
nor U16590 (N_16590,N_16438,N_16263);
or U16591 (N_16591,N_16472,N_16428);
nor U16592 (N_16592,N_16341,N_16253);
xnor U16593 (N_16593,N_16496,N_16466);
nor U16594 (N_16594,N_16288,N_16409);
xnor U16595 (N_16595,N_16323,N_16416);
nand U16596 (N_16596,N_16407,N_16421);
xor U16597 (N_16597,N_16445,N_16306);
or U16598 (N_16598,N_16320,N_16252);
and U16599 (N_16599,N_16346,N_16441);
and U16600 (N_16600,N_16431,N_16370);
xor U16601 (N_16601,N_16398,N_16272);
nor U16602 (N_16602,N_16267,N_16289);
or U16603 (N_16603,N_16276,N_16291);
nand U16604 (N_16604,N_16422,N_16447);
and U16605 (N_16605,N_16329,N_16287);
or U16606 (N_16606,N_16379,N_16362);
nor U16607 (N_16607,N_16491,N_16486);
or U16608 (N_16608,N_16443,N_16497);
xor U16609 (N_16609,N_16458,N_16485);
nand U16610 (N_16610,N_16493,N_16498);
nand U16611 (N_16611,N_16345,N_16255);
nand U16612 (N_16612,N_16305,N_16349);
xor U16613 (N_16613,N_16477,N_16484);
or U16614 (N_16614,N_16279,N_16357);
nor U16615 (N_16615,N_16334,N_16456);
nand U16616 (N_16616,N_16453,N_16391);
nand U16617 (N_16617,N_16302,N_16475);
or U16618 (N_16618,N_16467,N_16499);
nand U16619 (N_16619,N_16299,N_16400);
and U16620 (N_16620,N_16278,N_16427);
or U16621 (N_16621,N_16490,N_16318);
nor U16622 (N_16622,N_16481,N_16488);
xnor U16623 (N_16623,N_16419,N_16372);
and U16624 (N_16624,N_16361,N_16366);
xor U16625 (N_16625,N_16464,N_16327);
nand U16626 (N_16626,N_16389,N_16367);
nor U16627 (N_16627,N_16487,N_16362);
and U16628 (N_16628,N_16486,N_16468);
nor U16629 (N_16629,N_16304,N_16409);
nand U16630 (N_16630,N_16354,N_16356);
and U16631 (N_16631,N_16365,N_16263);
and U16632 (N_16632,N_16425,N_16490);
or U16633 (N_16633,N_16476,N_16423);
xor U16634 (N_16634,N_16364,N_16292);
xnor U16635 (N_16635,N_16302,N_16396);
and U16636 (N_16636,N_16253,N_16319);
nand U16637 (N_16637,N_16303,N_16287);
or U16638 (N_16638,N_16352,N_16258);
nand U16639 (N_16639,N_16409,N_16470);
and U16640 (N_16640,N_16305,N_16364);
and U16641 (N_16641,N_16371,N_16437);
nand U16642 (N_16642,N_16455,N_16448);
xor U16643 (N_16643,N_16389,N_16277);
nand U16644 (N_16644,N_16391,N_16395);
nand U16645 (N_16645,N_16494,N_16428);
or U16646 (N_16646,N_16264,N_16383);
nor U16647 (N_16647,N_16419,N_16377);
nand U16648 (N_16648,N_16392,N_16476);
nand U16649 (N_16649,N_16282,N_16384);
and U16650 (N_16650,N_16449,N_16273);
xor U16651 (N_16651,N_16399,N_16279);
nor U16652 (N_16652,N_16389,N_16283);
and U16653 (N_16653,N_16338,N_16328);
nor U16654 (N_16654,N_16335,N_16487);
xnor U16655 (N_16655,N_16447,N_16461);
or U16656 (N_16656,N_16367,N_16301);
nand U16657 (N_16657,N_16462,N_16283);
nand U16658 (N_16658,N_16363,N_16320);
xnor U16659 (N_16659,N_16444,N_16493);
xor U16660 (N_16660,N_16399,N_16287);
nand U16661 (N_16661,N_16262,N_16351);
nand U16662 (N_16662,N_16384,N_16348);
nor U16663 (N_16663,N_16270,N_16299);
and U16664 (N_16664,N_16345,N_16290);
nor U16665 (N_16665,N_16339,N_16299);
nor U16666 (N_16666,N_16312,N_16375);
nand U16667 (N_16667,N_16388,N_16261);
nor U16668 (N_16668,N_16479,N_16406);
xnor U16669 (N_16669,N_16400,N_16390);
and U16670 (N_16670,N_16255,N_16271);
and U16671 (N_16671,N_16290,N_16413);
nor U16672 (N_16672,N_16300,N_16344);
nand U16673 (N_16673,N_16395,N_16332);
nor U16674 (N_16674,N_16357,N_16361);
and U16675 (N_16675,N_16446,N_16371);
or U16676 (N_16676,N_16255,N_16396);
xor U16677 (N_16677,N_16482,N_16368);
nand U16678 (N_16678,N_16401,N_16458);
nand U16679 (N_16679,N_16343,N_16434);
nand U16680 (N_16680,N_16431,N_16495);
xnor U16681 (N_16681,N_16332,N_16314);
or U16682 (N_16682,N_16459,N_16350);
or U16683 (N_16683,N_16283,N_16488);
xnor U16684 (N_16684,N_16256,N_16454);
xor U16685 (N_16685,N_16340,N_16281);
and U16686 (N_16686,N_16286,N_16481);
xnor U16687 (N_16687,N_16303,N_16264);
or U16688 (N_16688,N_16281,N_16353);
xnor U16689 (N_16689,N_16381,N_16490);
xnor U16690 (N_16690,N_16408,N_16297);
xor U16691 (N_16691,N_16348,N_16393);
nor U16692 (N_16692,N_16371,N_16364);
xor U16693 (N_16693,N_16410,N_16344);
and U16694 (N_16694,N_16301,N_16475);
and U16695 (N_16695,N_16377,N_16481);
xnor U16696 (N_16696,N_16382,N_16336);
or U16697 (N_16697,N_16353,N_16439);
nor U16698 (N_16698,N_16335,N_16350);
and U16699 (N_16699,N_16269,N_16487);
and U16700 (N_16700,N_16251,N_16429);
or U16701 (N_16701,N_16332,N_16347);
nand U16702 (N_16702,N_16468,N_16352);
and U16703 (N_16703,N_16498,N_16478);
and U16704 (N_16704,N_16285,N_16477);
and U16705 (N_16705,N_16386,N_16499);
and U16706 (N_16706,N_16403,N_16364);
nand U16707 (N_16707,N_16387,N_16410);
nand U16708 (N_16708,N_16460,N_16368);
and U16709 (N_16709,N_16346,N_16293);
xnor U16710 (N_16710,N_16463,N_16303);
xor U16711 (N_16711,N_16315,N_16450);
nor U16712 (N_16712,N_16350,N_16361);
and U16713 (N_16713,N_16315,N_16303);
xnor U16714 (N_16714,N_16492,N_16456);
nand U16715 (N_16715,N_16470,N_16369);
nor U16716 (N_16716,N_16253,N_16347);
xor U16717 (N_16717,N_16403,N_16357);
xnor U16718 (N_16718,N_16373,N_16357);
and U16719 (N_16719,N_16493,N_16433);
nand U16720 (N_16720,N_16286,N_16451);
and U16721 (N_16721,N_16287,N_16453);
or U16722 (N_16722,N_16479,N_16415);
nor U16723 (N_16723,N_16452,N_16322);
and U16724 (N_16724,N_16379,N_16279);
nor U16725 (N_16725,N_16460,N_16330);
and U16726 (N_16726,N_16485,N_16256);
or U16727 (N_16727,N_16459,N_16473);
xnor U16728 (N_16728,N_16440,N_16395);
and U16729 (N_16729,N_16348,N_16450);
xor U16730 (N_16730,N_16325,N_16350);
and U16731 (N_16731,N_16434,N_16368);
and U16732 (N_16732,N_16291,N_16402);
xnor U16733 (N_16733,N_16380,N_16404);
xor U16734 (N_16734,N_16375,N_16419);
nor U16735 (N_16735,N_16316,N_16454);
and U16736 (N_16736,N_16464,N_16380);
nor U16737 (N_16737,N_16380,N_16332);
and U16738 (N_16738,N_16383,N_16482);
nor U16739 (N_16739,N_16320,N_16376);
xor U16740 (N_16740,N_16485,N_16334);
and U16741 (N_16741,N_16444,N_16442);
nor U16742 (N_16742,N_16396,N_16313);
nor U16743 (N_16743,N_16343,N_16299);
nor U16744 (N_16744,N_16279,N_16476);
nor U16745 (N_16745,N_16425,N_16440);
or U16746 (N_16746,N_16263,N_16440);
nand U16747 (N_16747,N_16276,N_16448);
nor U16748 (N_16748,N_16392,N_16424);
or U16749 (N_16749,N_16427,N_16361);
and U16750 (N_16750,N_16660,N_16748);
or U16751 (N_16751,N_16522,N_16686);
nand U16752 (N_16752,N_16541,N_16519);
nor U16753 (N_16753,N_16558,N_16638);
or U16754 (N_16754,N_16551,N_16639);
and U16755 (N_16755,N_16653,N_16706);
or U16756 (N_16756,N_16526,N_16509);
and U16757 (N_16757,N_16596,N_16722);
or U16758 (N_16758,N_16560,N_16671);
xor U16759 (N_16759,N_16702,N_16635);
xnor U16760 (N_16760,N_16725,N_16520);
and U16761 (N_16761,N_16680,N_16586);
nor U16762 (N_16762,N_16574,N_16713);
nand U16763 (N_16763,N_16597,N_16705);
nor U16764 (N_16764,N_16624,N_16636);
nand U16765 (N_16765,N_16626,N_16731);
nand U16766 (N_16766,N_16552,N_16678);
and U16767 (N_16767,N_16559,N_16614);
nor U16768 (N_16768,N_16701,N_16728);
xor U16769 (N_16769,N_16581,N_16715);
and U16770 (N_16770,N_16562,N_16647);
xor U16771 (N_16771,N_16504,N_16601);
and U16772 (N_16772,N_16696,N_16576);
xnor U16773 (N_16773,N_16683,N_16511);
xnor U16774 (N_16774,N_16727,N_16641);
nor U16775 (N_16775,N_16501,N_16606);
and U16776 (N_16776,N_16735,N_16707);
xnor U16777 (N_16777,N_16632,N_16536);
nand U16778 (N_16778,N_16712,N_16615);
nor U16779 (N_16779,N_16719,N_16741);
nand U16780 (N_16780,N_16546,N_16568);
nor U16781 (N_16781,N_16506,N_16625);
and U16782 (N_16782,N_16721,N_16613);
xor U16783 (N_16783,N_16555,N_16543);
nor U16784 (N_16784,N_16618,N_16666);
nand U16785 (N_16785,N_16667,N_16580);
and U16786 (N_16786,N_16532,N_16736);
nor U16787 (N_16787,N_16659,N_16740);
and U16788 (N_16788,N_16587,N_16648);
and U16789 (N_16789,N_16556,N_16577);
or U16790 (N_16790,N_16502,N_16658);
and U16791 (N_16791,N_16644,N_16621);
and U16792 (N_16792,N_16662,N_16542);
xor U16793 (N_16793,N_16684,N_16585);
nand U16794 (N_16794,N_16651,N_16533);
or U16795 (N_16795,N_16523,N_16718);
xor U16796 (N_16796,N_16665,N_16564);
nor U16797 (N_16797,N_16553,N_16646);
xor U16798 (N_16798,N_16578,N_16595);
and U16799 (N_16799,N_16744,N_16623);
nor U16800 (N_16800,N_16730,N_16611);
nor U16801 (N_16801,N_16570,N_16612);
and U16802 (N_16802,N_16616,N_16567);
nand U16803 (N_16803,N_16689,N_16609);
or U16804 (N_16804,N_16742,N_16729);
or U16805 (N_16805,N_16539,N_16720);
and U16806 (N_16806,N_16594,N_16517);
nand U16807 (N_16807,N_16513,N_16547);
nand U16808 (N_16808,N_16565,N_16535);
nand U16809 (N_16809,N_16540,N_16743);
xor U16810 (N_16810,N_16525,N_16619);
nand U16811 (N_16811,N_16685,N_16732);
nand U16812 (N_16812,N_16711,N_16500);
nand U16813 (N_16813,N_16608,N_16697);
or U16814 (N_16814,N_16668,N_16672);
nand U16815 (N_16815,N_16602,N_16717);
nand U16816 (N_16816,N_16627,N_16737);
nor U16817 (N_16817,N_16710,N_16703);
or U16818 (N_16818,N_16663,N_16692);
or U16819 (N_16819,N_16507,N_16657);
nor U16820 (N_16820,N_16512,N_16550);
or U16821 (N_16821,N_16548,N_16529);
xor U16822 (N_16822,N_16584,N_16588);
and U16823 (N_16823,N_16695,N_16749);
and U16824 (N_16824,N_16637,N_16654);
or U16825 (N_16825,N_16537,N_16591);
and U16826 (N_16826,N_16561,N_16571);
nor U16827 (N_16827,N_16634,N_16709);
or U16828 (N_16828,N_16549,N_16642);
and U16829 (N_16829,N_16505,N_16569);
nand U16830 (N_16830,N_16600,N_16734);
nand U16831 (N_16831,N_16714,N_16593);
and U16832 (N_16832,N_16677,N_16733);
nor U16833 (N_16833,N_16589,N_16746);
nand U16834 (N_16834,N_16592,N_16664);
nor U16835 (N_16835,N_16688,N_16690);
nand U16836 (N_16836,N_16628,N_16518);
nor U16837 (N_16837,N_16704,N_16528);
or U16838 (N_16838,N_16563,N_16516);
nand U16839 (N_16839,N_16524,N_16620);
or U16840 (N_16840,N_16652,N_16649);
or U16841 (N_16841,N_16515,N_16699);
or U16842 (N_16842,N_16554,N_16700);
xnor U16843 (N_16843,N_16566,N_16573);
nand U16844 (N_16844,N_16631,N_16617);
xnor U16845 (N_16845,N_16681,N_16557);
and U16846 (N_16846,N_16538,N_16622);
nand U16847 (N_16847,N_16726,N_16598);
or U16848 (N_16848,N_16514,N_16745);
or U16849 (N_16849,N_16503,N_16673);
nand U16850 (N_16850,N_16643,N_16661);
or U16851 (N_16851,N_16682,N_16530);
nor U16852 (N_16852,N_16521,N_16691);
nor U16853 (N_16853,N_16716,N_16534);
or U16854 (N_16854,N_16723,N_16544);
xor U16855 (N_16855,N_16640,N_16510);
and U16856 (N_16856,N_16675,N_16629);
xnor U16857 (N_16857,N_16545,N_16693);
xor U16858 (N_16858,N_16724,N_16698);
and U16859 (N_16859,N_16676,N_16669);
nand U16860 (N_16860,N_16582,N_16599);
nand U16861 (N_16861,N_16610,N_16694);
and U16862 (N_16862,N_16572,N_16583);
and U16863 (N_16863,N_16603,N_16607);
xor U16864 (N_16864,N_16630,N_16650);
nand U16865 (N_16865,N_16679,N_16655);
xor U16866 (N_16866,N_16739,N_16633);
and U16867 (N_16867,N_16527,N_16747);
nor U16868 (N_16868,N_16670,N_16531);
and U16869 (N_16869,N_16508,N_16579);
nor U16870 (N_16870,N_16604,N_16674);
or U16871 (N_16871,N_16645,N_16575);
nor U16872 (N_16872,N_16590,N_16605);
nand U16873 (N_16873,N_16656,N_16708);
or U16874 (N_16874,N_16687,N_16738);
nor U16875 (N_16875,N_16607,N_16563);
xnor U16876 (N_16876,N_16733,N_16672);
and U16877 (N_16877,N_16707,N_16587);
or U16878 (N_16878,N_16670,N_16719);
xor U16879 (N_16879,N_16526,N_16713);
nor U16880 (N_16880,N_16549,N_16714);
and U16881 (N_16881,N_16671,N_16579);
and U16882 (N_16882,N_16537,N_16506);
xnor U16883 (N_16883,N_16749,N_16628);
nand U16884 (N_16884,N_16600,N_16511);
nand U16885 (N_16885,N_16581,N_16726);
nor U16886 (N_16886,N_16574,N_16530);
xor U16887 (N_16887,N_16609,N_16541);
nand U16888 (N_16888,N_16602,N_16585);
nand U16889 (N_16889,N_16595,N_16620);
xor U16890 (N_16890,N_16696,N_16708);
nor U16891 (N_16891,N_16591,N_16579);
nand U16892 (N_16892,N_16601,N_16716);
and U16893 (N_16893,N_16667,N_16630);
and U16894 (N_16894,N_16635,N_16710);
nor U16895 (N_16895,N_16725,N_16527);
nor U16896 (N_16896,N_16670,N_16599);
or U16897 (N_16897,N_16703,N_16552);
xor U16898 (N_16898,N_16544,N_16740);
or U16899 (N_16899,N_16658,N_16654);
nand U16900 (N_16900,N_16723,N_16605);
and U16901 (N_16901,N_16571,N_16642);
nor U16902 (N_16902,N_16618,N_16583);
or U16903 (N_16903,N_16677,N_16695);
nor U16904 (N_16904,N_16677,N_16655);
and U16905 (N_16905,N_16615,N_16544);
or U16906 (N_16906,N_16658,N_16593);
xor U16907 (N_16907,N_16634,N_16501);
or U16908 (N_16908,N_16515,N_16540);
and U16909 (N_16909,N_16565,N_16545);
xor U16910 (N_16910,N_16645,N_16624);
and U16911 (N_16911,N_16621,N_16575);
or U16912 (N_16912,N_16521,N_16685);
nor U16913 (N_16913,N_16578,N_16606);
and U16914 (N_16914,N_16524,N_16715);
nor U16915 (N_16915,N_16573,N_16512);
xnor U16916 (N_16916,N_16690,N_16549);
xnor U16917 (N_16917,N_16588,N_16583);
nand U16918 (N_16918,N_16738,N_16740);
nor U16919 (N_16919,N_16580,N_16745);
or U16920 (N_16920,N_16707,N_16651);
nand U16921 (N_16921,N_16639,N_16734);
or U16922 (N_16922,N_16655,N_16641);
xnor U16923 (N_16923,N_16663,N_16681);
xor U16924 (N_16924,N_16722,N_16694);
nor U16925 (N_16925,N_16693,N_16618);
or U16926 (N_16926,N_16505,N_16586);
nand U16927 (N_16927,N_16614,N_16611);
xor U16928 (N_16928,N_16631,N_16684);
nand U16929 (N_16929,N_16619,N_16727);
nor U16930 (N_16930,N_16635,N_16603);
or U16931 (N_16931,N_16517,N_16748);
or U16932 (N_16932,N_16694,N_16506);
xnor U16933 (N_16933,N_16740,N_16624);
xor U16934 (N_16934,N_16712,N_16663);
or U16935 (N_16935,N_16508,N_16562);
or U16936 (N_16936,N_16629,N_16581);
nand U16937 (N_16937,N_16554,N_16605);
nand U16938 (N_16938,N_16563,N_16582);
or U16939 (N_16939,N_16529,N_16681);
nor U16940 (N_16940,N_16726,N_16545);
and U16941 (N_16941,N_16599,N_16568);
xor U16942 (N_16942,N_16593,N_16560);
nor U16943 (N_16943,N_16590,N_16712);
nand U16944 (N_16944,N_16587,N_16615);
nand U16945 (N_16945,N_16523,N_16697);
nand U16946 (N_16946,N_16519,N_16538);
xor U16947 (N_16947,N_16557,N_16599);
nor U16948 (N_16948,N_16520,N_16746);
and U16949 (N_16949,N_16704,N_16525);
or U16950 (N_16950,N_16708,N_16709);
xor U16951 (N_16951,N_16509,N_16691);
xnor U16952 (N_16952,N_16566,N_16631);
or U16953 (N_16953,N_16718,N_16740);
and U16954 (N_16954,N_16513,N_16717);
xor U16955 (N_16955,N_16605,N_16561);
xor U16956 (N_16956,N_16537,N_16511);
nor U16957 (N_16957,N_16724,N_16584);
nor U16958 (N_16958,N_16549,N_16534);
nor U16959 (N_16959,N_16505,N_16549);
nor U16960 (N_16960,N_16501,N_16516);
nand U16961 (N_16961,N_16737,N_16684);
and U16962 (N_16962,N_16533,N_16716);
nor U16963 (N_16963,N_16663,N_16710);
xnor U16964 (N_16964,N_16635,N_16723);
and U16965 (N_16965,N_16719,N_16575);
or U16966 (N_16966,N_16533,N_16722);
xnor U16967 (N_16967,N_16535,N_16674);
or U16968 (N_16968,N_16686,N_16597);
and U16969 (N_16969,N_16739,N_16647);
and U16970 (N_16970,N_16608,N_16664);
nand U16971 (N_16971,N_16626,N_16534);
nor U16972 (N_16972,N_16665,N_16630);
and U16973 (N_16973,N_16644,N_16687);
or U16974 (N_16974,N_16740,N_16589);
nand U16975 (N_16975,N_16681,N_16589);
nor U16976 (N_16976,N_16698,N_16697);
and U16977 (N_16977,N_16571,N_16583);
nand U16978 (N_16978,N_16553,N_16569);
or U16979 (N_16979,N_16700,N_16694);
nor U16980 (N_16980,N_16575,N_16544);
or U16981 (N_16981,N_16514,N_16605);
or U16982 (N_16982,N_16596,N_16676);
nand U16983 (N_16983,N_16629,N_16556);
nor U16984 (N_16984,N_16608,N_16704);
xnor U16985 (N_16985,N_16745,N_16508);
xor U16986 (N_16986,N_16719,N_16697);
and U16987 (N_16987,N_16602,N_16640);
xor U16988 (N_16988,N_16705,N_16545);
and U16989 (N_16989,N_16645,N_16726);
nand U16990 (N_16990,N_16655,N_16552);
nor U16991 (N_16991,N_16521,N_16576);
or U16992 (N_16992,N_16715,N_16717);
xnor U16993 (N_16993,N_16743,N_16592);
and U16994 (N_16994,N_16616,N_16610);
xnor U16995 (N_16995,N_16734,N_16738);
or U16996 (N_16996,N_16647,N_16505);
nand U16997 (N_16997,N_16687,N_16697);
xor U16998 (N_16998,N_16655,N_16663);
nand U16999 (N_16999,N_16728,N_16746);
and U17000 (N_17000,N_16759,N_16909);
and U17001 (N_17001,N_16978,N_16793);
or U17002 (N_17002,N_16987,N_16828);
xnor U17003 (N_17003,N_16833,N_16961);
or U17004 (N_17004,N_16901,N_16964);
and U17005 (N_17005,N_16829,N_16836);
nand U17006 (N_17006,N_16857,N_16785);
nor U17007 (N_17007,N_16900,N_16954);
and U17008 (N_17008,N_16960,N_16826);
nand U17009 (N_17009,N_16962,N_16877);
or U17010 (N_17010,N_16896,N_16846);
nand U17011 (N_17011,N_16819,N_16848);
and U17012 (N_17012,N_16970,N_16878);
and U17013 (N_17013,N_16980,N_16963);
nand U17014 (N_17014,N_16973,N_16906);
xor U17015 (N_17015,N_16843,N_16860);
nand U17016 (N_17016,N_16788,N_16940);
or U17017 (N_17017,N_16864,N_16892);
or U17018 (N_17018,N_16879,N_16989);
or U17019 (N_17019,N_16902,N_16827);
nor U17020 (N_17020,N_16981,N_16983);
nand U17021 (N_17021,N_16991,N_16905);
and U17022 (N_17022,N_16830,N_16899);
or U17023 (N_17023,N_16801,N_16931);
xnor U17024 (N_17024,N_16894,N_16769);
or U17025 (N_17025,N_16756,N_16893);
nor U17026 (N_17026,N_16881,N_16768);
xnor U17027 (N_17027,N_16751,N_16849);
and U17028 (N_17028,N_16992,N_16985);
xnor U17029 (N_17029,N_16949,N_16758);
nor U17030 (N_17030,N_16867,N_16927);
xnor U17031 (N_17031,N_16763,N_16839);
or U17032 (N_17032,N_16783,N_16859);
or U17033 (N_17033,N_16886,N_16911);
nor U17034 (N_17034,N_16873,N_16802);
nor U17035 (N_17035,N_16854,N_16773);
or U17036 (N_17036,N_16972,N_16816);
nand U17037 (N_17037,N_16998,N_16798);
nor U17038 (N_17038,N_16988,N_16795);
nand U17039 (N_17039,N_16806,N_16786);
nor U17040 (N_17040,N_16967,N_16999);
nand U17041 (N_17041,N_16868,N_16946);
and U17042 (N_17042,N_16957,N_16823);
or U17043 (N_17043,N_16924,N_16841);
nor U17044 (N_17044,N_16914,N_16814);
and U17045 (N_17045,N_16767,N_16789);
xnor U17046 (N_17046,N_16923,N_16969);
nand U17047 (N_17047,N_16907,N_16752);
or U17048 (N_17048,N_16938,N_16755);
and U17049 (N_17049,N_16955,N_16762);
nor U17050 (N_17050,N_16872,N_16869);
xor U17051 (N_17051,N_16822,N_16974);
or U17052 (N_17052,N_16837,N_16966);
and U17053 (N_17053,N_16765,N_16809);
xor U17054 (N_17054,N_16908,N_16920);
or U17055 (N_17055,N_16791,N_16831);
nand U17056 (N_17056,N_16956,N_16936);
or U17057 (N_17057,N_16889,N_16958);
xnor U17058 (N_17058,N_16904,N_16932);
nand U17059 (N_17059,N_16929,N_16817);
or U17060 (N_17060,N_16875,N_16820);
nor U17061 (N_17061,N_16891,N_16754);
and U17062 (N_17062,N_16910,N_16951);
and U17063 (N_17063,N_16794,N_16805);
nand U17064 (N_17064,N_16945,N_16876);
nand U17065 (N_17065,N_16774,N_16764);
xor U17066 (N_17066,N_16852,N_16871);
nand U17067 (N_17067,N_16842,N_16807);
nand U17068 (N_17068,N_16847,N_16979);
or U17069 (N_17069,N_16890,N_16855);
nor U17070 (N_17070,N_16779,N_16930);
xor U17071 (N_17071,N_16866,N_16898);
xnor U17072 (N_17072,N_16760,N_16861);
nor U17073 (N_17073,N_16797,N_16885);
xor U17074 (N_17074,N_16995,N_16821);
nor U17075 (N_17075,N_16778,N_16919);
or U17076 (N_17076,N_16916,N_16935);
nor U17077 (N_17077,N_16982,N_16853);
nand U17078 (N_17078,N_16825,N_16844);
nand U17079 (N_17079,N_16941,N_16968);
xnor U17080 (N_17080,N_16934,N_16813);
xnor U17081 (N_17081,N_16850,N_16766);
nor U17082 (N_17082,N_16921,N_16784);
nor U17083 (N_17083,N_16810,N_16808);
and U17084 (N_17084,N_16952,N_16928);
or U17085 (N_17085,N_16888,N_16942);
xnor U17086 (N_17086,N_16799,N_16757);
and U17087 (N_17087,N_16824,N_16753);
xor U17088 (N_17088,N_16917,N_16950);
or U17089 (N_17089,N_16939,N_16845);
nor U17090 (N_17090,N_16780,N_16965);
xor U17091 (N_17091,N_16777,N_16792);
xnor U17092 (N_17092,N_16947,N_16926);
xnor U17093 (N_17093,N_16975,N_16997);
and U17094 (N_17094,N_16986,N_16884);
or U17095 (N_17095,N_16770,N_16863);
xor U17096 (N_17096,N_16913,N_16925);
nand U17097 (N_17097,N_16787,N_16977);
nor U17098 (N_17098,N_16874,N_16856);
and U17099 (N_17099,N_16918,N_16944);
and U17100 (N_17100,N_16990,N_16771);
nand U17101 (N_17101,N_16761,N_16996);
nand U17102 (N_17102,N_16903,N_16840);
nor U17103 (N_17103,N_16976,N_16943);
nand U17104 (N_17104,N_16834,N_16804);
and U17105 (N_17105,N_16895,N_16796);
nand U17106 (N_17106,N_16959,N_16994);
nand U17107 (N_17107,N_16933,N_16912);
nand U17108 (N_17108,N_16835,N_16937);
xor U17109 (N_17109,N_16775,N_16811);
nor U17110 (N_17110,N_16915,N_16812);
xnor U17111 (N_17111,N_16897,N_16984);
nor U17112 (N_17112,N_16772,N_16815);
and U17113 (N_17113,N_16880,N_16858);
nand U17114 (N_17114,N_16971,N_16922);
nor U17115 (N_17115,N_16803,N_16782);
xor U17116 (N_17116,N_16832,N_16851);
nor U17117 (N_17117,N_16887,N_16781);
and U17118 (N_17118,N_16865,N_16993);
and U17119 (N_17119,N_16953,N_16838);
xnor U17120 (N_17120,N_16750,N_16800);
and U17121 (N_17121,N_16790,N_16870);
nand U17122 (N_17122,N_16883,N_16862);
or U17123 (N_17123,N_16882,N_16776);
nor U17124 (N_17124,N_16948,N_16818);
nand U17125 (N_17125,N_16782,N_16897);
or U17126 (N_17126,N_16988,N_16758);
xor U17127 (N_17127,N_16871,N_16937);
xor U17128 (N_17128,N_16885,N_16947);
nor U17129 (N_17129,N_16817,N_16824);
xor U17130 (N_17130,N_16780,N_16978);
nand U17131 (N_17131,N_16935,N_16839);
and U17132 (N_17132,N_16783,N_16812);
or U17133 (N_17133,N_16827,N_16967);
and U17134 (N_17134,N_16750,N_16994);
nand U17135 (N_17135,N_16959,N_16873);
and U17136 (N_17136,N_16971,N_16936);
nand U17137 (N_17137,N_16997,N_16813);
nand U17138 (N_17138,N_16913,N_16928);
nor U17139 (N_17139,N_16828,N_16901);
and U17140 (N_17140,N_16858,N_16983);
nand U17141 (N_17141,N_16892,N_16972);
nor U17142 (N_17142,N_16992,N_16903);
nand U17143 (N_17143,N_16978,N_16899);
xnor U17144 (N_17144,N_16780,N_16793);
nor U17145 (N_17145,N_16853,N_16838);
nand U17146 (N_17146,N_16909,N_16894);
and U17147 (N_17147,N_16772,N_16788);
nand U17148 (N_17148,N_16951,N_16780);
nand U17149 (N_17149,N_16756,N_16845);
nor U17150 (N_17150,N_16770,N_16812);
or U17151 (N_17151,N_16768,N_16806);
and U17152 (N_17152,N_16792,N_16880);
and U17153 (N_17153,N_16957,N_16880);
or U17154 (N_17154,N_16816,N_16990);
and U17155 (N_17155,N_16985,N_16806);
nor U17156 (N_17156,N_16965,N_16875);
xor U17157 (N_17157,N_16923,N_16993);
nand U17158 (N_17158,N_16774,N_16783);
nor U17159 (N_17159,N_16970,N_16984);
and U17160 (N_17160,N_16772,N_16896);
and U17161 (N_17161,N_16950,N_16992);
xnor U17162 (N_17162,N_16852,N_16985);
and U17163 (N_17163,N_16832,N_16776);
nand U17164 (N_17164,N_16931,N_16943);
nor U17165 (N_17165,N_16831,N_16865);
xor U17166 (N_17166,N_16917,N_16862);
nand U17167 (N_17167,N_16761,N_16976);
or U17168 (N_17168,N_16943,N_16923);
xnor U17169 (N_17169,N_16958,N_16897);
nor U17170 (N_17170,N_16805,N_16781);
or U17171 (N_17171,N_16874,N_16933);
nor U17172 (N_17172,N_16754,N_16805);
nor U17173 (N_17173,N_16762,N_16999);
or U17174 (N_17174,N_16760,N_16933);
or U17175 (N_17175,N_16971,N_16965);
nand U17176 (N_17176,N_16953,N_16994);
or U17177 (N_17177,N_16833,N_16790);
or U17178 (N_17178,N_16885,N_16777);
xnor U17179 (N_17179,N_16843,N_16812);
nand U17180 (N_17180,N_16768,N_16940);
xor U17181 (N_17181,N_16757,N_16838);
and U17182 (N_17182,N_16763,N_16817);
or U17183 (N_17183,N_16785,N_16893);
or U17184 (N_17184,N_16902,N_16786);
nor U17185 (N_17185,N_16959,N_16853);
or U17186 (N_17186,N_16960,N_16840);
or U17187 (N_17187,N_16927,N_16959);
nor U17188 (N_17188,N_16967,N_16862);
xor U17189 (N_17189,N_16776,N_16761);
nor U17190 (N_17190,N_16768,N_16847);
and U17191 (N_17191,N_16882,N_16778);
or U17192 (N_17192,N_16795,N_16827);
and U17193 (N_17193,N_16985,N_16796);
or U17194 (N_17194,N_16997,N_16885);
xnor U17195 (N_17195,N_16951,N_16895);
and U17196 (N_17196,N_16887,N_16814);
nor U17197 (N_17197,N_16811,N_16864);
or U17198 (N_17198,N_16852,N_16836);
xor U17199 (N_17199,N_16895,N_16885);
nor U17200 (N_17200,N_16991,N_16869);
nor U17201 (N_17201,N_16961,N_16872);
xnor U17202 (N_17202,N_16770,N_16768);
xnor U17203 (N_17203,N_16762,N_16802);
nor U17204 (N_17204,N_16778,N_16993);
and U17205 (N_17205,N_16948,N_16849);
nand U17206 (N_17206,N_16897,N_16975);
or U17207 (N_17207,N_16962,N_16967);
nor U17208 (N_17208,N_16886,N_16897);
nor U17209 (N_17209,N_16839,N_16863);
nand U17210 (N_17210,N_16796,N_16967);
nor U17211 (N_17211,N_16927,N_16947);
or U17212 (N_17212,N_16820,N_16853);
nand U17213 (N_17213,N_16854,N_16804);
and U17214 (N_17214,N_16775,N_16881);
or U17215 (N_17215,N_16825,N_16870);
and U17216 (N_17216,N_16886,N_16869);
nor U17217 (N_17217,N_16764,N_16979);
or U17218 (N_17218,N_16893,N_16833);
xor U17219 (N_17219,N_16813,N_16840);
or U17220 (N_17220,N_16829,N_16765);
nor U17221 (N_17221,N_16797,N_16953);
or U17222 (N_17222,N_16809,N_16891);
and U17223 (N_17223,N_16994,N_16951);
and U17224 (N_17224,N_16824,N_16764);
and U17225 (N_17225,N_16918,N_16928);
or U17226 (N_17226,N_16873,N_16962);
or U17227 (N_17227,N_16947,N_16804);
and U17228 (N_17228,N_16771,N_16925);
nor U17229 (N_17229,N_16963,N_16824);
nor U17230 (N_17230,N_16871,N_16848);
xor U17231 (N_17231,N_16947,N_16875);
and U17232 (N_17232,N_16947,N_16774);
nand U17233 (N_17233,N_16801,N_16924);
or U17234 (N_17234,N_16835,N_16983);
nand U17235 (N_17235,N_16919,N_16997);
and U17236 (N_17236,N_16930,N_16951);
xnor U17237 (N_17237,N_16997,N_16939);
nor U17238 (N_17238,N_16797,N_16848);
xor U17239 (N_17239,N_16751,N_16801);
nand U17240 (N_17240,N_16819,N_16953);
or U17241 (N_17241,N_16904,N_16902);
nand U17242 (N_17242,N_16870,N_16876);
and U17243 (N_17243,N_16814,N_16926);
xor U17244 (N_17244,N_16998,N_16878);
or U17245 (N_17245,N_16848,N_16980);
or U17246 (N_17246,N_16763,N_16879);
xnor U17247 (N_17247,N_16837,N_16857);
nor U17248 (N_17248,N_16831,N_16839);
or U17249 (N_17249,N_16842,N_16880);
nor U17250 (N_17250,N_17212,N_17012);
or U17251 (N_17251,N_17067,N_17209);
xor U17252 (N_17252,N_17243,N_17110);
and U17253 (N_17253,N_17004,N_17213);
and U17254 (N_17254,N_17094,N_17093);
nor U17255 (N_17255,N_17127,N_17028);
or U17256 (N_17256,N_17027,N_17114);
nand U17257 (N_17257,N_17052,N_17011);
nor U17258 (N_17258,N_17246,N_17106);
or U17259 (N_17259,N_17161,N_17136);
nand U17260 (N_17260,N_17063,N_17192);
nor U17261 (N_17261,N_17201,N_17214);
xnor U17262 (N_17262,N_17097,N_17072);
and U17263 (N_17263,N_17156,N_17245);
xnor U17264 (N_17264,N_17037,N_17077);
nand U17265 (N_17265,N_17112,N_17162);
nand U17266 (N_17266,N_17157,N_17155);
and U17267 (N_17267,N_17002,N_17150);
nor U17268 (N_17268,N_17239,N_17064);
nand U17269 (N_17269,N_17166,N_17070);
or U17270 (N_17270,N_17198,N_17111);
and U17271 (N_17271,N_17169,N_17146);
nand U17272 (N_17272,N_17230,N_17038);
nor U17273 (N_17273,N_17147,N_17091);
nor U17274 (N_17274,N_17119,N_17164);
nand U17275 (N_17275,N_17120,N_17102);
and U17276 (N_17276,N_17231,N_17203);
and U17277 (N_17277,N_17202,N_17086);
nor U17278 (N_17278,N_17189,N_17075);
nor U17279 (N_17279,N_17184,N_17177);
or U17280 (N_17280,N_17179,N_17148);
or U17281 (N_17281,N_17051,N_17099);
xnor U17282 (N_17282,N_17124,N_17207);
and U17283 (N_17283,N_17158,N_17024);
and U17284 (N_17284,N_17188,N_17105);
nand U17285 (N_17285,N_17168,N_17226);
or U17286 (N_17286,N_17137,N_17000);
or U17287 (N_17287,N_17204,N_17020);
xnor U17288 (N_17288,N_17101,N_17187);
and U17289 (N_17289,N_17066,N_17088);
and U17290 (N_17290,N_17109,N_17060);
nor U17291 (N_17291,N_17013,N_17001);
nor U17292 (N_17292,N_17030,N_17056);
nand U17293 (N_17293,N_17173,N_17135);
xnor U17294 (N_17294,N_17039,N_17116);
nand U17295 (N_17295,N_17005,N_17041);
nand U17296 (N_17296,N_17095,N_17074);
nand U17297 (N_17297,N_17160,N_17082);
nor U17298 (N_17298,N_17191,N_17104);
xor U17299 (N_17299,N_17218,N_17145);
or U17300 (N_17300,N_17085,N_17062);
xnor U17301 (N_17301,N_17032,N_17089);
xnor U17302 (N_17302,N_17221,N_17194);
nand U17303 (N_17303,N_17108,N_17199);
xor U17304 (N_17304,N_17205,N_17174);
or U17305 (N_17305,N_17073,N_17240);
or U17306 (N_17306,N_17176,N_17033);
and U17307 (N_17307,N_17183,N_17244);
and U17308 (N_17308,N_17196,N_17087);
or U17309 (N_17309,N_17128,N_17165);
nand U17310 (N_17310,N_17236,N_17098);
nand U17311 (N_17311,N_17009,N_17149);
and U17312 (N_17312,N_17055,N_17058);
nor U17313 (N_17313,N_17241,N_17224);
nor U17314 (N_17314,N_17131,N_17080);
or U17315 (N_17315,N_17228,N_17197);
xnor U17316 (N_17316,N_17132,N_17078);
nand U17317 (N_17317,N_17076,N_17185);
and U17318 (N_17318,N_17068,N_17096);
nor U17319 (N_17319,N_17152,N_17171);
xor U17320 (N_17320,N_17031,N_17061);
and U17321 (N_17321,N_17172,N_17021);
or U17322 (N_17322,N_17159,N_17014);
and U17323 (N_17323,N_17181,N_17222);
and U17324 (N_17324,N_17071,N_17069);
or U17325 (N_17325,N_17059,N_17232);
nand U17326 (N_17326,N_17193,N_17170);
xnor U17327 (N_17327,N_17216,N_17090);
and U17328 (N_17328,N_17122,N_17035);
xor U17329 (N_17329,N_17023,N_17040);
or U17330 (N_17330,N_17050,N_17123);
xnor U17331 (N_17331,N_17208,N_17019);
or U17332 (N_17332,N_17100,N_17084);
nor U17333 (N_17333,N_17010,N_17154);
xnor U17334 (N_17334,N_17219,N_17129);
nor U17335 (N_17335,N_17190,N_17015);
and U17336 (N_17336,N_17141,N_17107);
nor U17337 (N_17337,N_17079,N_17210);
and U17338 (N_17338,N_17235,N_17054);
nor U17339 (N_17339,N_17242,N_17036);
xnor U17340 (N_17340,N_17126,N_17034);
or U17341 (N_17341,N_17139,N_17217);
or U17342 (N_17342,N_17134,N_17045);
or U17343 (N_17343,N_17140,N_17048);
and U17344 (N_17344,N_17229,N_17081);
nor U17345 (N_17345,N_17225,N_17121);
and U17346 (N_17346,N_17180,N_17057);
and U17347 (N_17347,N_17065,N_17238);
and U17348 (N_17348,N_17003,N_17115);
xnor U17349 (N_17349,N_17133,N_17182);
nor U17350 (N_17350,N_17008,N_17223);
and U17351 (N_17351,N_17007,N_17206);
and U17352 (N_17352,N_17103,N_17200);
and U17353 (N_17353,N_17142,N_17248);
xor U17354 (N_17354,N_17049,N_17167);
nor U17355 (N_17355,N_17237,N_17227);
nor U17356 (N_17356,N_17022,N_17211);
and U17357 (N_17357,N_17153,N_17186);
or U17358 (N_17358,N_17025,N_17018);
nor U17359 (N_17359,N_17083,N_17195);
and U17360 (N_17360,N_17130,N_17151);
and U17361 (N_17361,N_17113,N_17016);
or U17362 (N_17362,N_17053,N_17117);
nand U17363 (N_17363,N_17006,N_17043);
nand U17364 (N_17364,N_17118,N_17215);
nor U17365 (N_17365,N_17178,N_17144);
or U17366 (N_17366,N_17175,N_17247);
or U17367 (N_17367,N_17092,N_17249);
nor U17368 (N_17368,N_17163,N_17044);
nor U17369 (N_17369,N_17042,N_17047);
nand U17370 (N_17370,N_17143,N_17220);
xnor U17371 (N_17371,N_17029,N_17046);
and U17372 (N_17372,N_17125,N_17138);
xnor U17373 (N_17373,N_17233,N_17017);
nand U17374 (N_17374,N_17026,N_17234);
nor U17375 (N_17375,N_17211,N_17075);
or U17376 (N_17376,N_17019,N_17030);
or U17377 (N_17377,N_17019,N_17189);
nand U17378 (N_17378,N_17098,N_17101);
nor U17379 (N_17379,N_17135,N_17094);
and U17380 (N_17380,N_17183,N_17115);
and U17381 (N_17381,N_17058,N_17232);
or U17382 (N_17382,N_17011,N_17061);
and U17383 (N_17383,N_17116,N_17155);
xor U17384 (N_17384,N_17082,N_17064);
or U17385 (N_17385,N_17177,N_17081);
and U17386 (N_17386,N_17174,N_17122);
or U17387 (N_17387,N_17085,N_17160);
xnor U17388 (N_17388,N_17128,N_17191);
xor U17389 (N_17389,N_17187,N_17097);
nand U17390 (N_17390,N_17127,N_17109);
or U17391 (N_17391,N_17121,N_17124);
xor U17392 (N_17392,N_17136,N_17179);
and U17393 (N_17393,N_17006,N_17215);
nand U17394 (N_17394,N_17071,N_17149);
nor U17395 (N_17395,N_17080,N_17114);
nor U17396 (N_17396,N_17002,N_17156);
nor U17397 (N_17397,N_17117,N_17061);
nor U17398 (N_17398,N_17095,N_17244);
and U17399 (N_17399,N_17031,N_17105);
nor U17400 (N_17400,N_17119,N_17171);
xnor U17401 (N_17401,N_17048,N_17043);
and U17402 (N_17402,N_17038,N_17078);
nor U17403 (N_17403,N_17203,N_17047);
xor U17404 (N_17404,N_17096,N_17023);
and U17405 (N_17405,N_17155,N_17196);
xor U17406 (N_17406,N_17020,N_17178);
and U17407 (N_17407,N_17127,N_17032);
nor U17408 (N_17408,N_17013,N_17022);
nor U17409 (N_17409,N_17033,N_17184);
xor U17410 (N_17410,N_17222,N_17057);
or U17411 (N_17411,N_17206,N_17171);
nor U17412 (N_17412,N_17078,N_17226);
or U17413 (N_17413,N_17189,N_17176);
xor U17414 (N_17414,N_17025,N_17170);
nor U17415 (N_17415,N_17181,N_17170);
or U17416 (N_17416,N_17068,N_17067);
or U17417 (N_17417,N_17052,N_17182);
nand U17418 (N_17418,N_17035,N_17055);
and U17419 (N_17419,N_17248,N_17035);
or U17420 (N_17420,N_17048,N_17142);
or U17421 (N_17421,N_17186,N_17041);
or U17422 (N_17422,N_17155,N_17043);
or U17423 (N_17423,N_17081,N_17237);
and U17424 (N_17424,N_17106,N_17030);
nor U17425 (N_17425,N_17184,N_17021);
nor U17426 (N_17426,N_17207,N_17144);
nand U17427 (N_17427,N_17200,N_17184);
xor U17428 (N_17428,N_17133,N_17223);
nand U17429 (N_17429,N_17034,N_17157);
xnor U17430 (N_17430,N_17212,N_17040);
nor U17431 (N_17431,N_17106,N_17157);
and U17432 (N_17432,N_17199,N_17135);
or U17433 (N_17433,N_17113,N_17230);
and U17434 (N_17434,N_17090,N_17056);
or U17435 (N_17435,N_17184,N_17104);
or U17436 (N_17436,N_17113,N_17220);
nor U17437 (N_17437,N_17090,N_17045);
or U17438 (N_17438,N_17226,N_17202);
xor U17439 (N_17439,N_17142,N_17136);
and U17440 (N_17440,N_17049,N_17115);
xnor U17441 (N_17441,N_17035,N_17185);
nor U17442 (N_17442,N_17054,N_17001);
nand U17443 (N_17443,N_17042,N_17054);
xor U17444 (N_17444,N_17080,N_17036);
xor U17445 (N_17445,N_17150,N_17151);
or U17446 (N_17446,N_17088,N_17126);
or U17447 (N_17447,N_17223,N_17119);
or U17448 (N_17448,N_17025,N_17080);
or U17449 (N_17449,N_17088,N_17120);
and U17450 (N_17450,N_17085,N_17153);
nor U17451 (N_17451,N_17045,N_17220);
xnor U17452 (N_17452,N_17234,N_17220);
nor U17453 (N_17453,N_17074,N_17104);
and U17454 (N_17454,N_17087,N_17068);
xnor U17455 (N_17455,N_17080,N_17054);
xor U17456 (N_17456,N_17231,N_17187);
nand U17457 (N_17457,N_17229,N_17177);
nor U17458 (N_17458,N_17206,N_17112);
or U17459 (N_17459,N_17156,N_17198);
nand U17460 (N_17460,N_17061,N_17087);
and U17461 (N_17461,N_17171,N_17009);
nor U17462 (N_17462,N_17220,N_17069);
xnor U17463 (N_17463,N_17172,N_17202);
nor U17464 (N_17464,N_17089,N_17222);
or U17465 (N_17465,N_17231,N_17216);
nand U17466 (N_17466,N_17209,N_17154);
nand U17467 (N_17467,N_17134,N_17026);
nand U17468 (N_17468,N_17023,N_17140);
and U17469 (N_17469,N_17222,N_17041);
nand U17470 (N_17470,N_17020,N_17233);
xor U17471 (N_17471,N_17037,N_17057);
or U17472 (N_17472,N_17094,N_17197);
or U17473 (N_17473,N_17077,N_17055);
nand U17474 (N_17474,N_17187,N_17201);
nor U17475 (N_17475,N_17247,N_17125);
or U17476 (N_17476,N_17211,N_17192);
and U17477 (N_17477,N_17085,N_17017);
xor U17478 (N_17478,N_17231,N_17225);
and U17479 (N_17479,N_17018,N_17223);
nor U17480 (N_17480,N_17014,N_17004);
nor U17481 (N_17481,N_17229,N_17030);
nor U17482 (N_17482,N_17138,N_17131);
nor U17483 (N_17483,N_17012,N_17240);
or U17484 (N_17484,N_17028,N_17247);
nor U17485 (N_17485,N_17235,N_17036);
xnor U17486 (N_17486,N_17177,N_17090);
nand U17487 (N_17487,N_17183,N_17235);
nand U17488 (N_17488,N_17133,N_17245);
nand U17489 (N_17489,N_17039,N_17082);
xnor U17490 (N_17490,N_17228,N_17198);
nand U17491 (N_17491,N_17022,N_17120);
and U17492 (N_17492,N_17210,N_17165);
or U17493 (N_17493,N_17031,N_17106);
nand U17494 (N_17494,N_17183,N_17140);
or U17495 (N_17495,N_17232,N_17147);
nor U17496 (N_17496,N_17135,N_17218);
nor U17497 (N_17497,N_17217,N_17200);
nor U17498 (N_17498,N_17143,N_17058);
xnor U17499 (N_17499,N_17118,N_17069);
xor U17500 (N_17500,N_17453,N_17334);
nor U17501 (N_17501,N_17486,N_17492);
xnor U17502 (N_17502,N_17276,N_17488);
nand U17503 (N_17503,N_17274,N_17422);
or U17504 (N_17504,N_17489,N_17449);
nand U17505 (N_17505,N_17436,N_17407);
xnor U17506 (N_17506,N_17278,N_17440);
nand U17507 (N_17507,N_17356,N_17326);
nand U17508 (N_17508,N_17448,N_17458);
and U17509 (N_17509,N_17343,N_17471);
and U17510 (N_17510,N_17462,N_17271);
nand U17511 (N_17511,N_17312,N_17338);
or U17512 (N_17512,N_17497,N_17258);
and U17513 (N_17513,N_17473,N_17275);
xnor U17514 (N_17514,N_17269,N_17266);
or U17515 (N_17515,N_17267,N_17482);
xnor U17516 (N_17516,N_17465,N_17369);
nor U17517 (N_17517,N_17336,N_17409);
and U17518 (N_17518,N_17364,N_17307);
nor U17519 (N_17519,N_17367,N_17273);
xor U17520 (N_17520,N_17253,N_17498);
or U17521 (N_17521,N_17260,N_17366);
nor U17522 (N_17522,N_17263,N_17328);
nand U17523 (N_17523,N_17353,N_17428);
or U17524 (N_17524,N_17327,N_17420);
or U17525 (N_17525,N_17375,N_17318);
or U17526 (N_17526,N_17388,N_17337);
nand U17527 (N_17527,N_17270,N_17329);
nor U17528 (N_17528,N_17426,N_17305);
nand U17529 (N_17529,N_17454,N_17324);
nand U17530 (N_17530,N_17401,N_17333);
and U17531 (N_17531,N_17394,N_17371);
nor U17532 (N_17532,N_17391,N_17309);
and U17533 (N_17533,N_17374,N_17279);
or U17534 (N_17534,N_17376,N_17405);
xnor U17535 (N_17535,N_17429,N_17325);
nor U17536 (N_17536,N_17302,N_17386);
xor U17537 (N_17537,N_17495,N_17250);
nor U17538 (N_17538,N_17413,N_17287);
or U17539 (N_17539,N_17314,N_17456);
nand U17540 (N_17540,N_17381,N_17423);
or U17541 (N_17541,N_17320,N_17424);
or U17542 (N_17542,N_17406,N_17351);
nand U17543 (N_17543,N_17444,N_17352);
or U17544 (N_17544,N_17288,N_17400);
and U17545 (N_17545,N_17331,N_17300);
or U17546 (N_17546,N_17304,N_17459);
and U17547 (N_17547,N_17355,N_17452);
and U17548 (N_17548,N_17340,N_17323);
nand U17549 (N_17549,N_17319,N_17435);
xor U17550 (N_17550,N_17335,N_17265);
nand U17551 (N_17551,N_17251,N_17468);
nor U17552 (N_17552,N_17308,N_17442);
or U17553 (N_17553,N_17280,N_17350);
xor U17554 (N_17554,N_17484,N_17354);
nand U17555 (N_17555,N_17349,N_17427);
nor U17556 (N_17556,N_17445,N_17430);
xnor U17557 (N_17557,N_17399,N_17415);
xnor U17558 (N_17558,N_17476,N_17363);
and U17559 (N_17559,N_17437,N_17293);
or U17560 (N_17560,N_17410,N_17358);
or U17561 (N_17561,N_17347,N_17262);
nand U17562 (N_17562,N_17383,N_17297);
nor U17563 (N_17563,N_17491,N_17438);
and U17564 (N_17564,N_17475,N_17342);
nand U17565 (N_17565,N_17461,N_17295);
and U17566 (N_17566,N_17480,N_17457);
and U17567 (N_17567,N_17421,N_17360);
or U17568 (N_17568,N_17313,N_17361);
and U17569 (N_17569,N_17447,N_17431);
nor U17570 (N_17570,N_17490,N_17306);
and U17571 (N_17571,N_17290,N_17433);
or U17572 (N_17572,N_17291,N_17359);
xnor U17573 (N_17573,N_17397,N_17432);
and U17574 (N_17574,N_17467,N_17344);
xor U17575 (N_17575,N_17402,N_17357);
or U17576 (N_17576,N_17483,N_17348);
nor U17577 (N_17577,N_17339,N_17418);
or U17578 (N_17578,N_17485,N_17494);
and U17579 (N_17579,N_17477,N_17254);
or U17580 (N_17580,N_17384,N_17256);
or U17581 (N_17581,N_17298,N_17463);
nor U17582 (N_17582,N_17434,N_17398);
or U17583 (N_17583,N_17368,N_17416);
and U17584 (N_17584,N_17332,N_17396);
or U17585 (N_17585,N_17460,N_17292);
or U17586 (N_17586,N_17479,N_17282);
xor U17587 (N_17587,N_17481,N_17439);
nand U17588 (N_17588,N_17496,N_17284);
nand U17589 (N_17589,N_17377,N_17310);
or U17590 (N_17590,N_17289,N_17277);
nand U17591 (N_17591,N_17255,N_17382);
xnor U17592 (N_17592,N_17311,N_17362);
or U17593 (N_17593,N_17372,N_17315);
nor U17594 (N_17594,N_17499,N_17330);
xnor U17595 (N_17595,N_17261,N_17487);
nor U17596 (N_17596,N_17451,N_17425);
nand U17597 (N_17597,N_17478,N_17268);
nor U17598 (N_17598,N_17294,N_17373);
xnor U17599 (N_17599,N_17419,N_17408);
nor U17600 (N_17600,N_17341,N_17412);
nand U17601 (N_17601,N_17301,N_17404);
and U17602 (N_17602,N_17286,N_17411);
nand U17603 (N_17603,N_17392,N_17464);
or U17604 (N_17604,N_17466,N_17321);
and U17605 (N_17605,N_17272,N_17414);
and U17606 (N_17606,N_17316,N_17252);
nand U17607 (N_17607,N_17296,N_17285);
xor U17608 (N_17608,N_17395,N_17303);
and U17609 (N_17609,N_17446,N_17469);
nand U17610 (N_17610,N_17387,N_17379);
nor U17611 (N_17611,N_17299,N_17470);
nand U17612 (N_17612,N_17389,N_17365);
and U17613 (N_17613,N_17370,N_17259);
xor U17614 (N_17614,N_17346,N_17443);
nor U17615 (N_17615,N_17317,N_17378);
xnor U17616 (N_17616,N_17385,N_17264);
or U17617 (N_17617,N_17345,N_17257);
xnor U17618 (N_17618,N_17281,N_17390);
and U17619 (N_17619,N_17441,N_17455);
nand U17620 (N_17620,N_17393,N_17472);
nor U17621 (N_17621,N_17380,N_17417);
and U17622 (N_17622,N_17450,N_17322);
and U17623 (N_17623,N_17403,N_17474);
xor U17624 (N_17624,N_17283,N_17493);
nor U17625 (N_17625,N_17409,N_17322);
nand U17626 (N_17626,N_17397,N_17481);
or U17627 (N_17627,N_17318,N_17301);
xnor U17628 (N_17628,N_17343,N_17392);
nand U17629 (N_17629,N_17253,N_17328);
xor U17630 (N_17630,N_17386,N_17337);
nor U17631 (N_17631,N_17385,N_17260);
nand U17632 (N_17632,N_17412,N_17371);
xnor U17633 (N_17633,N_17365,N_17452);
and U17634 (N_17634,N_17485,N_17460);
and U17635 (N_17635,N_17458,N_17433);
nand U17636 (N_17636,N_17454,N_17449);
xor U17637 (N_17637,N_17396,N_17470);
or U17638 (N_17638,N_17324,N_17458);
xor U17639 (N_17639,N_17258,N_17388);
and U17640 (N_17640,N_17404,N_17323);
nand U17641 (N_17641,N_17299,N_17252);
nand U17642 (N_17642,N_17318,N_17465);
nor U17643 (N_17643,N_17434,N_17481);
nand U17644 (N_17644,N_17279,N_17454);
nand U17645 (N_17645,N_17273,N_17296);
nor U17646 (N_17646,N_17258,N_17353);
nand U17647 (N_17647,N_17475,N_17378);
nand U17648 (N_17648,N_17250,N_17356);
or U17649 (N_17649,N_17476,N_17289);
xor U17650 (N_17650,N_17297,N_17406);
and U17651 (N_17651,N_17425,N_17334);
and U17652 (N_17652,N_17324,N_17280);
xnor U17653 (N_17653,N_17315,N_17429);
and U17654 (N_17654,N_17428,N_17324);
and U17655 (N_17655,N_17469,N_17367);
xor U17656 (N_17656,N_17385,N_17363);
nor U17657 (N_17657,N_17269,N_17337);
nor U17658 (N_17658,N_17310,N_17272);
and U17659 (N_17659,N_17344,N_17276);
xor U17660 (N_17660,N_17371,N_17434);
nand U17661 (N_17661,N_17416,N_17315);
or U17662 (N_17662,N_17309,N_17317);
nor U17663 (N_17663,N_17291,N_17311);
xnor U17664 (N_17664,N_17410,N_17388);
xnor U17665 (N_17665,N_17347,N_17429);
or U17666 (N_17666,N_17408,N_17386);
xor U17667 (N_17667,N_17376,N_17399);
nor U17668 (N_17668,N_17387,N_17456);
nor U17669 (N_17669,N_17397,N_17280);
nand U17670 (N_17670,N_17279,N_17464);
and U17671 (N_17671,N_17281,N_17289);
xor U17672 (N_17672,N_17333,N_17319);
or U17673 (N_17673,N_17339,N_17320);
nand U17674 (N_17674,N_17317,N_17492);
and U17675 (N_17675,N_17326,N_17350);
xor U17676 (N_17676,N_17498,N_17371);
or U17677 (N_17677,N_17456,N_17349);
nand U17678 (N_17678,N_17277,N_17446);
and U17679 (N_17679,N_17329,N_17324);
nor U17680 (N_17680,N_17261,N_17447);
xor U17681 (N_17681,N_17470,N_17289);
nand U17682 (N_17682,N_17273,N_17396);
nor U17683 (N_17683,N_17355,N_17458);
and U17684 (N_17684,N_17371,N_17496);
xnor U17685 (N_17685,N_17292,N_17372);
and U17686 (N_17686,N_17253,N_17286);
xnor U17687 (N_17687,N_17422,N_17388);
or U17688 (N_17688,N_17447,N_17429);
nor U17689 (N_17689,N_17289,N_17304);
nand U17690 (N_17690,N_17280,N_17490);
and U17691 (N_17691,N_17416,N_17348);
and U17692 (N_17692,N_17337,N_17492);
and U17693 (N_17693,N_17458,N_17380);
or U17694 (N_17694,N_17315,N_17473);
nand U17695 (N_17695,N_17339,N_17318);
nor U17696 (N_17696,N_17288,N_17377);
nand U17697 (N_17697,N_17262,N_17415);
nor U17698 (N_17698,N_17266,N_17284);
nor U17699 (N_17699,N_17473,N_17365);
and U17700 (N_17700,N_17442,N_17394);
and U17701 (N_17701,N_17456,N_17461);
nand U17702 (N_17702,N_17352,N_17445);
nor U17703 (N_17703,N_17496,N_17392);
nand U17704 (N_17704,N_17279,N_17476);
and U17705 (N_17705,N_17476,N_17342);
nor U17706 (N_17706,N_17450,N_17382);
or U17707 (N_17707,N_17317,N_17497);
or U17708 (N_17708,N_17456,N_17324);
xnor U17709 (N_17709,N_17308,N_17401);
or U17710 (N_17710,N_17415,N_17449);
and U17711 (N_17711,N_17386,N_17373);
nand U17712 (N_17712,N_17376,N_17425);
nand U17713 (N_17713,N_17325,N_17321);
or U17714 (N_17714,N_17436,N_17366);
xnor U17715 (N_17715,N_17271,N_17441);
nor U17716 (N_17716,N_17287,N_17483);
nor U17717 (N_17717,N_17471,N_17491);
or U17718 (N_17718,N_17349,N_17373);
nand U17719 (N_17719,N_17482,N_17346);
and U17720 (N_17720,N_17480,N_17388);
and U17721 (N_17721,N_17283,N_17482);
nand U17722 (N_17722,N_17266,N_17364);
or U17723 (N_17723,N_17447,N_17340);
nand U17724 (N_17724,N_17448,N_17384);
and U17725 (N_17725,N_17253,N_17259);
nor U17726 (N_17726,N_17270,N_17376);
xor U17727 (N_17727,N_17329,N_17354);
and U17728 (N_17728,N_17370,N_17415);
or U17729 (N_17729,N_17468,N_17265);
or U17730 (N_17730,N_17352,N_17254);
nor U17731 (N_17731,N_17371,N_17435);
nand U17732 (N_17732,N_17283,N_17253);
or U17733 (N_17733,N_17381,N_17443);
nand U17734 (N_17734,N_17341,N_17458);
and U17735 (N_17735,N_17360,N_17402);
or U17736 (N_17736,N_17360,N_17451);
nand U17737 (N_17737,N_17415,N_17405);
and U17738 (N_17738,N_17298,N_17466);
or U17739 (N_17739,N_17434,N_17290);
and U17740 (N_17740,N_17360,N_17383);
and U17741 (N_17741,N_17453,N_17388);
nor U17742 (N_17742,N_17387,N_17293);
xor U17743 (N_17743,N_17456,N_17444);
or U17744 (N_17744,N_17384,N_17424);
or U17745 (N_17745,N_17338,N_17259);
and U17746 (N_17746,N_17332,N_17421);
or U17747 (N_17747,N_17443,N_17476);
nor U17748 (N_17748,N_17259,N_17464);
and U17749 (N_17749,N_17471,N_17295);
nand U17750 (N_17750,N_17560,N_17717);
nor U17751 (N_17751,N_17625,N_17604);
xnor U17752 (N_17752,N_17571,N_17714);
nor U17753 (N_17753,N_17684,N_17616);
nor U17754 (N_17754,N_17622,N_17748);
and U17755 (N_17755,N_17536,N_17510);
nand U17756 (N_17756,N_17583,N_17648);
nand U17757 (N_17757,N_17600,N_17634);
nand U17758 (N_17758,N_17698,N_17561);
and U17759 (N_17759,N_17655,N_17525);
or U17760 (N_17760,N_17647,N_17545);
and U17761 (N_17761,N_17703,N_17578);
or U17762 (N_17762,N_17518,N_17743);
nand U17763 (N_17763,N_17738,N_17638);
nand U17764 (N_17764,N_17620,N_17736);
nor U17765 (N_17765,N_17547,N_17678);
xor U17766 (N_17766,N_17594,N_17606);
and U17767 (N_17767,N_17595,N_17500);
xnor U17768 (N_17768,N_17591,N_17696);
nand U17769 (N_17769,N_17633,N_17552);
xnor U17770 (N_17770,N_17701,N_17713);
and U17771 (N_17771,N_17746,N_17715);
nor U17772 (N_17772,N_17544,N_17687);
nand U17773 (N_17773,N_17659,N_17563);
nor U17774 (N_17774,N_17593,N_17501);
nand U17775 (N_17775,N_17601,N_17689);
nand U17776 (N_17776,N_17611,N_17586);
and U17777 (N_17777,N_17666,N_17677);
nand U17778 (N_17778,N_17539,N_17749);
nor U17779 (N_17779,N_17630,N_17671);
nand U17780 (N_17780,N_17619,N_17697);
or U17781 (N_17781,N_17681,N_17734);
nor U17782 (N_17782,N_17589,N_17683);
nor U17783 (N_17783,N_17679,N_17556);
or U17784 (N_17784,N_17688,N_17721);
or U17785 (N_17785,N_17641,N_17651);
or U17786 (N_17786,N_17657,N_17546);
and U17787 (N_17787,N_17555,N_17708);
or U17788 (N_17788,N_17632,N_17694);
and U17789 (N_17789,N_17509,N_17669);
xnor U17790 (N_17790,N_17613,N_17598);
and U17791 (N_17791,N_17540,N_17650);
xor U17792 (N_17792,N_17532,N_17720);
nor U17793 (N_17793,N_17605,N_17585);
nor U17794 (N_17794,N_17637,N_17596);
nand U17795 (N_17795,N_17513,N_17635);
or U17796 (N_17796,N_17549,N_17692);
and U17797 (N_17797,N_17642,N_17618);
nor U17798 (N_17798,N_17504,N_17639);
nand U17799 (N_17799,N_17723,N_17672);
nand U17800 (N_17800,N_17658,N_17534);
xnor U17801 (N_17801,N_17685,N_17514);
or U17802 (N_17802,N_17537,N_17739);
or U17803 (N_17803,N_17629,N_17624);
xnor U17804 (N_17804,N_17574,N_17573);
or U17805 (N_17805,N_17668,N_17542);
or U17806 (N_17806,N_17718,N_17538);
and U17807 (N_17807,N_17569,N_17654);
nor U17808 (N_17808,N_17646,N_17524);
or U17809 (N_17809,N_17680,N_17614);
or U17810 (N_17810,N_17609,N_17660);
or U17811 (N_17811,N_17568,N_17674);
nor U17812 (N_17812,N_17709,N_17607);
and U17813 (N_17813,N_17682,N_17732);
xor U17814 (N_17814,N_17516,N_17512);
nand U17815 (N_17815,N_17693,N_17575);
or U17816 (N_17816,N_17597,N_17704);
xnor U17817 (N_17817,N_17729,N_17554);
and U17818 (N_17818,N_17615,N_17608);
nand U17819 (N_17819,N_17565,N_17737);
nand U17820 (N_17820,N_17652,N_17640);
nor U17821 (N_17821,N_17588,N_17686);
xor U17822 (N_17822,N_17550,N_17741);
xnor U17823 (N_17823,N_17558,N_17747);
nand U17824 (N_17824,N_17725,N_17508);
nand U17825 (N_17825,N_17533,N_17735);
and U17826 (N_17826,N_17644,N_17699);
nand U17827 (N_17827,N_17645,N_17621);
nand U17828 (N_17828,N_17528,N_17700);
and U17829 (N_17829,N_17521,N_17522);
or U17830 (N_17830,N_17580,N_17590);
nor U17831 (N_17831,N_17502,N_17535);
xnor U17832 (N_17832,N_17527,N_17626);
and U17833 (N_17833,N_17530,N_17636);
nand U17834 (N_17834,N_17710,N_17567);
or U17835 (N_17835,N_17745,N_17690);
nand U17836 (N_17836,N_17531,N_17553);
xnor U17837 (N_17837,N_17592,N_17730);
xnor U17838 (N_17838,N_17662,N_17603);
nand U17839 (N_17839,N_17731,N_17551);
nor U17840 (N_17840,N_17577,N_17582);
nor U17841 (N_17841,N_17543,N_17566);
or U17842 (N_17842,N_17711,N_17503);
and U17843 (N_17843,N_17517,N_17726);
and U17844 (N_17844,N_17599,N_17649);
and U17845 (N_17845,N_17548,N_17612);
xor U17846 (N_17846,N_17673,N_17617);
nor U17847 (N_17847,N_17706,N_17520);
and U17848 (N_17848,N_17670,N_17695);
or U17849 (N_17849,N_17664,N_17505);
and U17850 (N_17850,N_17564,N_17665);
xnor U17851 (N_17851,N_17602,N_17661);
or U17852 (N_17852,N_17728,N_17722);
nand U17853 (N_17853,N_17576,N_17623);
nand U17854 (N_17854,N_17663,N_17707);
nand U17855 (N_17855,N_17572,N_17587);
nand U17856 (N_17856,N_17667,N_17702);
and U17857 (N_17857,N_17506,N_17643);
or U17858 (N_17858,N_17584,N_17740);
or U17859 (N_17859,N_17507,N_17742);
and U17860 (N_17860,N_17653,N_17719);
or U17861 (N_17861,N_17570,N_17511);
xor U17862 (N_17862,N_17676,N_17744);
nor U17863 (N_17863,N_17628,N_17581);
and U17864 (N_17864,N_17656,N_17529);
nor U17865 (N_17865,N_17557,N_17627);
xnor U17866 (N_17866,N_17675,N_17610);
xnor U17867 (N_17867,N_17515,N_17579);
nor U17868 (N_17868,N_17712,N_17562);
or U17869 (N_17869,N_17523,N_17631);
nor U17870 (N_17870,N_17519,N_17541);
nor U17871 (N_17871,N_17716,N_17733);
nor U17872 (N_17872,N_17559,N_17724);
nor U17873 (N_17873,N_17691,N_17727);
and U17874 (N_17874,N_17705,N_17526);
or U17875 (N_17875,N_17662,N_17743);
or U17876 (N_17876,N_17687,N_17606);
nand U17877 (N_17877,N_17676,N_17584);
nor U17878 (N_17878,N_17648,N_17724);
or U17879 (N_17879,N_17582,N_17627);
xnor U17880 (N_17880,N_17643,N_17714);
nor U17881 (N_17881,N_17748,N_17666);
nor U17882 (N_17882,N_17575,N_17551);
nor U17883 (N_17883,N_17636,N_17668);
xnor U17884 (N_17884,N_17530,N_17505);
or U17885 (N_17885,N_17575,N_17579);
and U17886 (N_17886,N_17533,N_17651);
nor U17887 (N_17887,N_17546,N_17715);
xor U17888 (N_17888,N_17636,N_17535);
and U17889 (N_17889,N_17726,N_17709);
xor U17890 (N_17890,N_17599,N_17717);
nor U17891 (N_17891,N_17736,N_17749);
xor U17892 (N_17892,N_17745,N_17709);
nand U17893 (N_17893,N_17506,N_17507);
nor U17894 (N_17894,N_17696,N_17726);
xnor U17895 (N_17895,N_17631,N_17567);
and U17896 (N_17896,N_17617,N_17588);
and U17897 (N_17897,N_17544,N_17625);
and U17898 (N_17898,N_17520,N_17656);
or U17899 (N_17899,N_17652,N_17585);
xor U17900 (N_17900,N_17534,N_17607);
nor U17901 (N_17901,N_17721,N_17640);
and U17902 (N_17902,N_17668,N_17622);
and U17903 (N_17903,N_17544,N_17657);
xor U17904 (N_17904,N_17639,N_17619);
and U17905 (N_17905,N_17707,N_17617);
or U17906 (N_17906,N_17609,N_17508);
nor U17907 (N_17907,N_17628,N_17724);
and U17908 (N_17908,N_17692,N_17531);
and U17909 (N_17909,N_17664,N_17550);
or U17910 (N_17910,N_17588,N_17723);
nand U17911 (N_17911,N_17530,N_17621);
or U17912 (N_17912,N_17519,N_17616);
xor U17913 (N_17913,N_17597,N_17552);
xor U17914 (N_17914,N_17582,N_17541);
and U17915 (N_17915,N_17589,N_17617);
xor U17916 (N_17916,N_17589,N_17516);
nor U17917 (N_17917,N_17684,N_17748);
and U17918 (N_17918,N_17557,N_17620);
xnor U17919 (N_17919,N_17732,N_17585);
and U17920 (N_17920,N_17548,N_17528);
or U17921 (N_17921,N_17697,N_17595);
nand U17922 (N_17922,N_17726,N_17539);
xnor U17923 (N_17923,N_17535,N_17675);
nand U17924 (N_17924,N_17641,N_17506);
and U17925 (N_17925,N_17543,N_17624);
xor U17926 (N_17926,N_17612,N_17637);
or U17927 (N_17927,N_17516,N_17652);
or U17928 (N_17928,N_17669,N_17696);
nand U17929 (N_17929,N_17636,N_17680);
nand U17930 (N_17930,N_17524,N_17702);
and U17931 (N_17931,N_17617,N_17700);
nand U17932 (N_17932,N_17719,N_17605);
and U17933 (N_17933,N_17709,N_17738);
xor U17934 (N_17934,N_17738,N_17556);
nor U17935 (N_17935,N_17684,N_17646);
xor U17936 (N_17936,N_17730,N_17707);
xor U17937 (N_17937,N_17641,N_17672);
and U17938 (N_17938,N_17652,N_17725);
nor U17939 (N_17939,N_17719,N_17671);
and U17940 (N_17940,N_17700,N_17689);
nor U17941 (N_17941,N_17689,N_17708);
or U17942 (N_17942,N_17690,N_17686);
xor U17943 (N_17943,N_17579,N_17696);
and U17944 (N_17944,N_17537,N_17702);
and U17945 (N_17945,N_17669,N_17629);
xor U17946 (N_17946,N_17579,N_17527);
nand U17947 (N_17947,N_17678,N_17588);
or U17948 (N_17948,N_17605,N_17681);
nand U17949 (N_17949,N_17733,N_17600);
nor U17950 (N_17950,N_17539,N_17705);
and U17951 (N_17951,N_17639,N_17643);
nor U17952 (N_17952,N_17566,N_17541);
or U17953 (N_17953,N_17539,N_17521);
and U17954 (N_17954,N_17645,N_17571);
nand U17955 (N_17955,N_17588,N_17630);
or U17956 (N_17956,N_17542,N_17533);
nor U17957 (N_17957,N_17693,N_17594);
nand U17958 (N_17958,N_17695,N_17529);
and U17959 (N_17959,N_17739,N_17727);
or U17960 (N_17960,N_17726,N_17523);
and U17961 (N_17961,N_17721,N_17534);
or U17962 (N_17962,N_17656,N_17508);
xor U17963 (N_17963,N_17540,N_17572);
xnor U17964 (N_17964,N_17675,N_17564);
xor U17965 (N_17965,N_17538,N_17501);
nor U17966 (N_17966,N_17508,N_17551);
or U17967 (N_17967,N_17537,N_17647);
nor U17968 (N_17968,N_17551,N_17737);
nand U17969 (N_17969,N_17721,N_17741);
nor U17970 (N_17970,N_17515,N_17548);
and U17971 (N_17971,N_17723,N_17557);
or U17972 (N_17972,N_17654,N_17531);
nand U17973 (N_17973,N_17542,N_17700);
xor U17974 (N_17974,N_17599,N_17511);
and U17975 (N_17975,N_17718,N_17672);
or U17976 (N_17976,N_17705,N_17746);
nor U17977 (N_17977,N_17700,N_17597);
nor U17978 (N_17978,N_17723,N_17687);
or U17979 (N_17979,N_17507,N_17650);
xor U17980 (N_17980,N_17566,N_17669);
nand U17981 (N_17981,N_17676,N_17555);
nand U17982 (N_17982,N_17591,N_17535);
nand U17983 (N_17983,N_17748,N_17626);
xnor U17984 (N_17984,N_17614,N_17601);
or U17985 (N_17985,N_17664,N_17615);
xor U17986 (N_17986,N_17637,N_17638);
nor U17987 (N_17987,N_17542,N_17717);
nand U17988 (N_17988,N_17547,N_17717);
xor U17989 (N_17989,N_17669,N_17641);
and U17990 (N_17990,N_17639,N_17600);
or U17991 (N_17991,N_17543,N_17713);
and U17992 (N_17992,N_17569,N_17560);
or U17993 (N_17993,N_17696,N_17748);
and U17994 (N_17994,N_17527,N_17703);
xnor U17995 (N_17995,N_17575,N_17743);
nor U17996 (N_17996,N_17736,N_17530);
xor U17997 (N_17997,N_17584,N_17529);
xnor U17998 (N_17998,N_17535,N_17651);
xnor U17999 (N_17999,N_17576,N_17684);
or U18000 (N_18000,N_17929,N_17756);
and U18001 (N_18001,N_17826,N_17880);
nand U18002 (N_18002,N_17981,N_17940);
nand U18003 (N_18003,N_17989,N_17785);
xnor U18004 (N_18004,N_17824,N_17985);
nor U18005 (N_18005,N_17829,N_17848);
or U18006 (N_18006,N_17791,N_17978);
xor U18007 (N_18007,N_17926,N_17953);
nand U18008 (N_18008,N_17818,N_17762);
nor U18009 (N_18009,N_17997,N_17776);
and U18010 (N_18010,N_17781,N_17951);
or U18011 (N_18011,N_17778,N_17758);
or U18012 (N_18012,N_17918,N_17806);
nand U18013 (N_18013,N_17939,N_17982);
xor U18014 (N_18014,N_17830,N_17854);
or U18015 (N_18015,N_17761,N_17919);
nand U18016 (N_18016,N_17901,N_17965);
and U18017 (N_18017,N_17960,N_17879);
xor U18018 (N_18018,N_17902,N_17899);
and U18019 (N_18019,N_17796,N_17755);
and U18020 (N_18020,N_17890,N_17921);
nand U18021 (N_18021,N_17937,N_17786);
and U18022 (N_18022,N_17993,N_17999);
or U18023 (N_18023,N_17764,N_17843);
and U18024 (N_18024,N_17840,N_17851);
and U18025 (N_18025,N_17831,N_17979);
xor U18026 (N_18026,N_17819,N_17892);
nand U18027 (N_18027,N_17842,N_17906);
or U18028 (N_18028,N_17910,N_17948);
nor U18029 (N_18029,N_17904,N_17774);
nand U18030 (N_18030,N_17907,N_17779);
or U18031 (N_18031,N_17784,N_17964);
and U18032 (N_18032,N_17752,N_17810);
nor U18033 (N_18033,N_17980,N_17945);
or U18034 (N_18034,N_17827,N_17861);
nand U18035 (N_18035,N_17967,N_17805);
xor U18036 (N_18036,N_17927,N_17911);
xor U18037 (N_18037,N_17971,N_17941);
nand U18038 (N_18038,N_17789,N_17994);
or U18039 (N_18039,N_17894,N_17828);
or U18040 (N_18040,N_17770,N_17913);
xnor U18041 (N_18041,N_17923,N_17874);
and U18042 (N_18042,N_17962,N_17991);
and U18043 (N_18043,N_17782,N_17849);
xnor U18044 (N_18044,N_17969,N_17812);
xnor U18045 (N_18045,N_17920,N_17833);
and U18046 (N_18046,N_17869,N_17792);
nand U18047 (N_18047,N_17825,N_17814);
nand U18048 (N_18048,N_17905,N_17817);
xnor U18049 (N_18049,N_17775,N_17928);
or U18050 (N_18050,N_17803,N_17832);
xor U18051 (N_18051,N_17959,N_17887);
xor U18052 (N_18052,N_17858,N_17820);
xnor U18053 (N_18053,N_17790,N_17875);
and U18054 (N_18054,N_17877,N_17788);
and U18055 (N_18055,N_17798,N_17841);
nor U18056 (N_18056,N_17772,N_17963);
or U18057 (N_18057,N_17915,N_17973);
nand U18058 (N_18058,N_17765,N_17942);
xor U18059 (N_18059,N_17751,N_17924);
nor U18060 (N_18060,N_17768,N_17972);
nor U18061 (N_18061,N_17816,N_17996);
nand U18062 (N_18062,N_17931,N_17783);
nand U18063 (N_18063,N_17836,N_17896);
and U18064 (N_18064,N_17865,N_17970);
and U18065 (N_18065,N_17864,N_17780);
xnor U18066 (N_18066,N_17850,N_17838);
and U18067 (N_18067,N_17860,N_17800);
xor U18068 (N_18068,N_17955,N_17922);
xor U18069 (N_18069,N_17908,N_17898);
and U18070 (N_18070,N_17797,N_17794);
xor U18071 (N_18071,N_17844,N_17799);
and U18072 (N_18072,N_17750,N_17754);
or U18073 (N_18073,N_17958,N_17807);
nor U18074 (N_18074,N_17802,N_17900);
and U18075 (N_18075,N_17847,N_17975);
nand U18076 (N_18076,N_17916,N_17938);
nand U18077 (N_18077,N_17866,N_17852);
xnor U18078 (N_18078,N_17873,N_17884);
and U18079 (N_18079,N_17809,N_17952);
or U18080 (N_18080,N_17863,N_17995);
or U18081 (N_18081,N_17871,N_17855);
and U18082 (N_18082,N_17769,N_17897);
xnor U18083 (N_18083,N_17823,N_17974);
nor U18084 (N_18084,N_17808,N_17881);
nor U18085 (N_18085,N_17857,N_17815);
nand U18086 (N_18086,N_17976,N_17932);
xor U18087 (N_18087,N_17757,N_17767);
nand U18088 (N_18088,N_17990,N_17947);
xor U18089 (N_18089,N_17912,N_17771);
nand U18090 (N_18090,N_17867,N_17956);
nand U18091 (N_18091,N_17760,N_17853);
or U18092 (N_18092,N_17801,N_17903);
nor U18093 (N_18093,N_17773,N_17883);
and U18094 (N_18094,N_17998,N_17862);
and U18095 (N_18095,N_17968,N_17909);
or U18096 (N_18096,N_17984,N_17944);
and U18097 (N_18097,N_17961,N_17804);
xor U18098 (N_18098,N_17917,N_17846);
nor U18099 (N_18099,N_17845,N_17914);
xor U18100 (N_18100,N_17885,N_17868);
and U18101 (N_18101,N_17886,N_17950);
nor U18102 (N_18102,N_17895,N_17856);
nor U18103 (N_18103,N_17777,N_17787);
or U18104 (N_18104,N_17763,N_17793);
nand U18105 (N_18105,N_17878,N_17966);
nor U18106 (N_18106,N_17925,N_17766);
and U18107 (N_18107,N_17891,N_17949);
nand U18108 (N_18108,N_17882,N_17933);
nand U18109 (N_18109,N_17834,N_17977);
nand U18110 (N_18110,N_17813,N_17943);
or U18111 (N_18111,N_17986,N_17839);
nor U18112 (N_18112,N_17837,N_17889);
xnor U18113 (N_18113,N_17821,N_17753);
and U18114 (N_18114,N_17893,N_17936);
nand U18115 (N_18115,N_17988,N_17888);
xnor U18116 (N_18116,N_17930,N_17957);
and U18117 (N_18117,N_17946,N_17876);
xnor U18118 (N_18118,N_17992,N_17835);
nor U18119 (N_18119,N_17872,N_17759);
xor U18120 (N_18120,N_17987,N_17822);
and U18121 (N_18121,N_17811,N_17935);
nand U18122 (N_18122,N_17983,N_17934);
xor U18123 (N_18123,N_17859,N_17795);
or U18124 (N_18124,N_17870,N_17954);
nor U18125 (N_18125,N_17756,N_17900);
nand U18126 (N_18126,N_17910,N_17822);
nand U18127 (N_18127,N_17908,N_17888);
nand U18128 (N_18128,N_17820,N_17904);
nor U18129 (N_18129,N_17847,N_17878);
or U18130 (N_18130,N_17841,N_17760);
or U18131 (N_18131,N_17975,N_17972);
xor U18132 (N_18132,N_17992,N_17883);
nor U18133 (N_18133,N_17900,N_17933);
nand U18134 (N_18134,N_17751,N_17756);
nor U18135 (N_18135,N_17913,N_17988);
xor U18136 (N_18136,N_17821,N_17951);
and U18137 (N_18137,N_17906,N_17775);
xor U18138 (N_18138,N_17817,N_17956);
nand U18139 (N_18139,N_17978,N_17927);
and U18140 (N_18140,N_17902,N_17950);
nand U18141 (N_18141,N_17981,N_17909);
and U18142 (N_18142,N_17776,N_17846);
nor U18143 (N_18143,N_17853,N_17996);
xor U18144 (N_18144,N_17930,N_17984);
or U18145 (N_18145,N_17889,N_17954);
xnor U18146 (N_18146,N_17824,N_17797);
and U18147 (N_18147,N_17936,N_17945);
nand U18148 (N_18148,N_17991,N_17957);
or U18149 (N_18149,N_17908,N_17837);
or U18150 (N_18150,N_17814,N_17990);
nor U18151 (N_18151,N_17914,N_17878);
nand U18152 (N_18152,N_17791,N_17971);
and U18153 (N_18153,N_17915,N_17867);
and U18154 (N_18154,N_17755,N_17788);
nand U18155 (N_18155,N_17863,N_17969);
xnor U18156 (N_18156,N_17882,N_17957);
xnor U18157 (N_18157,N_17958,N_17756);
xnor U18158 (N_18158,N_17891,N_17850);
xnor U18159 (N_18159,N_17932,N_17879);
xnor U18160 (N_18160,N_17891,N_17907);
and U18161 (N_18161,N_17801,N_17930);
nor U18162 (N_18162,N_17888,N_17781);
and U18163 (N_18163,N_17899,N_17924);
or U18164 (N_18164,N_17877,N_17967);
and U18165 (N_18165,N_17826,N_17913);
and U18166 (N_18166,N_17901,N_17983);
nand U18167 (N_18167,N_17829,N_17921);
xnor U18168 (N_18168,N_17830,N_17792);
nand U18169 (N_18169,N_17754,N_17920);
nand U18170 (N_18170,N_17874,N_17886);
nand U18171 (N_18171,N_17875,N_17827);
or U18172 (N_18172,N_17821,N_17960);
nand U18173 (N_18173,N_17865,N_17906);
nand U18174 (N_18174,N_17830,N_17819);
nand U18175 (N_18175,N_17879,N_17939);
and U18176 (N_18176,N_17948,N_17813);
or U18177 (N_18177,N_17789,N_17828);
and U18178 (N_18178,N_17899,N_17962);
nor U18179 (N_18179,N_17788,N_17921);
xor U18180 (N_18180,N_17777,N_17830);
or U18181 (N_18181,N_17979,N_17752);
nand U18182 (N_18182,N_17838,N_17845);
or U18183 (N_18183,N_17827,N_17803);
or U18184 (N_18184,N_17973,N_17982);
and U18185 (N_18185,N_17829,N_17940);
nor U18186 (N_18186,N_17863,N_17845);
nand U18187 (N_18187,N_17789,N_17901);
nor U18188 (N_18188,N_17794,N_17848);
xnor U18189 (N_18189,N_17983,N_17894);
or U18190 (N_18190,N_17879,N_17816);
xor U18191 (N_18191,N_17808,N_17929);
nor U18192 (N_18192,N_17770,N_17782);
or U18193 (N_18193,N_17955,N_17993);
or U18194 (N_18194,N_17811,N_17861);
nor U18195 (N_18195,N_17898,N_17792);
nand U18196 (N_18196,N_17934,N_17793);
nor U18197 (N_18197,N_17916,N_17885);
or U18198 (N_18198,N_17973,N_17882);
nand U18199 (N_18199,N_17751,N_17801);
nand U18200 (N_18200,N_17967,N_17917);
and U18201 (N_18201,N_17897,N_17779);
or U18202 (N_18202,N_17886,N_17949);
nand U18203 (N_18203,N_17793,N_17832);
or U18204 (N_18204,N_17907,N_17875);
and U18205 (N_18205,N_17902,N_17904);
and U18206 (N_18206,N_17796,N_17847);
or U18207 (N_18207,N_17894,N_17897);
xor U18208 (N_18208,N_17991,N_17770);
xnor U18209 (N_18209,N_17758,N_17845);
xnor U18210 (N_18210,N_17901,N_17803);
and U18211 (N_18211,N_17949,N_17888);
nor U18212 (N_18212,N_17912,N_17897);
xnor U18213 (N_18213,N_17801,N_17967);
and U18214 (N_18214,N_17852,N_17972);
and U18215 (N_18215,N_17761,N_17769);
xnor U18216 (N_18216,N_17777,N_17835);
nand U18217 (N_18217,N_17872,N_17851);
nor U18218 (N_18218,N_17885,N_17784);
nand U18219 (N_18219,N_17892,N_17859);
or U18220 (N_18220,N_17925,N_17818);
and U18221 (N_18221,N_17954,N_17794);
and U18222 (N_18222,N_17977,N_17774);
or U18223 (N_18223,N_17807,N_17968);
nand U18224 (N_18224,N_17797,N_17948);
xor U18225 (N_18225,N_17971,N_17767);
or U18226 (N_18226,N_17896,N_17840);
nand U18227 (N_18227,N_17970,N_17916);
nand U18228 (N_18228,N_17998,N_17880);
xor U18229 (N_18229,N_17838,N_17996);
xnor U18230 (N_18230,N_17968,N_17804);
xnor U18231 (N_18231,N_17983,N_17862);
and U18232 (N_18232,N_17765,N_17884);
or U18233 (N_18233,N_17808,N_17965);
nor U18234 (N_18234,N_17765,N_17866);
nand U18235 (N_18235,N_17870,N_17780);
and U18236 (N_18236,N_17828,N_17854);
nor U18237 (N_18237,N_17906,N_17952);
nor U18238 (N_18238,N_17894,N_17886);
nor U18239 (N_18239,N_17907,N_17766);
and U18240 (N_18240,N_17832,N_17787);
and U18241 (N_18241,N_17974,N_17987);
nor U18242 (N_18242,N_17998,N_17889);
or U18243 (N_18243,N_17940,N_17901);
xor U18244 (N_18244,N_17835,N_17934);
or U18245 (N_18245,N_17802,N_17826);
nor U18246 (N_18246,N_17864,N_17753);
nor U18247 (N_18247,N_17780,N_17954);
and U18248 (N_18248,N_17783,N_17894);
nand U18249 (N_18249,N_17943,N_17759);
xor U18250 (N_18250,N_18108,N_18103);
or U18251 (N_18251,N_18219,N_18195);
or U18252 (N_18252,N_18058,N_18085);
nor U18253 (N_18253,N_18158,N_18107);
nor U18254 (N_18254,N_18201,N_18057);
nor U18255 (N_18255,N_18050,N_18032);
nand U18256 (N_18256,N_18213,N_18168);
and U18257 (N_18257,N_18084,N_18088);
and U18258 (N_18258,N_18031,N_18020);
or U18259 (N_18259,N_18115,N_18000);
nor U18260 (N_18260,N_18045,N_18124);
xor U18261 (N_18261,N_18118,N_18191);
or U18262 (N_18262,N_18221,N_18049);
xor U18263 (N_18263,N_18178,N_18038);
or U18264 (N_18264,N_18006,N_18003);
and U18265 (N_18265,N_18225,N_18034);
nand U18266 (N_18266,N_18017,N_18236);
and U18267 (N_18267,N_18206,N_18153);
nor U18268 (N_18268,N_18177,N_18184);
nor U18269 (N_18269,N_18069,N_18146);
xor U18270 (N_18270,N_18217,N_18144);
and U18271 (N_18271,N_18176,N_18162);
nand U18272 (N_18272,N_18052,N_18222);
or U18273 (N_18273,N_18143,N_18133);
nand U18274 (N_18274,N_18248,N_18102);
nor U18275 (N_18275,N_18029,N_18033);
xor U18276 (N_18276,N_18012,N_18204);
nand U18277 (N_18277,N_18190,N_18086);
nand U18278 (N_18278,N_18099,N_18189);
nand U18279 (N_18279,N_18185,N_18224);
nor U18280 (N_18280,N_18125,N_18170);
nor U18281 (N_18281,N_18130,N_18200);
xnor U18282 (N_18282,N_18030,N_18087);
or U18283 (N_18283,N_18209,N_18041);
nand U18284 (N_18284,N_18002,N_18043);
xnor U18285 (N_18285,N_18132,N_18167);
and U18286 (N_18286,N_18244,N_18098);
nand U18287 (N_18287,N_18120,N_18110);
xor U18288 (N_18288,N_18181,N_18090);
xnor U18289 (N_18289,N_18059,N_18161);
and U18290 (N_18290,N_18060,N_18121);
xnor U18291 (N_18291,N_18051,N_18235);
and U18292 (N_18292,N_18216,N_18066);
nor U18293 (N_18293,N_18027,N_18117);
nor U18294 (N_18294,N_18054,N_18021);
or U18295 (N_18295,N_18135,N_18089);
and U18296 (N_18296,N_18065,N_18123);
or U18297 (N_18297,N_18242,N_18077);
and U18298 (N_18298,N_18180,N_18228);
xor U18299 (N_18299,N_18232,N_18005);
or U18300 (N_18300,N_18151,N_18068);
or U18301 (N_18301,N_18009,N_18053);
xor U18302 (N_18302,N_18091,N_18014);
and U18303 (N_18303,N_18187,N_18172);
xor U18304 (N_18304,N_18202,N_18067);
xnor U18305 (N_18305,N_18212,N_18138);
nor U18306 (N_18306,N_18198,N_18171);
nand U18307 (N_18307,N_18223,N_18105);
nand U18308 (N_18308,N_18145,N_18082);
nand U18309 (N_18309,N_18131,N_18015);
xor U18310 (N_18310,N_18055,N_18197);
xor U18311 (N_18311,N_18156,N_18239);
and U18312 (N_18312,N_18079,N_18164);
xor U18313 (N_18313,N_18016,N_18022);
and U18314 (N_18314,N_18104,N_18147);
nand U18315 (N_18315,N_18010,N_18205);
nand U18316 (N_18316,N_18095,N_18196);
and U18317 (N_18317,N_18136,N_18100);
or U18318 (N_18318,N_18119,N_18234);
and U18319 (N_18319,N_18063,N_18149);
nand U18320 (N_18320,N_18193,N_18159);
and U18321 (N_18321,N_18246,N_18064);
and U18322 (N_18322,N_18179,N_18194);
or U18323 (N_18323,N_18163,N_18062);
xnor U18324 (N_18324,N_18243,N_18019);
nand U18325 (N_18325,N_18111,N_18046);
nand U18326 (N_18326,N_18109,N_18192);
and U18327 (N_18327,N_18230,N_18044);
or U18328 (N_18328,N_18233,N_18011);
xor U18329 (N_18329,N_18070,N_18214);
xor U18330 (N_18330,N_18116,N_18028);
and U18331 (N_18331,N_18227,N_18231);
and U18332 (N_18332,N_18139,N_18238);
xnor U18333 (N_18333,N_18078,N_18083);
nand U18334 (N_18334,N_18249,N_18160);
nand U18335 (N_18335,N_18157,N_18126);
nor U18336 (N_18336,N_18148,N_18025);
or U18337 (N_18337,N_18026,N_18101);
xor U18338 (N_18338,N_18007,N_18226);
nand U18339 (N_18339,N_18106,N_18004);
nand U18340 (N_18340,N_18142,N_18048);
xnor U18341 (N_18341,N_18129,N_18073);
nor U18342 (N_18342,N_18097,N_18040);
nand U18343 (N_18343,N_18199,N_18218);
or U18344 (N_18344,N_18237,N_18169);
nor U18345 (N_18345,N_18134,N_18210);
nor U18346 (N_18346,N_18080,N_18241);
or U18347 (N_18347,N_18093,N_18018);
nand U18348 (N_18348,N_18042,N_18154);
or U18349 (N_18349,N_18155,N_18186);
nand U18350 (N_18350,N_18188,N_18165);
and U18351 (N_18351,N_18074,N_18183);
and U18352 (N_18352,N_18035,N_18072);
nand U18353 (N_18353,N_18076,N_18013);
nor U18354 (N_18354,N_18008,N_18096);
or U18355 (N_18355,N_18208,N_18245);
or U18356 (N_18356,N_18113,N_18207);
xnor U18357 (N_18357,N_18037,N_18061);
nand U18358 (N_18358,N_18220,N_18166);
or U18359 (N_18359,N_18229,N_18173);
xor U18360 (N_18360,N_18175,N_18140);
xnor U18361 (N_18361,N_18240,N_18211);
nor U18362 (N_18362,N_18094,N_18039);
and U18363 (N_18363,N_18001,N_18215);
xnor U18364 (N_18364,N_18150,N_18203);
nor U18365 (N_18365,N_18127,N_18128);
or U18366 (N_18366,N_18071,N_18047);
or U18367 (N_18367,N_18137,N_18174);
nor U18368 (N_18368,N_18247,N_18081);
nand U18369 (N_18369,N_18114,N_18122);
nor U18370 (N_18370,N_18075,N_18141);
xnor U18371 (N_18371,N_18092,N_18112);
or U18372 (N_18372,N_18152,N_18023);
and U18373 (N_18373,N_18036,N_18024);
nand U18374 (N_18374,N_18182,N_18056);
or U18375 (N_18375,N_18236,N_18093);
nor U18376 (N_18376,N_18028,N_18164);
nand U18377 (N_18377,N_18079,N_18105);
nand U18378 (N_18378,N_18022,N_18106);
or U18379 (N_18379,N_18181,N_18207);
xor U18380 (N_18380,N_18195,N_18191);
and U18381 (N_18381,N_18138,N_18233);
and U18382 (N_18382,N_18095,N_18167);
or U18383 (N_18383,N_18070,N_18217);
or U18384 (N_18384,N_18199,N_18043);
nand U18385 (N_18385,N_18022,N_18238);
xnor U18386 (N_18386,N_18013,N_18105);
nor U18387 (N_18387,N_18039,N_18104);
nand U18388 (N_18388,N_18146,N_18152);
xnor U18389 (N_18389,N_18094,N_18200);
xor U18390 (N_18390,N_18208,N_18120);
nand U18391 (N_18391,N_18036,N_18137);
or U18392 (N_18392,N_18190,N_18216);
nand U18393 (N_18393,N_18133,N_18064);
nand U18394 (N_18394,N_18035,N_18094);
nor U18395 (N_18395,N_18227,N_18013);
xor U18396 (N_18396,N_18035,N_18118);
xnor U18397 (N_18397,N_18194,N_18006);
nor U18398 (N_18398,N_18246,N_18134);
or U18399 (N_18399,N_18068,N_18182);
nor U18400 (N_18400,N_18248,N_18155);
nor U18401 (N_18401,N_18150,N_18076);
nor U18402 (N_18402,N_18020,N_18118);
nand U18403 (N_18403,N_18055,N_18079);
or U18404 (N_18404,N_18068,N_18191);
nand U18405 (N_18405,N_18206,N_18228);
nor U18406 (N_18406,N_18016,N_18148);
or U18407 (N_18407,N_18131,N_18073);
nor U18408 (N_18408,N_18167,N_18032);
nand U18409 (N_18409,N_18048,N_18238);
nor U18410 (N_18410,N_18141,N_18003);
and U18411 (N_18411,N_18040,N_18159);
xor U18412 (N_18412,N_18151,N_18041);
xor U18413 (N_18413,N_18122,N_18111);
and U18414 (N_18414,N_18235,N_18065);
or U18415 (N_18415,N_18142,N_18003);
nand U18416 (N_18416,N_18047,N_18192);
and U18417 (N_18417,N_18080,N_18121);
nand U18418 (N_18418,N_18221,N_18090);
nand U18419 (N_18419,N_18206,N_18030);
nand U18420 (N_18420,N_18022,N_18128);
or U18421 (N_18421,N_18196,N_18217);
and U18422 (N_18422,N_18113,N_18249);
or U18423 (N_18423,N_18225,N_18147);
nor U18424 (N_18424,N_18123,N_18106);
xor U18425 (N_18425,N_18085,N_18176);
nor U18426 (N_18426,N_18144,N_18197);
or U18427 (N_18427,N_18053,N_18055);
nor U18428 (N_18428,N_18124,N_18031);
or U18429 (N_18429,N_18102,N_18197);
xnor U18430 (N_18430,N_18066,N_18045);
nand U18431 (N_18431,N_18185,N_18074);
nor U18432 (N_18432,N_18002,N_18139);
nand U18433 (N_18433,N_18059,N_18018);
and U18434 (N_18434,N_18217,N_18162);
nor U18435 (N_18435,N_18084,N_18130);
and U18436 (N_18436,N_18107,N_18225);
xor U18437 (N_18437,N_18212,N_18149);
nand U18438 (N_18438,N_18110,N_18212);
or U18439 (N_18439,N_18066,N_18245);
or U18440 (N_18440,N_18149,N_18191);
and U18441 (N_18441,N_18005,N_18099);
nand U18442 (N_18442,N_18045,N_18209);
nand U18443 (N_18443,N_18229,N_18118);
nor U18444 (N_18444,N_18213,N_18064);
or U18445 (N_18445,N_18053,N_18211);
and U18446 (N_18446,N_18085,N_18218);
and U18447 (N_18447,N_18098,N_18118);
nand U18448 (N_18448,N_18174,N_18031);
nor U18449 (N_18449,N_18021,N_18246);
nand U18450 (N_18450,N_18080,N_18108);
nor U18451 (N_18451,N_18162,N_18101);
xnor U18452 (N_18452,N_18029,N_18042);
nand U18453 (N_18453,N_18115,N_18187);
or U18454 (N_18454,N_18033,N_18201);
or U18455 (N_18455,N_18147,N_18022);
nor U18456 (N_18456,N_18155,N_18046);
xor U18457 (N_18457,N_18143,N_18200);
nor U18458 (N_18458,N_18036,N_18184);
xor U18459 (N_18459,N_18124,N_18211);
xnor U18460 (N_18460,N_18054,N_18029);
or U18461 (N_18461,N_18019,N_18000);
and U18462 (N_18462,N_18019,N_18094);
xor U18463 (N_18463,N_18098,N_18224);
nor U18464 (N_18464,N_18011,N_18039);
nor U18465 (N_18465,N_18035,N_18042);
nor U18466 (N_18466,N_18014,N_18161);
nand U18467 (N_18467,N_18022,N_18073);
and U18468 (N_18468,N_18207,N_18045);
or U18469 (N_18469,N_18066,N_18063);
and U18470 (N_18470,N_18175,N_18050);
and U18471 (N_18471,N_18151,N_18169);
or U18472 (N_18472,N_18058,N_18243);
or U18473 (N_18473,N_18185,N_18098);
nor U18474 (N_18474,N_18038,N_18204);
nor U18475 (N_18475,N_18022,N_18244);
or U18476 (N_18476,N_18121,N_18107);
nand U18477 (N_18477,N_18088,N_18111);
or U18478 (N_18478,N_18032,N_18197);
nor U18479 (N_18479,N_18180,N_18089);
nand U18480 (N_18480,N_18056,N_18061);
or U18481 (N_18481,N_18060,N_18236);
xnor U18482 (N_18482,N_18041,N_18108);
nor U18483 (N_18483,N_18014,N_18120);
xor U18484 (N_18484,N_18140,N_18240);
xor U18485 (N_18485,N_18153,N_18058);
and U18486 (N_18486,N_18194,N_18105);
and U18487 (N_18487,N_18239,N_18146);
nand U18488 (N_18488,N_18014,N_18013);
nor U18489 (N_18489,N_18136,N_18230);
or U18490 (N_18490,N_18015,N_18220);
and U18491 (N_18491,N_18220,N_18058);
and U18492 (N_18492,N_18200,N_18108);
nor U18493 (N_18493,N_18123,N_18226);
or U18494 (N_18494,N_18081,N_18135);
nand U18495 (N_18495,N_18033,N_18188);
xnor U18496 (N_18496,N_18142,N_18089);
and U18497 (N_18497,N_18213,N_18089);
or U18498 (N_18498,N_18238,N_18107);
xnor U18499 (N_18499,N_18057,N_18058);
nand U18500 (N_18500,N_18477,N_18261);
and U18501 (N_18501,N_18281,N_18280);
and U18502 (N_18502,N_18384,N_18371);
or U18503 (N_18503,N_18328,N_18480);
nor U18504 (N_18504,N_18494,N_18315);
and U18505 (N_18505,N_18283,N_18346);
or U18506 (N_18506,N_18333,N_18256);
or U18507 (N_18507,N_18367,N_18471);
xor U18508 (N_18508,N_18478,N_18262);
and U18509 (N_18509,N_18474,N_18433);
or U18510 (N_18510,N_18303,N_18291);
nand U18511 (N_18511,N_18387,N_18286);
nand U18512 (N_18512,N_18373,N_18360);
or U18513 (N_18513,N_18296,N_18440);
nor U18514 (N_18514,N_18421,N_18419);
or U18515 (N_18515,N_18329,N_18452);
or U18516 (N_18516,N_18332,N_18415);
nand U18517 (N_18517,N_18405,N_18472);
and U18518 (N_18518,N_18284,N_18279);
nor U18519 (N_18519,N_18325,N_18492);
nand U18520 (N_18520,N_18330,N_18495);
xor U18521 (N_18521,N_18355,N_18410);
or U18522 (N_18522,N_18382,N_18409);
or U18523 (N_18523,N_18344,N_18251);
xnor U18524 (N_18524,N_18431,N_18352);
nand U18525 (N_18525,N_18372,N_18427);
nand U18526 (N_18526,N_18422,N_18458);
nand U18527 (N_18527,N_18450,N_18392);
nor U18528 (N_18528,N_18308,N_18377);
nor U18529 (N_18529,N_18309,N_18314);
or U18530 (N_18530,N_18311,N_18271);
and U18531 (N_18531,N_18435,N_18374);
xnor U18532 (N_18532,N_18368,N_18453);
and U18533 (N_18533,N_18423,N_18445);
nor U18534 (N_18534,N_18408,N_18297);
nand U18535 (N_18535,N_18499,N_18335);
xnor U18536 (N_18536,N_18305,N_18481);
xor U18537 (N_18537,N_18337,N_18420);
nand U18538 (N_18538,N_18430,N_18389);
nand U18539 (N_18539,N_18488,N_18414);
xnor U18540 (N_18540,N_18424,N_18270);
nand U18541 (N_18541,N_18380,N_18353);
nand U18542 (N_18542,N_18340,N_18259);
nor U18543 (N_18543,N_18407,N_18432);
xnor U18544 (N_18544,N_18267,N_18482);
nand U18545 (N_18545,N_18266,N_18348);
xor U18546 (N_18546,N_18293,N_18300);
xnor U18547 (N_18547,N_18253,N_18304);
xor U18548 (N_18548,N_18274,N_18277);
or U18549 (N_18549,N_18307,N_18317);
and U18550 (N_18550,N_18456,N_18475);
and U18551 (N_18551,N_18276,N_18418);
or U18552 (N_18552,N_18349,N_18463);
xnor U18553 (N_18553,N_18461,N_18285);
or U18554 (N_18554,N_18447,N_18275);
and U18555 (N_18555,N_18393,N_18264);
xnor U18556 (N_18556,N_18292,N_18263);
or U18557 (N_18557,N_18400,N_18468);
nand U18558 (N_18558,N_18252,N_18250);
nor U18559 (N_18559,N_18294,N_18483);
nor U18560 (N_18560,N_18396,N_18361);
nor U18561 (N_18561,N_18470,N_18404);
or U18562 (N_18562,N_18341,N_18364);
nand U18563 (N_18563,N_18269,N_18306);
nor U18564 (N_18564,N_18473,N_18365);
and U18565 (N_18565,N_18376,N_18397);
and U18566 (N_18566,N_18487,N_18370);
nor U18567 (N_18567,N_18287,N_18464);
and U18568 (N_18568,N_18282,N_18466);
nand U18569 (N_18569,N_18278,N_18493);
nor U18570 (N_18570,N_18441,N_18467);
nor U18571 (N_18571,N_18402,N_18322);
or U18572 (N_18572,N_18255,N_18485);
nor U18573 (N_18573,N_18381,N_18316);
nor U18574 (N_18574,N_18358,N_18497);
nand U18575 (N_18575,N_18327,N_18448);
and U18576 (N_18576,N_18417,N_18439);
nand U18577 (N_18577,N_18290,N_18394);
nor U18578 (N_18578,N_18398,N_18268);
xnor U18579 (N_18579,N_18460,N_18442);
nor U18580 (N_18580,N_18390,N_18496);
nand U18581 (N_18581,N_18336,N_18257);
or U18582 (N_18582,N_18265,N_18359);
nand U18583 (N_18583,N_18298,N_18258);
xor U18584 (N_18584,N_18366,N_18416);
and U18585 (N_18585,N_18446,N_18498);
nor U18586 (N_18586,N_18383,N_18342);
nand U18587 (N_18587,N_18288,N_18323);
or U18588 (N_18588,N_18338,N_18331);
nand U18589 (N_18589,N_18484,N_18443);
nor U18590 (N_18590,N_18476,N_18391);
nand U18591 (N_18591,N_18313,N_18462);
nor U18592 (N_18592,N_18406,N_18491);
or U18593 (N_18593,N_18299,N_18388);
nand U18594 (N_18594,N_18479,N_18345);
or U18595 (N_18595,N_18438,N_18362);
xor U18596 (N_18596,N_18490,N_18395);
nor U18597 (N_18597,N_18451,N_18434);
xor U18598 (N_18598,N_18310,N_18334);
or U18599 (N_18599,N_18302,N_18357);
nor U18600 (N_18600,N_18457,N_18375);
nor U18601 (N_18601,N_18403,N_18319);
xnor U18602 (N_18602,N_18312,N_18379);
nor U18603 (N_18603,N_18326,N_18455);
xor U18604 (N_18604,N_18489,N_18385);
and U18605 (N_18605,N_18428,N_18324);
and U18606 (N_18606,N_18401,N_18413);
or U18607 (N_18607,N_18386,N_18339);
nor U18608 (N_18608,N_18436,N_18378);
nor U18609 (N_18609,N_18273,N_18363);
or U18610 (N_18610,N_18343,N_18321);
nor U18611 (N_18611,N_18437,N_18369);
nand U18612 (N_18612,N_18260,N_18449);
xnor U18613 (N_18613,N_18426,N_18454);
nand U18614 (N_18614,N_18318,N_18351);
xor U18615 (N_18615,N_18412,N_18295);
nor U18616 (N_18616,N_18459,N_18354);
and U18617 (N_18617,N_18301,N_18254);
nand U18618 (N_18618,N_18350,N_18320);
nor U18619 (N_18619,N_18399,N_18356);
or U18620 (N_18620,N_18465,N_18289);
and U18621 (N_18621,N_18411,N_18486);
or U18622 (N_18622,N_18444,N_18429);
nand U18623 (N_18623,N_18347,N_18469);
xnor U18624 (N_18624,N_18425,N_18272);
nor U18625 (N_18625,N_18449,N_18284);
xor U18626 (N_18626,N_18266,N_18472);
nand U18627 (N_18627,N_18385,N_18313);
or U18628 (N_18628,N_18496,N_18276);
nand U18629 (N_18629,N_18437,N_18331);
or U18630 (N_18630,N_18456,N_18443);
xnor U18631 (N_18631,N_18405,N_18433);
and U18632 (N_18632,N_18391,N_18415);
xor U18633 (N_18633,N_18377,N_18419);
and U18634 (N_18634,N_18389,N_18481);
or U18635 (N_18635,N_18464,N_18349);
and U18636 (N_18636,N_18298,N_18309);
and U18637 (N_18637,N_18473,N_18337);
nand U18638 (N_18638,N_18481,N_18349);
and U18639 (N_18639,N_18339,N_18456);
or U18640 (N_18640,N_18353,N_18469);
or U18641 (N_18641,N_18267,N_18289);
nor U18642 (N_18642,N_18359,N_18358);
xor U18643 (N_18643,N_18347,N_18388);
nand U18644 (N_18644,N_18315,N_18393);
or U18645 (N_18645,N_18315,N_18412);
or U18646 (N_18646,N_18338,N_18370);
nor U18647 (N_18647,N_18486,N_18408);
xnor U18648 (N_18648,N_18425,N_18381);
nor U18649 (N_18649,N_18268,N_18391);
xnor U18650 (N_18650,N_18275,N_18313);
nor U18651 (N_18651,N_18293,N_18256);
xor U18652 (N_18652,N_18329,N_18278);
xor U18653 (N_18653,N_18327,N_18252);
nand U18654 (N_18654,N_18393,N_18460);
nand U18655 (N_18655,N_18446,N_18447);
nor U18656 (N_18656,N_18297,N_18392);
nor U18657 (N_18657,N_18409,N_18266);
and U18658 (N_18658,N_18320,N_18333);
xnor U18659 (N_18659,N_18351,N_18444);
nor U18660 (N_18660,N_18381,N_18440);
nand U18661 (N_18661,N_18414,N_18483);
and U18662 (N_18662,N_18413,N_18486);
nor U18663 (N_18663,N_18442,N_18264);
or U18664 (N_18664,N_18487,N_18302);
nand U18665 (N_18665,N_18283,N_18294);
or U18666 (N_18666,N_18283,N_18301);
xnor U18667 (N_18667,N_18272,N_18499);
or U18668 (N_18668,N_18300,N_18259);
and U18669 (N_18669,N_18366,N_18393);
and U18670 (N_18670,N_18484,N_18416);
or U18671 (N_18671,N_18421,N_18453);
nand U18672 (N_18672,N_18302,N_18284);
nor U18673 (N_18673,N_18430,N_18281);
and U18674 (N_18674,N_18348,N_18440);
nor U18675 (N_18675,N_18321,N_18474);
xor U18676 (N_18676,N_18476,N_18424);
xnor U18677 (N_18677,N_18467,N_18453);
or U18678 (N_18678,N_18437,N_18406);
nor U18679 (N_18679,N_18362,N_18409);
xnor U18680 (N_18680,N_18275,N_18281);
nor U18681 (N_18681,N_18417,N_18490);
and U18682 (N_18682,N_18317,N_18336);
nand U18683 (N_18683,N_18306,N_18332);
and U18684 (N_18684,N_18472,N_18377);
nand U18685 (N_18685,N_18349,N_18451);
or U18686 (N_18686,N_18488,N_18428);
nand U18687 (N_18687,N_18498,N_18403);
xnor U18688 (N_18688,N_18452,N_18489);
nor U18689 (N_18689,N_18414,N_18277);
and U18690 (N_18690,N_18384,N_18410);
or U18691 (N_18691,N_18320,N_18343);
nor U18692 (N_18692,N_18361,N_18480);
or U18693 (N_18693,N_18286,N_18439);
xor U18694 (N_18694,N_18385,N_18412);
and U18695 (N_18695,N_18376,N_18255);
nand U18696 (N_18696,N_18412,N_18393);
and U18697 (N_18697,N_18351,N_18368);
and U18698 (N_18698,N_18379,N_18338);
and U18699 (N_18699,N_18374,N_18455);
nor U18700 (N_18700,N_18275,N_18386);
or U18701 (N_18701,N_18277,N_18322);
nand U18702 (N_18702,N_18394,N_18381);
xnor U18703 (N_18703,N_18291,N_18360);
or U18704 (N_18704,N_18309,N_18344);
and U18705 (N_18705,N_18350,N_18468);
nand U18706 (N_18706,N_18475,N_18423);
xnor U18707 (N_18707,N_18262,N_18311);
nand U18708 (N_18708,N_18301,N_18417);
nor U18709 (N_18709,N_18276,N_18351);
xnor U18710 (N_18710,N_18250,N_18486);
and U18711 (N_18711,N_18406,N_18345);
xnor U18712 (N_18712,N_18471,N_18319);
xnor U18713 (N_18713,N_18409,N_18312);
or U18714 (N_18714,N_18419,N_18356);
and U18715 (N_18715,N_18379,N_18322);
nand U18716 (N_18716,N_18429,N_18395);
and U18717 (N_18717,N_18485,N_18444);
nor U18718 (N_18718,N_18427,N_18259);
xnor U18719 (N_18719,N_18484,N_18458);
nand U18720 (N_18720,N_18374,N_18497);
nor U18721 (N_18721,N_18404,N_18312);
nand U18722 (N_18722,N_18403,N_18411);
or U18723 (N_18723,N_18460,N_18467);
and U18724 (N_18724,N_18497,N_18307);
or U18725 (N_18725,N_18310,N_18261);
and U18726 (N_18726,N_18344,N_18316);
nor U18727 (N_18727,N_18413,N_18407);
or U18728 (N_18728,N_18433,N_18285);
nand U18729 (N_18729,N_18303,N_18375);
or U18730 (N_18730,N_18470,N_18416);
nand U18731 (N_18731,N_18300,N_18390);
and U18732 (N_18732,N_18367,N_18473);
nand U18733 (N_18733,N_18337,N_18470);
or U18734 (N_18734,N_18369,N_18374);
and U18735 (N_18735,N_18275,N_18490);
and U18736 (N_18736,N_18357,N_18394);
and U18737 (N_18737,N_18328,N_18361);
nand U18738 (N_18738,N_18486,N_18340);
nand U18739 (N_18739,N_18336,N_18348);
and U18740 (N_18740,N_18276,N_18428);
xor U18741 (N_18741,N_18250,N_18450);
nand U18742 (N_18742,N_18442,N_18417);
nor U18743 (N_18743,N_18434,N_18279);
xnor U18744 (N_18744,N_18292,N_18469);
nor U18745 (N_18745,N_18384,N_18492);
or U18746 (N_18746,N_18262,N_18404);
nand U18747 (N_18747,N_18459,N_18362);
nor U18748 (N_18748,N_18366,N_18376);
nand U18749 (N_18749,N_18270,N_18423);
xnor U18750 (N_18750,N_18629,N_18719);
or U18751 (N_18751,N_18730,N_18624);
or U18752 (N_18752,N_18502,N_18570);
nor U18753 (N_18753,N_18585,N_18533);
xnor U18754 (N_18754,N_18690,N_18732);
nand U18755 (N_18755,N_18577,N_18616);
nand U18756 (N_18756,N_18634,N_18595);
and U18757 (N_18757,N_18584,N_18644);
and U18758 (N_18758,N_18664,N_18564);
and U18759 (N_18759,N_18687,N_18503);
nor U18760 (N_18760,N_18523,N_18515);
xnor U18761 (N_18761,N_18548,N_18642);
nor U18762 (N_18762,N_18610,N_18683);
xnor U18763 (N_18763,N_18622,N_18703);
or U18764 (N_18764,N_18551,N_18505);
and U18765 (N_18765,N_18611,N_18547);
or U18766 (N_18766,N_18630,N_18580);
nand U18767 (N_18767,N_18617,N_18534);
xnor U18768 (N_18768,N_18678,N_18623);
nand U18769 (N_18769,N_18602,N_18597);
nand U18770 (N_18770,N_18699,N_18576);
nand U18771 (N_18771,N_18528,N_18641);
or U18772 (N_18772,N_18681,N_18676);
xnor U18773 (N_18773,N_18532,N_18635);
nand U18774 (N_18774,N_18621,N_18579);
nor U18775 (N_18775,N_18725,N_18536);
or U18776 (N_18776,N_18514,N_18631);
nor U18777 (N_18777,N_18707,N_18513);
nand U18778 (N_18778,N_18521,N_18662);
nor U18779 (N_18779,N_18645,N_18705);
or U18780 (N_18780,N_18625,N_18729);
xor U18781 (N_18781,N_18566,N_18658);
nand U18782 (N_18782,N_18659,N_18511);
nand U18783 (N_18783,N_18501,N_18557);
and U18784 (N_18784,N_18748,N_18587);
nor U18785 (N_18785,N_18620,N_18558);
or U18786 (N_18786,N_18731,N_18565);
xnor U18787 (N_18787,N_18582,N_18650);
nor U18788 (N_18788,N_18727,N_18749);
nor U18789 (N_18789,N_18575,N_18594);
and U18790 (N_18790,N_18668,N_18607);
nand U18791 (N_18791,N_18737,N_18667);
or U18792 (N_18792,N_18603,N_18590);
nor U18793 (N_18793,N_18684,N_18663);
xnor U18794 (N_18794,N_18546,N_18696);
nand U18795 (N_18795,N_18531,N_18688);
xnor U18796 (N_18796,N_18578,N_18518);
or U18797 (N_18797,N_18540,N_18706);
and U18798 (N_18798,N_18504,N_18653);
or U18799 (N_18799,N_18553,N_18626);
or U18800 (N_18800,N_18649,N_18637);
and U18801 (N_18801,N_18717,N_18581);
nor U18802 (N_18802,N_18652,N_18702);
nand U18803 (N_18803,N_18686,N_18685);
xnor U18804 (N_18804,N_18525,N_18657);
nor U18805 (N_18805,N_18700,N_18526);
xor U18806 (N_18806,N_18710,N_18651);
or U18807 (N_18807,N_18606,N_18601);
and U18808 (N_18808,N_18713,N_18643);
nand U18809 (N_18809,N_18704,N_18638);
nor U18810 (N_18810,N_18512,N_18561);
xor U18811 (N_18811,N_18520,N_18596);
nor U18812 (N_18812,N_18735,N_18605);
and U18813 (N_18813,N_18543,N_18556);
and U18814 (N_18814,N_18583,N_18682);
nor U18815 (N_18815,N_18695,N_18655);
xor U18816 (N_18816,N_18656,N_18591);
or U18817 (N_18817,N_18573,N_18720);
or U18818 (N_18818,N_18742,N_18692);
nand U18819 (N_18819,N_18508,N_18734);
nand U18820 (N_18820,N_18571,N_18640);
and U18821 (N_18821,N_18627,N_18673);
or U18822 (N_18822,N_18509,N_18661);
xor U18823 (N_18823,N_18527,N_18599);
xnor U18824 (N_18824,N_18746,N_18697);
and U18825 (N_18825,N_18745,N_18669);
xnor U18826 (N_18826,N_18545,N_18500);
nor U18827 (N_18827,N_18554,N_18672);
and U18828 (N_18828,N_18524,N_18743);
nand U18829 (N_18829,N_18537,N_18738);
xor U18830 (N_18830,N_18708,N_18636);
nor U18831 (N_18831,N_18588,N_18600);
xor U18832 (N_18832,N_18613,N_18718);
nor U18833 (N_18833,N_18541,N_18522);
nor U18834 (N_18834,N_18721,N_18715);
or U18835 (N_18835,N_18677,N_18550);
nor U18836 (N_18836,N_18724,N_18549);
and U18837 (N_18837,N_18618,N_18608);
nor U18838 (N_18838,N_18563,N_18593);
or U18839 (N_18839,N_18740,N_18728);
and U18840 (N_18840,N_18701,N_18654);
xnor U18841 (N_18841,N_18598,N_18538);
and U18842 (N_18842,N_18555,N_18712);
nand U18843 (N_18843,N_18716,N_18741);
xnor U18844 (N_18844,N_18559,N_18666);
and U18845 (N_18845,N_18674,N_18529);
and U18846 (N_18846,N_18747,N_18744);
nand U18847 (N_18847,N_18698,N_18660);
or U18848 (N_18848,N_18711,N_18680);
xnor U18849 (N_18849,N_18736,N_18568);
nand U18850 (N_18850,N_18648,N_18609);
or U18851 (N_18851,N_18665,N_18693);
nand U18852 (N_18852,N_18723,N_18510);
or U18853 (N_18853,N_18679,N_18560);
and U18854 (N_18854,N_18619,N_18506);
xnor U18855 (N_18855,N_18572,N_18589);
and U18856 (N_18856,N_18647,N_18542);
and U18857 (N_18857,N_18604,N_18507);
or U18858 (N_18858,N_18691,N_18675);
nor U18859 (N_18859,N_18567,N_18535);
xnor U18860 (N_18860,N_18614,N_18562);
xor U18861 (N_18861,N_18689,N_18639);
and U18862 (N_18862,N_18592,N_18628);
and U18863 (N_18863,N_18574,N_18615);
or U18864 (N_18864,N_18516,N_18519);
or U18865 (N_18865,N_18733,N_18612);
xor U18866 (N_18866,N_18646,N_18670);
xor U18867 (N_18867,N_18586,N_18739);
or U18868 (N_18868,N_18633,N_18722);
and U18869 (N_18869,N_18517,N_18714);
nand U18870 (N_18870,N_18552,N_18694);
xor U18871 (N_18871,N_18632,N_18569);
or U18872 (N_18872,N_18671,N_18726);
or U18873 (N_18873,N_18539,N_18530);
nand U18874 (N_18874,N_18544,N_18709);
nor U18875 (N_18875,N_18515,N_18685);
or U18876 (N_18876,N_18653,N_18622);
nand U18877 (N_18877,N_18605,N_18671);
or U18878 (N_18878,N_18639,N_18550);
xor U18879 (N_18879,N_18718,N_18579);
xor U18880 (N_18880,N_18723,N_18741);
or U18881 (N_18881,N_18633,N_18735);
nand U18882 (N_18882,N_18717,N_18634);
xnor U18883 (N_18883,N_18717,N_18594);
nand U18884 (N_18884,N_18574,N_18596);
nand U18885 (N_18885,N_18690,N_18566);
xnor U18886 (N_18886,N_18589,N_18709);
and U18887 (N_18887,N_18632,N_18508);
and U18888 (N_18888,N_18675,N_18655);
nand U18889 (N_18889,N_18512,N_18597);
or U18890 (N_18890,N_18580,N_18540);
or U18891 (N_18891,N_18614,N_18555);
or U18892 (N_18892,N_18643,N_18692);
xnor U18893 (N_18893,N_18543,N_18561);
or U18894 (N_18894,N_18734,N_18535);
xnor U18895 (N_18895,N_18677,N_18646);
or U18896 (N_18896,N_18686,N_18737);
or U18897 (N_18897,N_18667,N_18714);
xnor U18898 (N_18898,N_18543,N_18566);
nand U18899 (N_18899,N_18725,N_18619);
or U18900 (N_18900,N_18509,N_18652);
or U18901 (N_18901,N_18606,N_18516);
or U18902 (N_18902,N_18649,N_18696);
nor U18903 (N_18903,N_18574,N_18693);
xnor U18904 (N_18904,N_18505,N_18626);
nor U18905 (N_18905,N_18599,N_18718);
or U18906 (N_18906,N_18505,N_18514);
nand U18907 (N_18907,N_18606,N_18569);
nand U18908 (N_18908,N_18573,N_18721);
nor U18909 (N_18909,N_18609,N_18701);
nand U18910 (N_18910,N_18510,N_18585);
or U18911 (N_18911,N_18612,N_18584);
nand U18912 (N_18912,N_18595,N_18575);
nand U18913 (N_18913,N_18520,N_18506);
and U18914 (N_18914,N_18718,N_18720);
nand U18915 (N_18915,N_18663,N_18577);
nand U18916 (N_18916,N_18593,N_18678);
and U18917 (N_18917,N_18581,N_18664);
nor U18918 (N_18918,N_18714,N_18562);
or U18919 (N_18919,N_18527,N_18523);
or U18920 (N_18920,N_18719,N_18740);
and U18921 (N_18921,N_18700,N_18680);
and U18922 (N_18922,N_18597,N_18573);
nor U18923 (N_18923,N_18636,N_18590);
xor U18924 (N_18924,N_18746,N_18514);
xor U18925 (N_18925,N_18572,N_18692);
nand U18926 (N_18926,N_18599,N_18556);
or U18927 (N_18927,N_18560,N_18747);
and U18928 (N_18928,N_18538,N_18555);
nand U18929 (N_18929,N_18538,N_18549);
or U18930 (N_18930,N_18527,N_18684);
and U18931 (N_18931,N_18519,N_18551);
or U18932 (N_18932,N_18522,N_18635);
nand U18933 (N_18933,N_18588,N_18551);
and U18934 (N_18934,N_18679,N_18723);
or U18935 (N_18935,N_18656,N_18607);
and U18936 (N_18936,N_18603,N_18610);
nor U18937 (N_18937,N_18574,N_18538);
or U18938 (N_18938,N_18699,N_18635);
xor U18939 (N_18939,N_18534,N_18718);
and U18940 (N_18940,N_18668,N_18575);
nor U18941 (N_18941,N_18517,N_18675);
or U18942 (N_18942,N_18723,N_18591);
xor U18943 (N_18943,N_18639,N_18712);
xor U18944 (N_18944,N_18594,N_18504);
xor U18945 (N_18945,N_18649,N_18646);
and U18946 (N_18946,N_18703,N_18593);
xnor U18947 (N_18947,N_18727,N_18547);
xnor U18948 (N_18948,N_18672,N_18600);
nand U18949 (N_18949,N_18633,N_18594);
nand U18950 (N_18950,N_18672,N_18579);
nor U18951 (N_18951,N_18614,N_18646);
nor U18952 (N_18952,N_18617,N_18630);
or U18953 (N_18953,N_18524,N_18749);
nor U18954 (N_18954,N_18685,N_18522);
nor U18955 (N_18955,N_18672,N_18515);
and U18956 (N_18956,N_18522,N_18642);
and U18957 (N_18957,N_18652,N_18656);
and U18958 (N_18958,N_18744,N_18542);
or U18959 (N_18959,N_18603,N_18608);
nand U18960 (N_18960,N_18569,N_18578);
nor U18961 (N_18961,N_18698,N_18612);
xnor U18962 (N_18962,N_18713,N_18714);
or U18963 (N_18963,N_18536,N_18502);
and U18964 (N_18964,N_18713,N_18519);
or U18965 (N_18965,N_18521,N_18567);
nor U18966 (N_18966,N_18712,N_18659);
xor U18967 (N_18967,N_18620,N_18730);
nand U18968 (N_18968,N_18666,N_18724);
or U18969 (N_18969,N_18536,N_18520);
and U18970 (N_18970,N_18533,N_18545);
nor U18971 (N_18971,N_18566,N_18626);
or U18972 (N_18972,N_18504,N_18674);
or U18973 (N_18973,N_18522,N_18598);
and U18974 (N_18974,N_18728,N_18567);
nor U18975 (N_18975,N_18637,N_18523);
xnor U18976 (N_18976,N_18645,N_18644);
nor U18977 (N_18977,N_18577,N_18720);
nand U18978 (N_18978,N_18624,N_18747);
nor U18979 (N_18979,N_18639,N_18744);
xor U18980 (N_18980,N_18717,N_18545);
nor U18981 (N_18981,N_18665,N_18519);
and U18982 (N_18982,N_18620,N_18667);
and U18983 (N_18983,N_18520,N_18721);
and U18984 (N_18984,N_18651,N_18677);
nor U18985 (N_18985,N_18568,N_18527);
and U18986 (N_18986,N_18612,N_18705);
and U18987 (N_18987,N_18713,N_18695);
nand U18988 (N_18988,N_18702,N_18620);
nand U18989 (N_18989,N_18662,N_18540);
xnor U18990 (N_18990,N_18695,N_18609);
or U18991 (N_18991,N_18727,N_18575);
xor U18992 (N_18992,N_18717,N_18651);
nand U18993 (N_18993,N_18583,N_18653);
nand U18994 (N_18994,N_18589,N_18604);
nor U18995 (N_18995,N_18699,N_18698);
nor U18996 (N_18996,N_18599,N_18691);
and U18997 (N_18997,N_18700,N_18536);
or U18998 (N_18998,N_18632,N_18515);
nor U18999 (N_18999,N_18604,N_18734);
nor U19000 (N_19000,N_18792,N_18985);
nor U19001 (N_19001,N_18760,N_18877);
nand U19002 (N_19002,N_18777,N_18898);
nand U19003 (N_19003,N_18962,N_18788);
nor U19004 (N_19004,N_18933,N_18847);
nor U19005 (N_19005,N_18955,N_18977);
nand U19006 (N_19006,N_18758,N_18757);
nor U19007 (N_19007,N_18887,N_18826);
and U19008 (N_19008,N_18867,N_18773);
nand U19009 (N_19009,N_18993,N_18850);
nand U19010 (N_19010,N_18912,N_18827);
nand U19011 (N_19011,N_18840,N_18774);
nand U19012 (N_19012,N_18916,N_18771);
and U19013 (N_19013,N_18872,N_18852);
nor U19014 (N_19014,N_18837,N_18811);
or U19015 (N_19015,N_18886,N_18915);
xor U19016 (N_19016,N_18945,N_18791);
nor U19017 (N_19017,N_18804,N_18823);
nand U19018 (N_19018,N_18973,N_18842);
nor U19019 (N_19019,N_18839,N_18941);
nand U19020 (N_19020,N_18810,N_18772);
nor U19021 (N_19021,N_18753,N_18902);
nand U19022 (N_19022,N_18950,N_18861);
xnor U19023 (N_19023,N_18942,N_18853);
nand U19024 (N_19024,N_18963,N_18974);
or U19025 (N_19025,N_18883,N_18935);
xor U19026 (N_19026,N_18889,N_18809);
xnor U19027 (N_19027,N_18800,N_18854);
and U19028 (N_19028,N_18863,N_18938);
xor U19029 (N_19029,N_18756,N_18778);
nand U19030 (N_19030,N_18754,N_18891);
and U19031 (N_19031,N_18799,N_18903);
and U19032 (N_19032,N_18980,N_18992);
or U19033 (N_19033,N_18875,N_18957);
and U19034 (N_19034,N_18901,N_18948);
and U19035 (N_19035,N_18989,N_18798);
nor U19036 (N_19036,N_18899,N_18905);
or U19037 (N_19037,N_18943,N_18768);
nor U19038 (N_19038,N_18932,N_18914);
xnor U19039 (N_19039,N_18986,N_18865);
nor U19040 (N_19040,N_18919,N_18881);
nor U19041 (N_19041,N_18940,N_18953);
or U19042 (N_19042,N_18892,N_18924);
xor U19043 (N_19043,N_18824,N_18880);
or U19044 (N_19044,N_18911,N_18780);
nor U19045 (N_19045,N_18781,N_18838);
nand U19046 (N_19046,N_18815,N_18830);
nor U19047 (N_19047,N_18906,N_18949);
xor U19048 (N_19048,N_18990,N_18779);
nand U19049 (N_19049,N_18923,N_18834);
or U19050 (N_19050,N_18995,N_18856);
nor U19051 (N_19051,N_18927,N_18767);
nor U19052 (N_19052,N_18972,N_18797);
nand U19053 (N_19053,N_18787,N_18818);
or U19054 (N_19054,N_18782,N_18936);
xnor U19055 (N_19055,N_18884,N_18864);
nand U19056 (N_19056,N_18984,N_18828);
xor U19057 (N_19057,N_18983,N_18954);
nor U19058 (N_19058,N_18930,N_18775);
and U19059 (N_19059,N_18969,N_18848);
and U19060 (N_19060,N_18752,N_18843);
xnor U19061 (N_19061,N_18965,N_18956);
and U19062 (N_19062,N_18803,N_18960);
or U19063 (N_19063,N_18894,N_18808);
xor U19064 (N_19064,N_18866,N_18964);
or U19065 (N_19065,N_18802,N_18829);
nor U19066 (N_19066,N_18776,N_18825);
nor U19067 (N_19067,N_18999,N_18893);
xnor U19068 (N_19068,N_18944,N_18789);
xnor U19069 (N_19069,N_18766,N_18762);
nand U19070 (N_19070,N_18836,N_18925);
and U19071 (N_19071,N_18784,N_18988);
xor U19072 (N_19072,N_18907,N_18939);
or U19073 (N_19073,N_18857,N_18759);
xnor U19074 (N_19074,N_18910,N_18982);
xnor U19075 (N_19075,N_18822,N_18796);
nor U19076 (N_19076,N_18952,N_18859);
or U19077 (N_19077,N_18967,N_18868);
nor U19078 (N_19078,N_18975,N_18918);
nor U19079 (N_19079,N_18994,N_18998);
nor U19080 (N_19080,N_18817,N_18846);
nand U19081 (N_19081,N_18959,N_18874);
or U19082 (N_19082,N_18885,N_18761);
xnor U19083 (N_19083,N_18921,N_18770);
xor U19084 (N_19084,N_18801,N_18991);
xnor U19085 (N_19085,N_18805,N_18896);
nor U19086 (N_19086,N_18831,N_18812);
and U19087 (N_19087,N_18764,N_18819);
xnor U19088 (N_19088,N_18844,N_18968);
xnor U19089 (N_19089,N_18928,N_18904);
and U19090 (N_19090,N_18979,N_18851);
or U19091 (N_19091,N_18858,N_18786);
and U19092 (N_19092,N_18997,N_18821);
nand U19093 (N_19093,N_18849,N_18946);
nor U19094 (N_19094,N_18862,N_18934);
nor U19095 (N_19095,N_18793,N_18922);
nor U19096 (N_19096,N_18755,N_18832);
or U19097 (N_19097,N_18947,N_18845);
nand U19098 (N_19098,N_18981,N_18814);
nor U19099 (N_19099,N_18895,N_18900);
and U19100 (N_19100,N_18931,N_18794);
nand U19101 (N_19101,N_18855,N_18795);
xor U19102 (N_19102,N_18929,N_18870);
nor U19103 (N_19103,N_18790,N_18890);
nand U19104 (N_19104,N_18835,N_18813);
nor U19105 (N_19105,N_18882,N_18917);
or U19106 (N_19106,N_18970,N_18833);
nand U19107 (N_19107,N_18765,N_18971);
or U19108 (N_19108,N_18987,N_18878);
or U19109 (N_19109,N_18966,N_18873);
and U19110 (N_19110,N_18961,N_18751);
nand U19111 (N_19111,N_18978,N_18820);
nand U19112 (N_19112,N_18807,N_18937);
nand U19113 (N_19113,N_18816,N_18951);
nand U19114 (N_19114,N_18888,N_18879);
or U19115 (N_19115,N_18750,N_18783);
and U19116 (N_19116,N_18763,N_18869);
or U19117 (N_19117,N_18769,N_18913);
xor U19118 (N_19118,N_18806,N_18841);
xnor U19119 (N_19119,N_18909,N_18908);
and U19120 (N_19120,N_18897,N_18871);
or U19121 (N_19121,N_18958,N_18860);
and U19122 (N_19122,N_18920,N_18926);
and U19123 (N_19123,N_18876,N_18996);
nor U19124 (N_19124,N_18785,N_18976);
nor U19125 (N_19125,N_18855,N_18776);
nor U19126 (N_19126,N_18985,N_18930);
or U19127 (N_19127,N_18805,N_18789);
or U19128 (N_19128,N_18913,N_18855);
and U19129 (N_19129,N_18988,N_18896);
and U19130 (N_19130,N_18907,N_18948);
or U19131 (N_19131,N_18985,N_18863);
or U19132 (N_19132,N_18896,N_18794);
nand U19133 (N_19133,N_18882,N_18977);
and U19134 (N_19134,N_18852,N_18859);
or U19135 (N_19135,N_18976,N_18926);
or U19136 (N_19136,N_18939,N_18777);
xor U19137 (N_19137,N_18977,N_18908);
and U19138 (N_19138,N_18813,N_18997);
or U19139 (N_19139,N_18794,N_18852);
xnor U19140 (N_19140,N_18785,N_18954);
nor U19141 (N_19141,N_18897,N_18778);
nand U19142 (N_19142,N_18888,N_18819);
or U19143 (N_19143,N_18966,N_18859);
xor U19144 (N_19144,N_18803,N_18805);
or U19145 (N_19145,N_18910,N_18936);
xor U19146 (N_19146,N_18824,N_18852);
and U19147 (N_19147,N_18804,N_18827);
xnor U19148 (N_19148,N_18883,N_18945);
or U19149 (N_19149,N_18774,N_18941);
nand U19150 (N_19150,N_18920,N_18952);
or U19151 (N_19151,N_18947,N_18889);
and U19152 (N_19152,N_18918,N_18904);
or U19153 (N_19153,N_18992,N_18988);
nand U19154 (N_19154,N_18809,N_18980);
nor U19155 (N_19155,N_18839,N_18757);
xor U19156 (N_19156,N_18786,N_18916);
nor U19157 (N_19157,N_18906,N_18974);
and U19158 (N_19158,N_18771,N_18911);
or U19159 (N_19159,N_18978,N_18983);
nand U19160 (N_19160,N_18930,N_18959);
or U19161 (N_19161,N_18922,N_18809);
or U19162 (N_19162,N_18854,N_18848);
nor U19163 (N_19163,N_18806,N_18922);
nand U19164 (N_19164,N_18860,N_18983);
or U19165 (N_19165,N_18809,N_18987);
nor U19166 (N_19166,N_18989,N_18981);
and U19167 (N_19167,N_18811,N_18967);
nand U19168 (N_19168,N_18818,N_18806);
or U19169 (N_19169,N_18896,N_18965);
xor U19170 (N_19170,N_18938,N_18955);
or U19171 (N_19171,N_18914,N_18799);
nor U19172 (N_19172,N_18924,N_18898);
and U19173 (N_19173,N_18874,N_18947);
xor U19174 (N_19174,N_18946,N_18750);
xor U19175 (N_19175,N_18950,N_18841);
xor U19176 (N_19176,N_18938,N_18796);
nor U19177 (N_19177,N_18978,N_18830);
xor U19178 (N_19178,N_18982,N_18797);
nor U19179 (N_19179,N_18802,N_18847);
and U19180 (N_19180,N_18958,N_18902);
xor U19181 (N_19181,N_18977,N_18844);
and U19182 (N_19182,N_18970,N_18961);
and U19183 (N_19183,N_18934,N_18848);
and U19184 (N_19184,N_18969,N_18785);
nand U19185 (N_19185,N_18960,N_18948);
and U19186 (N_19186,N_18803,N_18840);
xor U19187 (N_19187,N_18836,N_18823);
nor U19188 (N_19188,N_18951,N_18834);
nand U19189 (N_19189,N_18905,N_18980);
or U19190 (N_19190,N_18873,N_18993);
nor U19191 (N_19191,N_18833,N_18760);
nand U19192 (N_19192,N_18885,N_18823);
xor U19193 (N_19193,N_18771,N_18752);
or U19194 (N_19194,N_18901,N_18871);
or U19195 (N_19195,N_18830,N_18751);
nor U19196 (N_19196,N_18949,N_18899);
xor U19197 (N_19197,N_18859,N_18919);
xnor U19198 (N_19198,N_18831,N_18885);
nand U19199 (N_19199,N_18752,N_18988);
and U19200 (N_19200,N_18820,N_18863);
nor U19201 (N_19201,N_18805,N_18878);
xor U19202 (N_19202,N_18928,N_18982);
nand U19203 (N_19203,N_18894,N_18837);
or U19204 (N_19204,N_18965,N_18876);
and U19205 (N_19205,N_18885,N_18778);
nand U19206 (N_19206,N_18795,N_18852);
or U19207 (N_19207,N_18901,N_18885);
xnor U19208 (N_19208,N_18923,N_18775);
nor U19209 (N_19209,N_18792,N_18835);
or U19210 (N_19210,N_18993,N_18843);
nor U19211 (N_19211,N_18964,N_18896);
xnor U19212 (N_19212,N_18765,N_18787);
or U19213 (N_19213,N_18830,N_18960);
xor U19214 (N_19214,N_18924,N_18830);
xor U19215 (N_19215,N_18912,N_18843);
nand U19216 (N_19216,N_18860,N_18961);
xor U19217 (N_19217,N_18817,N_18919);
and U19218 (N_19218,N_18852,N_18998);
nor U19219 (N_19219,N_18829,N_18892);
and U19220 (N_19220,N_18838,N_18819);
or U19221 (N_19221,N_18815,N_18834);
nand U19222 (N_19222,N_18838,N_18921);
nand U19223 (N_19223,N_18785,N_18814);
nand U19224 (N_19224,N_18850,N_18833);
and U19225 (N_19225,N_18948,N_18921);
xor U19226 (N_19226,N_18918,N_18869);
and U19227 (N_19227,N_18865,N_18834);
nor U19228 (N_19228,N_18938,N_18962);
xor U19229 (N_19229,N_18995,N_18821);
xnor U19230 (N_19230,N_18974,N_18888);
and U19231 (N_19231,N_18772,N_18898);
nor U19232 (N_19232,N_18959,N_18833);
nand U19233 (N_19233,N_18895,N_18754);
nor U19234 (N_19234,N_18790,N_18827);
nand U19235 (N_19235,N_18859,N_18954);
and U19236 (N_19236,N_18856,N_18878);
and U19237 (N_19237,N_18855,N_18920);
nand U19238 (N_19238,N_18899,N_18840);
nor U19239 (N_19239,N_18939,N_18784);
xor U19240 (N_19240,N_18751,N_18969);
or U19241 (N_19241,N_18792,N_18908);
and U19242 (N_19242,N_18789,N_18840);
nand U19243 (N_19243,N_18928,N_18756);
nand U19244 (N_19244,N_18831,N_18782);
nand U19245 (N_19245,N_18963,N_18831);
or U19246 (N_19246,N_18932,N_18784);
or U19247 (N_19247,N_18992,N_18837);
nor U19248 (N_19248,N_18782,N_18788);
nor U19249 (N_19249,N_18915,N_18856);
or U19250 (N_19250,N_19212,N_19054);
or U19251 (N_19251,N_19150,N_19248);
nand U19252 (N_19252,N_19091,N_19053);
and U19253 (N_19253,N_19083,N_19061);
and U19254 (N_19254,N_19160,N_19206);
or U19255 (N_19255,N_19186,N_19159);
or U19256 (N_19256,N_19030,N_19217);
and U19257 (N_19257,N_19190,N_19137);
nor U19258 (N_19258,N_19135,N_19022);
xor U19259 (N_19259,N_19068,N_19020);
and U19260 (N_19260,N_19066,N_19173);
nor U19261 (N_19261,N_19152,N_19191);
nand U19262 (N_19262,N_19187,N_19034);
xor U19263 (N_19263,N_19193,N_19236);
and U19264 (N_19264,N_19126,N_19218);
and U19265 (N_19265,N_19085,N_19154);
or U19266 (N_19266,N_19112,N_19049);
nand U19267 (N_19267,N_19077,N_19165);
nand U19268 (N_19268,N_19104,N_19094);
or U19269 (N_19269,N_19241,N_19003);
nand U19270 (N_19270,N_19016,N_19011);
nor U19271 (N_19271,N_19082,N_19175);
nand U19272 (N_19272,N_19174,N_19099);
or U19273 (N_19273,N_19079,N_19111);
xor U19274 (N_19274,N_19025,N_19050);
nor U19275 (N_19275,N_19227,N_19007);
and U19276 (N_19276,N_19044,N_19105);
nand U19277 (N_19277,N_19033,N_19101);
or U19278 (N_19278,N_19113,N_19151);
and U19279 (N_19279,N_19225,N_19219);
nand U19280 (N_19280,N_19235,N_19169);
and U19281 (N_19281,N_19214,N_19084);
nor U19282 (N_19282,N_19095,N_19089);
and U19283 (N_19283,N_19189,N_19170);
and U19284 (N_19284,N_19001,N_19162);
and U19285 (N_19285,N_19223,N_19032);
xnor U19286 (N_19286,N_19136,N_19010);
nand U19287 (N_19287,N_19167,N_19243);
xnor U19288 (N_19288,N_19177,N_19188);
nor U19289 (N_19289,N_19209,N_19004);
or U19290 (N_19290,N_19106,N_19100);
nor U19291 (N_19291,N_19201,N_19071);
nor U19292 (N_19292,N_19140,N_19141);
or U19293 (N_19293,N_19143,N_19005);
xnor U19294 (N_19294,N_19184,N_19081);
nor U19295 (N_19295,N_19233,N_19014);
or U19296 (N_19296,N_19074,N_19045);
and U19297 (N_19297,N_19012,N_19062);
xor U19298 (N_19298,N_19072,N_19220);
and U19299 (N_19299,N_19052,N_19231);
or U19300 (N_19300,N_19164,N_19125);
and U19301 (N_19301,N_19073,N_19000);
and U19302 (N_19302,N_19192,N_19098);
nand U19303 (N_19303,N_19117,N_19148);
nor U19304 (N_19304,N_19119,N_19041);
nor U19305 (N_19305,N_19246,N_19158);
nand U19306 (N_19306,N_19021,N_19103);
nor U19307 (N_19307,N_19060,N_19096);
nor U19308 (N_19308,N_19038,N_19182);
xor U19309 (N_19309,N_19092,N_19240);
nor U19310 (N_19310,N_19087,N_19031);
nor U19311 (N_19311,N_19131,N_19245);
xnor U19312 (N_19312,N_19035,N_19069);
nand U19313 (N_19313,N_19207,N_19180);
or U19314 (N_19314,N_19139,N_19238);
nand U19315 (N_19315,N_19063,N_19161);
nor U19316 (N_19316,N_19056,N_19093);
nor U19317 (N_19317,N_19157,N_19009);
nor U19318 (N_19318,N_19055,N_19226);
and U19319 (N_19319,N_19086,N_19115);
nand U19320 (N_19320,N_19224,N_19121);
nand U19321 (N_19321,N_19002,N_19181);
xor U19322 (N_19322,N_19120,N_19039);
and U19323 (N_19323,N_19216,N_19163);
nor U19324 (N_19324,N_19183,N_19075);
nor U19325 (N_19325,N_19202,N_19067);
or U19326 (N_19326,N_19065,N_19208);
nor U19327 (N_19327,N_19176,N_19026);
or U19328 (N_19328,N_19048,N_19019);
and U19329 (N_19329,N_19229,N_19059);
or U19330 (N_19330,N_19239,N_19203);
or U19331 (N_19331,N_19211,N_19051);
or U19332 (N_19332,N_19128,N_19168);
nand U19333 (N_19333,N_19097,N_19197);
and U19334 (N_19334,N_19130,N_19247);
or U19335 (N_19335,N_19185,N_19123);
nand U19336 (N_19336,N_19043,N_19057);
nor U19337 (N_19337,N_19042,N_19204);
nand U19338 (N_19338,N_19027,N_19155);
or U19339 (N_19339,N_19237,N_19018);
nor U19340 (N_19340,N_19200,N_19198);
and U19341 (N_19341,N_19078,N_19144);
xor U19342 (N_19342,N_19156,N_19194);
nand U19343 (N_19343,N_19008,N_19088);
or U19344 (N_19344,N_19107,N_19172);
and U19345 (N_19345,N_19017,N_19047);
nor U19346 (N_19346,N_19064,N_19040);
nand U19347 (N_19347,N_19058,N_19110);
or U19348 (N_19348,N_19199,N_19195);
xor U19349 (N_19349,N_19171,N_19179);
or U19350 (N_19350,N_19132,N_19228);
xor U19351 (N_19351,N_19232,N_19178);
xor U19352 (N_19352,N_19127,N_19244);
or U19353 (N_19353,N_19210,N_19102);
and U19354 (N_19354,N_19114,N_19146);
xnor U19355 (N_19355,N_19076,N_19023);
or U19356 (N_19356,N_19129,N_19133);
xnor U19357 (N_19357,N_19138,N_19036);
or U19358 (N_19358,N_19221,N_19013);
and U19359 (N_19359,N_19145,N_19108);
nand U19360 (N_19360,N_19015,N_19090);
or U19361 (N_19361,N_19213,N_19142);
nand U19362 (N_19362,N_19028,N_19134);
nor U19363 (N_19363,N_19249,N_19122);
nand U19364 (N_19364,N_19109,N_19196);
nor U19365 (N_19365,N_19006,N_19124);
nor U19366 (N_19366,N_19205,N_19166);
nand U19367 (N_19367,N_19147,N_19024);
or U19368 (N_19368,N_19222,N_19149);
xnor U19369 (N_19369,N_19215,N_19242);
nor U19370 (N_19370,N_19230,N_19080);
and U19371 (N_19371,N_19037,N_19153);
and U19372 (N_19372,N_19234,N_19116);
xnor U19373 (N_19373,N_19118,N_19046);
and U19374 (N_19374,N_19029,N_19070);
nor U19375 (N_19375,N_19114,N_19157);
and U19376 (N_19376,N_19020,N_19057);
nand U19377 (N_19377,N_19061,N_19118);
xor U19378 (N_19378,N_19043,N_19167);
nand U19379 (N_19379,N_19172,N_19201);
or U19380 (N_19380,N_19166,N_19116);
nor U19381 (N_19381,N_19049,N_19092);
and U19382 (N_19382,N_19110,N_19001);
or U19383 (N_19383,N_19113,N_19234);
xor U19384 (N_19384,N_19027,N_19146);
or U19385 (N_19385,N_19001,N_19071);
nand U19386 (N_19386,N_19046,N_19060);
or U19387 (N_19387,N_19001,N_19187);
xnor U19388 (N_19388,N_19140,N_19039);
xnor U19389 (N_19389,N_19155,N_19214);
nand U19390 (N_19390,N_19172,N_19004);
and U19391 (N_19391,N_19149,N_19035);
or U19392 (N_19392,N_19182,N_19103);
nand U19393 (N_19393,N_19149,N_19153);
and U19394 (N_19394,N_19115,N_19042);
nor U19395 (N_19395,N_19010,N_19146);
nor U19396 (N_19396,N_19058,N_19031);
nand U19397 (N_19397,N_19128,N_19100);
and U19398 (N_19398,N_19106,N_19237);
nor U19399 (N_19399,N_19004,N_19061);
and U19400 (N_19400,N_19153,N_19245);
and U19401 (N_19401,N_19014,N_19167);
or U19402 (N_19402,N_19203,N_19148);
xor U19403 (N_19403,N_19051,N_19182);
and U19404 (N_19404,N_19078,N_19189);
xnor U19405 (N_19405,N_19161,N_19123);
nor U19406 (N_19406,N_19083,N_19020);
nand U19407 (N_19407,N_19113,N_19190);
xnor U19408 (N_19408,N_19237,N_19085);
xor U19409 (N_19409,N_19192,N_19171);
xor U19410 (N_19410,N_19094,N_19041);
and U19411 (N_19411,N_19179,N_19127);
nor U19412 (N_19412,N_19178,N_19020);
nor U19413 (N_19413,N_19240,N_19140);
nand U19414 (N_19414,N_19180,N_19106);
xor U19415 (N_19415,N_19225,N_19244);
nand U19416 (N_19416,N_19122,N_19129);
nor U19417 (N_19417,N_19166,N_19021);
nor U19418 (N_19418,N_19039,N_19172);
nor U19419 (N_19419,N_19014,N_19211);
and U19420 (N_19420,N_19039,N_19035);
xor U19421 (N_19421,N_19134,N_19071);
and U19422 (N_19422,N_19001,N_19163);
and U19423 (N_19423,N_19225,N_19140);
and U19424 (N_19424,N_19095,N_19229);
or U19425 (N_19425,N_19107,N_19211);
nand U19426 (N_19426,N_19135,N_19232);
nor U19427 (N_19427,N_19026,N_19090);
or U19428 (N_19428,N_19080,N_19175);
or U19429 (N_19429,N_19009,N_19160);
or U19430 (N_19430,N_19064,N_19134);
nor U19431 (N_19431,N_19159,N_19014);
xor U19432 (N_19432,N_19147,N_19083);
nor U19433 (N_19433,N_19001,N_19116);
nand U19434 (N_19434,N_19126,N_19069);
nor U19435 (N_19435,N_19172,N_19092);
nor U19436 (N_19436,N_19211,N_19013);
or U19437 (N_19437,N_19085,N_19136);
and U19438 (N_19438,N_19208,N_19172);
xnor U19439 (N_19439,N_19153,N_19045);
or U19440 (N_19440,N_19072,N_19104);
nor U19441 (N_19441,N_19133,N_19104);
nand U19442 (N_19442,N_19111,N_19158);
and U19443 (N_19443,N_19002,N_19241);
nand U19444 (N_19444,N_19095,N_19216);
and U19445 (N_19445,N_19103,N_19119);
xor U19446 (N_19446,N_19073,N_19127);
or U19447 (N_19447,N_19007,N_19098);
and U19448 (N_19448,N_19107,N_19090);
xor U19449 (N_19449,N_19216,N_19031);
and U19450 (N_19450,N_19171,N_19041);
and U19451 (N_19451,N_19061,N_19181);
xnor U19452 (N_19452,N_19009,N_19144);
and U19453 (N_19453,N_19169,N_19180);
nand U19454 (N_19454,N_19238,N_19183);
nand U19455 (N_19455,N_19158,N_19039);
or U19456 (N_19456,N_19106,N_19181);
and U19457 (N_19457,N_19046,N_19033);
or U19458 (N_19458,N_19006,N_19159);
xor U19459 (N_19459,N_19188,N_19058);
and U19460 (N_19460,N_19191,N_19068);
nand U19461 (N_19461,N_19143,N_19204);
or U19462 (N_19462,N_19166,N_19192);
or U19463 (N_19463,N_19238,N_19040);
or U19464 (N_19464,N_19009,N_19013);
and U19465 (N_19465,N_19065,N_19136);
nand U19466 (N_19466,N_19011,N_19164);
nor U19467 (N_19467,N_19205,N_19001);
xnor U19468 (N_19468,N_19211,N_19199);
xnor U19469 (N_19469,N_19014,N_19150);
and U19470 (N_19470,N_19034,N_19097);
xor U19471 (N_19471,N_19153,N_19100);
or U19472 (N_19472,N_19038,N_19235);
or U19473 (N_19473,N_19143,N_19116);
nand U19474 (N_19474,N_19198,N_19041);
nand U19475 (N_19475,N_19217,N_19050);
nand U19476 (N_19476,N_19070,N_19117);
xnor U19477 (N_19477,N_19049,N_19119);
nor U19478 (N_19478,N_19225,N_19025);
xnor U19479 (N_19479,N_19161,N_19133);
nor U19480 (N_19480,N_19036,N_19090);
and U19481 (N_19481,N_19157,N_19225);
and U19482 (N_19482,N_19191,N_19224);
nor U19483 (N_19483,N_19118,N_19105);
xor U19484 (N_19484,N_19032,N_19091);
and U19485 (N_19485,N_19108,N_19135);
nor U19486 (N_19486,N_19101,N_19201);
nor U19487 (N_19487,N_19093,N_19205);
nor U19488 (N_19488,N_19016,N_19208);
or U19489 (N_19489,N_19096,N_19038);
nor U19490 (N_19490,N_19088,N_19012);
or U19491 (N_19491,N_19110,N_19123);
nor U19492 (N_19492,N_19058,N_19052);
nand U19493 (N_19493,N_19128,N_19030);
or U19494 (N_19494,N_19235,N_19157);
nand U19495 (N_19495,N_19095,N_19118);
or U19496 (N_19496,N_19233,N_19166);
and U19497 (N_19497,N_19080,N_19121);
nand U19498 (N_19498,N_19000,N_19059);
or U19499 (N_19499,N_19038,N_19202);
nand U19500 (N_19500,N_19416,N_19371);
and U19501 (N_19501,N_19403,N_19455);
nor U19502 (N_19502,N_19389,N_19339);
nor U19503 (N_19503,N_19362,N_19357);
and U19504 (N_19504,N_19493,N_19476);
and U19505 (N_19505,N_19361,N_19359);
nor U19506 (N_19506,N_19278,N_19288);
nand U19507 (N_19507,N_19481,N_19447);
nand U19508 (N_19508,N_19282,N_19445);
nor U19509 (N_19509,N_19304,N_19433);
nand U19510 (N_19510,N_19457,N_19489);
nand U19511 (N_19511,N_19353,N_19270);
nand U19512 (N_19512,N_19318,N_19471);
nand U19513 (N_19513,N_19292,N_19460);
and U19514 (N_19514,N_19423,N_19297);
nor U19515 (N_19515,N_19451,N_19442);
nor U19516 (N_19516,N_19355,N_19333);
nand U19517 (N_19517,N_19364,N_19388);
or U19518 (N_19518,N_19310,N_19443);
nand U19519 (N_19519,N_19492,N_19430);
nand U19520 (N_19520,N_19463,N_19474);
nand U19521 (N_19521,N_19321,N_19348);
or U19522 (N_19522,N_19345,N_19448);
nor U19523 (N_19523,N_19346,N_19324);
and U19524 (N_19524,N_19486,N_19274);
nand U19525 (N_19525,N_19295,N_19382);
or U19526 (N_19526,N_19257,N_19342);
and U19527 (N_19527,N_19432,N_19469);
and U19528 (N_19528,N_19290,N_19478);
and U19529 (N_19529,N_19465,N_19289);
xnor U19530 (N_19530,N_19287,N_19259);
nor U19531 (N_19531,N_19250,N_19347);
xnor U19532 (N_19532,N_19373,N_19407);
nor U19533 (N_19533,N_19490,N_19496);
xnor U19534 (N_19534,N_19296,N_19273);
nor U19535 (N_19535,N_19375,N_19285);
or U19536 (N_19536,N_19323,N_19360);
xnor U19537 (N_19537,N_19409,N_19459);
nor U19538 (N_19538,N_19365,N_19383);
xnor U19539 (N_19539,N_19390,N_19370);
or U19540 (N_19540,N_19330,N_19434);
nor U19541 (N_19541,N_19425,N_19293);
nand U19542 (N_19542,N_19488,N_19284);
and U19543 (N_19543,N_19462,N_19393);
nor U19544 (N_19544,N_19429,N_19435);
nor U19545 (N_19545,N_19438,N_19466);
nand U19546 (N_19546,N_19379,N_19439);
nor U19547 (N_19547,N_19441,N_19475);
and U19548 (N_19548,N_19483,N_19453);
nand U19549 (N_19549,N_19314,N_19252);
nand U19550 (N_19550,N_19413,N_19408);
or U19551 (N_19551,N_19341,N_19380);
xnor U19552 (N_19552,N_19258,N_19385);
or U19553 (N_19553,N_19377,N_19480);
nor U19554 (N_19554,N_19387,N_19251);
nor U19555 (N_19555,N_19271,N_19300);
nor U19556 (N_19556,N_19283,N_19395);
and U19557 (N_19557,N_19322,N_19326);
nor U19558 (N_19558,N_19454,N_19349);
xor U19559 (N_19559,N_19468,N_19325);
nor U19560 (N_19560,N_19410,N_19456);
xnor U19561 (N_19561,N_19461,N_19277);
xor U19562 (N_19562,N_19320,N_19394);
nand U19563 (N_19563,N_19266,N_19426);
nor U19564 (N_19564,N_19263,N_19372);
or U19565 (N_19565,N_19446,N_19291);
nor U19566 (N_19566,N_19437,N_19401);
or U19567 (N_19567,N_19419,N_19449);
or U19568 (N_19568,N_19444,N_19422);
or U19569 (N_19569,N_19335,N_19491);
and U19570 (N_19570,N_19332,N_19298);
and U19571 (N_19571,N_19305,N_19269);
or U19572 (N_19572,N_19398,N_19315);
xor U19573 (N_19573,N_19399,N_19268);
and U19574 (N_19574,N_19427,N_19309);
and U19575 (N_19575,N_19458,N_19363);
and U19576 (N_19576,N_19344,N_19440);
and U19577 (N_19577,N_19487,N_19262);
and U19578 (N_19578,N_19436,N_19368);
nand U19579 (N_19579,N_19265,N_19261);
or U19580 (N_19580,N_19400,N_19473);
and U19581 (N_19581,N_19338,N_19350);
and U19582 (N_19582,N_19497,N_19319);
xor U19583 (N_19583,N_19358,N_19303);
xor U19584 (N_19584,N_19386,N_19470);
and U19585 (N_19585,N_19412,N_19381);
or U19586 (N_19586,N_19260,N_19498);
or U19587 (N_19587,N_19307,N_19331);
or U19588 (N_19588,N_19495,N_19391);
nand U19589 (N_19589,N_19316,N_19327);
and U19590 (N_19590,N_19313,N_19286);
or U19591 (N_19591,N_19351,N_19484);
and U19592 (N_19592,N_19255,N_19482);
xor U19593 (N_19593,N_19254,N_19450);
nor U19594 (N_19594,N_19276,N_19367);
or U19595 (N_19595,N_19421,N_19485);
nor U19596 (N_19596,N_19280,N_19317);
and U19597 (N_19597,N_19374,N_19301);
xnor U19598 (N_19598,N_19464,N_19376);
xnor U19599 (N_19599,N_19340,N_19329);
xor U19600 (N_19600,N_19499,N_19369);
nor U19601 (N_19601,N_19281,N_19431);
or U19602 (N_19602,N_19299,N_19334);
and U19603 (N_19603,N_19311,N_19272);
or U19604 (N_19604,N_19479,N_19253);
or U19605 (N_19605,N_19418,N_19343);
xor U19606 (N_19606,N_19414,N_19392);
or U19607 (N_19607,N_19396,N_19294);
or U19608 (N_19608,N_19306,N_19424);
nand U19609 (N_19609,N_19477,N_19302);
nand U19610 (N_19610,N_19402,N_19420);
xnor U19611 (N_19611,N_19452,N_19494);
or U19612 (N_19612,N_19354,N_19356);
nand U19613 (N_19613,N_19308,N_19279);
and U19614 (N_19614,N_19397,N_19472);
and U19615 (N_19615,N_19415,N_19352);
or U19616 (N_19616,N_19312,N_19467);
xor U19617 (N_19617,N_19406,N_19328);
nor U19618 (N_19618,N_19417,N_19337);
nand U19619 (N_19619,N_19336,N_19378);
or U19620 (N_19620,N_19275,N_19405);
nand U19621 (N_19621,N_19264,N_19256);
or U19622 (N_19622,N_19411,N_19366);
nand U19623 (N_19623,N_19428,N_19267);
or U19624 (N_19624,N_19404,N_19384);
or U19625 (N_19625,N_19302,N_19489);
xnor U19626 (N_19626,N_19431,N_19363);
nor U19627 (N_19627,N_19280,N_19338);
xnor U19628 (N_19628,N_19436,N_19353);
or U19629 (N_19629,N_19467,N_19485);
xnor U19630 (N_19630,N_19390,N_19379);
nor U19631 (N_19631,N_19450,N_19348);
or U19632 (N_19632,N_19426,N_19297);
nor U19633 (N_19633,N_19476,N_19339);
nor U19634 (N_19634,N_19332,N_19340);
or U19635 (N_19635,N_19262,N_19351);
and U19636 (N_19636,N_19266,N_19289);
or U19637 (N_19637,N_19382,N_19473);
and U19638 (N_19638,N_19316,N_19409);
and U19639 (N_19639,N_19334,N_19294);
nor U19640 (N_19640,N_19449,N_19488);
xor U19641 (N_19641,N_19317,N_19391);
nand U19642 (N_19642,N_19376,N_19399);
xor U19643 (N_19643,N_19427,N_19416);
and U19644 (N_19644,N_19478,N_19491);
nor U19645 (N_19645,N_19413,N_19271);
or U19646 (N_19646,N_19301,N_19278);
nand U19647 (N_19647,N_19337,N_19430);
nand U19648 (N_19648,N_19335,N_19251);
or U19649 (N_19649,N_19441,N_19439);
nand U19650 (N_19650,N_19377,N_19320);
nand U19651 (N_19651,N_19252,N_19380);
nand U19652 (N_19652,N_19398,N_19474);
and U19653 (N_19653,N_19429,N_19399);
and U19654 (N_19654,N_19360,N_19448);
nand U19655 (N_19655,N_19292,N_19429);
xor U19656 (N_19656,N_19483,N_19492);
nor U19657 (N_19657,N_19465,N_19453);
or U19658 (N_19658,N_19284,N_19471);
nand U19659 (N_19659,N_19345,N_19317);
or U19660 (N_19660,N_19374,N_19343);
and U19661 (N_19661,N_19296,N_19399);
xor U19662 (N_19662,N_19471,N_19267);
xnor U19663 (N_19663,N_19426,N_19490);
xnor U19664 (N_19664,N_19273,N_19366);
nand U19665 (N_19665,N_19306,N_19429);
xor U19666 (N_19666,N_19343,N_19298);
xor U19667 (N_19667,N_19491,N_19350);
and U19668 (N_19668,N_19270,N_19478);
nand U19669 (N_19669,N_19276,N_19475);
and U19670 (N_19670,N_19265,N_19459);
nor U19671 (N_19671,N_19455,N_19329);
nand U19672 (N_19672,N_19390,N_19441);
and U19673 (N_19673,N_19423,N_19446);
nor U19674 (N_19674,N_19369,N_19398);
and U19675 (N_19675,N_19471,N_19333);
and U19676 (N_19676,N_19401,N_19490);
or U19677 (N_19677,N_19432,N_19456);
or U19678 (N_19678,N_19267,N_19404);
and U19679 (N_19679,N_19400,N_19346);
nand U19680 (N_19680,N_19455,N_19292);
or U19681 (N_19681,N_19367,N_19492);
xnor U19682 (N_19682,N_19327,N_19392);
xor U19683 (N_19683,N_19486,N_19363);
nand U19684 (N_19684,N_19300,N_19351);
nand U19685 (N_19685,N_19375,N_19302);
nand U19686 (N_19686,N_19462,N_19471);
and U19687 (N_19687,N_19477,N_19333);
nor U19688 (N_19688,N_19381,N_19394);
or U19689 (N_19689,N_19447,N_19317);
or U19690 (N_19690,N_19383,N_19340);
xor U19691 (N_19691,N_19296,N_19348);
nor U19692 (N_19692,N_19352,N_19360);
xnor U19693 (N_19693,N_19341,N_19388);
or U19694 (N_19694,N_19321,N_19265);
nand U19695 (N_19695,N_19350,N_19374);
nor U19696 (N_19696,N_19374,N_19329);
nor U19697 (N_19697,N_19422,N_19309);
nand U19698 (N_19698,N_19406,N_19382);
or U19699 (N_19699,N_19284,N_19250);
xnor U19700 (N_19700,N_19315,N_19378);
nor U19701 (N_19701,N_19291,N_19267);
xnor U19702 (N_19702,N_19303,N_19384);
nand U19703 (N_19703,N_19433,N_19307);
xnor U19704 (N_19704,N_19380,N_19464);
nand U19705 (N_19705,N_19398,N_19308);
nand U19706 (N_19706,N_19498,N_19495);
xor U19707 (N_19707,N_19367,N_19410);
nand U19708 (N_19708,N_19302,N_19306);
xnor U19709 (N_19709,N_19346,N_19291);
xor U19710 (N_19710,N_19439,N_19408);
nor U19711 (N_19711,N_19479,N_19302);
nand U19712 (N_19712,N_19251,N_19334);
or U19713 (N_19713,N_19423,N_19453);
and U19714 (N_19714,N_19327,N_19376);
xor U19715 (N_19715,N_19362,N_19441);
and U19716 (N_19716,N_19412,N_19489);
nor U19717 (N_19717,N_19493,N_19400);
or U19718 (N_19718,N_19407,N_19316);
or U19719 (N_19719,N_19308,N_19484);
or U19720 (N_19720,N_19443,N_19307);
and U19721 (N_19721,N_19376,N_19322);
and U19722 (N_19722,N_19392,N_19273);
nor U19723 (N_19723,N_19353,N_19393);
or U19724 (N_19724,N_19449,N_19412);
nor U19725 (N_19725,N_19296,N_19395);
and U19726 (N_19726,N_19275,N_19430);
and U19727 (N_19727,N_19406,N_19280);
xor U19728 (N_19728,N_19388,N_19483);
xnor U19729 (N_19729,N_19280,N_19360);
nand U19730 (N_19730,N_19400,N_19290);
and U19731 (N_19731,N_19339,N_19498);
or U19732 (N_19732,N_19330,N_19485);
or U19733 (N_19733,N_19323,N_19274);
or U19734 (N_19734,N_19491,N_19325);
xnor U19735 (N_19735,N_19271,N_19317);
xor U19736 (N_19736,N_19361,N_19435);
or U19737 (N_19737,N_19475,N_19499);
nand U19738 (N_19738,N_19382,N_19398);
or U19739 (N_19739,N_19342,N_19356);
or U19740 (N_19740,N_19335,N_19294);
nor U19741 (N_19741,N_19483,N_19265);
nand U19742 (N_19742,N_19385,N_19443);
and U19743 (N_19743,N_19261,N_19365);
nand U19744 (N_19744,N_19348,N_19353);
nor U19745 (N_19745,N_19375,N_19424);
and U19746 (N_19746,N_19334,N_19353);
xnor U19747 (N_19747,N_19465,N_19425);
and U19748 (N_19748,N_19403,N_19435);
and U19749 (N_19749,N_19389,N_19348);
and U19750 (N_19750,N_19546,N_19533);
nand U19751 (N_19751,N_19604,N_19559);
xor U19752 (N_19752,N_19625,N_19588);
or U19753 (N_19753,N_19608,N_19566);
and U19754 (N_19754,N_19662,N_19554);
and U19755 (N_19755,N_19666,N_19603);
nor U19756 (N_19756,N_19563,N_19636);
xnor U19757 (N_19757,N_19530,N_19702);
nor U19758 (N_19758,N_19526,N_19631);
nand U19759 (N_19759,N_19722,N_19705);
nand U19760 (N_19760,N_19502,N_19508);
xor U19761 (N_19761,N_19657,N_19744);
nand U19762 (N_19762,N_19684,N_19735);
nand U19763 (N_19763,N_19598,N_19544);
nor U19764 (N_19764,N_19585,N_19632);
or U19765 (N_19765,N_19556,N_19540);
and U19766 (N_19766,N_19504,N_19527);
xnor U19767 (N_19767,N_19561,N_19635);
or U19768 (N_19768,N_19541,N_19693);
and U19769 (N_19769,N_19673,N_19731);
nor U19770 (N_19770,N_19729,N_19738);
and U19771 (N_19771,N_19617,N_19507);
xnor U19772 (N_19772,N_19615,N_19688);
or U19773 (N_19773,N_19686,N_19601);
nand U19774 (N_19774,N_19647,N_19741);
or U19775 (N_19775,N_19536,N_19614);
nor U19776 (N_19776,N_19624,N_19745);
and U19777 (N_19777,N_19720,N_19558);
or U19778 (N_19778,N_19668,N_19611);
xor U19779 (N_19779,N_19574,N_19512);
nor U19780 (N_19780,N_19732,N_19648);
nor U19781 (N_19781,N_19630,N_19733);
xnor U19782 (N_19782,N_19743,N_19538);
or U19783 (N_19783,N_19710,N_19695);
xnor U19784 (N_19784,N_19620,N_19643);
xor U19785 (N_19785,N_19580,N_19728);
and U19786 (N_19786,N_19618,N_19523);
nand U19787 (N_19787,N_19678,N_19597);
and U19788 (N_19788,N_19547,N_19716);
or U19789 (N_19789,N_19736,N_19609);
nand U19790 (N_19790,N_19665,N_19641);
and U19791 (N_19791,N_19714,N_19582);
nor U19792 (N_19792,N_19669,N_19542);
and U19793 (N_19793,N_19687,N_19593);
or U19794 (N_19794,N_19658,N_19555);
nand U19795 (N_19795,N_19596,N_19589);
nand U19796 (N_19796,N_19592,N_19653);
nor U19797 (N_19797,N_19740,N_19590);
or U19798 (N_19798,N_19660,N_19628);
and U19799 (N_19799,N_19683,N_19664);
and U19800 (N_19800,N_19500,N_19637);
or U19801 (N_19801,N_19706,N_19699);
xor U19802 (N_19802,N_19537,N_19517);
xnor U19803 (N_19803,N_19676,N_19513);
xnor U19804 (N_19804,N_19718,N_19511);
nand U19805 (N_19805,N_19654,N_19514);
or U19806 (N_19806,N_19655,N_19713);
xnor U19807 (N_19807,N_19642,N_19534);
and U19808 (N_19808,N_19570,N_19501);
xnor U19809 (N_19809,N_19646,N_19724);
and U19810 (N_19810,N_19562,N_19606);
nor U19811 (N_19811,N_19553,N_19730);
or U19812 (N_19812,N_19616,N_19605);
nand U19813 (N_19813,N_19645,N_19583);
nor U19814 (N_19814,N_19633,N_19519);
or U19815 (N_19815,N_19564,N_19712);
or U19816 (N_19816,N_19667,N_19621);
nand U19817 (N_19817,N_19721,N_19602);
nand U19818 (N_19818,N_19515,N_19539);
or U19819 (N_19819,N_19595,N_19685);
nand U19820 (N_19820,N_19650,N_19579);
or U19821 (N_19821,N_19652,N_19619);
and U19822 (N_19822,N_19516,N_19677);
and U19823 (N_19823,N_19622,N_19510);
and U19824 (N_19824,N_19569,N_19709);
or U19825 (N_19825,N_19734,N_19529);
nand U19826 (N_19826,N_19679,N_19656);
nand U19827 (N_19827,N_19726,N_19692);
nand U19828 (N_19828,N_19703,N_19551);
nor U19829 (N_19829,N_19575,N_19557);
nand U19830 (N_19830,N_19661,N_19587);
xor U19831 (N_19831,N_19638,N_19649);
or U19832 (N_19832,N_19503,N_19531);
nand U19833 (N_19833,N_19576,N_19634);
nand U19834 (N_19834,N_19535,N_19629);
nor U19835 (N_19835,N_19715,N_19675);
xor U19836 (N_19836,N_19701,N_19690);
xnor U19837 (N_19837,N_19742,N_19543);
nor U19838 (N_19838,N_19600,N_19567);
nor U19839 (N_19839,N_19613,N_19651);
nand U19840 (N_19840,N_19694,N_19505);
and U19841 (N_19841,N_19626,N_19689);
or U19842 (N_19842,N_19640,N_19571);
nor U19843 (N_19843,N_19581,N_19627);
and U19844 (N_19844,N_19698,N_19739);
nand U19845 (N_19845,N_19568,N_19548);
nand U19846 (N_19846,N_19607,N_19696);
and U19847 (N_19847,N_19521,N_19525);
or U19848 (N_19848,N_19680,N_19719);
nor U19849 (N_19849,N_19746,N_19747);
nand U19850 (N_19850,N_19586,N_19725);
nand U19851 (N_19851,N_19578,N_19599);
or U19852 (N_19852,N_19520,N_19584);
nor U19853 (N_19853,N_19727,N_19681);
or U19854 (N_19854,N_19623,N_19691);
nand U19855 (N_19855,N_19708,N_19672);
nor U19856 (N_19856,N_19524,N_19572);
nor U19857 (N_19857,N_19545,N_19518);
nand U19858 (N_19858,N_19549,N_19552);
xnor U19859 (N_19859,N_19697,N_19573);
nor U19860 (N_19860,N_19700,N_19612);
nor U19861 (N_19861,N_19682,N_19594);
nor U19862 (N_19862,N_19748,N_19528);
xor U19863 (N_19863,N_19717,N_19670);
nor U19864 (N_19864,N_19737,N_19711);
nand U19865 (N_19865,N_19639,N_19610);
nor U19866 (N_19866,N_19707,N_19674);
nand U19867 (N_19867,N_19671,N_19659);
and U19868 (N_19868,N_19532,N_19644);
xor U19869 (N_19869,N_19749,N_19509);
nor U19870 (N_19870,N_19704,N_19560);
xnor U19871 (N_19871,N_19663,N_19565);
nor U19872 (N_19872,N_19591,N_19550);
nand U19873 (N_19873,N_19522,N_19577);
or U19874 (N_19874,N_19506,N_19723);
xnor U19875 (N_19875,N_19619,N_19507);
nand U19876 (N_19876,N_19511,N_19669);
xnor U19877 (N_19877,N_19640,N_19732);
xor U19878 (N_19878,N_19737,N_19503);
nand U19879 (N_19879,N_19647,N_19607);
xor U19880 (N_19880,N_19526,N_19609);
xor U19881 (N_19881,N_19665,N_19656);
nor U19882 (N_19882,N_19577,N_19520);
or U19883 (N_19883,N_19680,N_19599);
and U19884 (N_19884,N_19505,N_19562);
nor U19885 (N_19885,N_19539,N_19584);
xor U19886 (N_19886,N_19644,N_19727);
xnor U19887 (N_19887,N_19622,N_19625);
nand U19888 (N_19888,N_19652,N_19515);
or U19889 (N_19889,N_19560,N_19702);
nor U19890 (N_19890,N_19678,N_19558);
nor U19891 (N_19891,N_19570,N_19678);
nand U19892 (N_19892,N_19553,N_19530);
nand U19893 (N_19893,N_19601,N_19572);
nand U19894 (N_19894,N_19588,N_19728);
or U19895 (N_19895,N_19735,N_19604);
nand U19896 (N_19896,N_19637,N_19701);
nor U19897 (N_19897,N_19723,N_19573);
nand U19898 (N_19898,N_19532,N_19639);
nor U19899 (N_19899,N_19574,N_19552);
xor U19900 (N_19900,N_19537,N_19500);
nor U19901 (N_19901,N_19609,N_19652);
nor U19902 (N_19902,N_19652,N_19529);
and U19903 (N_19903,N_19652,N_19575);
or U19904 (N_19904,N_19668,N_19613);
or U19905 (N_19905,N_19528,N_19709);
and U19906 (N_19906,N_19650,N_19696);
nand U19907 (N_19907,N_19635,N_19535);
or U19908 (N_19908,N_19722,N_19736);
or U19909 (N_19909,N_19608,N_19613);
nand U19910 (N_19910,N_19667,N_19674);
and U19911 (N_19911,N_19546,N_19628);
or U19912 (N_19912,N_19601,N_19505);
nor U19913 (N_19913,N_19551,N_19573);
nand U19914 (N_19914,N_19610,N_19570);
nor U19915 (N_19915,N_19543,N_19557);
and U19916 (N_19916,N_19553,N_19557);
and U19917 (N_19917,N_19650,N_19631);
or U19918 (N_19918,N_19680,N_19706);
and U19919 (N_19919,N_19647,N_19700);
nand U19920 (N_19920,N_19535,N_19608);
and U19921 (N_19921,N_19655,N_19690);
nor U19922 (N_19922,N_19548,N_19739);
xnor U19923 (N_19923,N_19607,N_19636);
nor U19924 (N_19924,N_19684,N_19670);
xor U19925 (N_19925,N_19519,N_19569);
and U19926 (N_19926,N_19605,N_19510);
xnor U19927 (N_19927,N_19573,N_19580);
and U19928 (N_19928,N_19599,N_19604);
and U19929 (N_19929,N_19739,N_19675);
or U19930 (N_19930,N_19580,N_19741);
and U19931 (N_19931,N_19713,N_19542);
and U19932 (N_19932,N_19616,N_19533);
and U19933 (N_19933,N_19702,N_19719);
or U19934 (N_19934,N_19715,N_19658);
or U19935 (N_19935,N_19657,N_19536);
or U19936 (N_19936,N_19581,N_19555);
nand U19937 (N_19937,N_19686,N_19623);
and U19938 (N_19938,N_19630,N_19702);
nor U19939 (N_19939,N_19582,N_19617);
and U19940 (N_19940,N_19732,N_19662);
nand U19941 (N_19941,N_19647,N_19676);
and U19942 (N_19942,N_19537,N_19552);
nor U19943 (N_19943,N_19530,N_19740);
or U19944 (N_19944,N_19563,N_19543);
nor U19945 (N_19945,N_19597,N_19540);
xor U19946 (N_19946,N_19551,N_19745);
or U19947 (N_19947,N_19570,N_19542);
and U19948 (N_19948,N_19556,N_19631);
nor U19949 (N_19949,N_19724,N_19634);
nor U19950 (N_19950,N_19620,N_19520);
nor U19951 (N_19951,N_19572,N_19641);
nor U19952 (N_19952,N_19740,N_19661);
or U19953 (N_19953,N_19630,N_19601);
or U19954 (N_19954,N_19517,N_19632);
xor U19955 (N_19955,N_19531,N_19616);
nand U19956 (N_19956,N_19723,N_19530);
xor U19957 (N_19957,N_19537,N_19748);
nor U19958 (N_19958,N_19558,N_19510);
xor U19959 (N_19959,N_19726,N_19538);
xnor U19960 (N_19960,N_19620,N_19604);
xnor U19961 (N_19961,N_19677,N_19644);
nand U19962 (N_19962,N_19685,N_19612);
nor U19963 (N_19963,N_19683,N_19515);
or U19964 (N_19964,N_19723,N_19729);
nand U19965 (N_19965,N_19663,N_19562);
and U19966 (N_19966,N_19530,N_19677);
and U19967 (N_19967,N_19638,N_19730);
and U19968 (N_19968,N_19542,N_19575);
xor U19969 (N_19969,N_19509,N_19614);
nand U19970 (N_19970,N_19652,N_19597);
and U19971 (N_19971,N_19728,N_19704);
and U19972 (N_19972,N_19648,N_19599);
nor U19973 (N_19973,N_19603,N_19547);
nand U19974 (N_19974,N_19579,N_19687);
xnor U19975 (N_19975,N_19590,N_19557);
or U19976 (N_19976,N_19504,N_19741);
nor U19977 (N_19977,N_19748,N_19686);
nand U19978 (N_19978,N_19563,N_19677);
nor U19979 (N_19979,N_19630,N_19692);
and U19980 (N_19980,N_19708,N_19657);
or U19981 (N_19981,N_19576,N_19525);
and U19982 (N_19982,N_19696,N_19663);
nor U19983 (N_19983,N_19713,N_19676);
or U19984 (N_19984,N_19679,N_19544);
or U19985 (N_19985,N_19682,N_19509);
and U19986 (N_19986,N_19531,N_19508);
nand U19987 (N_19987,N_19520,N_19749);
or U19988 (N_19988,N_19558,N_19636);
nand U19989 (N_19989,N_19556,N_19590);
nor U19990 (N_19990,N_19550,N_19510);
and U19991 (N_19991,N_19544,N_19717);
nor U19992 (N_19992,N_19713,N_19548);
or U19993 (N_19993,N_19558,N_19666);
nand U19994 (N_19994,N_19610,N_19749);
or U19995 (N_19995,N_19502,N_19740);
or U19996 (N_19996,N_19513,N_19565);
xor U19997 (N_19997,N_19668,N_19582);
nor U19998 (N_19998,N_19716,N_19524);
and U19999 (N_19999,N_19658,N_19688);
and UO_0 (O_0,N_19949,N_19920);
nor UO_1 (O_1,N_19753,N_19944);
nor UO_2 (O_2,N_19890,N_19881);
xor UO_3 (O_3,N_19819,N_19948);
and UO_4 (O_4,N_19969,N_19817);
nor UO_5 (O_5,N_19932,N_19763);
or UO_6 (O_6,N_19853,N_19955);
or UO_7 (O_7,N_19901,N_19892);
nor UO_8 (O_8,N_19906,N_19918);
xor UO_9 (O_9,N_19751,N_19876);
nand UO_10 (O_10,N_19985,N_19992);
or UO_11 (O_11,N_19778,N_19858);
xor UO_12 (O_12,N_19889,N_19841);
and UO_13 (O_13,N_19910,N_19830);
and UO_14 (O_14,N_19986,N_19801);
nor UO_15 (O_15,N_19759,N_19800);
or UO_16 (O_16,N_19884,N_19869);
xnor UO_17 (O_17,N_19839,N_19861);
nand UO_18 (O_18,N_19963,N_19996);
and UO_19 (O_19,N_19849,N_19882);
nor UO_20 (O_20,N_19850,N_19950);
xnor UO_21 (O_21,N_19919,N_19938);
nor UO_22 (O_22,N_19872,N_19810);
and UO_23 (O_23,N_19905,N_19788);
nand UO_24 (O_24,N_19897,N_19988);
nand UO_25 (O_25,N_19979,N_19762);
nand UO_26 (O_26,N_19870,N_19842);
nand UO_27 (O_27,N_19931,N_19991);
and UO_28 (O_28,N_19813,N_19898);
and UO_29 (O_29,N_19832,N_19798);
nor UO_30 (O_30,N_19771,N_19846);
or UO_31 (O_31,N_19895,N_19868);
nand UO_32 (O_32,N_19930,N_19886);
nor UO_33 (O_33,N_19761,N_19987);
or UO_34 (O_34,N_19780,N_19767);
nor UO_35 (O_35,N_19785,N_19903);
or UO_36 (O_36,N_19925,N_19994);
and UO_37 (O_37,N_19779,N_19885);
nor UO_38 (O_38,N_19777,N_19834);
and UO_39 (O_39,N_19847,N_19999);
nand UO_40 (O_40,N_19860,N_19917);
xor UO_41 (O_41,N_19758,N_19899);
xor UO_42 (O_42,N_19995,N_19790);
nor UO_43 (O_43,N_19802,N_19833);
nand UO_44 (O_44,N_19808,N_19928);
and UO_45 (O_45,N_19964,N_19970);
nand UO_46 (O_46,N_19982,N_19936);
nor UO_47 (O_47,N_19806,N_19826);
and UO_48 (O_48,N_19803,N_19824);
xor UO_49 (O_49,N_19837,N_19854);
xor UO_50 (O_50,N_19939,N_19945);
nor UO_51 (O_51,N_19768,N_19909);
nand UO_52 (O_52,N_19941,N_19975);
xnor UO_53 (O_53,N_19840,N_19951);
and UO_54 (O_54,N_19937,N_19794);
xor UO_55 (O_55,N_19760,N_19815);
xnor UO_56 (O_56,N_19913,N_19754);
xor UO_57 (O_57,N_19998,N_19864);
or UO_58 (O_58,N_19799,N_19835);
nor UO_59 (O_59,N_19923,N_19980);
and UO_60 (O_60,N_19770,N_19848);
nand UO_61 (O_61,N_19829,N_19862);
xor UO_62 (O_62,N_19844,N_19871);
or UO_63 (O_63,N_19878,N_19933);
nand UO_64 (O_64,N_19879,N_19900);
and UO_65 (O_65,N_19911,N_19797);
or UO_66 (O_66,N_19765,N_19965);
nor UO_67 (O_67,N_19877,N_19859);
and UO_68 (O_68,N_19784,N_19821);
xor UO_69 (O_69,N_19880,N_19831);
or UO_70 (O_70,N_19775,N_19855);
or UO_71 (O_71,N_19795,N_19883);
and UO_72 (O_72,N_19845,N_19791);
or UO_73 (O_73,N_19953,N_19971);
or UO_74 (O_74,N_19894,N_19968);
nor UO_75 (O_75,N_19907,N_19764);
and UO_76 (O_76,N_19924,N_19921);
nor UO_77 (O_77,N_19960,N_19787);
and UO_78 (O_78,N_19789,N_19843);
nor UO_79 (O_79,N_19954,N_19772);
and UO_80 (O_80,N_19774,N_19974);
nor UO_81 (O_81,N_19927,N_19926);
or UO_82 (O_82,N_19782,N_19958);
nor UO_83 (O_83,N_19750,N_19993);
nand UO_84 (O_84,N_19793,N_19783);
or UO_85 (O_85,N_19755,N_19989);
nand UO_86 (O_86,N_19873,N_19896);
and UO_87 (O_87,N_19916,N_19922);
nor UO_88 (O_88,N_19786,N_19792);
and UO_89 (O_89,N_19856,N_19959);
or UO_90 (O_90,N_19891,N_19934);
nand UO_91 (O_91,N_19947,N_19943);
or UO_92 (O_92,N_19972,N_19887);
nor UO_93 (O_93,N_19807,N_19940);
nand UO_94 (O_94,N_19852,N_19966);
nor UO_95 (O_95,N_19838,N_19804);
or UO_96 (O_96,N_19820,N_19981);
and UO_97 (O_97,N_19851,N_19956);
or UO_98 (O_98,N_19863,N_19866);
and UO_99 (O_99,N_19978,N_19822);
nor UO_100 (O_100,N_19756,N_19912);
nor UO_101 (O_101,N_19888,N_19962);
nand UO_102 (O_102,N_19961,N_19929);
nor UO_103 (O_103,N_19990,N_19752);
xnor UO_104 (O_104,N_19997,N_19893);
nand UO_105 (O_105,N_19874,N_19828);
nor UO_106 (O_106,N_19812,N_19823);
xnor UO_107 (O_107,N_19816,N_19867);
nor UO_108 (O_108,N_19857,N_19757);
xor UO_109 (O_109,N_19827,N_19952);
nor UO_110 (O_110,N_19976,N_19904);
or UO_111 (O_111,N_19984,N_19865);
or UO_112 (O_112,N_19957,N_19946);
and UO_113 (O_113,N_19942,N_19796);
or UO_114 (O_114,N_19983,N_19809);
xnor UO_115 (O_115,N_19776,N_19805);
xor UO_116 (O_116,N_19814,N_19902);
nand UO_117 (O_117,N_19773,N_19977);
xor UO_118 (O_118,N_19811,N_19875);
and UO_119 (O_119,N_19818,N_19973);
xnor UO_120 (O_120,N_19836,N_19967);
nor UO_121 (O_121,N_19908,N_19825);
or UO_122 (O_122,N_19935,N_19766);
or UO_123 (O_123,N_19915,N_19781);
and UO_124 (O_124,N_19914,N_19769);
or UO_125 (O_125,N_19925,N_19833);
and UO_126 (O_126,N_19781,N_19972);
nand UO_127 (O_127,N_19835,N_19827);
nor UO_128 (O_128,N_19922,N_19783);
nand UO_129 (O_129,N_19969,N_19991);
xor UO_130 (O_130,N_19897,N_19839);
nor UO_131 (O_131,N_19882,N_19902);
nand UO_132 (O_132,N_19957,N_19884);
or UO_133 (O_133,N_19911,N_19906);
nor UO_134 (O_134,N_19957,N_19878);
nand UO_135 (O_135,N_19875,N_19939);
and UO_136 (O_136,N_19770,N_19984);
nor UO_137 (O_137,N_19953,N_19818);
xnor UO_138 (O_138,N_19964,N_19974);
and UO_139 (O_139,N_19946,N_19893);
or UO_140 (O_140,N_19825,N_19982);
or UO_141 (O_141,N_19882,N_19925);
nor UO_142 (O_142,N_19760,N_19820);
nand UO_143 (O_143,N_19809,N_19970);
and UO_144 (O_144,N_19914,N_19779);
xnor UO_145 (O_145,N_19750,N_19828);
xnor UO_146 (O_146,N_19753,N_19856);
nor UO_147 (O_147,N_19777,N_19931);
nor UO_148 (O_148,N_19786,N_19827);
and UO_149 (O_149,N_19891,N_19828);
nand UO_150 (O_150,N_19956,N_19762);
and UO_151 (O_151,N_19769,N_19973);
nand UO_152 (O_152,N_19760,N_19838);
xor UO_153 (O_153,N_19877,N_19891);
and UO_154 (O_154,N_19889,N_19799);
xor UO_155 (O_155,N_19923,N_19786);
nand UO_156 (O_156,N_19867,N_19945);
xor UO_157 (O_157,N_19782,N_19929);
or UO_158 (O_158,N_19754,N_19967);
nor UO_159 (O_159,N_19930,N_19952);
nor UO_160 (O_160,N_19922,N_19886);
and UO_161 (O_161,N_19929,N_19899);
nand UO_162 (O_162,N_19765,N_19848);
nand UO_163 (O_163,N_19847,N_19932);
and UO_164 (O_164,N_19902,N_19916);
or UO_165 (O_165,N_19910,N_19834);
or UO_166 (O_166,N_19844,N_19828);
xor UO_167 (O_167,N_19816,N_19916);
and UO_168 (O_168,N_19888,N_19940);
nand UO_169 (O_169,N_19812,N_19929);
xor UO_170 (O_170,N_19908,N_19932);
nand UO_171 (O_171,N_19881,N_19822);
nand UO_172 (O_172,N_19916,N_19898);
nand UO_173 (O_173,N_19818,N_19967);
nand UO_174 (O_174,N_19853,N_19937);
and UO_175 (O_175,N_19799,N_19896);
and UO_176 (O_176,N_19842,N_19989);
nand UO_177 (O_177,N_19947,N_19850);
xor UO_178 (O_178,N_19931,N_19781);
xor UO_179 (O_179,N_19888,N_19904);
nor UO_180 (O_180,N_19872,N_19946);
nand UO_181 (O_181,N_19763,N_19916);
nand UO_182 (O_182,N_19808,N_19932);
and UO_183 (O_183,N_19803,N_19843);
nand UO_184 (O_184,N_19804,N_19979);
or UO_185 (O_185,N_19767,N_19925);
nor UO_186 (O_186,N_19942,N_19814);
or UO_187 (O_187,N_19833,N_19969);
nor UO_188 (O_188,N_19946,N_19944);
xor UO_189 (O_189,N_19798,N_19845);
nand UO_190 (O_190,N_19892,N_19816);
and UO_191 (O_191,N_19964,N_19779);
nand UO_192 (O_192,N_19871,N_19881);
or UO_193 (O_193,N_19823,N_19972);
nand UO_194 (O_194,N_19969,N_19836);
nand UO_195 (O_195,N_19893,N_19856);
nand UO_196 (O_196,N_19915,N_19862);
nand UO_197 (O_197,N_19859,N_19923);
and UO_198 (O_198,N_19974,N_19950);
xnor UO_199 (O_199,N_19977,N_19771);
nor UO_200 (O_200,N_19968,N_19950);
xor UO_201 (O_201,N_19975,N_19820);
xnor UO_202 (O_202,N_19882,N_19762);
or UO_203 (O_203,N_19960,N_19785);
nor UO_204 (O_204,N_19758,N_19836);
xnor UO_205 (O_205,N_19923,N_19982);
xor UO_206 (O_206,N_19944,N_19847);
nand UO_207 (O_207,N_19758,N_19973);
xor UO_208 (O_208,N_19866,N_19884);
xnor UO_209 (O_209,N_19845,N_19776);
nand UO_210 (O_210,N_19824,N_19906);
nor UO_211 (O_211,N_19784,N_19834);
nor UO_212 (O_212,N_19864,N_19777);
nand UO_213 (O_213,N_19888,N_19953);
and UO_214 (O_214,N_19817,N_19991);
xnor UO_215 (O_215,N_19952,N_19838);
xnor UO_216 (O_216,N_19950,N_19960);
nand UO_217 (O_217,N_19962,N_19936);
and UO_218 (O_218,N_19890,N_19984);
xor UO_219 (O_219,N_19782,N_19809);
nand UO_220 (O_220,N_19979,N_19777);
xor UO_221 (O_221,N_19789,N_19892);
or UO_222 (O_222,N_19871,N_19795);
xnor UO_223 (O_223,N_19903,N_19970);
or UO_224 (O_224,N_19787,N_19982);
nor UO_225 (O_225,N_19792,N_19820);
nand UO_226 (O_226,N_19754,N_19785);
or UO_227 (O_227,N_19757,N_19922);
or UO_228 (O_228,N_19917,N_19931);
xor UO_229 (O_229,N_19822,N_19863);
nand UO_230 (O_230,N_19819,N_19871);
and UO_231 (O_231,N_19900,N_19850);
or UO_232 (O_232,N_19788,N_19883);
xnor UO_233 (O_233,N_19993,N_19890);
nand UO_234 (O_234,N_19813,N_19893);
nand UO_235 (O_235,N_19866,N_19811);
nand UO_236 (O_236,N_19753,N_19813);
nand UO_237 (O_237,N_19988,N_19809);
xor UO_238 (O_238,N_19836,N_19817);
xnor UO_239 (O_239,N_19777,N_19858);
nand UO_240 (O_240,N_19802,N_19987);
and UO_241 (O_241,N_19988,N_19806);
nand UO_242 (O_242,N_19987,N_19778);
or UO_243 (O_243,N_19869,N_19779);
and UO_244 (O_244,N_19937,N_19993);
and UO_245 (O_245,N_19766,N_19980);
nor UO_246 (O_246,N_19988,N_19778);
nand UO_247 (O_247,N_19801,N_19859);
and UO_248 (O_248,N_19863,N_19988);
nor UO_249 (O_249,N_19785,N_19871);
and UO_250 (O_250,N_19939,N_19979);
nor UO_251 (O_251,N_19869,N_19907);
xnor UO_252 (O_252,N_19846,N_19777);
xor UO_253 (O_253,N_19961,N_19886);
nand UO_254 (O_254,N_19902,N_19841);
and UO_255 (O_255,N_19846,N_19934);
nand UO_256 (O_256,N_19917,N_19820);
or UO_257 (O_257,N_19954,N_19883);
and UO_258 (O_258,N_19751,N_19818);
xor UO_259 (O_259,N_19818,N_19898);
nand UO_260 (O_260,N_19919,N_19923);
nand UO_261 (O_261,N_19919,N_19904);
nand UO_262 (O_262,N_19793,N_19817);
nor UO_263 (O_263,N_19988,N_19850);
xnor UO_264 (O_264,N_19878,N_19851);
or UO_265 (O_265,N_19984,N_19912);
or UO_266 (O_266,N_19755,N_19981);
nand UO_267 (O_267,N_19936,N_19755);
and UO_268 (O_268,N_19940,N_19948);
or UO_269 (O_269,N_19834,N_19906);
or UO_270 (O_270,N_19944,N_19788);
nor UO_271 (O_271,N_19816,N_19868);
nand UO_272 (O_272,N_19979,N_19941);
or UO_273 (O_273,N_19836,N_19915);
and UO_274 (O_274,N_19795,N_19813);
nand UO_275 (O_275,N_19872,N_19847);
nand UO_276 (O_276,N_19827,N_19780);
nand UO_277 (O_277,N_19841,N_19941);
or UO_278 (O_278,N_19756,N_19865);
and UO_279 (O_279,N_19933,N_19809);
nor UO_280 (O_280,N_19872,N_19881);
xor UO_281 (O_281,N_19899,N_19884);
nor UO_282 (O_282,N_19752,N_19860);
xnor UO_283 (O_283,N_19962,N_19951);
or UO_284 (O_284,N_19795,N_19875);
or UO_285 (O_285,N_19807,N_19802);
and UO_286 (O_286,N_19796,N_19853);
nor UO_287 (O_287,N_19867,N_19961);
xnor UO_288 (O_288,N_19817,N_19895);
nand UO_289 (O_289,N_19962,N_19817);
xnor UO_290 (O_290,N_19822,N_19763);
nand UO_291 (O_291,N_19848,N_19972);
or UO_292 (O_292,N_19890,N_19808);
nor UO_293 (O_293,N_19960,N_19859);
and UO_294 (O_294,N_19870,N_19990);
and UO_295 (O_295,N_19897,N_19860);
xnor UO_296 (O_296,N_19774,N_19981);
xor UO_297 (O_297,N_19969,N_19916);
and UO_298 (O_298,N_19868,N_19812);
nor UO_299 (O_299,N_19970,N_19888);
nand UO_300 (O_300,N_19943,N_19876);
and UO_301 (O_301,N_19979,N_19797);
xor UO_302 (O_302,N_19990,N_19867);
nand UO_303 (O_303,N_19893,N_19783);
nor UO_304 (O_304,N_19821,N_19881);
nor UO_305 (O_305,N_19908,N_19970);
xor UO_306 (O_306,N_19810,N_19820);
and UO_307 (O_307,N_19931,N_19926);
xnor UO_308 (O_308,N_19986,N_19871);
xor UO_309 (O_309,N_19944,N_19769);
xor UO_310 (O_310,N_19934,N_19755);
and UO_311 (O_311,N_19908,N_19991);
and UO_312 (O_312,N_19765,N_19989);
or UO_313 (O_313,N_19763,N_19843);
xor UO_314 (O_314,N_19815,N_19820);
and UO_315 (O_315,N_19896,N_19956);
or UO_316 (O_316,N_19892,N_19904);
nand UO_317 (O_317,N_19926,N_19756);
or UO_318 (O_318,N_19970,N_19776);
or UO_319 (O_319,N_19889,N_19810);
xor UO_320 (O_320,N_19765,N_19781);
or UO_321 (O_321,N_19989,N_19859);
xnor UO_322 (O_322,N_19923,N_19915);
xor UO_323 (O_323,N_19934,N_19841);
xnor UO_324 (O_324,N_19837,N_19862);
or UO_325 (O_325,N_19980,N_19833);
and UO_326 (O_326,N_19778,N_19997);
nand UO_327 (O_327,N_19947,N_19752);
nor UO_328 (O_328,N_19822,N_19811);
or UO_329 (O_329,N_19982,N_19898);
or UO_330 (O_330,N_19864,N_19817);
and UO_331 (O_331,N_19959,N_19801);
or UO_332 (O_332,N_19845,N_19931);
or UO_333 (O_333,N_19862,N_19854);
or UO_334 (O_334,N_19932,N_19790);
nor UO_335 (O_335,N_19759,N_19967);
xnor UO_336 (O_336,N_19961,N_19906);
xnor UO_337 (O_337,N_19912,N_19998);
nand UO_338 (O_338,N_19763,N_19955);
nor UO_339 (O_339,N_19976,N_19936);
or UO_340 (O_340,N_19971,N_19754);
and UO_341 (O_341,N_19985,N_19864);
and UO_342 (O_342,N_19800,N_19781);
nand UO_343 (O_343,N_19764,N_19791);
xor UO_344 (O_344,N_19811,N_19908);
xor UO_345 (O_345,N_19983,N_19771);
xnor UO_346 (O_346,N_19776,N_19905);
nor UO_347 (O_347,N_19758,N_19965);
and UO_348 (O_348,N_19919,N_19893);
nor UO_349 (O_349,N_19956,N_19874);
or UO_350 (O_350,N_19871,N_19995);
and UO_351 (O_351,N_19878,N_19783);
nand UO_352 (O_352,N_19855,N_19946);
nand UO_353 (O_353,N_19976,N_19873);
xnor UO_354 (O_354,N_19936,N_19814);
xnor UO_355 (O_355,N_19877,N_19903);
or UO_356 (O_356,N_19760,N_19919);
and UO_357 (O_357,N_19830,N_19884);
xnor UO_358 (O_358,N_19757,N_19920);
nor UO_359 (O_359,N_19752,N_19842);
nand UO_360 (O_360,N_19987,N_19763);
nand UO_361 (O_361,N_19771,N_19819);
and UO_362 (O_362,N_19900,N_19946);
nand UO_363 (O_363,N_19970,N_19864);
nor UO_364 (O_364,N_19839,N_19850);
or UO_365 (O_365,N_19891,N_19838);
nor UO_366 (O_366,N_19933,N_19936);
and UO_367 (O_367,N_19755,N_19882);
or UO_368 (O_368,N_19773,N_19772);
and UO_369 (O_369,N_19827,N_19751);
or UO_370 (O_370,N_19778,N_19862);
nand UO_371 (O_371,N_19804,N_19999);
or UO_372 (O_372,N_19936,N_19849);
and UO_373 (O_373,N_19766,N_19848);
or UO_374 (O_374,N_19935,N_19964);
nand UO_375 (O_375,N_19900,N_19763);
nand UO_376 (O_376,N_19976,N_19909);
nor UO_377 (O_377,N_19823,N_19990);
or UO_378 (O_378,N_19777,N_19773);
nor UO_379 (O_379,N_19936,N_19840);
xor UO_380 (O_380,N_19771,N_19912);
nand UO_381 (O_381,N_19795,N_19977);
nor UO_382 (O_382,N_19759,N_19867);
xor UO_383 (O_383,N_19855,N_19798);
nor UO_384 (O_384,N_19913,N_19903);
and UO_385 (O_385,N_19803,N_19982);
xor UO_386 (O_386,N_19927,N_19832);
nand UO_387 (O_387,N_19895,N_19905);
nor UO_388 (O_388,N_19799,N_19794);
and UO_389 (O_389,N_19759,N_19786);
nand UO_390 (O_390,N_19983,N_19949);
nand UO_391 (O_391,N_19976,N_19785);
nor UO_392 (O_392,N_19924,N_19816);
nor UO_393 (O_393,N_19810,N_19992);
and UO_394 (O_394,N_19924,N_19943);
xnor UO_395 (O_395,N_19753,N_19912);
xnor UO_396 (O_396,N_19912,N_19796);
nand UO_397 (O_397,N_19868,N_19869);
and UO_398 (O_398,N_19974,N_19978);
xnor UO_399 (O_399,N_19895,N_19910);
and UO_400 (O_400,N_19955,N_19930);
or UO_401 (O_401,N_19994,N_19968);
nor UO_402 (O_402,N_19959,N_19819);
nand UO_403 (O_403,N_19796,N_19906);
or UO_404 (O_404,N_19842,N_19792);
nor UO_405 (O_405,N_19778,N_19787);
and UO_406 (O_406,N_19782,N_19948);
or UO_407 (O_407,N_19962,N_19756);
nor UO_408 (O_408,N_19849,N_19875);
nand UO_409 (O_409,N_19876,N_19788);
nor UO_410 (O_410,N_19797,N_19937);
xor UO_411 (O_411,N_19979,N_19878);
xor UO_412 (O_412,N_19858,N_19936);
nor UO_413 (O_413,N_19919,N_19843);
or UO_414 (O_414,N_19943,N_19910);
nand UO_415 (O_415,N_19764,N_19995);
xor UO_416 (O_416,N_19967,N_19965);
or UO_417 (O_417,N_19771,N_19837);
xnor UO_418 (O_418,N_19810,N_19783);
xor UO_419 (O_419,N_19935,N_19807);
nor UO_420 (O_420,N_19762,N_19851);
or UO_421 (O_421,N_19940,N_19935);
or UO_422 (O_422,N_19780,N_19757);
nor UO_423 (O_423,N_19853,N_19799);
xor UO_424 (O_424,N_19779,N_19958);
and UO_425 (O_425,N_19960,N_19892);
and UO_426 (O_426,N_19803,N_19866);
nor UO_427 (O_427,N_19967,N_19993);
nor UO_428 (O_428,N_19976,N_19890);
xnor UO_429 (O_429,N_19918,N_19983);
and UO_430 (O_430,N_19995,N_19925);
nand UO_431 (O_431,N_19930,N_19750);
xor UO_432 (O_432,N_19836,N_19978);
nor UO_433 (O_433,N_19834,N_19902);
or UO_434 (O_434,N_19781,N_19943);
or UO_435 (O_435,N_19751,N_19920);
nand UO_436 (O_436,N_19929,N_19879);
nor UO_437 (O_437,N_19974,N_19998);
nor UO_438 (O_438,N_19783,N_19953);
and UO_439 (O_439,N_19810,N_19811);
and UO_440 (O_440,N_19847,N_19911);
and UO_441 (O_441,N_19760,N_19880);
and UO_442 (O_442,N_19887,N_19927);
and UO_443 (O_443,N_19866,N_19822);
or UO_444 (O_444,N_19855,N_19884);
xnor UO_445 (O_445,N_19995,N_19785);
or UO_446 (O_446,N_19888,N_19752);
xor UO_447 (O_447,N_19756,N_19792);
xnor UO_448 (O_448,N_19942,N_19751);
or UO_449 (O_449,N_19984,N_19883);
xor UO_450 (O_450,N_19986,N_19972);
and UO_451 (O_451,N_19993,N_19923);
and UO_452 (O_452,N_19807,N_19951);
or UO_453 (O_453,N_19929,N_19760);
nor UO_454 (O_454,N_19971,N_19820);
and UO_455 (O_455,N_19762,N_19948);
xnor UO_456 (O_456,N_19958,N_19994);
or UO_457 (O_457,N_19791,N_19754);
and UO_458 (O_458,N_19828,N_19995);
or UO_459 (O_459,N_19894,N_19982);
nand UO_460 (O_460,N_19957,N_19816);
xor UO_461 (O_461,N_19795,N_19810);
and UO_462 (O_462,N_19980,N_19844);
or UO_463 (O_463,N_19830,N_19866);
and UO_464 (O_464,N_19987,N_19843);
or UO_465 (O_465,N_19938,N_19789);
xnor UO_466 (O_466,N_19903,N_19888);
or UO_467 (O_467,N_19875,N_19812);
or UO_468 (O_468,N_19958,N_19841);
nor UO_469 (O_469,N_19805,N_19780);
nor UO_470 (O_470,N_19872,N_19888);
nand UO_471 (O_471,N_19986,N_19802);
and UO_472 (O_472,N_19949,N_19937);
xnor UO_473 (O_473,N_19833,N_19977);
or UO_474 (O_474,N_19916,N_19795);
or UO_475 (O_475,N_19789,N_19820);
nor UO_476 (O_476,N_19824,N_19823);
xnor UO_477 (O_477,N_19968,N_19809);
nor UO_478 (O_478,N_19794,N_19976);
and UO_479 (O_479,N_19813,N_19931);
and UO_480 (O_480,N_19834,N_19950);
or UO_481 (O_481,N_19994,N_19855);
nand UO_482 (O_482,N_19833,N_19995);
xnor UO_483 (O_483,N_19878,N_19934);
nand UO_484 (O_484,N_19756,N_19790);
xor UO_485 (O_485,N_19769,N_19952);
nor UO_486 (O_486,N_19848,N_19845);
xor UO_487 (O_487,N_19848,N_19948);
nand UO_488 (O_488,N_19851,N_19767);
or UO_489 (O_489,N_19773,N_19800);
nor UO_490 (O_490,N_19996,N_19787);
and UO_491 (O_491,N_19760,N_19979);
nor UO_492 (O_492,N_19761,N_19791);
xor UO_493 (O_493,N_19772,N_19817);
nor UO_494 (O_494,N_19815,N_19862);
xnor UO_495 (O_495,N_19772,N_19802);
and UO_496 (O_496,N_19945,N_19958);
nand UO_497 (O_497,N_19806,N_19778);
and UO_498 (O_498,N_19900,N_19956);
nand UO_499 (O_499,N_19825,N_19770);
or UO_500 (O_500,N_19900,N_19820);
and UO_501 (O_501,N_19775,N_19944);
xor UO_502 (O_502,N_19766,N_19868);
nor UO_503 (O_503,N_19782,N_19807);
or UO_504 (O_504,N_19886,N_19817);
nor UO_505 (O_505,N_19762,N_19872);
xnor UO_506 (O_506,N_19892,N_19935);
xnor UO_507 (O_507,N_19754,N_19990);
xor UO_508 (O_508,N_19879,N_19957);
and UO_509 (O_509,N_19892,N_19879);
nand UO_510 (O_510,N_19781,N_19898);
nor UO_511 (O_511,N_19751,N_19900);
nor UO_512 (O_512,N_19973,N_19992);
nor UO_513 (O_513,N_19754,N_19838);
xnor UO_514 (O_514,N_19976,N_19778);
or UO_515 (O_515,N_19911,N_19820);
nor UO_516 (O_516,N_19790,N_19971);
and UO_517 (O_517,N_19804,N_19830);
or UO_518 (O_518,N_19994,N_19803);
and UO_519 (O_519,N_19993,N_19771);
nand UO_520 (O_520,N_19772,N_19964);
or UO_521 (O_521,N_19789,N_19763);
nor UO_522 (O_522,N_19822,N_19852);
and UO_523 (O_523,N_19766,N_19810);
or UO_524 (O_524,N_19804,N_19819);
xor UO_525 (O_525,N_19931,N_19791);
xnor UO_526 (O_526,N_19910,N_19865);
nand UO_527 (O_527,N_19877,N_19838);
nand UO_528 (O_528,N_19975,N_19794);
nand UO_529 (O_529,N_19897,N_19981);
xor UO_530 (O_530,N_19954,N_19990);
nand UO_531 (O_531,N_19939,N_19878);
nor UO_532 (O_532,N_19826,N_19768);
nand UO_533 (O_533,N_19990,N_19934);
and UO_534 (O_534,N_19971,N_19845);
nor UO_535 (O_535,N_19765,N_19950);
nand UO_536 (O_536,N_19752,N_19960);
nor UO_537 (O_537,N_19782,N_19857);
and UO_538 (O_538,N_19874,N_19759);
xnor UO_539 (O_539,N_19917,N_19836);
nand UO_540 (O_540,N_19842,N_19775);
nor UO_541 (O_541,N_19911,N_19995);
xnor UO_542 (O_542,N_19812,N_19853);
nand UO_543 (O_543,N_19756,N_19921);
nand UO_544 (O_544,N_19885,N_19797);
nand UO_545 (O_545,N_19821,N_19916);
nor UO_546 (O_546,N_19963,N_19802);
or UO_547 (O_547,N_19819,N_19908);
and UO_548 (O_548,N_19891,N_19909);
nor UO_549 (O_549,N_19767,N_19968);
xor UO_550 (O_550,N_19903,N_19879);
nor UO_551 (O_551,N_19995,N_19953);
nor UO_552 (O_552,N_19888,N_19928);
xnor UO_553 (O_553,N_19798,N_19807);
xor UO_554 (O_554,N_19981,N_19786);
and UO_555 (O_555,N_19982,N_19829);
or UO_556 (O_556,N_19982,N_19798);
xor UO_557 (O_557,N_19755,N_19896);
nor UO_558 (O_558,N_19776,N_19791);
nor UO_559 (O_559,N_19792,N_19921);
xor UO_560 (O_560,N_19949,N_19750);
and UO_561 (O_561,N_19952,N_19774);
xor UO_562 (O_562,N_19835,N_19860);
nor UO_563 (O_563,N_19883,N_19901);
xnor UO_564 (O_564,N_19829,N_19891);
and UO_565 (O_565,N_19853,N_19974);
and UO_566 (O_566,N_19942,N_19829);
nor UO_567 (O_567,N_19976,N_19808);
and UO_568 (O_568,N_19955,N_19801);
xnor UO_569 (O_569,N_19766,N_19918);
or UO_570 (O_570,N_19954,N_19754);
xor UO_571 (O_571,N_19789,N_19946);
nor UO_572 (O_572,N_19769,N_19995);
or UO_573 (O_573,N_19895,N_19863);
or UO_574 (O_574,N_19933,N_19900);
or UO_575 (O_575,N_19941,N_19902);
nand UO_576 (O_576,N_19873,N_19961);
or UO_577 (O_577,N_19868,N_19917);
and UO_578 (O_578,N_19969,N_19800);
nand UO_579 (O_579,N_19863,N_19899);
and UO_580 (O_580,N_19809,N_19772);
nand UO_581 (O_581,N_19954,N_19970);
nand UO_582 (O_582,N_19857,N_19823);
and UO_583 (O_583,N_19914,N_19751);
xnor UO_584 (O_584,N_19977,N_19776);
or UO_585 (O_585,N_19814,N_19890);
nand UO_586 (O_586,N_19800,N_19814);
or UO_587 (O_587,N_19961,N_19870);
and UO_588 (O_588,N_19967,N_19936);
xnor UO_589 (O_589,N_19857,N_19947);
or UO_590 (O_590,N_19865,N_19796);
xnor UO_591 (O_591,N_19779,N_19900);
and UO_592 (O_592,N_19858,N_19825);
and UO_593 (O_593,N_19869,N_19822);
and UO_594 (O_594,N_19786,N_19925);
nand UO_595 (O_595,N_19956,N_19939);
nand UO_596 (O_596,N_19894,N_19812);
or UO_597 (O_597,N_19924,N_19985);
or UO_598 (O_598,N_19867,N_19861);
xnor UO_599 (O_599,N_19985,N_19968);
nand UO_600 (O_600,N_19753,N_19846);
or UO_601 (O_601,N_19879,N_19972);
xor UO_602 (O_602,N_19965,N_19834);
and UO_603 (O_603,N_19876,N_19804);
or UO_604 (O_604,N_19795,N_19766);
and UO_605 (O_605,N_19997,N_19796);
nand UO_606 (O_606,N_19799,N_19810);
or UO_607 (O_607,N_19754,N_19957);
or UO_608 (O_608,N_19856,N_19977);
nor UO_609 (O_609,N_19994,N_19811);
nand UO_610 (O_610,N_19839,N_19859);
nand UO_611 (O_611,N_19826,N_19973);
or UO_612 (O_612,N_19961,N_19815);
nand UO_613 (O_613,N_19860,N_19968);
or UO_614 (O_614,N_19870,N_19796);
and UO_615 (O_615,N_19992,N_19780);
or UO_616 (O_616,N_19965,N_19862);
nand UO_617 (O_617,N_19865,N_19951);
and UO_618 (O_618,N_19922,N_19921);
nand UO_619 (O_619,N_19920,N_19778);
and UO_620 (O_620,N_19864,N_19944);
xor UO_621 (O_621,N_19997,N_19843);
nor UO_622 (O_622,N_19864,N_19829);
nor UO_623 (O_623,N_19891,N_19809);
nor UO_624 (O_624,N_19818,N_19781);
nand UO_625 (O_625,N_19921,N_19913);
nor UO_626 (O_626,N_19753,N_19796);
and UO_627 (O_627,N_19898,N_19885);
or UO_628 (O_628,N_19767,N_19994);
and UO_629 (O_629,N_19953,N_19761);
xor UO_630 (O_630,N_19801,N_19946);
xnor UO_631 (O_631,N_19952,N_19753);
nand UO_632 (O_632,N_19958,N_19991);
or UO_633 (O_633,N_19897,N_19834);
or UO_634 (O_634,N_19782,N_19893);
xor UO_635 (O_635,N_19910,N_19824);
and UO_636 (O_636,N_19857,N_19938);
and UO_637 (O_637,N_19934,N_19971);
xnor UO_638 (O_638,N_19942,N_19813);
or UO_639 (O_639,N_19999,N_19820);
or UO_640 (O_640,N_19762,N_19764);
nor UO_641 (O_641,N_19848,N_19782);
nand UO_642 (O_642,N_19945,N_19797);
nand UO_643 (O_643,N_19914,N_19870);
or UO_644 (O_644,N_19976,N_19914);
xnor UO_645 (O_645,N_19987,N_19955);
and UO_646 (O_646,N_19766,N_19835);
nor UO_647 (O_647,N_19865,N_19993);
and UO_648 (O_648,N_19839,N_19905);
nand UO_649 (O_649,N_19911,N_19926);
xor UO_650 (O_650,N_19848,N_19847);
xor UO_651 (O_651,N_19962,N_19902);
or UO_652 (O_652,N_19823,N_19864);
xor UO_653 (O_653,N_19802,N_19980);
xor UO_654 (O_654,N_19968,N_19836);
xor UO_655 (O_655,N_19926,N_19775);
nand UO_656 (O_656,N_19880,N_19858);
xor UO_657 (O_657,N_19789,N_19797);
and UO_658 (O_658,N_19973,N_19760);
xor UO_659 (O_659,N_19926,N_19840);
or UO_660 (O_660,N_19830,N_19848);
nor UO_661 (O_661,N_19952,N_19811);
nand UO_662 (O_662,N_19799,N_19809);
or UO_663 (O_663,N_19856,N_19869);
nor UO_664 (O_664,N_19934,N_19969);
xor UO_665 (O_665,N_19977,N_19839);
and UO_666 (O_666,N_19852,N_19828);
and UO_667 (O_667,N_19967,N_19937);
xnor UO_668 (O_668,N_19863,N_19956);
and UO_669 (O_669,N_19948,N_19913);
and UO_670 (O_670,N_19998,N_19962);
xnor UO_671 (O_671,N_19953,N_19848);
xor UO_672 (O_672,N_19908,N_19756);
nand UO_673 (O_673,N_19755,N_19996);
nand UO_674 (O_674,N_19911,N_19781);
or UO_675 (O_675,N_19945,N_19843);
or UO_676 (O_676,N_19842,N_19817);
nand UO_677 (O_677,N_19805,N_19884);
xnor UO_678 (O_678,N_19817,N_19921);
nor UO_679 (O_679,N_19765,N_19981);
and UO_680 (O_680,N_19867,N_19973);
xnor UO_681 (O_681,N_19802,N_19832);
xor UO_682 (O_682,N_19850,N_19763);
and UO_683 (O_683,N_19886,N_19970);
xnor UO_684 (O_684,N_19879,N_19975);
nor UO_685 (O_685,N_19762,N_19900);
and UO_686 (O_686,N_19893,N_19934);
nand UO_687 (O_687,N_19779,N_19797);
or UO_688 (O_688,N_19818,N_19815);
and UO_689 (O_689,N_19780,N_19894);
or UO_690 (O_690,N_19903,N_19883);
nor UO_691 (O_691,N_19876,N_19762);
nand UO_692 (O_692,N_19864,N_19880);
and UO_693 (O_693,N_19779,N_19784);
xnor UO_694 (O_694,N_19893,N_19905);
and UO_695 (O_695,N_19774,N_19860);
nand UO_696 (O_696,N_19806,N_19852);
and UO_697 (O_697,N_19992,N_19860);
nor UO_698 (O_698,N_19816,N_19869);
xnor UO_699 (O_699,N_19844,N_19881);
nor UO_700 (O_700,N_19840,N_19777);
or UO_701 (O_701,N_19929,N_19845);
and UO_702 (O_702,N_19793,N_19762);
nand UO_703 (O_703,N_19950,N_19975);
or UO_704 (O_704,N_19888,N_19892);
and UO_705 (O_705,N_19783,N_19979);
xor UO_706 (O_706,N_19991,N_19875);
xor UO_707 (O_707,N_19751,N_19960);
nand UO_708 (O_708,N_19781,N_19872);
nand UO_709 (O_709,N_19883,N_19983);
or UO_710 (O_710,N_19950,N_19888);
nand UO_711 (O_711,N_19977,N_19941);
and UO_712 (O_712,N_19914,N_19878);
nand UO_713 (O_713,N_19823,N_19930);
and UO_714 (O_714,N_19776,N_19848);
nor UO_715 (O_715,N_19902,N_19837);
nor UO_716 (O_716,N_19856,N_19805);
and UO_717 (O_717,N_19753,N_19949);
xnor UO_718 (O_718,N_19901,N_19965);
xor UO_719 (O_719,N_19842,N_19932);
nand UO_720 (O_720,N_19896,N_19894);
nor UO_721 (O_721,N_19922,N_19819);
nor UO_722 (O_722,N_19782,N_19810);
xor UO_723 (O_723,N_19794,N_19784);
nand UO_724 (O_724,N_19918,N_19871);
xnor UO_725 (O_725,N_19754,N_19834);
nand UO_726 (O_726,N_19978,N_19772);
and UO_727 (O_727,N_19767,N_19923);
xor UO_728 (O_728,N_19772,N_19932);
nor UO_729 (O_729,N_19752,N_19987);
or UO_730 (O_730,N_19900,N_19979);
nor UO_731 (O_731,N_19808,N_19780);
nand UO_732 (O_732,N_19819,N_19765);
nor UO_733 (O_733,N_19769,N_19963);
nand UO_734 (O_734,N_19921,N_19892);
or UO_735 (O_735,N_19876,N_19968);
and UO_736 (O_736,N_19991,N_19840);
xor UO_737 (O_737,N_19859,N_19855);
or UO_738 (O_738,N_19781,N_19819);
xor UO_739 (O_739,N_19788,N_19904);
and UO_740 (O_740,N_19798,N_19835);
nor UO_741 (O_741,N_19934,N_19840);
xor UO_742 (O_742,N_19905,N_19891);
or UO_743 (O_743,N_19771,N_19770);
nand UO_744 (O_744,N_19802,N_19997);
xor UO_745 (O_745,N_19813,N_19764);
nor UO_746 (O_746,N_19969,N_19750);
xor UO_747 (O_747,N_19922,N_19917);
nand UO_748 (O_748,N_19983,N_19862);
nand UO_749 (O_749,N_19945,N_19750);
xor UO_750 (O_750,N_19885,N_19864);
and UO_751 (O_751,N_19830,N_19809);
and UO_752 (O_752,N_19788,N_19770);
and UO_753 (O_753,N_19884,N_19769);
nand UO_754 (O_754,N_19897,N_19950);
nor UO_755 (O_755,N_19862,N_19844);
xnor UO_756 (O_756,N_19959,N_19986);
nor UO_757 (O_757,N_19845,N_19780);
and UO_758 (O_758,N_19770,N_19962);
or UO_759 (O_759,N_19954,N_19867);
or UO_760 (O_760,N_19866,N_19858);
and UO_761 (O_761,N_19964,N_19931);
xor UO_762 (O_762,N_19845,N_19818);
or UO_763 (O_763,N_19838,N_19892);
xor UO_764 (O_764,N_19871,N_19982);
and UO_765 (O_765,N_19885,N_19927);
or UO_766 (O_766,N_19939,N_19776);
and UO_767 (O_767,N_19865,N_19992);
xnor UO_768 (O_768,N_19913,N_19897);
nand UO_769 (O_769,N_19815,N_19883);
and UO_770 (O_770,N_19842,N_19927);
xnor UO_771 (O_771,N_19890,N_19765);
and UO_772 (O_772,N_19894,N_19752);
and UO_773 (O_773,N_19924,N_19990);
nor UO_774 (O_774,N_19821,N_19921);
and UO_775 (O_775,N_19992,N_19784);
xor UO_776 (O_776,N_19929,N_19973);
xor UO_777 (O_777,N_19868,N_19855);
xnor UO_778 (O_778,N_19811,N_19979);
and UO_779 (O_779,N_19804,N_19980);
and UO_780 (O_780,N_19781,N_19878);
xnor UO_781 (O_781,N_19772,N_19784);
and UO_782 (O_782,N_19763,N_19925);
or UO_783 (O_783,N_19903,N_19914);
xor UO_784 (O_784,N_19971,N_19939);
or UO_785 (O_785,N_19778,N_19847);
and UO_786 (O_786,N_19832,N_19931);
xor UO_787 (O_787,N_19916,N_19864);
xor UO_788 (O_788,N_19772,N_19750);
or UO_789 (O_789,N_19918,N_19862);
nand UO_790 (O_790,N_19960,N_19755);
or UO_791 (O_791,N_19838,N_19833);
nor UO_792 (O_792,N_19839,N_19894);
xor UO_793 (O_793,N_19786,N_19960);
and UO_794 (O_794,N_19861,N_19757);
xnor UO_795 (O_795,N_19976,N_19979);
xor UO_796 (O_796,N_19847,N_19795);
xor UO_797 (O_797,N_19878,N_19992);
xnor UO_798 (O_798,N_19753,N_19859);
nor UO_799 (O_799,N_19976,N_19986);
and UO_800 (O_800,N_19917,N_19950);
or UO_801 (O_801,N_19783,N_19824);
xnor UO_802 (O_802,N_19757,N_19946);
nor UO_803 (O_803,N_19899,N_19880);
or UO_804 (O_804,N_19819,N_19855);
nand UO_805 (O_805,N_19775,N_19933);
xnor UO_806 (O_806,N_19977,N_19980);
xnor UO_807 (O_807,N_19884,N_19881);
and UO_808 (O_808,N_19912,N_19944);
xnor UO_809 (O_809,N_19983,N_19969);
and UO_810 (O_810,N_19929,N_19846);
and UO_811 (O_811,N_19981,N_19910);
or UO_812 (O_812,N_19987,N_19951);
and UO_813 (O_813,N_19865,N_19897);
nand UO_814 (O_814,N_19878,N_19928);
or UO_815 (O_815,N_19758,N_19858);
and UO_816 (O_816,N_19885,N_19994);
nor UO_817 (O_817,N_19848,N_19833);
nand UO_818 (O_818,N_19773,N_19971);
xnor UO_819 (O_819,N_19909,N_19946);
nand UO_820 (O_820,N_19770,N_19863);
or UO_821 (O_821,N_19771,N_19800);
or UO_822 (O_822,N_19990,N_19865);
or UO_823 (O_823,N_19909,N_19760);
nor UO_824 (O_824,N_19785,N_19800);
nand UO_825 (O_825,N_19957,N_19847);
nand UO_826 (O_826,N_19890,N_19948);
nor UO_827 (O_827,N_19941,N_19942);
and UO_828 (O_828,N_19948,N_19917);
or UO_829 (O_829,N_19917,N_19938);
xor UO_830 (O_830,N_19927,N_19815);
xnor UO_831 (O_831,N_19781,N_19958);
and UO_832 (O_832,N_19984,N_19997);
or UO_833 (O_833,N_19848,N_19913);
nor UO_834 (O_834,N_19999,N_19845);
nand UO_835 (O_835,N_19778,N_19914);
or UO_836 (O_836,N_19923,N_19774);
and UO_837 (O_837,N_19830,N_19900);
nor UO_838 (O_838,N_19763,N_19991);
and UO_839 (O_839,N_19872,N_19750);
nand UO_840 (O_840,N_19914,N_19985);
nand UO_841 (O_841,N_19825,N_19981);
xnor UO_842 (O_842,N_19796,N_19826);
or UO_843 (O_843,N_19964,N_19796);
nor UO_844 (O_844,N_19906,N_19884);
xor UO_845 (O_845,N_19916,N_19873);
nand UO_846 (O_846,N_19956,N_19976);
nor UO_847 (O_847,N_19760,N_19886);
nand UO_848 (O_848,N_19815,N_19834);
nand UO_849 (O_849,N_19958,N_19961);
and UO_850 (O_850,N_19818,N_19779);
nand UO_851 (O_851,N_19868,N_19814);
nor UO_852 (O_852,N_19887,N_19840);
xnor UO_853 (O_853,N_19920,N_19836);
xnor UO_854 (O_854,N_19894,N_19825);
nor UO_855 (O_855,N_19895,N_19951);
xnor UO_856 (O_856,N_19839,N_19987);
or UO_857 (O_857,N_19885,N_19988);
nor UO_858 (O_858,N_19905,N_19955);
nor UO_859 (O_859,N_19802,N_19783);
nand UO_860 (O_860,N_19989,N_19920);
nor UO_861 (O_861,N_19931,N_19826);
nand UO_862 (O_862,N_19787,N_19754);
nand UO_863 (O_863,N_19808,N_19859);
xnor UO_864 (O_864,N_19844,N_19903);
or UO_865 (O_865,N_19968,N_19889);
nor UO_866 (O_866,N_19879,N_19992);
or UO_867 (O_867,N_19938,N_19827);
xor UO_868 (O_868,N_19794,N_19926);
or UO_869 (O_869,N_19952,N_19808);
nand UO_870 (O_870,N_19869,N_19788);
xor UO_871 (O_871,N_19956,N_19763);
and UO_872 (O_872,N_19759,N_19845);
or UO_873 (O_873,N_19939,N_19839);
xnor UO_874 (O_874,N_19943,N_19884);
nand UO_875 (O_875,N_19858,N_19784);
nand UO_876 (O_876,N_19889,N_19948);
nand UO_877 (O_877,N_19839,N_19990);
nor UO_878 (O_878,N_19888,N_19852);
and UO_879 (O_879,N_19940,N_19761);
nand UO_880 (O_880,N_19937,N_19939);
nor UO_881 (O_881,N_19758,N_19826);
and UO_882 (O_882,N_19836,N_19861);
and UO_883 (O_883,N_19946,N_19780);
xnor UO_884 (O_884,N_19837,N_19829);
nand UO_885 (O_885,N_19897,N_19962);
and UO_886 (O_886,N_19989,N_19996);
nor UO_887 (O_887,N_19948,N_19805);
nand UO_888 (O_888,N_19780,N_19846);
and UO_889 (O_889,N_19798,N_19867);
xor UO_890 (O_890,N_19922,N_19798);
xor UO_891 (O_891,N_19850,N_19809);
xnor UO_892 (O_892,N_19813,N_19761);
or UO_893 (O_893,N_19818,N_19876);
and UO_894 (O_894,N_19819,N_19829);
and UO_895 (O_895,N_19780,N_19755);
nand UO_896 (O_896,N_19868,N_19808);
nand UO_897 (O_897,N_19820,N_19772);
and UO_898 (O_898,N_19989,N_19905);
and UO_899 (O_899,N_19998,N_19818);
xnor UO_900 (O_900,N_19950,N_19846);
nand UO_901 (O_901,N_19967,N_19758);
nor UO_902 (O_902,N_19849,N_19767);
nand UO_903 (O_903,N_19874,N_19961);
nand UO_904 (O_904,N_19955,N_19843);
nor UO_905 (O_905,N_19886,N_19977);
xnor UO_906 (O_906,N_19804,N_19778);
nand UO_907 (O_907,N_19904,N_19833);
or UO_908 (O_908,N_19885,N_19818);
nor UO_909 (O_909,N_19972,N_19792);
and UO_910 (O_910,N_19831,N_19912);
nor UO_911 (O_911,N_19974,N_19934);
nor UO_912 (O_912,N_19912,N_19752);
xor UO_913 (O_913,N_19788,N_19993);
and UO_914 (O_914,N_19995,N_19771);
and UO_915 (O_915,N_19985,N_19893);
nor UO_916 (O_916,N_19784,N_19819);
nor UO_917 (O_917,N_19757,N_19773);
or UO_918 (O_918,N_19957,N_19858);
or UO_919 (O_919,N_19977,N_19931);
nor UO_920 (O_920,N_19858,N_19976);
nand UO_921 (O_921,N_19767,N_19861);
xnor UO_922 (O_922,N_19914,N_19814);
and UO_923 (O_923,N_19818,N_19960);
and UO_924 (O_924,N_19944,N_19940);
or UO_925 (O_925,N_19959,N_19869);
nand UO_926 (O_926,N_19875,N_19824);
nor UO_927 (O_927,N_19751,N_19757);
nor UO_928 (O_928,N_19898,N_19949);
or UO_929 (O_929,N_19958,N_19813);
xor UO_930 (O_930,N_19903,N_19906);
nor UO_931 (O_931,N_19844,N_19849);
xnor UO_932 (O_932,N_19984,N_19951);
nor UO_933 (O_933,N_19780,N_19856);
nand UO_934 (O_934,N_19825,N_19929);
and UO_935 (O_935,N_19802,N_19795);
and UO_936 (O_936,N_19973,N_19934);
nor UO_937 (O_937,N_19825,N_19980);
and UO_938 (O_938,N_19812,N_19928);
xnor UO_939 (O_939,N_19964,N_19926);
nand UO_940 (O_940,N_19990,N_19999);
nand UO_941 (O_941,N_19811,N_19761);
or UO_942 (O_942,N_19940,N_19836);
nor UO_943 (O_943,N_19884,N_19940);
xor UO_944 (O_944,N_19885,N_19821);
xnor UO_945 (O_945,N_19763,N_19924);
nand UO_946 (O_946,N_19919,N_19930);
nor UO_947 (O_947,N_19944,N_19792);
nand UO_948 (O_948,N_19978,N_19787);
nand UO_949 (O_949,N_19964,N_19877);
and UO_950 (O_950,N_19872,N_19899);
or UO_951 (O_951,N_19864,N_19786);
xnor UO_952 (O_952,N_19752,N_19964);
nor UO_953 (O_953,N_19945,N_19923);
nor UO_954 (O_954,N_19980,N_19965);
nor UO_955 (O_955,N_19987,N_19969);
or UO_956 (O_956,N_19968,N_19982);
and UO_957 (O_957,N_19961,N_19761);
nand UO_958 (O_958,N_19765,N_19996);
xnor UO_959 (O_959,N_19887,N_19809);
nor UO_960 (O_960,N_19892,N_19787);
and UO_961 (O_961,N_19882,N_19922);
xor UO_962 (O_962,N_19790,N_19913);
and UO_963 (O_963,N_19865,N_19944);
xnor UO_964 (O_964,N_19910,N_19828);
or UO_965 (O_965,N_19922,N_19883);
nor UO_966 (O_966,N_19887,N_19807);
nor UO_967 (O_967,N_19961,N_19752);
nand UO_968 (O_968,N_19827,N_19937);
and UO_969 (O_969,N_19955,N_19830);
and UO_970 (O_970,N_19764,N_19796);
and UO_971 (O_971,N_19869,N_19794);
or UO_972 (O_972,N_19993,N_19872);
xor UO_973 (O_973,N_19924,N_19911);
xnor UO_974 (O_974,N_19834,N_19766);
xor UO_975 (O_975,N_19840,N_19828);
or UO_976 (O_976,N_19978,N_19810);
nor UO_977 (O_977,N_19803,N_19805);
nor UO_978 (O_978,N_19834,N_19842);
nor UO_979 (O_979,N_19961,N_19853);
nor UO_980 (O_980,N_19916,N_19860);
and UO_981 (O_981,N_19938,N_19931);
xor UO_982 (O_982,N_19852,N_19833);
nand UO_983 (O_983,N_19948,N_19887);
or UO_984 (O_984,N_19985,N_19791);
xnor UO_985 (O_985,N_19806,N_19782);
xor UO_986 (O_986,N_19838,N_19934);
and UO_987 (O_987,N_19887,N_19890);
or UO_988 (O_988,N_19916,N_19909);
and UO_989 (O_989,N_19811,N_19934);
xor UO_990 (O_990,N_19837,N_19818);
nor UO_991 (O_991,N_19823,N_19891);
or UO_992 (O_992,N_19947,N_19779);
or UO_993 (O_993,N_19755,N_19893);
nand UO_994 (O_994,N_19859,N_19996);
xnor UO_995 (O_995,N_19941,N_19937);
xnor UO_996 (O_996,N_19811,N_19893);
and UO_997 (O_997,N_19795,N_19784);
nand UO_998 (O_998,N_19776,N_19797);
nor UO_999 (O_999,N_19798,N_19805);
xor UO_1000 (O_1000,N_19803,N_19942);
nand UO_1001 (O_1001,N_19926,N_19953);
nand UO_1002 (O_1002,N_19852,N_19766);
nor UO_1003 (O_1003,N_19762,N_19996);
xnor UO_1004 (O_1004,N_19833,N_19992);
or UO_1005 (O_1005,N_19870,N_19772);
xor UO_1006 (O_1006,N_19780,N_19904);
or UO_1007 (O_1007,N_19751,N_19980);
nor UO_1008 (O_1008,N_19806,N_19797);
and UO_1009 (O_1009,N_19861,N_19956);
xnor UO_1010 (O_1010,N_19911,N_19877);
nor UO_1011 (O_1011,N_19996,N_19843);
nand UO_1012 (O_1012,N_19989,N_19929);
xor UO_1013 (O_1013,N_19816,N_19980);
xnor UO_1014 (O_1014,N_19834,N_19918);
xor UO_1015 (O_1015,N_19940,N_19947);
nand UO_1016 (O_1016,N_19788,N_19766);
or UO_1017 (O_1017,N_19964,N_19813);
nor UO_1018 (O_1018,N_19774,N_19967);
nand UO_1019 (O_1019,N_19901,N_19983);
nand UO_1020 (O_1020,N_19992,N_19866);
nor UO_1021 (O_1021,N_19890,N_19902);
xor UO_1022 (O_1022,N_19882,N_19916);
nor UO_1023 (O_1023,N_19918,N_19827);
and UO_1024 (O_1024,N_19929,N_19854);
nor UO_1025 (O_1025,N_19969,N_19933);
nand UO_1026 (O_1026,N_19912,N_19893);
xor UO_1027 (O_1027,N_19903,N_19796);
or UO_1028 (O_1028,N_19876,N_19753);
nand UO_1029 (O_1029,N_19819,N_19752);
and UO_1030 (O_1030,N_19878,N_19940);
and UO_1031 (O_1031,N_19896,N_19782);
or UO_1032 (O_1032,N_19815,N_19775);
xnor UO_1033 (O_1033,N_19973,N_19962);
nor UO_1034 (O_1034,N_19883,N_19917);
xor UO_1035 (O_1035,N_19830,N_19974);
nor UO_1036 (O_1036,N_19992,N_19956);
and UO_1037 (O_1037,N_19793,N_19849);
or UO_1038 (O_1038,N_19755,N_19926);
or UO_1039 (O_1039,N_19903,N_19832);
nor UO_1040 (O_1040,N_19999,N_19762);
xnor UO_1041 (O_1041,N_19899,N_19861);
nand UO_1042 (O_1042,N_19974,N_19884);
and UO_1043 (O_1043,N_19764,N_19835);
and UO_1044 (O_1044,N_19928,N_19851);
and UO_1045 (O_1045,N_19799,N_19752);
xor UO_1046 (O_1046,N_19788,N_19862);
or UO_1047 (O_1047,N_19850,N_19787);
nor UO_1048 (O_1048,N_19942,N_19793);
nand UO_1049 (O_1049,N_19807,N_19838);
or UO_1050 (O_1050,N_19826,N_19799);
nand UO_1051 (O_1051,N_19807,N_19931);
xor UO_1052 (O_1052,N_19927,N_19838);
nor UO_1053 (O_1053,N_19765,N_19986);
nor UO_1054 (O_1054,N_19934,N_19945);
nand UO_1055 (O_1055,N_19859,N_19983);
nand UO_1056 (O_1056,N_19949,N_19833);
xor UO_1057 (O_1057,N_19945,N_19769);
and UO_1058 (O_1058,N_19780,N_19978);
nor UO_1059 (O_1059,N_19835,N_19875);
nor UO_1060 (O_1060,N_19982,N_19797);
nor UO_1061 (O_1061,N_19986,N_19916);
and UO_1062 (O_1062,N_19801,N_19832);
or UO_1063 (O_1063,N_19973,N_19945);
nor UO_1064 (O_1064,N_19851,N_19919);
nor UO_1065 (O_1065,N_19822,N_19868);
and UO_1066 (O_1066,N_19759,N_19810);
nand UO_1067 (O_1067,N_19882,N_19968);
xnor UO_1068 (O_1068,N_19829,N_19908);
and UO_1069 (O_1069,N_19923,N_19991);
nor UO_1070 (O_1070,N_19835,N_19780);
nor UO_1071 (O_1071,N_19955,N_19947);
or UO_1072 (O_1072,N_19870,N_19776);
and UO_1073 (O_1073,N_19888,N_19926);
nand UO_1074 (O_1074,N_19808,N_19806);
xor UO_1075 (O_1075,N_19878,N_19937);
xor UO_1076 (O_1076,N_19982,N_19990);
xnor UO_1077 (O_1077,N_19792,N_19834);
nor UO_1078 (O_1078,N_19977,N_19831);
xor UO_1079 (O_1079,N_19757,N_19779);
nor UO_1080 (O_1080,N_19926,N_19793);
and UO_1081 (O_1081,N_19847,N_19825);
nor UO_1082 (O_1082,N_19768,N_19927);
or UO_1083 (O_1083,N_19937,N_19875);
or UO_1084 (O_1084,N_19837,N_19821);
xor UO_1085 (O_1085,N_19852,N_19943);
or UO_1086 (O_1086,N_19918,N_19879);
nor UO_1087 (O_1087,N_19755,N_19812);
and UO_1088 (O_1088,N_19917,N_19990);
xnor UO_1089 (O_1089,N_19963,N_19905);
or UO_1090 (O_1090,N_19833,N_19882);
or UO_1091 (O_1091,N_19836,N_19970);
nand UO_1092 (O_1092,N_19845,N_19921);
or UO_1093 (O_1093,N_19838,N_19788);
or UO_1094 (O_1094,N_19935,N_19898);
nand UO_1095 (O_1095,N_19834,N_19783);
nor UO_1096 (O_1096,N_19750,N_19811);
nor UO_1097 (O_1097,N_19858,N_19889);
nor UO_1098 (O_1098,N_19942,N_19774);
and UO_1099 (O_1099,N_19909,N_19842);
nor UO_1100 (O_1100,N_19812,N_19932);
and UO_1101 (O_1101,N_19820,N_19972);
and UO_1102 (O_1102,N_19929,N_19931);
xnor UO_1103 (O_1103,N_19944,N_19960);
or UO_1104 (O_1104,N_19956,N_19797);
nand UO_1105 (O_1105,N_19876,N_19838);
nor UO_1106 (O_1106,N_19933,N_19971);
nor UO_1107 (O_1107,N_19992,N_19946);
and UO_1108 (O_1108,N_19952,N_19915);
nand UO_1109 (O_1109,N_19852,N_19941);
and UO_1110 (O_1110,N_19909,N_19837);
nor UO_1111 (O_1111,N_19961,N_19833);
nand UO_1112 (O_1112,N_19867,N_19982);
and UO_1113 (O_1113,N_19800,N_19884);
nand UO_1114 (O_1114,N_19861,N_19825);
nand UO_1115 (O_1115,N_19937,N_19978);
and UO_1116 (O_1116,N_19914,N_19949);
xnor UO_1117 (O_1117,N_19983,N_19762);
xnor UO_1118 (O_1118,N_19891,N_19866);
nand UO_1119 (O_1119,N_19996,N_19887);
or UO_1120 (O_1120,N_19852,N_19909);
or UO_1121 (O_1121,N_19987,N_19800);
and UO_1122 (O_1122,N_19817,N_19835);
nor UO_1123 (O_1123,N_19870,N_19941);
nand UO_1124 (O_1124,N_19841,N_19947);
and UO_1125 (O_1125,N_19987,N_19826);
or UO_1126 (O_1126,N_19993,N_19780);
nand UO_1127 (O_1127,N_19833,N_19829);
nor UO_1128 (O_1128,N_19780,N_19893);
or UO_1129 (O_1129,N_19968,N_19918);
and UO_1130 (O_1130,N_19956,N_19759);
and UO_1131 (O_1131,N_19882,N_19963);
or UO_1132 (O_1132,N_19887,N_19946);
nor UO_1133 (O_1133,N_19759,N_19847);
nand UO_1134 (O_1134,N_19782,N_19803);
nor UO_1135 (O_1135,N_19801,N_19841);
nand UO_1136 (O_1136,N_19873,N_19951);
nor UO_1137 (O_1137,N_19776,N_19847);
xnor UO_1138 (O_1138,N_19834,N_19991);
nor UO_1139 (O_1139,N_19899,N_19855);
and UO_1140 (O_1140,N_19963,N_19792);
xor UO_1141 (O_1141,N_19776,N_19803);
and UO_1142 (O_1142,N_19852,N_19890);
nor UO_1143 (O_1143,N_19922,N_19859);
nor UO_1144 (O_1144,N_19830,N_19854);
and UO_1145 (O_1145,N_19826,N_19765);
xnor UO_1146 (O_1146,N_19943,N_19772);
and UO_1147 (O_1147,N_19997,N_19974);
xnor UO_1148 (O_1148,N_19844,N_19887);
or UO_1149 (O_1149,N_19758,N_19827);
nor UO_1150 (O_1150,N_19977,N_19794);
and UO_1151 (O_1151,N_19867,N_19951);
or UO_1152 (O_1152,N_19920,N_19894);
nand UO_1153 (O_1153,N_19940,N_19828);
nor UO_1154 (O_1154,N_19758,N_19990);
nand UO_1155 (O_1155,N_19916,N_19771);
and UO_1156 (O_1156,N_19955,N_19923);
xor UO_1157 (O_1157,N_19821,N_19859);
nand UO_1158 (O_1158,N_19996,N_19999);
nand UO_1159 (O_1159,N_19978,N_19851);
xor UO_1160 (O_1160,N_19923,N_19962);
nand UO_1161 (O_1161,N_19792,N_19930);
nor UO_1162 (O_1162,N_19972,N_19804);
xor UO_1163 (O_1163,N_19898,N_19994);
nand UO_1164 (O_1164,N_19865,N_19873);
nand UO_1165 (O_1165,N_19834,N_19829);
nand UO_1166 (O_1166,N_19855,N_19989);
or UO_1167 (O_1167,N_19993,N_19947);
and UO_1168 (O_1168,N_19999,N_19800);
nand UO_1169 (O_1169,N_19965,N_19993);
nor UO_1170 (O_1170,N_19869,N_19921);
and UO_1171 (O_1171,N_19786,N_19913);
or UO_1172 (O_1172,N_19828,N_19939);
and UO_1173 (O_1173,N_19775,N_19810);
xor UO_1174 (O_1174,N_19787,N_19887);
xor UO_1175 (O_1175,N_19963,N_19956);
xnor UO_1176 (O_1176,N_19750,N_19884);
and UO_1177 (O_1177,N_19755,N_19974);
or UO_1178 (O_1178,N_19935,N_19934);
and UO_1179 (O_1179,N_19987,N_19860);
xor UO_1180 (O_1180,N_19909,N_19957);
and UO_1181 (O_1181,N_19874,N_19900);
nor UO_1182 (O_1182,N_19887,N_19839);
and UO_1183 (O_1183,N_19995,N_19787);
and UO_1184 (O_1184,N_19854,N_19937);
nand UO_1185 (O_1185,N_19891,N_19773);
nor UO_1186 (O_1186,N_19785,N_19769);
xor UO_1187 (O_1187,N_19860,N_19972);
nor UO_1188 (O_1188,N_19880,N_19926);
xor UO_1189 (O_1189,N_19899,N_19859);
nor UO_1190 (O_1190,N_19783,N_19762);
nor UO_1191 (O_1191,N_19781,N_19919);
xnor UO_1192 (O_1192,N_19999,N_19895);
and UO_1193 (O_1193,N_19817,N_19846);
xnor UO_1194 (O_1194,N_19939,N_19829);
xnor UO_1195 (O_1195,N_19788,N_19960);
or UO_1196 (O_1196,N_19975,N_19786);
or UO_1197 (O_1197,N_19860,N_19984);
or UO_1198 (O_1198,N_19896,N_19757);
xnor UO_1199 (O_1199,N_19793,N_19799);
nand UO_1200 (O_1200,N_19968,N_19804);
or UO_1201 (O_1201,N_19821,N_19774);
nand UO_1202 (O_1202,N_19966,N_19869);
xnor UO_1203 (O_1203,N_19823,N_19772);
xor UO_1204 (O_1204,N_19944,N_19863);
xnor UO_1205 (O_1205,N_19887,N_19903);
nand UO_1206 (O_1206,N_19803,N_19875);
or UO_1207 (O_1207,N_19810,N_19961);
nand UO_1208 (O_1208,N_19762,N_19801);
or UO_1209 (O_1209,N_19854,N_19807);
xnor UO_1210 (O_1210,N_19913,N_19766);
xnor UO_1211 (O_1211,N_19818,N_19986);
nand UO_1212 (O_1212,N_19854,N_19932);
nand UO_1213 (O_1213,N_19813,N_19791);
and UO_1214 (O_1214,N_19836,N_19900);
and UO_1215 (O_1215,N_19928,N_19825);
and UO_1216 (O_1216,N_19785,N_19763);
or UO_1217 (O_1217,N_19930,N_19752);
nor UO_1218 (O_1218,N_19955,N_19917);
xnor UO_1219 (O_1219,N_19945,N_19858);
xor UO_1220 (O_1220,N_19911,N_19818);
nor UO_1221 (O_1221,N_19861,N_19754);
nand UO_1222 (O_1222,N_19955,N_19814);
nor UO_1223 (O_1223,N_19833,N_19784);
xor UO_1224 (O_1224,N_19922,N_19802);
nand UO_1225 (O_1225,N_19832,N_19756);
xnor UO_1226 (O_1226,N_19800,N_19806);
nor UO_1227 (O_1227,N_19859,N_19976);
and UO_1228 (O_1228,N_19936,N_19866);
nand UO_1229 (O_1229,N_19960,N_19988);
nor UO_1230 (O_1230,N_19792,N_19975);
or UO_1231 (O_1231,N_19931,N_19902);
nand UO_1232 (O_1232,N_19946,N_19899);
or UO_1233 (O_1233,N_19750,N_19916);
xor UO_1234 (O_1234,N_19862,N_19806);
or UO_1235 (O_1235,N_19963,N_19883);
and UO_1236 (O_1236,N_19909,N_19855);
or UO_1237 (O_1237,N_19753,N_19783);
nor UO_1238 (O_1238,N_19836,N_19857);
xnor UO_1239 (O_1239,N_19777,N_19910);
and UO_1240 (O_1240,N_19903,N_19994);
nor UO_1241 (O_1241,N_19922,N_19866);
nor UO_1242 (O_1242,N_19858,N_19927);
xnor UO_1243 (O_1243,N_19897,N_19900);
nand UO_1244 (O_1244,N_19965,N_19949);
xnor UO_1245 (O_1245,N_19975,N_19848);
nor UO_1246 (O_1246,N_19763,N_19775);
nor UO_1247 (O_1247,N_19853,N_19788);
or UO_1248 (O_1248,N_19937,N_19823);
nor UO_1249 (O_1249,N_19775,N_19903);
xnor UO_1250 (O_1250,N_19786,N_19978);
xnor UO_1251 (O_1251,N_19905,N_19879);
and UO_1252 (O_1252,N_19832,N_19912);
and UO_1253 (O_1253,N_19802,N_19752);
and UO_1254 (O_1254,N_19876,N_19987);
and UO_1255 (O_1255,N_19995,N_19922);
nand UO_1256 (O_1256,N_19792,N_19754);
nor UO_1257 (O_1257,N_19827,N_19940);
or UO_1258 (O_1258,N_19885,N_19841);
xnor UO_1259 (O_1259,N_19797,N_19823);
xnor UO_1260 (O_1260,N_19899,N_19791);
nor UO_1261 (O_1261,N_19982,N_19801);
or UO_1262 (O_1262,N_19970,N_19858);
nor UO_1263 (O_1263,N_19776,N_19832);
nor UO_1264 (O_1264,N_19927,N_19912);
or UO_1265 (O_1265,N_19962,N_19840);
xnor UO_1266 (O_1266,N_19997,N_19962);
xor UO_1267 (O_1267,N_19952,N_19794);
or UO_1268 (O_1268,N_19968,N_19770);
or UO_1269 (O_1269,N_19766,N_19758);
nor UO_1270 (O_1270,N_19885,N_19773);
nor UO_1271 (O_1271,N_19768,N_19894);
nor UO_1272 (O_1272,N_19835,N_19797);
nand UO_1273 (O_1273,N_19808,N_19896);
or UO_1274 (O_1274,N_19969,N_19878);
xnor UO_1275 (O_1275,N_19903,N_19964);
nand UO_1276 (O_1276,N_19937,N_19948);
nor UO_1277 (O_1277,N_19817,N_19881);
or UO_1278 (O_1278,N_19797,N_19943);
and UO_1279 (O_1279,N_19999,N_19991);
xnor UO_1280 (O_1280,N_19763,N_19918);
xnor UO_1281 (O_1281,N_19939,N_19916);
xor UO_1282 (O_1282,N_19953,N_19922);
nand UO_1283 (O_1283,N_19836,N_19933);
nand UO_1284 (O_1284,N_19985,N_19781);
or UO_1285 (O_1285,N_19853,N_19927);
nand UO_1286 (O_1286,N_19768,N_19842);
xor UO_1287 (O_1287,N_19877,N_19872);
or UO_1288 (O_1288,N_19791,N_19904);
nor UO_1289 (O_1289,N_19782,N_19963);
nor UO_1290 (O_1290,N_19765,N_19843);
and UO_1291 (O_1291,N_19950,N_19763);
and UO_1292 (O_1292,N_19874,N_19814);
or UO_1293 (O_1293,N_19976,N_19815);
nand UO_1294 (O_1294,N_19839,N_19952);
nor UO_1295 (O_1295,N_19763,N_19957);
nand UO_1296 (O_1296,N_19980,N_19798);
xnor UO_1297 (O_1297,N_19981,N_19756);
nand UO_1298 (O_1298,N_19898,N_19871);
nor UO_1299 (O_1299,N_19961,N_19980);
and UO_1300 (O_1300,N_19862,N_19997);
xnor UO_1301 (O_1301,N_19785,N_19986);
xnor UO_1302 (O_1302,N_19760,N_19938);
and UO_1303 (O_1303,N_19923,N_19793);
nand UO_1304 (O_1304,N_19874,N_19987);
or UO_1305 (O_1305,N_19894,N_19927);
nand UO_1306 (O_1306,N_19974,N_19815);
or UO_1307 (O_1307,N_19815,N_19808);
nand UO_1308 (O_1308,N_19959,N_19771);
nor UO_1309 (O_1309,N_19815,N_19879);
xnor UO_1310 (O_1310,N_19780,N_19951);
or UO_1311 (O_1311,N_19856,N_19953);
nand UO_1312 (O_1312,N_19792,N_19771);
and UO_1313 (O_1313,N_19829,N_19988);
and UO_1314 (O_1314,N_19831,N_19871);
or UO_1315 (O_1315,N_19899,N_19847);
or UO_1316 (O_1316,N_19887,N_19767);
nor UO_1317 (O_1317,N_19758,N_19831);
xnor UO_1318 (O_1318,N_19837,N_19767);
and UO_1319 (O_1319,N_19975,N_19771);
xor UO_1320 (O_1320,N_19925,N_19997);
xor UO_1321 (O_1321,N_19878,N_19899);
xnor UO_1322 (O_1322,N_19931,N_19776);
or UO_1323 (O_1323,N_19796,N_19830);
and UO_1324 (O_1324,N_19788,N_19909);
nand UO_1325 (O_1325,N_19889,N_19769);
or UO_1326 (O_1326,N_19888,N_19834);
nand UO_1327 (O_1327,N_19797,N_19960);
nand UO_1328 (O_1328,N_19986,N_19847);
nand UO_1329 (O_1329,N_19962,N_19790);
and UO_1330 (O_1330,N_19863,N_19760);
nor UO_1331 (O_1331,N_19793,N_19920);
nor UO_1332 (O_1332,N_19888,N_19968);
and UO_1333 (O_1333,N_19771,N_19826);
nand UO_1334 (O_1334,N_19886,N_19803);
xnor UO_1335 (O_1335,N_19812,N_19833);
xor UO_1336 (O_1336,N_19783,N_19963);
and UO_1337 (O_1337,N_19900,N_19981);
nor UO_1338 (O_1338,N_19777,N_19862);
and UO_1339 (O_1339,N_19906,N_19929);
nor UO_1340 (O_1340,N_19937,N_19958);
nor UO_1341 (O_1341,N_19918,N_19771);
and UO_1342 (O_1342,N_19817,N_19910);
and UO_1343 (O_1343,N_19798,N_19960);
or UO_1344 (O_1344,N_19836,N_19856);
and UO_1345 (O_1345,N_19815,N_19759);
and UO_1346 (O_1346,N_19820,N_19832);
xor UO_1347 (O_1347,N_19885,N_19986);
nor UO_1348 (O_1348,N_19890,N_19756);
nand UO_1349 (O_1349,N_19789,N_19986);
xor UO_1350 (O_1350,N_19931,N_19918);
or UO_1351 (O_1351,N_19782,N_19831);
xnor UO_1352 (O_1352,N_19902,N_19752);
xor UO_1353 (O_1353,N_19972,N_19939);
and UO_1354 (O_1354,N_19802,N_19824);
nor UO_1355 (O_1355,N_19805,N_19854);
nor UO_1356 (O_1356,N_19750,N_19897);
nand UO_1357 (O_1357,N_19972,N_19956);
nor UO_1358 (O_1358,N_19943,N_19900);
and UO_1359 (O_1359,N_19959,N_19963);
nor UO_1360 (O_1360,N_19879,N_19931);
xnor UO_1361 (O_1361,N_19925,N_19810);
xor UO_1362 (O_1362,N_19992,N_19863);
and UO_1363 (O_1363,N_19943,N_19859);
nor UO_1364 (O_1364,N_19955,N_19878);
nand UO_1365 (O_1365,N_19829,N_19990);
xnor UO_1366 (O_1366,N_19912,N_19863);
or UO_1367 (O_1367,N_19878,N_19871);
or UO_1368 (O_1368,N_19921,N_19791);
nor UO_1369 (O_1369,N_19918,N_19943);
and UO_1370 (O_1370,N_19809,N_19972);
xor UO_1371 (O_1371,N_19908,N_19868);
or UO_1372 (O_1372,N_19852,N_19841);
and UO_1373 (O_1373,N_19789,N_19937);
nor UO_1374 (O_1374,N_19772,N_19752);
and UO_1375 (O_1375,N_19901,N_19772);
nand UO_1376 (O_1376,N_19825,N_19867);
nor UO_1377 (O_1377,N_19772,N_19791);
or UO_1378 (O_1378,N_19911,N_19943);
and UO_1379 (O_1379,N_19854,N_19995);
nand UO_1380 (O_1380,N_19832,N_19848);
nor UO_1381 (O_1381,N_19904,N_19828);
or UO_1382 (O_1382,N_19817,N_19963);
and UO_1383 (O_1383,N_19773,N_19934);
and UO_1384 (O_1384,N_19948,N_19947);
nand UO_1385 (O_1385,N_19968,N_19933);
nand UO_1386 (O_1386,N_19767,N_19800);
and UO_1387 (O_1387,N_19863,N_19875);
nand UO_1388 (O_1388,N_19807,N_19953);
nor UO_1389 (O_1389,N_19970,N_19794);
nor UO_1390 (O_1390,N_19980,N_19945);
nand UO_1391 (O_1391,N_19855,N_19975);
and UO_1392 (O_1392,N_19873,N_19856);
nand UO_1393 (O_1393,N_19791,N_19765);
nor UO_1394 (O_1394,N_19994,N_19832);
nand UO_1395 (O_1395,N_19992,N_19952);
and UO_1396 (O_1396,N_19752,N_19956);
or UO_1397 (O_1397,N_19949,N_19876);
xor UO_1398 (O_1398,N_19846,N_19899);
and UO_1399 (O_1399,N_19919,N_19755);
or UO_1400 (O_1400,N_19914,N_19893);
nor UO_1401 (O_1401,N_19886,N_19976);
and UO_1402 (O_1402,N_19924,N_19794);
and UO_1403 (O_1403,N_19929,N_19892);
nor UO_1404 (O_1404,N_19935,N_19792);
and UO_1405 (O_1405,N_19841,N_19978);
nor UO_1406 (O_1406,N_19841,N_19884);
xnor UO_1407 (O_1407,N_19894,N_19851);
xnor UO_1408 (O_1408,N_19781,N_19838);
nor UO_1409 (O_1409,N_19850,N_19785);
nor UO_1410 (O_1410,N_19855,N_19986);
nor UO_1411 (O_1411,N_19986,N_19879);
xor UO_1412 (O_1412,N_19845,N_19904);
xor UO_1413 (O_1413,N_19989,N_19806);
and UO_1414 (O_1414,N_19955,N_19842);
xor UO_1415 (O_1415,N_19833,N_19810);
or UO_1416 (O_1416,N_19846,N_19874);
xor UO_1417 (O_1417,N_19940,N_19981);
and UO_1418 (O_1418,N_19944,N_19763);
or UO_1419 (O_1419,N_19977,N_19881);
nor UO_1420 (O_1420,N_19895,N_19962);
nand UO_1421 (O_1421,N_19940,N_19995);
and UO_1422 (O_1422,N_19977,N_19937);
or UO_1423 (O_1423,N_19769,N_19969);
nand UO_1424 (O_1424,N_19838,N_19998);
nand UO_1425 (O_1425,N_19885,N_19758);
nor UO_1426 (O_1426,N_19915,N_19882);
nor UO_1427 (O_1427,N_19765,N_19766);
nor UO_1428 (O_1428,N_19896,N_19854);
xnor UO_1429 (O_1429,N_19812,N_19940);
and UO_1430 (O_1430,N_19782,N_19915);
and UO_1431 (O_1431,N_19933,N_19921);
or UO_1432 (O_1432,N_19965,N_19923);
and UO_1433 (O_1433,N_19921,N_19880);
nand UO_1434 (O_1434,N_19953,N_19808);
nor UO_1435 (O_1435,N_19861,N_19950);
nor UO_1436 (O_1436,N_19991,N_19772);
nor UO_1437 (O_1437,N_19800,N_19941);
or UO_1438 (O_1438,N_19952,N_19929);
xnor UO_1439 (O_1439,N_19940,N_19915);
or UO_1440 (O_1440,N_19904,N_19887);
nor UO_1441 (O_1441,N_19846,N_19960);
nor UO_1442 (O_1442,N_19937,N_19769);
nor UO_1443 (O_1443,N_19886,N_19994);
xor UO_1444 (O_1444,N_19894,N_19902);
xor UO_1445 (O_1445,N_19811,N_19805);
and UO_1446 (O_1446,N_19904,N_19882);
or UO_1447 (O_1447,N_19849,N_19796);
xnor UO_1448 (O_1448,N_19785,N_19864);
xor UO_1449 (O_1449,N_19985,N_19997);
or UO_1450 (O_1450,N_19991,N_19752);
nand UO_1451 (O_1451,N_19799,N_19941);
nor UO_1452 (O_1452,N_19920,N_19934);
nand UO_1453 (O_1453,N_19849,N_19917);
nand UO_1454 (O_1454,N_19878,N_19900);
and UO_1455 (O_1455,N_19997,N_19826);
nand UO_1456 (O_1456,N_19778,N_19762);
xor UO_1457 (O_1457,N_19825,N_19789);
or UO_1458 (O_1458,N_19950,N_19832);
or UO_1459 (O_1459,N_19969,N_19822);
nand UO_1460 (O_1460,N_19764,N_19771);
or UO_1461 (O_1461,N_19771,N_19905);
nand UO_1462 (O_1462,N_19767,N_19881);
nand UO_1463 (O_1463,N_19961,N_19803);
or UO_1464 (O_1464,N_19964,N_19957);
nor UO_1465 (O_1465,N_19879,N_19966);
xnor UO_1466 (O_1466,N_19817,N_19815);
or UO_1467 (O_1467,N_19920,N_19866);
nand UO_1468 (O_1468,N_19879,N_19842);
nand UO_1469 (O_1469,N_19778,N_19923);
nand UO_1470 (O_1470,N_19940,N_19802);
nor UO_1471 (O_1471,N_19851,N_19784);
nor UO_1472 (O_1472,N_19984,N_19988);
nor UO_1473 (O_1473,N_19799,N_19933);
xor UO_1474 (O_1474,N_19967,N_19868);
or UO_1475 (O_1475,N_19782,N_19914);
and UO_1476 (O_1476,N_19964,N_19983);
xor UO_1477 (O_1477,N_19889,N_19956);
nor UO_1478 (O_1478,N_19829,N_19756);
and UO_1479 (O_1479,N_19919,N_19966);
or UO_1480 (O_1480,N_19906,N_19904);
or UO_1481 (O_1481,N_19776,N_19808);
xnor UO_1482 (O_1482,N_19942,N_19954);
xnor UO_1483 (O_1483,N_19827,N_19776);
nand UO_1484 (O_1484,N_19871,N_19835);
or UO_1485 (O_1485,N_19785,N_19831);
nand UO_1486 (O_1486,N_19777,N_19835);
nand UO_1487 (O_1487,N_19773,N_19864);
nor UO_1488 (O_1488,N_19863,N_19845);
or UO_1489 (O_1489,N_19848,N_19928);
nor UO_1490 (O_1490,N_19965,N_19870);
or UO_1491 (O_1491,N_19777,N_19969);
and UO_1492 (O_1492,N_19767,N_19827);
or UO_1493 (O_1493,N_19879,N_19880);
nor UO_1494 (O_1494,N_19834,N_19879);
and UO_1495 (O_1495,N_19882,N_19754);
and UO_1496 (O_1496,N_19870,N_19792);
and UO_1497 (O_1497,N_19922,N_19865);
nor UO_1498 (O_1498,N_19981,N_19835);
or UO_1499 (O_1499,N_19796,N_19931);
xor UO_1500 (O_1500,N_19903,N_19780);
nand UO_1501 (O_1501,N_19889,N_19833);
xnor UO_1502 (O_1502,N_19872,N_19953);
or UO_1503 (O_1503,N_19951,N_19917);
xor UO_1504 (O_1504,N_19923,N_19862);
xnor UO_1505 (O_1505,N_19789,N_19954);
nor UO_1506 (O_1506,N_19830,N_19754);
nand UO_1507 (O_1507,N_19951,N_19909);
or UO_1508 (O_1508,N_19939,N_19864);
nand UO_1509 (O_1509,N_19900,N_19826);
xnor UO_1510 (O_1510,N_19919,N_19784);
and UO_1511 (O_1511,N_19751,N_19897);
nand UO_1512 (O_1512,N_19899,N_19942);
xor UO_1513 (O_1513,N_19961,N_19797);
nand UO_1514 (O_1514,N_19921,N_19917);
nand UO_1515 (O_1515,N_19844,N_19770);
nand UO_1516 (O_1516,N_19920,N_19988);
and UO_1517 (O_1517,N_19925,N_19873);
nand UO_1518 (O_1518,N_19867,N_19860);
or UO_1519 (O_1519,N_19800,N_19919);
nand UO_1520 (O_1520,N_19900,N_19884);
nand UO_1521 (O_1521,N_19800,N_19967);
or UO_1522 (O_1522,N_19869,N_19833);
nor UO_1523 (O_1523,N_19866,N_19913);
and UO_1524 (O_1524,N_19995,N_19933);
nand UO_1525 (O_1525,N_19980,N_19996);
and UO_1526 (O_1526,N_19811,N_19976);
or UO_1527 (O_1527,N_19892,N_19802);
xnor UO_1528 (O_1528,N_19980,N_19934);
xor UO_1529 (O_1529,N_19803,N_19853);
nand UO_1530 (O_1530,N_19886,N_19903);
xnor UO_1531 (O_1531,N_19861,N_19893);
nand UO_1532 (O_1532,N_19799,N_19985);
xor UO_1533 (O_1533,N_19810,N_19968);
nand UO_1534 (O_1534,N_19898,N_19858);
and UO_1535 (O_1535,N_19827,N_19850);
or UO_1536 (O_1536,N_19965,N_19904);
or UO_1537 (O_1537,N_19771,N_19871);
nor UO_1538 (O_1538,N_19790,N_19966);
xnor UO_1539 (O_1539,N_19866,N_19819);
nand UO_1540 (O_1540,N_19810,N_19974);
xor UO_1541 (O_1541,N_19826,N_19842);
and UO_1542 (O_1542,N_19956,N_19847);
nor UO_1543 (O_1543,N_19845,N_19974);
or UO_1544 (O_1544,N_19755,N_19766);
nor UO_1545 (O_1545,N_19977,N_19764);
and UO_1546 (O_1546,N_19766,N_19806);
nand UO_1547 (O_1547,N_19920,N_19933);
or UO_1548 (O_1548,N_19972,N_19850);
xnor UO_1549 (O_1549,N_19922,N_19931);
nor UO_1550 (O_1550,N_19826,N_19984);
xnor UO_1551 (O_1551,N_19866,N_19766);
and UO_1552 (O_1552,N_19886,N_19827);
nor UO_1553 (O_1553,N_19890,N_19981);
nand UO_1554 (O_1554,N_19971,N_19943);
nor UO_1555 (O_1555,N_19949,N_19926);
xnor UO_1556 (O_1556,N_19993,N_19914);
nor UO_1557 (O_1557,N_19927,N_19915);
or UO_1558 (O_1558,N_19826,N_19924);
or UO_1559 (O_1559,N_19776,N_19910);
nand UO_1560 (O_1560,N_19927,N_19799);
xnor UO_1561 (O_1561,N_19756,N_19891);
and UO_1562 (O_1562,N_19837,N_19896);
xor UO_1563 (O_1563,N_19996,N_19939);
nand UO_1564 (O_1564,N_19827,N_19956);
and UO_1565 (O_1565,N_19895,N_19787);
or UO_1566 (O_1566,N_19834,N_19885);
nor UO_1567 (O_1567,N_19811,N_19918);
nor UO_1568 (O_1568,N_19788,N_19970);
and UO_1569 (O_1569,N_19964,N_19878);
nor UO_1570 (O_1570,N_19829,N_19876);
or UO_1571 (O_1571,N_19973,N_19753);
or UO_1572 (O_1572,N_19764,N_19952);
or UO_1573 (O_1573,N_19825,N_19892);
nor UO_1574 (O_1574,N_19757,N_19756);
nand UO_1575 (O_1575,N_19826,N_19786);
xor UO_1576 (O_1576,N_19972,N_19876);
or UO_1577 (O_1577,N_19862,N_19764);
and UO_1578 (O_1578,N_19991,N_19785);
nand UO_1579 (O_1579,N_19800,N_19916);
nor UO_1580 (O_1580,N_19915,N_19848);
nand UO_1581 (O_1581,N_19756,N_19847);
nand UO_1582 (O_1582,N_19990,N_19803);
or UO_1583 (O_1583,N_19854,N_19802);
xor UO_1584 (O_1584,N_19996,N_19890);
nor UO_1585 (O_1585,N_19883,N_19772);
nand UO_1586 (O_1586,N_19996,N_19923);
nand UO_1587 (O_1587,N_19924,N_19830);
or UO_1588 (O_1588,N_19777,N_19971);
nor UO_1589 (O_1589,N_19989,N_19771);
or UO_1590 (O_1590,N_19864,N_19776);
nor UO_1591 (O_1591,N_19865,N_19842);
nor UO_1592 (O_1592,N_19945,N_19948);
or UO_1593 (O_1593,N_19782,N_19907);
and UO_1594 (O_1594,N_19783,N_19840);
nand UO_1595 (O_1595,N_19922,N_19911);
nand UO_1596 (O_1596,N_19801,N_19897);
xnor UO_1597 (O_1597,N_19929,N_19765);
nor UO_1598 (O_1598,N_19786,N_19915);
and UO_1599 (O_1599,N_19850,N_19967);
nor UO_1600 (O_1600,N_19772,N_19763);
xor UO_1601 (O_1601,N_19992,N_19761);
xor UO_1602 (O_1602,N_19866,N_19899);
nand UO_1603 (O_1603,N_19792,N_19854);
nor UO_1604 (O_1604,N_19998,N_19812);
nor UO_1605 (O_1605,N_19858,N_19906);
and UO_1606 (O_1606,N_19795,N_19791);
and UO_1607 (O_1607,N_19825,N_19886);
and UO_1608 (O_1608,N_19795,N_19980);
nand UO_1609 (O_1609,N_19947,N_19788);
nand UO_1610 (O_1610,N_19957,N_19965);
and UO_1611 (O_1611,N_19873,N_19802);
or UO_1612 (O_1612,N_19815,N_19755);
xor UO_1613 (O_1613,N_19827,N_19816);
nor UO_1614 (O_1614,N_19866,N_19783);
and UO_1615 (O_1615,N_19862,N_19977);
and UO_1616 (O_1616,N_19753,N_19820);
nand UO_1617 (O_1617,N_19920,N_19839);
or UO_1618 (O_1618,N_19854,N_19757);
and UO_1619 (O_1619,N_19951,N_19961);
and UO_1620 (O_1620,N_19839,N_19946);
and UO_1621 (O_1621,N_19984,N_19958);
xor UO_1622 (O_1622,N_19868,N_19842);
nand UO_1623 (O_1623,N_19806,N_19751);
xnor UO_1624 (O_1624,N_19866,N_19834);
nor UO_1625 (O_1625,N_19813,N_19837);
and UO_1626 (O_1626,N_19814,N_19957);
xnor UO_1627 (O_1627,N_19864,N_19974);
nor UO_1628 (O_1628,N_19940,N_19914);
nor UO_1629 (O_1629,N_19810,N_19995);
nand UO_1630 (O_1630,N_19987,N_19857);
or UO_1631 (O_1631,N_19956,N_19783);
xor UO_1632 (O_1632,N_19999,N_19757);
xnor UO_1633 (O_1633,N_19965,N_19821);
nand UO_1634 (O_1634,N_19767,N_19867);
xnor UO_1635 (O_1635,N_19809,N_19900);
and UO_1636 (O_1636,N_19972,N_19889);
nand UO_1637 (O_1637,N_19999,N_19827);
xor UO_1638 (O_1638,N_19753,N_19808);
or UO_1639 (O_1639,N_19790,N_19828);
nor UO_1640 (O_1640,N_19980,N_19957);
or UO_1641 (O_1641,N_19785,N_19818);
xnor UO_1642 (O_1642,N_19795,N_19764);
or UO_1643 (O_1643,N_19758,N_19909);
and UO_1644 (O_1644,N_19800,N_19991);
nand UO_1645 (O_1645,N_19905,N_19926);
xor UO_1646 (O_1646,N_19788,N_19804);
xor UO_1647 (O_1647,N_19968,N_19777);
nor UO_1648 (O_1648,N_19799,N_19878);
and UO_1649 (O_1649,N_19805,N_19756);
and UO_1650 (O_1650,N_19983,N_19806);
nor UO_1651 (O_1651,N_19822,N_19958);
and UO_1652 (O_1652,N_19864,N_19847);
nand UO_1653 (O_1653,N_19958,N_19765);
and UO_1654 (O_1654,N_19803,N_19848);
or UO_1655 (O_1655,N_19885,N_19853);
nor UO_1656 (O_1656,N_19953,N_19817);
and UO_1657 (O_1657,N_19859,N_19975);
xor UO_1658 (O_1658,N_19910,N_19957);
nand UO_1659 (O_1659,N_19782,N_19964);
nand UO_1660 (O_1660,N_19882,N_19879);
and UO_1661 (O_1661,N_19913,N_19886);
nand UO_1662 (O_1662,N_19917,N_19923);
nor UO_1663 (O_1663,N_19834,N_19798);
and UO_1664 (O_1664,N_19751,N_19786);
nand UO_1665 (O_1665,N_19986,N_19762);
or UO_1666 (O_1666,N_19830,N_19756);
and UO_1667 (O_1667,N_19774,N_19950);
or UO_1668 (O_1668,N_19849,N_19769);
nand UO_1669 (O_1669,N_19864,N_19981);
nand UO_1670 (O_1670,N_19971,N_19814);
nand UO_1671 (O_1671,N_19770,N_19852);
nand UO_1672 (O_1672,N_19915,N_19776);
or UO_1673 (O_1673,N_19892,N_19855);
xor UO_1674 (O_1674,N_19841,N_19933);
nor UO_1675 (O_1675,N_19837,N_19897);
and UO_1676 (O_1676,N_19839,N_19818);
xnor UO_1677 (O_1677,N_19913,N_19945);
nor UO_1678 (O_1678,N_19913,N_19990);
and UO_1679 (O_1679,N_19868,N_19752);
xor UO_1680 (O_1680,N_19911,N_19827);
and UO_1681 (O_1681,N_19787,N_19868);
nor UO_1682 (O_1682,N_19997,N_19959);
xor UO_1683 (O_1683,N_19811,N_19868);
and UO_1684 (O_1684,N_19752,N_19793);
nand UO_1685 (O_1685,N_19894,N_19876);
nand UO_1686 (O_1686,N_19971,N_19965);
xor UO_1687 (O_1687,N_19977,N_19783);
nor UO_1688 (O_1688,N_19774,N_19870);
and UO_1689 (O_1689,N_19867,N_19942);
nor UO_1690 (O_1690,N_19980,N_19982);
xnor UO_1691 (O_1691,N_19822,N_19827);
or UO_1692 (O_1692,N_19860,N_19799);
and UO_1693 (O_1693,N_19873,N_19973);
nor UO_1694 (O_1694,N_19920,N_19883);
nor UO_1695 (O_1695,N_19982,N_19875);
and UO_1696 (O_1696,N_19995,N_19757);
xnor UO_1697 (O_1697,N_19998,N_19931);
nand UO_1698 (O_1698,N_19813,N_19911);
xor UO_1699 (O_1699,N_19860,N_19884);
or UO_1700 (O_1700,N_19805,N_19885);
xnor UO_1701 (O_1701,N_19946,N_19856);
and UO_1702 (O_1702,N_19954,N_19846);
or UO_1703 (O_1703,N_19943,N_19892);
nand UO_1704 (O_1704,N_19989,N_19917);
and UO_1705 (O_1705,N_19812,N_19856);
and UO_1706 (O_1706,N_19844,N_19930);
and UO_1707 (O_1707,N_19871,N_19808);
and UO_1708 (O_1708,N_19990,N_19833);
nand UO_1709 (O_1709,N_19817,N_19752);
xnor UO_1710 (O_1710,N_19773,N_19814);
and UO_1711 (O_1711,N_19872,N_19766);
or UO_1712 (O_1712,N_19858,N_19952);
nor UO_1713 (O_1713,N_19994,N_19956);
xnor UO_1714 (O_1714,N_19900,N_19814);
nor UO_1715 (O_1715,N_19892,N_19987);
nand UO_1716 (O_1716,N_19881,N_19886);
nor UO_1717 (O_1717,N_19753,N_19892);
and UO_1718 (O_1718,N_19822,N_19860);
and UO_1719 (O_1719,N_19821,N_19900);
or UO_1720 (O_1720,N_19977,N_19791);
and UO_1721 (O_1721,N_19763,N_19986);
xnor UO_1722 (O_1722,N_19759,N_19824);
and UO_1723 (O_1723,N_19763,N_19824);
nand UO_1724 (O_1724,N_19916,N_19826);
or UO_1725 (O_1725,N_19802,N_19906);
and UO_1726 (O_1726,N_19833,N_19816);
nand UO_1727 (O_1727,N_19845,N_19819);
xnor UO_1728 (O_1728,N_19916,N_19790);
nand UO_1729 (O_1729,N_19943,N_19969);
and UO_1730 (O_1730,N_19981,N_19912);
nor UO_1731 (O_1731,N_19968,N_19912);
and UO_1732 (O_1732,N_19940,N_19991);
nand UO_1733 (O_1733,N_19847,N_19755);
and UO_1734 (O_1734,N_19928,N_19999);
and UO_1735 (O_1735,N_19910,N_19879);
nor UO_1736 (O_1736,N_19994,N_19900);
nor UO_1737 (O_1737,N_19878,N_19757);
or UO_1738 (O_1738,N_19989,N_19888);
and UO_1739 (O_1739,N_19840,N_19860);
or UO_1740 (O_1740,N_19852,N_19821);
and UO_1741 (O_1741,N_19932,N_19888);
nor UO_1742 (O_1742,N_19797,N_19889);
xor UO_1743 (O_1743,N_19971,N_19775);
or UO_1744 (O_1744,N_19921,N_19939);
xnor UO_1745 (O_1745,N_19813,N_19890);
nand UO_1746 (O_1746,N_19876,N_19939);
nor UO_1747 (O_1747,N_19917,N_19969);
xnor UO_1748 (O_1748,N_19973,N_19881);
xnor UO_1749 (O_1749,N_19997,N_19939);
nand UO_1750 (O_1750,N_19997,N_19970);
nor UO_1751 (O_1751,N_19915,N_19962);
and UO_1752 (O_1752,N_19980,N_19967);
and UO_1753 (O_1753,N_19990,N_19949);
nor UO_1754 (O_1754,N_19795,N_19917);
and UO_1755 (O_1755,N_19884,N_19788);
nand UO_1756 (O_1756,N_19951,N_19759);
or UO_1757 (O_1757,N_19917,N_19896);
or UO_1758 (O_1758,N_19954,N_19900);
nand UO_1759 (O_1759,N_19840,N_19984);
nor UO_1760 (O_1760,N_19804,N_19985);
and UO_1761 (O_1761,N_19782,N_19847);
and UO_1762 (O_1762,N_19892,N_19773);
or UO_1763 (O_1763,N_19790,N_19768);
nor UO_1764 (O_1764,N_19792,N_19773);
and UO_1765 (O_1765,N_19801,N_19932);
nor UO_1766 (O_1766,N_19765,N_19963);
nor UO_1767 (O_1767,N_19846,N_19985);
or UO_1768 (O_1768,N_19951,N_19882);
nand UO_1769 (O_1769,N_19756,N_19882);
or UO_1770 (O_1770,N_19751,N_19937);
xor UO_1771 (O_1771,N_19931,N_19849);
or UO_1772 (O_1772,N_19975,N_19885);
or UO_1773 (O_1773,N_19780,N_19758);
nand UO_1774 (O_1774,N_19786,N_19829);
xnor UO_1775 (O_1775,N_19827,N_19986);
nand UO_1776 (O_1776,N_19808,N_19818);
nand UO_1777 (O_1777,N_19916,N_19858);
or UO_1778 (O_1778,N_19982,N_19892);
or UO_1779 (O_1779,N_19989,N_19901);
and UO_1780 (O_1780,N_19884,N_19958);
and UO_1781 (O_1781,N_19752,N_19829);
nand UO_1782 (O_1782,N_19914,N_19766);
xor UO_1783 (O_1783,N_19908,N_19790);
nand UO_1784 (O_1784,N_19814,N_19770);
xnor UO_1785 (O_1785,N_19753,N_19898);
or UO_1786 (O_1786,N_19930,N_19793);
nand UO_1787 (O_1787,N_19903,N_19868);
xnor UO_1788 (O_1788,N_19810,N_19855);
or UO_1789 (O_1789,N_19908,N_19859);
and UO_1790 (O_1790,N_19788,N_19768);
nor UO_1791 (O_1791,N_19895,N_19928);
xnor UO_1792 (O_1792,N_19851,N_19957);
or UO_1793 (O_1793,N_19915,N_19840);
xnor UO_1794 (O_1794,N_19821,N_19973);
nor UO_1795 (O_1795,N_19978,N_19759);
nor UO_1796 (O_1796,N_19816,N_19902);
xor UO_1797 (O_1797,N_19848,N_19937);
and UO_1798 (O_1798,N_19964,N_19894);
xnor UO_1799 (O_1799,N_19928,N_19776);
xnor UO_1800 (O_1800,N_19955,N_19897);
nand UO_1801 (O_1801,N_19929,N_19927);
or UO_1802 (O_1802,N_19798,N_19761);
or UO_1803 (O_1803,N_19772,N_19847);
nor UO_1804 (O_1804,N_19988,N_19760);
nor UO_1805 (O_1805,N_19995,N_19899);
and UO_1806 (O_1806,N_19965,N_19754);
nand UO_1807 (O_1807,N_19773,N_19753);
and UO_1808 (O_1808,N_19943,N_19958);
or UO_1809 (O_1809,N_19847,N_19821);
nand UO_1810 (O_1810,N_19972,N_19950);
xor UO_1811 (O_1811,N_19956,N_19894);
nand UO_1812 (O_1812,N_19882,N_19910);
and UO_1813 (O_1813,N_19790,N_19987);
nor UO_1814 (O_1814,N_19764,N_19830);
and UO_1815 (O_1815,N_19985,N_19844);
xnor UO_1816 (O_1816,N_19751,N_19987);
and UO_1817 (O_1817,N_19931,N_19925);
nor UO_1818 (O_1818,N_19779,N_19830);
and UO_1819 (O_1819,N_19779,N_19970);
or UO_1820 (O_1820,N_19891,N_19821);
xnor UO_1821 (O_1821,N_19888,N_19811);
and UO_1822 (O_1822,N_19980,N_19783);
or UO_1823 (O_1823,N_19810,N_19788);
and UO_1824 (O_1824,N_19863,N_19846);
nor UO_1825 (O_1825,N_19916,N_19967);
nand UO_1826 (O_1826,N_19779,N_19949);
nand UO_1827 (O_1827,N_19972,N_19885);
or UO_1828 (O_1828,N_19802,N_19958);
or UO_1829 (O_1829,N_19869,N_19898);
and UO_1830 (O_1830,N_19803,N_19998);
xnor UO_1831 (O_1831,N_19962,N_19925);
and UO_1832 (O_1832,N_19942,N_19946);
or UO_1833 (O_1833,N_19886,N_19885);
and UO_1834 (O_1834,N_19862,N_19963);
or UO_1835 (O_1835,N_19984,N_19818);
or UO_1836 (O_1836,N_19750,N_19925);
or UO_1837 (O_1837,N_19863,N_19935);
nand UO_1838 (O_1838,N_19783,N_19826);
nor UO_1839 (O_1839,N_19931,N_19843);
or UO_1840 (O_1840,N_19823,N_19861);
nand UO_1841 (O_1841,N_19854,N_19926);
nand UO_1842 (O_1842,N_19890,N_19941);
or UO_1843 (O_1843,N_19857,N_19935);
and UO_1844 (O_1844,N_19852,N_19965);
nand UO_1845 (O_1845,N_19810,N_19918);
xnor UO_1846 (O_1846,N_19918,N_19751);
nand UO_1847 (O_1847,N_19895,N_19763);
nand UO_1848 (O_1848,N_19792,N_19781);
nor UO_1849 (O_1849,N_19802,N_19775);
xor UO_1850 (O_1850,N_19853,N_19916);
nor UO_1851 (O_1851,N_19767,N_19879);
or UO_1852 (O_1852,N_19957,N_19983);
or UO_1853 (O_1853,N_19795,N_19928);
or UO_1854 (O_1854,N_19972,N_19991);
or UO_1855 (O_1855,N_19990,N_19804);
or UO_1856 (O_1856,N_19950,N_19963);
nor UO_1857 (O_1857,N_19935,N_19959);
nor UO_1858 (O_1858,N_19828,N_19993);
or UO_1859 (O_1859,N_19817,N_19782);
nor UO_1860 (O_1860,N_19812,N_19993);
or UO_1861 (O_1861,N_19989,N_19865);
nand UO_1862 (O_1862,N_19778,N_19936);
nor UO_1863 (O_1863,N_19898,N_19806);
nor UO_1864 (O_1864,N_19954,N_19838);
nor UO_1865 (O_1865,N_19753,N_19825);
or UO_1866 (O_1866,N_19812,N_19902);
and UO_1867 (O_1867,N_19897,N_19995);
and UO_1868 (O_1868,N_19831,N_19850);
or UO_1869 (O_1869,N_19913,N_19915);
and UO_1870 (O_1870,N_19900,N_19910);
or UO_1871 (O_1871,N_19867,N_19796);
and UO_1872 (O_1872,N_19934,N_19837);
xnor UO_1873 (O_1873,N_19906,N_19933);
nor UO_1874 (O_1874,N_19772,N_19889);
and UO_1875 (O_1875,N_19781,N_19968);
nand UO_1876 (O_1876,N_19969,N_19901);
or UO_1877 (O_1877,N_19989,N_19998);
nor UO_1878 (O_1878,N_19801,N_19962);
nand UO_1879 (O_1879,N_19976,N_19800);
xnor UO_1880 (O_1880,N_19972,N_19973);
nor UO_1881 (O_1881,N_19811,N_19945);
and UO_1882 (O_1882,N_19819,N_19949);
xor UO_1883 (O_1883,N_19933,N_19853);
and UO_1884 (O_1884,N_19914,N_19888);
nand UO_1885 (O_1885,N_19838,N_19811);
nor UO_1886 (O_1886,N_19772,N_19987);
and UO_1887 (O_1887,N_19839,N_19959);
nor UO_1888 (O_1888,N_19992,N_19807);
nor UO_1889 (O_1889,N_19880,N_19750);
xnor UO_1890 (O_1890,N_19910,N_19812);
and UO_1891 (O_1891,N_19919,N_19880);
xor UO_1892 (O_1892,N_19935,N_19989);
xor UO_1893 (O_1893,N_19977,N_19945);
nand UO_1894 (O_1894,N_19814,N_19839);
xor UO_1895 (O_1895,N_19841,N_19963);
nand UO_1896 (O_1896,N_19937,N_19897);
xor UO_1897 (O_1897,N_19842,N_19789);
nand UO_1898 (O_1898,N_19836,N_19880);
nand UO_1899 (O_1899,N_19896,N_19798);
and UO_1900 (O_1900,N_19831,N_19878);
and UO_1901 (O_1901,N_19899,N_19798);
xor UO_1902 (O_1902,N_19753,N_19882);
and UO_1903 (O_1903,N_19872,N_19827);
nor UO_1904 (O_1904,N_19921,N_19993);
nand UO_1905 (O_1905,N_19837,N_19760);
and UO_1906 (O_1906,N_19882,N_19770);
and UO_1907 (O_1907,N_19756,N_19768);
and UO_1908 (O_1908,N_19839,N_19867);
and UO_1909 (O_1909,N_19822,N_19856);
and UO_1910 (O_1910,N_19764,N_19911);
nand UO_1911 (O_1911,N_19832,N_19971);
or UO_1912 (O_1912,N_19867,N_19795);
xnor UO_1913 (O_1913,N_19968,N_19800);
nor UO_1914 (O_1914,N_19889,N_19882);
or UO_1915 (O_1915,N_19945,N_19879);
nand UO_1916 (O_1916,N_19961,N_19965);
nand UO_1917 (O_1917,N_19971,N_19836);
or UO_1918 (O_1918,N_19845,N_19811);
nand UO_1919 (O_1919,N_19787,N_19912);
or UO_1920 (O_1920,N_19857,N_19846);
and UO_1921 (O_1921,N_19785,N_19902);
nor UO_1922 (O_1922,N_19755,N_19790);
or UO_1923 (O_1923,N_19851,N_19783);
and UO_1924 (O_1924,N_19941,N_19785);
nor UO_1925 (O_1925,N_19864,N_19909);
nor UO_1926 (O_1926,N_19917,N_19997);
nor UO_1927 (O_1927,N_19755,N_19963);
or UO_1928 (O_1928,N_19758,N_19833);
nor UO_1929 (O_1929,N_19975,N_19753);
and UO_1930 (O_1930,N_19792,N_19942);
and UO_1931 (O_1931,N_19891,N_19789);
or UO_1932 (O_1932,N_19977,N_19959);
nor UO_1933 (O_1933,N_19944,N_19767);
and UO_1934 (O_1934,N_19789,N_19851);
nand UO_1935 (O_1935,N_19932,N_19934);
or UO_1936 (O_1936,N_19917,N_19817);
xor UO_1937 (O_1937,N_19909,N_19997);
and UO_1938 (O_1938,N_19980,N_19794);
or UO_1939 (O_1939,N_19964,N_19828);
xnor UO_1940 (O_1940,N_19980,N_19763);
or UO_1941 (O_1941,N_19816,N_19970);
nand UO_1942 (O_1942,N_19854,N_19763);
xor UO_1943 (O_1943,N_19872,N_19919);
xnor UO_1944 (O_1944,N_19833,N_19915);
xor UO_1945 (O_1945,N_19999,N_19864);
and UO_1946 (O_1946,N_19841,N_19873);
and UO_1947 (O_1947,N_19985,N_19944);
nand UO_1948 (O_1948,N_19820,N_19941);
and UO_1949 (O_1949,N_19972,N_19988);
and UO_1950 (O_1950,N_19762,N_19946);
xor UO_1951 (O_1951,N_19764,N_19923);
xnor UO_1952 (O_1952,N_19971,N_19969);
nor UO_1953 (O_1953,N_19939,N_19798);
nand UO_1954 (O_1954,N_19793,N_19945);
nand UO_1955 (O_1955,N_19852,N_19883);
xor UO_1956 (O_1956,N_19866,N_19926);
xor UO_1957 (O_1957,N_19949,N_19798);
nor UO_1958 (O_1958,N_19764,N_19893);
nor UO_1959 (O_1959,N_19774,N_19800);
and UO_1960 (O_1960,N_19945,N_19947);
or UO_1961 (O_1961,N_19935,N_19902);
nand UO_1962 (O_1962,N_19759,N_19774);
nor UO_1963 (O_1963,N_19781,N_19978);
nand UO_1964 (O_1964,N_19935,N_19927);
or UO_1965 (O_1965,N_19797,N_19774);
nor UO_1966 (O_1966,N_19917,N_19873);
xnor UO_1967 (O_1967,N_19812,N_19798);
nor UO_1968 (O_1968,N_19768,N_19860);
or UO_1969 (O_1969,N_19896,N_19752);
xor UO_1970 (O_1970,N_19989,N_19778);
or UO_1971 (O_1971,N_19795,N_19863);
nand UO_1972 (O_1972,N_19848,N_19819);
xor UO_1973 (O_1973,N_19761,N_19814);
nor UO_1974 (O_1974,N_19982,N_19981);
nor UO_1975 (O_1975,N_19822,N_19823);
xor UO_1976 (O_1976,N_19954,N_19836);
nor UO_1977 (O_1977,N_19910,N_19850);
nand UO_1978 (O_1978,N_19938,N_19765);
nand UO_1979 (O_1979,N_19958,N_19851);
nor UO_1980 (O_1980,N_19761,N_19929);
and UO_1981 (O_1981,N_19905,N_19832);
or UO_1982 (O_1982,N_19798,N_19881);
or UO_1983 (O_1983,N_19783,N_19937);
or UO_1984 (O_1984,N_19985,N_19808);
or UO_1985 (O_1985,N_19988,N_19823);
xnor UO_1986 (O_1986,N_19806,N_19910);
or UO_1987 (O_1987,N_19903,N_19973);
xnor UO_1988 (O_1988,N_19808,N_19872);
xnor UO_1989 (O_1989,N_19951,N_19901);
nand UO_1990 (O_1990,N_19751,N_19969);
nand UO_1991 (O_1991,N_19950,N_19836);
nor UO_1992 (O_1992,N_19955,N_19993);
xnor UO_1993 (O_1993,N_19991,N_19788);
or UO_1994 (O_1994,N_19849,N_19877);
and UO_1995 (O_1995,N_19755,N_19774);
and UO_1996 (O_1996,N_19835,N_19982);
xor UO_1997 (O_1997,N_19816,N_19825);
and UO_1998 (O_1998,N_19904,N_19813);
nor UO_1999 (O_1999,N_19834,N_19836);
nand UO_2000 (O_2000,N_19933,N_19982);
and UO_2001 (O_2001,N_19908,N_19958);
nor UO_2002 (O_2002,N_19832,N_19864);
nand UO_2003 (O_2003,N_19758,N_19769);
nor UO_2004 (O_2004,N_19854,N_19801);
or UO_2005 (O_2005,N_19759,N_19949);
nand UO_2006 (O_2006,N_19938,N_19768);
nor UO_2007 (O_2007,N_19766,N_19870);
xnor UO_2008 (O_2008,N_19849,N_19833);
xnor UO_2009 (O_2009,N_19889,N_19892);
nor UO_2010 (O_2010,N_19961,N_19755);
and UO_2011 (O_2011,N_19846,N_19841);
nor UO_2012 (O_2012,N_19908,N_19917);
or UO_2013 (O_2013,N_19811,N_19881);
and UO_2014 (O_2014,N_19958,N_19796);
nand UO_2015 (O_2015,N_19805,N_19843);
nor UO_2016 (O_2016,N_19980,N_19978);
nor UO_2017 (O_2017,N_19963,N_19989);
xnor UO_2018 (O_2018,N_19849,N_19966);
nand UO_2019 (O_2019,N_19854,N_19833);
and UO_2020 (O_2020,N_19826,N_19870);
and UO_2021 (O_2021,N_19792,N_19941);
and UO_2022 (O_2022,N_19791,N_19923);
nor UO_2023 (O_2023,N_19811,N_19997);
xnor UO_2024 (O_2024,N_19831,N_19955);
and UO_2025 (O_2025,N_19835,N_19945);
and UO_2026 (O_2026,N_19800,N_19896);
or UO_2027 (O_2027,N_19925,N_19866);
xnor UO_2028 (O_2028,N_19947,N_19815);
or UO_2029 (O_2029,N_19789,N_19927);
nand UO_2030 (O_2030,N_19812,N_19758);
or UO_2031 (O_2031,N_19820,N_19794);
xor UO_2032 (O_2032,N_19992,N_19892);
xor UO_2033 (O_2033,N_19752,N_19874);
and UO_2034 (O_2034,N_19942,N_19910);
nand UO_2035 (O_2035,N_19923,N_19891);
or UO_2036 (O_2036,N_19784,N_19764);
xor UO_2037 (O_2037,N_19874,N_19785);
nand UO_2038 (O_2038,N_19906,N_19901);
nor UO_2039 (O_2039,N_19844,N_19806);
nor UO_2040 (O_2040,N_19861,N_19750);
nand UO_2041 (O_2041,N_19965,N_19839);
and UO_2042 (O_2042,N_19913,N_19833);
nor UO_2043 (O_2043,N_19790,N_19968);
nor UO_2044 (O_2044,N_19891,N_19998);
and UO_2045 (O_2045,N_19966,N_19917);
and UO_2046 (O_2046,N_19922,N_19833);
nor UO_2047 (O_2047,N_19919,N_19809);
xor UO_2048 (O_2048,N_19925,N_19803);
and UO_2049 (O_2049,N_19793,N_19773);
xnor UO_2050 (O_2050,N_19900,N_19942);
nor UO_2051 (O_2051,N_19842,N_19802);
or UO_2052 (O_2052,N_19848,N_19950);
nor UO_2053 (O_2053,N_19782,N_19939);
or UO_2054 (O_2054,N_19960,N_19967);
nor UO_2055 (O_2055,N_19823,N_19900);
or UO_2056 (O_2056,N_19912,N_19874);
nand UO_2057 (O_2057,N_19974,N_19977);
nand UO_2058 (O_2058,N_19840,N_19943);
xnor UO_2059 (O_2059,N_19793,N_19986);
nand UO_2060 (O_2060,N_19879,N_19869);
and UO_2061 (O_2061,N_19936,N_19777);
or UO_2062 (O_2062,N_19867,N_19788);
nand UO_2063 (O_2063,N_19882,N_19760);
nand UO_2064 (O_2064,N_19990,N_19783);
xnor UO_2065 (O_2065,N_19882,N_19975);
and UO_2066 (O_2066,N_19791,N_19783);
nand UO_2067 (O_2067,N_19781,N_19964);
nor UO_2068 (O_2068,N_19765,N_19756);
nand UO_2069 (O_2069,N_19913,N_19805);
and UO_2070 (O_2070,N_19856,N_19932);
and UO_2071 (O_2071,N_19794,N_19996);
or UO_2072 (O_2072,N_19826,N_19854);
nand UO_2073 (O_2073,N_19796,N_19787);
nor UO_2074 (O_2074,N_19951,N_19937);
nor UO_2075 (O_2075,N_19903,N_19968);
nor UO_2076 (O_2076,N_19838,N_19865);
xor UO_2077 (O_2077,N_19998,N_19795);
and UO_2078 (O_2078,N_19866,N_19842);
xnor UO_2079 (O_2079,N_19766,N_19819);
xnor UO_2080 (O_2080,N_19808,N_19960);
xnor UO_2081 (O_2081,N_19952,N_19833);
and UO_2082 (O_2082,N_19897,N_19797);
xor UO_2083 (O_2083,N_19859,N_19775);
and UO_2084 (O_2084,N_19886,N_19964);
or UO_2085 (O_2085,N_19800,N_19776);
or UO_2086 (O_2086,N_19756,N_19755);
xnor UO_2087 (O_2087,N_19784,N_19939);
xor UO_2088 (O_2088,N_19968,N_19999);
and UO_2089 (O_2089,N_19932,N_19977);
and UO_2090 (O_2090,N_19813,N_19840);
and UO_2091 (O_2091,N_19828,N_19936);
or UO_2092 (O_2092,N_19903,N_19889);
nor UO_2093 (O_2093,N_19766,N_19887);
nor UO_2094 (O_2094,N_19939,N_19807);
xor UO_2095 (O_2095,N_19837,N_19790);
nand UO_2096 (O_2096,N_19993,N_19879);
and UO_2097 (O_2097,N_19898,N_19862);
xnor UO_2098 (O_2098,N_19841,N_19786);
or UO_2099 (O_2099,N_19850,N_19943);
nand UO_2100 (O_2100,N_19931,N_19959);
and UO_2101 (O_2101,N_19998,N_19804);
nor UO_2102 (O_2102,N_19911,N_19990);
nor UO_2103 (O_2103,N_19825,N_19969);
xor UO_2104 (O_2104,N_19860,N_19779);
and UO_2105 (O_2105,N_19832,N_19873);
nor UO_2106 (O_2106,N_19802,N_19960);
xnor UO_2107 (O_2107,N_19787,N_19918);
nand UO_2108 (O_2108,N_19823,N_19938);
and UO_2109 (O_2109,N_19888,N_19795);
and UO_2110 (O_2110,N_19912,N_19926);
xnor UO_2111 (O_2111,N_19859,N_19861);
and UO_2112 (O_2112,N_19970,N_19780);
nand UO_2113 (O_2113,N_19888,N_19777);
and UO_2114 (O_2114,N_19856,N_19831);
and UO_2115 (O_2115,N_19944,N_19975);
nor UO_2116 (O_2116,N_19904,N_19862);
nor UO_2117 (O_2117,N_19816,N_19811);
nand UO_2118 (O_2118,N_19895,N_19835);
nor UO_2119 (O_2119,N_19875,N_19821);
nand UO_2120 (O_2120,N_19946,N_19791);
and UO_2121 (O_2121,N_19766,N_19799);
or UO_2122 (O_2122,N_19985,N_19780);
nand UO_2123 (O_2123,N_19780,N_19935);
and UO_2124 (O_2124,N_19841,N_19860);
xor UO_2125 (O_2125,N_19904,N_19863);
or UO_2126 (O_2126,N_19818,N_19761);
and UO_2127 (O_2127,N_19750,N_19798);
nor UO_2128 (O_2128,N_19867,N_19874);
and UO_2129 (O_2129,N_19930,N_19980);
nor UO_2130 (O_2130,N_19836,N_19982);
nor UO_2131 (O_2131,N_19811,N_19855);
and UO_2132 (O_2132,N_19970,N_19793);
nand UO_2133 (O_2133,N_19847,N_19953);
and UO_2134 (O_2134,N_19895,N_19754);
nor UO_2135 (O_2135,N_19879,N_19821);
or UO_2136 (O_2136,N_19941,N_19836);
nand UO_2137 (O_2137,N_19848,N_19981);
nand UO_2138 (O_2138,N_19961,N_19772);
or UO_2139 (O_2139,N_19766,N_19966);
nor UO_2140 (O_2140,N_19897,N_19905);
and UO_2141 (O_2141,N_19987,N_19786);
nand UO_2142 (O_2142,N_19894,N_19799);
xnor UO_2143 (O_2143,N_19880,N_19801);
nand UO_2144 (O_2144,N_19934,N_19962);
xnor UO_2145 (O_2145,N_19756,N_19894);
nor UO_2146 (O_2146,N_19975,N_19878);
nor UO_2147 (O_2147,N_19785,N_19936);
or UO_2148 (O_2148,N_19860,N_19956);
and UO_2149 (O_2149,N_19957,N_19815);
or UO_2150 (O_2150,N_19940,N_19867);
nor UO_2151 (O_2151,N_19886,N_19787);
xnor UO_2152 (O_2152,N_19929,N_19886);
and UO_2153 (O_2153,N_19817,N_19967);
xor UO_2154 (O_2154,N_19803,N_19800);
nor UO_2155 (O_2155,N_19884,N_19786);
xnor UO_2156 (O_2156,N_19943,N_19870);
nand UO_2157 (O_2157,N_19763,N_19766);
xnor UO_2158 (O_2158,N_19827,N_19893);
nand UO_2159 (O_2159,N_19828,N_19835);
nand UO_2160 (O_2160,N_19768,N_19957);
nor UO_2161 (O_2161,N_19776,N_19923);
nand UO_2162 (O_2162,N_19768,N_19808);
and UO_2163 (O_2163,N_19782,N_19927);
xnor UO_2164 (O_2164,N_19887,N_19987);
and UO_2165 (O_2165,N_19834,N_19979);
or UO_2166 (O_2166,N_19872,N_19870);
and UO_2167 (O_2167,N_19821,N_19824);
nand UO_2168 (O_2168,N_19811,N_19789);
nor UO_2169 (O_2169,N_19856,N_19885);
xnor UO_2170 (O_2170,N_19825,N_19977);
and UO_2171 (O_2171,N_19980,N_19812);
nor UO_2172 (O_2172,N_19954,N_19854);
or UO_2173 (O_2173,N_19821,N_19757);
and UO_2174 (O_2174,N_19935,N_19999);
and UO_2175 (O_2175,N_19796,N_19752);
nand UO_2176 (O_2176,N_19845,N_19989);
or UO_2177 (O_2177,N_19857,N_19974);
or UO_2178 (O_2178,N_19813,N_19823);
or UO_2179 (O_2179,N_19932,N_19988);
and UO_2180 (O_2180,N_19833,N_19928);
nor UO_2181 (O_2181,N_19753,N_19815);
and UO_2182 (O_2182,N_19863,N_19908);
nand UO_2183 (O_2183,N_19811,N_19974);
nor UO_2184 (O_2184,N_19876,N_19849);
nor UO_2185 (O_2185,N_19891,N_19911);
nand UO_2186 (O_2186,N_19758,N_19900);
nor UO_2187 (O_2187,N_19837,N_19937);
and UO_2188 (O_2188,N_19859,N_19755);
nand UO_2189 (O_2189,N_19909,N_19769);
nor UO_2190 (O_2190,N_19885,N_19770);
nand UO_2191 (O_2191,N_19950,N_19775);
xor UO_2192 (O_2192,N_19776,N_19994);
nor UO_2193 (O_2193,N_19989,N_19802);
nor UO_2194 (O_2194,N_19754,N_19860);
xnor UO_2195 (O_2195,N_19843,N_19884);
nor UO_2196 (O_2196,N_19876,N_19944);
xnor UO_2197 (O_2197,N_19865,N_19954);
xor UO_2198 (O_2198,N_19994,N_19990);
xor UO_2199 (O_2199,N_19857,N_19828);
nor UO_2200 (O_2200,N_19753,N_19817);
or UO_2201 (O_2201,N_19885,N_19954);
nand UO_2202 (O_2202,N_19811,N_19927);
nand UO_2203 (O_2203,N_19916,N_19974);
nand UO_2204 (O_2204,N_19868,N_19929);
or UO_2205 (O_2205,N_19787,N_19752);
and UO_2206 (O_2206,N_19992,N_19948);
nand UO_2207 (O_2207,N_19998,N_19944);
nor UO_2208 (O_2208,N_19781,N_19797);
or UO_2209 (O_2209,N_19782,N_19997);
xnor UO_2210 (O_2210,N_19875,N_19978);
nor UO_2211 (O_2211,N_19905,N_19772);
nor UO_2212 (O_2212,N_19796,N_19805);
xnor UO_2213 (O_2213,N_19935,N_19914);
or UO_2214 (O_2214,N_19753,N_19941);
nand UO_2215 (O_2215,N_19929,N_19803);
and UO_2216 (O_2216,N_19967,N_19921);
and UO_2217 (O_2217,N_19822,N_19759);
xnor UO_2218 (O_2218,N_19913,N_19774);
nand UO_2219 (O_2219,N_19880,N_19950);
nand UO_2220 (O_2220,N_19792,N_19770);
xor UO_2221 (O_2221,N_19803,N_19924);
nand UO_2222 (O_2222,N_19902,N_19930);
or UO_2223 (O_2223,N_19801,N_19863);
nor UO_2224 (O_2224,N_19778,N_19994);
xnor UO_2225 (O_2225,N_19919,N_19890);
nor UO_2226 (O_2226,N_19893,N_19883);
and UO_2227 (O_2227,N_19955,N_19873);
and UO_2228 (O_2228,N_19756,N_19861);
nor UO_2229 (O_2229,N_19964,N_19842);
xor UO_2230 (O_2230,N_19772,N_19769);
and UO_2231 (O_2231,N_19974,N_19806);
xor UO_2232 (O_2232,N_19850,N_19802);
and UO_2233 (O_2233,N_19949,N_19915);
and UO_2234 (O_2234,N_19939,N_19920);
xor UO_2235 (O_2235,N_19833,N_19948);
nand UO_2236 (O_2236,N_19860,N_19940);
nor UO_2237 (O_2237,N_19839,N_19957);
nand UO_2238 (O_2238,N_19991,N_19959);
nor UO_2239 (O_2239,N_19799,N_19767);
nand UO_2240 (O_2240,N_19882,N_19935);
or UO_2241 (O_2241,N_19765,N_19776);
or UO_2242 (O_2242,N_19935,N_19951);
xnor UO_2243 (O_2243,N_19816,N_19886);
xor UO_2244 (O_2244,N_19753,N_19919);
and UO_2245 (O_2245,N_19939,N_19770);
nor UO_2246 (O_2246,N_19895,N_19984);
xor UO_2247 (O_2247,N_19921,N_19900);
and UO_2248 (O_2248,N_19976,N_19969);
and UO_2249 (O_2249,N_19829,N_19879);
xor UO_2250 (O_2250,N_19772,N_19927);
nor UO_2251 (O_2251,N_19822,N_19831);
nor UO_2252 (O_2252,N_19817,N_19858);
and UO_2253 (O_2253,N_19800,N_19764);
nand UO_2254 (O_2254,N_19817,N_19809);
and UO_2255 (O_2255,N_19943,N_19827);
and UO_2256 (O_2256,N_19992,N_19798);
nand UO_2257 (O_2257,N_19815,N_19904);
and UO_2258 (O_2258,N_19922,N_19928);
xor UO_2259 (O_2259,N_19849,N_19890);
xnor UO_2260 (O_2260,N_19986,N_19905);
and UO_2261 (O_2261,N_19903,N_19865);
or UO_2262 (O_2262,N_19975,N_19890);
nand UO_2263 (O_2263,N_19841,N_19765);
or UO_2264 (O_2264,N_19918,N_19903);
or UO_2265 (O_2265,N_19756,N_19934);
nor UO_2266 (O_2266,N_19837,N_19765);
and UO_2267 (O_2267,N_19968,N_19920);
nand UO_2268 (O_2268,N_19922,N_19976);
nor UO_2269 (O_2269,N_19833,N_19766);
nor UO_2270 (O_2270,N_19948,N_19888);
nor UO_2271 (O_2271,N_19788,N_19842);
nor UO_2272 (O_2272,N_19833,N_19930);
or UO_2273 (O_2273,N_19896,N_19796);
xor UO_2274 (O_2274,N_19860,N_19783);
nor UO_2275 (O_2275,N_19964,N_19895);
nand UO_2276 (O_2276,N_19902,N_19969);
xnor UO_2277 (O_2277,N_19992,N_19785);
nor UO_2278 (O_2278,N_19912,N_19782);
nor UO_2279 (O_2279,N_19848,N_19958);
xnor UO_2280 (O_2280,N_19993,N_19881);
or UO_2281 (O_2281,N_19971,N_19861);
nor UO_2282 (O_2282,N_19949,N_19796);
nor UO_2283 (O_2283,N_19898,N_19911);
nor UO_2284 (O_2284,N_19940,N_19932);
and UO_2285 (O_2285,N_19848,N_19969);
nand UO_2286 (O_2286,N_19765,N_19960);
nor UO_2287 (O_2287,N_19844,N_19902);
or UO_2288 (O_2288,N_19872,N_19958);
nor UO_2289 (O_2289,N_19835,N_19918);
xor UO_2290 (O_2290,N_19977,N_19826);
nand UO_2291 (O_2291,N_19792,N_19782);
nor UO_2292 (O_2292,N_19818,N_19789);
nand UO_2293 (O_2293,N_19988,N_19874);
and UO_2294 (O_2294,N_19830,N_19801);
nand UO_2295 (O_2295,N_19959,N_19857);
xor UO_2296 (O_2296,N_19953,N_19881);
and UO_2297 (O_2297,N_19889,N_19987);
nor UO_2298 (O_2298,N_19830,N_19871);
xnor UO_2299 (O_2299,N_19881,N_19829);
nand UO_2300 (O_2300,N_19966,N_19856);
xor UO_2301 (O_2301,N_19973,N_19864);
or UO_2302 (O_2302,N_19805,N_19879);
or UO_2303 (O_2303,N_19946,N_19853);
xnor UO_2304 (O_2304,N_19972,N_19963);
nand UO_2305 (O_2305,N_19827,N_19777);
nand UO_2306 (O_2306,N_19782,N_19794);
xnor UO_2307 (O_2307,N_19948,N_19769);
or UO_2308 (O_2308,N_19807,N_19787);
nor UO_2309 (O_2309,N_19961,N_19774);
xor UO_2310 (O_2310,N_19815,N_19843);
and UO_2311 (O_2311,N_19958,N_19771);
nor UO_2312 (O_2312,N_19815,N_19795);
and UO_2313 (O_2313,N_19914,N_19790);
xnor UO_2314 (O_2314,N_19985,N_19947);
nor UO_2315 (O_2315,N_19977,N_19981);
and UO_2316 (O_2316,N_19764,N_19786);
nand UO_2317 (O_2317,N_19882,N_19872);
and UO_2318 (O_2318,N_19972,N_19858);
nor UO_2319 (O_2319,N_19987,N_19956);
nor UO_2320 (O_2320,N_19873,N_19893);
and UO_2321 (O_2321,N_19933,N_19925);
nand UO_2322 (O_2322,N_19755,N_19857);
and UO_2323 (O_2323,N_19965,N_19918);
nor UO_2324 (O_2324,N_19762,N_19824);
or UO_2325 (O_2325,N_19760,N_19892);
or UO_2326 (O_2326,N_19972,N_19911);
and UO_2327 (O_2327,N_19833,N_19851);
xnor UO_2328 (O_2328,N_19762,N_19847);
or UO_2329 (O_2329,N_19961,N_19862);
nand UO_2330 (O_2330,N_19758,N_19898);
or UO_2331 (O_2331,N_19751,N_19947);
xor UO_2332 (O_2332,N_19825,N_19944);
nor UO_2333 (O_2333,N_19896,N_19825);
or UO_2334 (O_2334,N_19908,N_19929);
or UO_2335 (O_2335,N_19987,N_19978);
and UO_2336 (O_2336,N_19760,N_19915);
nand UO_2337 (O_2337,N_19892,N_19872);
nor UO_2338 (O_2338,N_19766,N_19953);
and UO_2339 (O_2339,N_19892,N_19866);
nor UO_2340 (O_2340,N_19883,N_19791);
or UO_2341 (O_2341,N_19977,N_19947);
and UO_2342 (O_2342,N_19999,N_19763);
nand UO_2343 (O_2343,N_19876,N_19970);
nor UO_2344 (O_2344,N_19758,N_19902);
or UO_2345 (O_2345,N_19983,N_19811);
and UO_2346 (O_2346,N_19823,N_19965);
and UO_2347 (O_2347,N_19933,N_19926);
or UO_2348 (O_2348,N_19916,N_19803);
xor UO_2349 (O_2349,N_19995,N_19759);
nor UO_2350 (O_2350,N_19770,N_19791);
or UO_2351 (O_2351,N_19859,N_19871);
nand UO_2352 (O_2352,N_19937,N_19796);
xnor UO_2353 (O_2353,N_19774,N_19782);
xor UO_2354 (O_2354,N_19888,N_19890);
nor UO_2355 (O_2355,N_19859,N_19769);
nand UO_2356 (O_2356,N_19877,N_19895);
nand UO_2357 (O_2357,N_19983,N_19962);
nand UO_2358 (O_2358,N_19930,N_19908);
or UO_2359 (O_2359,N_19959,N_19901);
or UO_2360 (O_2360,N_19772,N_19912);
xor UO_2361 (O_2361,N_19790,N_19894);
or UO_2362 (O_2362,N_19910,N_19758);
and UO_2363 (O_2363,N_19998,N_19793);
nand UO_2364 (O_2364,N_19926,N_19835);
xor UO_2365 (O_2365,N_19934,N_19908);
or UO_2366 (O_2366,N_19811,N_19861);
nand UO_2367 (O_2367,N_19982,N_19772);
nand UO_2368 (O_2368,N_19920,N_19991);
and UO_2369 (O_2369,N_19999,N_19857);
and UO_2370 (O_2370,N_19992,N_19804);
nand UO_2371 (O_2371,N_19912,N_19817);
and UO_2372 (O_2372,N_19835,N_19752);
and UO_2373 (O_2373,N_19867,N_19894);
or UO_2374 (O_2374,N_19886,N_19901);
and UO_2375 (O_2375,N_19853,N_19809);
and UO_2376 (O_2376,N_19907,N_19995);
and UO_2377 (O_2377,N_19821,N_19976);
nor UO_2378 (O_2378,N_19831,N_19796);
xor UO_2379 (O_2379,N_19896,N_19851);
or UO_2380 (O_2380,N_19808,N_19888);
and UO_2381 (O_2381,N_19840,N_19901);
nor UO_2382 (O_2382,N_19860,N_19762);
and UO_2383 (O_2383,N_19859,N_19764);
nand UO_2384 (O_2384,N_19979,N_19864);
nor UO_2385 (O_2385,N_19896,N_19959);
nor UO_2386 (O_2386,N_19997,N_19853);
nand UO_2387 (O_2387,N_19833,N_19986);
xnor UO_2388 (O_2388,N_19939,N_19928);
nand UO_2389 (O_2389,N_19843,N_19844);
xor UO_2390 (O_2390,N_19888,N_19916);
xor UO_2391 (O_2391,N_19903,N_19985);
or UO_2392 (O_2392,N_19967,N_19897);
nand UO_2393 (O_2393,N_19867,N_19992);
or UO_2394 (O_2394,N_19907,N_19922);
xnor UO_2395 (O_2395,N_19990,N_19841);
and UO_2396 (O_2396,N_19777,N_19757);
and UO_2397 (O_2397,N_19803,N_19893);
nor UO_2398 (O_2398,N_19962,N_19833);
or UO_2399 (O_2399,N_19863,N_19979);
nand UO_2400 (O_2400,N_19784,N_19802);
and UO_2401 (O_2401,N_19835,N_19956);
and UO_2402 (O_2402,N_19931,N_19878);
nor UO_2403 (O_2403,N_19904,N_19779);
nor UO_2404 (O_2404,N_19751,N_19803);
xnor UO_2405 (O_2405,N_19755,N_19902);
xnor UO_2406 (O_2406,N_19971,N_19847);
or UO_2407 (O_2407,N_19849,N_19872);
xnor UO_2408 (O_2408,N_19917,N_19837);
and UO_2409 (O_2409,N_19824,N_19952);
xor UO_2410 (O_2410,N_19758,N_19810);
nor UO_2411 (O_2411,N_19836,N_19958);
or UO_2412 (O_2412,N_19849,N_19819);
nand UO_2413 (O_2413,N_19859,N_19991);
nand UO_2414 (O_2414,N_19951,N_19884);
nor UO_2415 (O_2415,N_19786,N_19879);
nor UO_2416 (O_2416,N_19820,N_19993);
and UO_2417 (O_2417,N_19784,N_19905);
xnor UO_2418 (O_2418,N_19847,N_19942);
xnor UO_2419 (O_2419,N_19867,N_19972);
nand UO_2420 (O_2420,N_19859,N_19760);
and UO_2421 (O_2421,N_19841,N_19843);
and UO_2422 (O_2422,N_19994,N_19870);
nand UO_2423 (O_2423,N_19884,N_19852);
and UO_2424 (O_2424,N_19834,N_19851);
nor UO_2425 (O_2425,N_19834,N_19765);
or UO_2426 (O_2426,N_19825,N_19875);
xnor UO_2427 (O_2427,N_19943,N_19934);
or UO_2428 (O_2428,N_19766,N_19951);
xnor UO_2429 (O_2429,N_19901,N_19954);
xor UO_2430 (O_2430,N_19873,N_19861);
and UO_2431 (O_2431,N_19789,N_19795);
nor UO_2432 (O_2432,N_19985,N_19872);
or UO_2433 (O_2433,N_19872,N_19823);
xor UO_2434 (O_2434,N_19937,N_19954);
nor UO_2435 (O_2435,N_19873,N_19756);
or UO_2436 (O_2436,N_19913,N_19902);
nand UO_2437 (O_2437,N_19854,N_19811);
xor UO_2438 (O_2438,N_19881,N_19930);
nor UO_2439 (O_2439,N_19932,N_19805);
nor UO_2440 (O_2440,N_19961,N_19921);
nand UO_2441 (O_2441,N_19868,N_19845);
nand UO_2442 (O_2442,N_19783,N_19844);
and UO_2443 (O_2443,N_19820,N_19949);
and UO_2444 (O_2444,N_19750,N_19823);
nor UO_2445 (O_2445,N_19764,N_19944);
nor UO_2446 (O_2446,N_19884,N_19991);
and UO_2447 (O_2447,N_19815,N_19773);
xor UO_2448 (O_2448,N_19897,N_19795);
and UO_2449 (O_2449,N_19820,N_19859);
nand UO_2450 (O_2450,N_19830,N_19864);
nand UO_2451 (O_2451,N_19908,N_19989);
nand UO_2452 (O_2452,N_19954,N_19780);
nand UO_2453 (O_2453,N_19846,N_19976);
xnor UO_2454 (O_2454,N_19936,N_19768);
nand UO_2455 (O_2455,N_19971,N_19867);
nor UO_2456 (O_2456,N_19754,N_19898);
or UO_2457 (O_2457,N_19925,N_19943);
xnor UO_2458 (O_2458,N_19922,N_19876);
nand UO_2459 (O_2459,N_19992,N_19904);
and UO_2460 (O_2460,N_19979,N_19857);
nand UO_2461 (O_2461,N_19907,N_19825);
or UO_2462 (O_2462,N_19924,N_19821);
nand UO_2463 (O_2463,N_19970,N_19968);
xnor UO_2464 (O_2464,N_19971,N_19838);
xor UO_2465 (O_2465,N_19924,N_19906);
and UO_2466 (O_2466,N_19908,N_19913);
nand UO_2467 (O_2467,N_19884,N_19959);
xor UO_2468 (O_2468,N_19788,N_19771);
xnor UO_2469 (O_2469,N_19876,N_19930);
and UO_2470 (O_2470,N_19937,N_19982);
nand UO_2471 (O_2471,N_19901,N_19999);
nor UO_2472 (O_2472,N_19948,N_19938);
or UO_2473 (O_2473,N_19899,N_19958);
xor UO_2474 (O_2474,N_19964,N_19865);
or UO_2475 (O_2475,N_19916,N_19996);
or UO_2476 (O_2476,N_19878,N_19918);
nand UO_2477 (O_2477,N_19954,N_19825);
and UO_2478 (O_2478,N_19943,N_19883);
and UO_2479 (O_2479,N_19822,N_19810);
nor UO_2480 (O_2480,N_19824,N_19857);
and UO_2481 (O_2481,N_19873,N_19923);
nor UO_2482 (O_2482,N_19858,N_19759);
or UO_2483 (O_2483,N_19959,N_19995);
nand UO_2484 (O_2484,N_19952,N_19754);
and UO_2485 (O_2485,N_19997,N_19892);
xor UO_2486 (O_2486,N_19800,N_19753);
xor UO_2487 (O_2487,N_19931,N_19839);
xor UO_2488 (O_2488,N_19972,N_19951);
and UO_2489 (O_2489,N_19795,N_19849);
nor UO_2490 (O_2490,N_19767,N_19826);
nor UO_2491 (O_2491,N_19891,N_19886);
nand UO_2492 (O_2492,N_19801,N_19819);
or UO_2493 (O_2493,N_19967,N_19795);
nor UO_2494 (O_2494,N_19916,N_19757);
nor UO_2495 (O_2495,N_19945,N_19908);
xor UO_2496 (O_2496,N_19997,N_19816);
nor UO_2497 (O_2497,N_19986,N_19943);
and UO_2498 (O_2498,N_19803,N_19980);
xor UO_2499 (O_2499,N_19855,N_19992);
endmodule