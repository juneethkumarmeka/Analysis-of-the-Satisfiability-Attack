module basic_1000_10000_1500_4_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_700,In_955);
nor U1 (N_1,In_637,In_361);
or U2 (N_2,In_522,In_925);
and U3 (N_3,In_885,In_452);
nor U4 (N_4,In_870,In_586);
nand U5 (N_5,In_904,In_158);
xnor U6 (N_6,In_227,In_910);
or U7 (N_7,In_430,In_901);
nor U8 (N_8,In_839,In_914);
and U9 (N_9,In_105,In_622);
nor U10 (N_10,In_768,In_36);
nor U11 (N_11,In_970,In_296);
xnor U12 (N_12,In_916,In_936);
nand U13 (N_13,In_715,In_193);
nand U14 (N_14,In_370,In_462);
nand U15 (N_15,In_742,In_170);
nand U16 (N_16,In_770,In_849);
nor U17 (N_17,In_418,In_345);
nand U18 (N_18,In_859,In_927);
or U19 (N_19,In_29,In_226);
xor U20 (N_20,In_455,In_617);
nor U21 (N_21,In_315,In_539);
nor U22 (N_22,In_15,In_546);
xnor U23 (N_23,In_640,In_777);
xnor U24 (N_24,In_673,In_479);
nand U25 (N_25,In_393,In_188);
xnor U26 (N_26,In_699,In_271);
xnor U27 (N_27,In_671,In_446);
nor U28 (N_28,In_390,In_367);
or U29 (N_29,In_391,In_382);
xor U30 (N_30,In_667,In_864);
xor U31 (N_31,In_93,In_938);
or U32 (N_32,In_662,In_820);
nand U33 (N_33,In_248,In_114);
and U34 (N_34,In_596,In_396);
xnor U35 (N_35,In_273,In_620);
nand U36 (N_36,In_74,In_321);
nor U37 (N_37,In_674,In_965);
nand U38 (N_38,In_990,In_817);
xnor U39 (N_39,In_894,In_77);
or U40 (N_40,In_854,In_788);
xnor U41 (N_41,In_184,In_363);
nand U42 (N_42,In_364,In_792);
or U43 (N_43,In_497,In_574);
nor U44 (N_44,In_134,In_840);
nor U45 (N_45,In_565,In_723);
and U46 (N_46,In_51,In_569);
nand U47 (N_47,In_576,In_478);
or U48 (N_48,In_948,In_877);
xor U49 (N_49,In_317,In_692);
xnor U50 (N_50,In_991,In_567);
or U51 (N_51,In_313,In_174);
nor U52 (N_52,In_491,In_428);
nor U53 (N_53,In_504,In_39);
nand U54 (N_54,In_470,In_500);
nand U55 (N_55,In_719,In_215);
xor U56 (N_56,In_848,In_985);
and U57 (N_57,In_149,In_251);
nand U58 (N_58,In_694,In_59);
nor U59 (N_59,In_460,In_505);
and U60 (N_60,In_49,In_544);
nand U61 (N_61,In_703,In_453);
and U62 (N_62,In_300,In_454);
and U63 (N_63,In_579,In_526);
nand U64 (N_64,In_135,In_809);
nand U65 (N_65,In_638,In_766);
nand U66 (N_66,In_443,In_228);
xnor U67 (N_67,In_989,In_326);
nand U68 (N_68,In_536,In_297);
or U69 (N_69,In_844,In_767);
nand U70 (N_70,In_305,In_669);
nand U71 (N_71,In_590,In_385);
and U72 (N_72,In_535,In_434);
nor U73 (N_73,In_823,In_529);
nor U74 (N_74,In_55,In_431);
xnor U75 (N_75,In_775,In_868);
nand U76 (N_76,In_38,In_758);
xnor U77 (N_77,In_352,In_132);
or U78 (N_78,In_162,In_451);
and U79 (N_79,In_912,In_474);
or U80 (N_80,In_639,In_140);
and U81 (N_81,In_90,In_69);
nand U82 (N_82,In_577,In_436);
xor U83 (N_83,In_602,In_865);
nand U84 (N_84,In_392,In_138);
or U85 (N_85,In_724,In_249);
xnor U86 (N_86,In_371,In_102);
xnor U87 (N_87,In_561,In_164);
xnor U88 (N_88,In_483,In_882);
xnor U89 (N_89,In_861,In_879);
or U90 (N_90,In_730,In_616);
nor U91 (N_91,In_769,In_66);
and U92 (N_92,In_476,In_417);
nor U93 (N_93,In_112,In_624);
nor U94 (N_94,In_83,In_172);
nand U95 (N_95,In_759,In_900);
or U96 (N_96,In_855,In_626);
xnor U97 (N_97,In_270,In_498);
or U98 (N_98,In_33,In_757);
nand U99 (N_99,In_869,In_377);
nor U100 (N_100,In_922,In_963);
nand U101 (N_101,In_531,In_24);
and U102 (N_102,In_409,In_661);
nand U103 (N_103,In_503,In_266);
nand U104 (N_104,In_813,In_182);
or U105 (N_105,In_831,In_276);
or U106 (N_106,In_580,In_22);
or U107 (N_107,In_939,In_427);
xnor U108 (N_108,In_27,In_736);
nor U109 (N_109,In_48,In_772);
xnor U110 (N_110,In_347,In_212);
and U111 (N_111,In_492,In_816);
nand U112 (N_112,In_244,In_945);
nand U113 (N_113,In_304,In_294);
nor U114 (N_114,In_734,In_560);
nand U115 (N_115,In_549,In_629);
or U116 (N_116,In_89,In_225);
and U117 (N_117,In_686,In_623);
and U118 (N_118,In_255,In_309);
or U119 (N_119,In_201,In_136);
xor U120 (N_120,In_538,In_811);
nand U121 (N_121,In_510,In_630);
nand U122 (N_122,In_883,In_429);
and U123 (N_123,In_433,In_835);
nor U124 (N_124,In_359,In_310);
and U125 (N_125,In_977,In_269);
nor U126 (N_126,In_5,In_351);
nand U127 (N_127,In_941,In_80);
and U128 (N_128,In_12,In_973);
xnor U129 (N_129,In_113,In_252);
or U130 (N_130,In_987,In_913);
nor U131 (N_131,In_44,In_950);
and U132 (N_132,In_964,In_87);
xor U133 (N_133,In_484,In_808);
xnor U134 (N_134,In_979,In_204);
or U135 (N_135,In_0,In_378);
nand U136 (N_136,In_655,In_488);
and U137 (N_137,In_551,In_822);
nor U138 (N_138,In_717,In_889);
and U139 (N_139,In_402,In_461);
or U140 (N_140,In_250,In_75);
and U141 (N_141,In_415,In_599);
nand U142 (N_142,In_236,In_895);
nor U143 (N_143,In_502,In_383);
or U144 (N_144,In_63,In_600);
nand U145 (N_145,In_85,In_545);
nor U146 (N_146,In_125,In_718);
nor U147 (N_147,In_40,In_419);
and U148 (N_148,In_70,In_542);
nor U149 (N_149,In_668,In_918);
nand U150 (N_150,In_217,In_589);
xor U151 (N_151,In_103,In_258);
nor U152 (N_152,In_106,In_46);
nand U153 (N_153,In_235,In_288);
and U154 (N_154,In_693,In_110);
nand U155 (N_155,In_156,In_108);
xor U156 (N_156,In_550,In_421);
and U157 (N_157,In_53,In_814);
nand U158 (N_158,In_213,In_776);
xor U159 (N_159,In_986,In_389);
and U160 (N_160,In_173,In_76);
and U161 (N_161,In_521,In_928);
or U162 (N_162,In_711,In_400);
nor U163 (N_163,In_548,In_358);
nand U164 (N_164,In_760,In_468);
nor U165 (N_165,In_657,In_564);
or U166 (N_166,In_96,In_971);
or U167 (N_167,In_17,In_680);
xor U168 (N_168,In_672,In_118);
and U169 (N_169,In_357,In_122);
and U170 (N_170,In_967,In_292);
or U171 (N_171,In_159,In_745);
nor U172 (N_172,In_449,In_802);
or U173 (N_173,In_954,In_641);
or U174 (N_174,In_805,In_993);
nor U175 (N_175,In_903,In_61);
nor U176 (N_176,In_525,In_314);
or U177 (N_177,In_785,In_746);
and U178 (N_178,In_395,In_853);
nor U179 (N_179,In_563,In_341);
or U180 (N_180,In_501,In_26);
nor U181 (N_181,In_308,In_681);
nand U182 (N_182,In_588,In_219);
or U183 (N_183,In_841,In_123);
nor U184 (N_184,In_19,In_253);
or U185 (N_185,In_243,In_239);
and U186 (N_186,In_482,In_54);
and U187 (N_187,In_177,In_131);
nand U188 (N_188,In_665,In_790);
nor U189 (N_189,In_334,In_753);
nor U190 (N_190,In_685,In_73);
or U191 (N_191,In_917,In_978);
nand U192 (N_192,In_603,In_871);
xnor U193 (N_193,In_604,In_984);
or U194 (N_194,In_755,In_435);
and U195 (N_195,In_793,In_824);
nor U196 (N_196,In_553,In_475);
xor U197 (N_197,In_71,In_466);
or U198 (N_198,In_163,In_1);
or U199 (N_199,In_6,In_423);
xor U200 (N_200,In_58,In_591);
nand U201 (N_201,In_56,In_151);
or U202 (N_202,In_952,In_930);
and U203 (N_203,In_789,In_860);
nand U204 (N_204,In_166,In_981);
xor U205 (N_205,In_884,In_289);
xor U206 (N_206,In_198,In_513);
xor U207 (N_207,In_473,In_797);
xnor U208 (N_208,In_281,In_306);
xor U209 (N_209,In_232,In_675);
nor U210 (N_210,In_448,In_739);
or U211 (N_211,In_330,In_366);
nor U212 (N_212,In_908,In_202);
nand U213 (N_213,In_495,In_842);
xnor U214 (N_214,In_893,In_931);
xor U215 (N_215,In_221,In_456);
nand U216 (N_216,In_187,In_552);
xor U217 (N_217,In_615,In_999);
xor U218 (N_218,In_799,In_386);
and U219 (N_219,In_688,In_146);
nand U220 (N_220,In_994,In_969);
nand U221 (N_221,In_459,In_741);
nand U222 (N_222,In_836,In_23);
xnor U223 (N_223,In_856,In_279);
and U224 (N_224,In_196,In_878);
nand U225 (N_225,In_101,In_594);
nor U226 (N_226,In_906,In_319);
or U227 (N_227,In_190,In_740);
and U228 (N_228,In_335,In_830);
nand U229 (N_229,In_566,In_690);
xor U230 (N_230,In_515,In_935);
and U231 (N_231,In_631,In_115);
or U232 (N_232,In_763,In_618);
nand U233 (N_233,In_988,In_783);
nand U234 (N_234,In_647,In_547);
nand U235 (N_235,In_958,In_157);
and U236 (N_236,In_169,In_832);
or U237 (N_237,In_11,In_465);
and U238 (N_238,In_154,In_205);
and U239 (N_239,In_178,In_88);
xor U240 (N_240,In_422,In_833);
or U241 (N_241,In_278,In_67);
or U242 (N_242,In_41,In_731);
xnor U243 (N_243,In_929,In_485);
and U244 (N_244,In_150,In_749);
or U245 (N_245,In_274,In_220);
or U246 (N_246,In_982,In_339);
and U247 (N_247,In_129,In_295);
xor U248 (N_248,In_152,In_408);
and U249 (N_249,In_233,In_713);
nand U250 (N_250,In_242,In_35);
and U251 (N_251,In_541,In_815);
nand U252 (N_252,In_354,In_593);
or U253 (N_253,In_953,In_705);
nand U254 (N_254,In_571,In_506);
and U255 (N_255,In_280,In_450);
xnor U256 (N_256,In_921,In_712);
nor U257 (N_257,In_206,In_773);
xnor U258 (N_258,In_168,In_956);
xnor U259 (N_259,In_704,In_818);
nor U260 (N_260,In_336,In_915);
nand U261 (N_261,In_237,In_99);
nand U262 (N_262,In_527,In_902);
or U263 (N_263,In_416,In_961);
xnor U264 (N_264,In_530,In_381);
nand U265 (N_265,In_645,In_697);
nor U266 (N_266,In_2,In_682);
or U267 (N_267,In_892,In_707);
or U268 (N_268,In_207,In_838);
and U269 (N_269,In_951,In_369);
or U270 (N_270,In_329,In_293);
nand U271 (N_271,In_562,In_720);
xnor U272 (N_272,In_520,In_656);
nand U273 (N_273,In_881,In_303);
xor U274 (N_274,In_607,In_86);
nand U275 (N_275,In_643,In_781);
nand U276 (N_276,In_282,In_494);
nor U277 (N_277,In_14,In_651);
nor U278 (N_278,In_664,In_160);
or U279 (N_279,In_998,In_683);
nand U280 (N_280,In_896,In_469);
nor U281 (N_281,In_866,In_437);
xnor U282 (N_282,In_532,In_947);
xor U283 (N_283,In_934,In_980);
xnor U284 (N_284,In_307,In_302);
xnor U285 (N_285,In_209,In_81);
nand U286 (N_286,In_199,In_612);
xor U287 (N_287,In_743,In_432);
nand U288 (N_288,In_283,In_570);
or U289 (N_289,In_666,In_897);
or U290 (N_290,In_846,In_144);
nand U291 (N_291,In_890,In_540);
and U292 (N_292,In_905,In_787);
or U293 (N_293,In_65,In_179);
xor U294 (N_294,In_62,In_50);
and U295 (N_295,In_353,In_175);
xor U296 (N_296,In_966,In_778);
and U297 (N_297,In_147,In_621);
or U298 (N_298,In_722,In_489);
nand U299 (N_299,In_197,In_441);
and U300 (N_300,In_13,In_124);
xor U301 (N_301,In_148,In_25);
nor U302 (N_302,In_275,In_609);
nand U303 (N_303,In_725,In_176);
nand U304 (N_304,In_234,In_957);
and U305 (N_305,In_333,In_750);
and U306 (N_306,In_874,In_9);
nand U307 (N_307,In_343,In_346);
nand U308 (N_308,In_677,In_262);
or U309 (N_309,In_272,In_754);
and U310 (N_310,In_43,In_405);
xnor U311 (N_311,In_937,In_764);
or U312 (N_312,In_509,In_97);
or U313 (N_313,In_791,In_208);
nand U314 (N_314,In_394,In_327);
or U315 (N_315,In_684,In_554);
xor U316 (N_316,In_133,In_907);
nand U317 (N_317,In_285,In_888);
nand U318 (N_318,In_803,In_246);
or U319 (N_319,In_825,In_194);
nand U320 (N_320,In_267,In_181);
xor U321 (N_321,In_399,In_557);
nor U322 (N_322,In_658,In_299);
nor U323 (N_323,In_847,In_57);
nor U324 (N_324,In_652,In_752);
nor U325 (N_325,In_398,In_404);
and U326 (N_326,In_128,In_349);
xor U327 (N_327,In_47,In_632);
or U328 (N_328,In_568,In_642);
nor U329 (N_329,In_200,In_247);
xor U330 (N_330,In_397,In_649);
xor U331 (N_331,In_932,In_804);
nor U332 (N_332,In_748,In_20);
or U333 (N_333,In_126,In_287);
nand U334 (N_334,In_635,In_801);
or U335 (N_335,In_942,In_241);
nand U336 (N_336,In_944,In_338);
and U337 (N_337,In_876,In_425);
nor U338 (N_338,In_862,In_872);
and U339 (N_339,In_45,In_438);
or U340 (N_340,In_121,In_143);
xor U341 (N_341,In_780,In_362);
nor U342 (N_342,In_614,In_880);
nand U343 (N_343,In_284,In_30);
xor U344 (N_344,In_611,In_414);
nor U345 (N_345,In_458,In_528);
nor U346 (N_346,In_442,In_139);
and U347 (N_347,In_507,In_16);
nor U348 (N_348,In_8,In_663);
nor U349 (N_349,In_222,In_898);
xor U350 (N_350,In_687,In_875);
or U351 (N_351,In_259,In_863);
or U352 (N_352,In_231,In_744);
or U353 (N_353,In_64,In_702);
xor U354 (N_354,In_411,In_608);
or U355 (N_355,In_606,In_650);
nor U356 (N_356,In_72,In_376);
or U357 (N_357,In_324,In_826);
xor U358 (N_358,In_779,In_678);
or U359 (N_359,In_845,In_762);
and U360 (N_360,In_486,In_32);
or U361 (N_361,In_737,In_192);
and U362 (N_362,In_514,In_534);
nand U363 (N_363,In_899,In_360);
nand U364 (N_364,In_613,In_95);
or U365 (N_365,In_245,In_130);
nand U366 (N_366,In_445,In_873);
xnor U367 (N_367,In_829,In_372);
nor U368 (N_368,In_229,In_240);
xor U369 (N_369,In_171,In_214);
nor U370 (N_370,In_496,In_924);
and U371 (N_371,In_426,In_867);
or U372 (N_372,In_940,In_806);
nand U373 (N_373,In_420,In_471);
nand U374 (N_374,In_379,In_508);
and U375 (N_375,In_595,In_518);
nand U376 (N_376,In_331,In_598);
or U377 (N_377,In_983,In_277);
nor U378 (N_378,In_765,In_583);
xnor U379 (N_379,In_412,In_256);
nand U380 (N_380,In_340,In_654);
xnor U381 (N_381,In_516,In_920);
nor U382 (N_382,In_582,In_524);
and U383 (N_383,In_111,In_633);
nand U384 (N_384,In_810,In_31);
or U385 (N_385,In_238,In_116);
xnor U386 (N_386,In_646,In_477);
nor U387 (N_387,In_344,In_365);
and U388 (N_388,In_676,In_78);
xnor U389 (N_389,In_79,In_943);
xor U390 (N_390,In_117,In_298);
xnor U391 (N_391,In_605,In_733);
nor U392 (N_392,In_726,In_578);
or U393 (N_393,In_68,In_493);
xor U394 (N_394,In_84,In_373);
nand U395 (N_395,In_992,In_328);
nor U396 (N_396,In_558,In_380);
or U397 (N_397,In_264,In_581);
or U398 (N_398,In_290,In_263);
xor U399 (N_399,In_843,In_537);
nor U400 (N_400,In_254,In_636);
nand U401 (N_401,In_210,In_301);
nand U402 (N_402,In_517,In_3);
and U403 (N_403,In_968,In_729);
xor U404 (N_404,In_751,In_960);
and U405 (N_405,In_974,In_721);
or U406 (N_406,In_10,In_710);
and U407 (N_407,In_782,In_962);
and U408 (N_408,In_559,In_996);
nand U409 (N_409,In_28,In_323);
xnor U410 (N_410,In_747,In_312);
nor U411 (N_411,In_698,In_909);
xnor U412 (N_412,In_104,In_52);
and U413 (N_413,In_342,In_679);
xnor U414 (N_414,In_857,In_191);
or U415 (N_415,In_774,In_186);
nand U416 (N_416,In_410,In_511);
nor U417 (N_417,In_320,In_512);
xnor U418 (N_418,In_689,In_127);
nor U419 (N_419,In_850,In_794);
and U420 (N_420,In_886,In_807);
nor U421 (N_421,In_42,In_738);
nand U422 (N_422,In_368,In_480);
or U423 (N_423,In_573,In_891);
or U424 (N_424,In_180,In_4);
xnor U425 (N_425,In_834,In_7);
nand U426 (N_426,In_837,In_523);
nand U427 (N_427,In_348,In_481);
or U428 (N_428,In_464,In_691);
xnor U429 (N_429,In_387,In_670);
nor U430 (N_430,In_555,In_644);
and U431 (N_431,In_660,In_141);
xor U432 (N_432,In_487,In_911);
or U433 (N_433,In_975,In_472);
and U434 (N_434,In_976,In_701);
nand U435 (N_435,In_355,In_919);
xnor U436 (N_436,In_318,In_107);
nand U437 (N_437,In_444,In_784);
xor U438 (N_438,In_796,In_519);
xnor U439 (N_439,In_424,In_619);
xnor U440 (N_440,In_21,In_332);
nand U441 (N_441,In_161,In_82);
nand U442 (N_442,In_634,In_735);
xnor U443 (N_443,In_972,In_627);
nand U444 (N_444,In_819,In_584);
xnor U445 (N_445,In_543,In_828);
or U446 (N_446,In_708,In_316);
and U447 (N_447,In_407,In_457);
and U448 (N_448,In_648,In_265);
or U449 (N_449,In_533,In_401);
nand U450 (N_450,In_575,In_167);
nor U451 (N_451,In_142,In_403);
xnor U452 (N_452,In_556,In_195);
and U453 (N_453,In_761,In_695);
nand U454 (N_454,In_933,In_356);
xnor U455 (N_455,In_812,In_311);
and U456 (N_456,In_463,In_800);
or U457 (N_457,In_261,In_727);
xnor U458 (N_458,In_291,In_572);
nand U459 (N_459,In_798,In_211);
nand U460 (N_460,In_587,In_145);
or U461 (N_461,In_659,In_447);
nor U462 (N_462,In_218,In_406);
and U463 (N_463,In_18,In_216);
and U464 (N_464,In_696,In_997);
xnor U465 (N_465,In_949,In_223);
or U466 (N_466,In_887,In_92);
xor U467 (N_467,In_337,In_467);
nor U468 (N_468,In_439,In_137);
nor U469 (N_469,In_786,In_375);
or U470 (N_470,In_268,In_490);
nor U471 (N_471,In_100,In_388);
and U472 (N_472,In_771,In_716);
xnor U473 (N_473,In_384,In_628);
or U474 (N_474,In_706,In_923);
or U475 (N_475,In_959,In_714);
nand U476 (N_476,In_827,In_585);
nor U477 (N_477,In_325,In_374);
nand U478 (N_478,In_946,In_153);
nor U479 (N_479,In_756,In_257);
or U480 (N_480,In_610,In_94);
nor U481 (N_481,In_499,In_165);
or U482 (N_482,In_260,In_185);
xnor U483 (N_483,In_795,In_34);
nand U484 (N_484,In_183,In_37);
nand U485 (N_485,In_625,In_91);
or U486 (N_486,In_224,In_120);
nor U487 (N_487,In_413,In_98);
xor U488 (N_488,In_732,In_852);
or U489 (N_489,In_858,In_155);
or U490 (N_490,In_601,In_60);
nor U491 (N_491,In_119,In_926);
or U492 (N_492,In_350,In_440);
xnor U493 (N_493,In_286,In_728);
or U494 (N_494,In_995,In_189);
and U495 (N_495,In_592,In_709);
nor U496 (N_496,In_821,In_109);
xnor U497 (N_497,In_851,In_322);
xor U498 (N_498,In_653,In_203);
xnor U499 (N_499,In_230,In_597);
nand U500 (N_500,In_21,In_924);
nor U501 (N_501,In_417,In_2);
and U502 (N_502,In_22,In_709);
nand U503 (N_503,In_505,In_335);
or U504 (N_504,In_519,In_663);
nand U505 (N_505,In_901,In_851);
nand U506 (N_506,In_848,In_816);
and U507 (N_507,In_317,In_234);
nand U508 (N_508,In_239,In_903);
nor U509 (N_509,In_328,In_371);
xor U510 (N_510,In_889,In_823);
or U511 (N_511,In_502,In_14);
nand U512 (N_512,In_4,In_247);
and U513 (N_513,In_460,In_647);
or U514 (N_514,In_894,In_737);
or U515 (N_515,In_890,In_889);
nor U516 (N_516,In_178,In_510);
nor U517 (N_517,In_743,In_507);
xnor U518 (N_518,In_74,In_715);
nand U519 (N_519,In_896,In_60);
nand U520 (N_520,In_947,In_909);
nor U521 (N_521,In_566,In_704);
and U522 (N_522,In_239,In_202);
nor U523 (N_523,In_833,In_506);
nor U524 (N_524,In_138,In_119);
nor U525 (N_525,In_787,In_488);
nand U526 (N_526,In_616,In_458);
xor U527 (N_527,In_548,In_265);
nand U528 (N_528,In_31,In_706);
and U529 (N_529,In_664,In_444);
xnor U530 (N_530,In_752,In_895);
and U531 (N_531,In_42,In_125);
nor U532 (N_532,In_18,In_258);
nand U533 (N_533,In_789,In_108);
and U534 (N_534,In_991,In_712);
and U535 (N_535,In_898,In_520);
xor U536 (N_536,In_31,In_490);
xor U537 (N_537,In_322,In_513);
nor U538 (N_538,In_877,In_387);
or U539 (N_539,In_208,In_513);
nand U540 (N_540,In_221,In_376);
xor U541 (N_541,In_198,In_72);
and U542 (N_542,In_90,In_334);
xnor U543 (N_543,In_41,In_430);
nand U544 (N_544,In_482,In_674);
and U545 (N_545,In_338,In_931);
xor U546 (N_546,In_35,In_385);
nor U547 (N_547,In_259,In_918);
and U548 (N_548,In_565,In_157);
and U549 (N_549,In_739,In_808);
xor U550 (N_550,In_833,In_834);
xnor U551 (N_551,In_922,In_26);
and U552 (N_552,In_36,In_205);
and U553 (N_553,In_711,In_712);
and U554 (N_554,In_343,In_392);
and U555 (N_555,In_734,In_517);
or U556 (N_556,In_694,In_790);
xnor U557 (N_557,In_64,In_56);
xnor U558 (N_558,In_309,In_703);
nor U559 (N_559,In_848,In_969);
nor U560 (N_560,In_44,In_79);
nand U561 (N_561,In_726,In_4);
and U562 (N_562,In_745,In_848);
and U563 (N_563,In_201,In_922);
nand U564 (N_564,In_897,In_341);
nand U565 (N_565,In_901,In_489);
nor U566 (N_566,In_530,In_534);
and U567 (N_567,In_854,In_510);
or U568 (N_568,In_235,In_329);
nor U569 (N_569,In_667,In_232);
and U570 (N_570,In_655,In_224);
xor U571 (N_571,In_972,In_47);
nor U572 (N_572,In_739,In_280);
nand U573 (N_573,In_305,In_905);
and U574 (N_574,In_267,In_11);
or U575 (N_575,In_754,In_686);
nor U576 (N_576,In_771,In_677);
xor U577 (N_577,In_374,In_94);
nand U578 (N_578,In_166,In_823);
and U579 (N_579,In_544,In_783);
and U580 (N_580,In_476,In_713);
and U581 (N_581,In_283,In_571);
and U582 (N_582,In_617,In_579);
nor U583 (N_583,In_766,In_483);
xor U584 (N_584,In_516,In_416);
nor U585 (N_585,In_244,In_944);
xor U586 (N_586,In_594,In_212);
nand U587 (N_587,In_421,In_457);
xor U588 (N_588,In_23,In_53);
nor U589 (N_589,In_791,In_166);
or U590 (N_590,In_327,In_722);
xnor U591 (N_591,In_684,In_200);
or U592 (N_592,In_516,In_927);
or U593 (N_593,In_554,In_238);
xnor U594 (N_594,In_527,In_74);
or U595 (N_595,In_713,In_606);
and U596 (N_596,In_213,In_956);
or U597 (N_597,In_534,In_133);
nand U598 (N_598,In_330,In_152);
nand U599 (N_599,In_16,In_953);
nand U600 (N_600,In_155,In_570);
or U601 (N_601,In_235,In_985);
xnor U602 (N_602,In_410,In_815);
nand U603 (N_603,In_740,In_899);
xnor U604 (N_604,In_886,In_452);
nand U605 (N_605,In_342,In_719);
and U606 (N_606,In_195,In_97);
and U607 (N_607,In_649,In_810);
and U608 (N_608,In_424,In_885);
and U609 (N_609,In_661,In_485);
or U610 (N_610,In_980,In_394);
nor U611 (N_611,In_273,In_556);
nand U612 (N_612,In_114,In_819);
or U613 (N_613,In_770,In_885);
nand U614 (N_614,In_352,In_834);
and U615 (N_615,In_446,In_650);
and U616 (N_616,In_917,In_439);
or U617 (N_617,In_478,In_933);
nor U618 (N_618,In_545,In_427);
nor U619 (N_619,In_367,In_812);
xnor U620 (N_620,In_609,In_212);
nor U621 (N_621,In_936,In_460);
or U622 (N_622,In_715,In_637);
nor U623 (N_623,In_688,In_9);
and U624 (N_624,In_626,In_790);
xnor U625 (N_625,In_705,In_295);
xnor U626 (N_626,In_697,In_753);
and U627 (N_627,In_242,In_102);
and U628 (N_628,In_911,In_93);
or U629 (N_629,In_574,In_657);
or U630 (N_630,In_810,In_0);
nor U631 (N_631,In_837,In_27);
and U632 (N_632,In_363,In_431);
nor U633 (N_633,In_258,In_856);
nor U634 (N_634,In_475,In_251);
nand U635 (N_635,In_868,In_202);
nor U636 (N_636,In_961,In_311);
or U637 (N_637,In_358,In_707);
or U638 (N_638,In_941,In_551);
xnor U639 (N_639,In_19,In_176);
nand U640 (N_640,In_825,In_132);
xnor U641 (N_641,In_703,In_934);
or U642 (N_642,In_633,In_579);
nand U643 (N_643,In_181,In_891);
or U644 (N_644,In_311,In_614);
and U645 (N_645,In_409,In_503);
or U646 (N_646,In_164,In_30);
xor U647 (N_647,In_129,In_240);
xor U648 (N_648,In_208,In_907);
xnor U649 (N_649,In_937,In_95);
nand U650 (N_650,In_548,In_605);
or U651 (N_651,In_282,In_920);
or U652 (N_652,In_394,In_123);
xnor U653 (N_653,In_365,In_24);
nor U654 (N_654,In_25,In_969);
and U655 (N_655,In_304,In_711);
nand U656 (N_656,In_554,In_423);
or U657 (N_657,In_100,In_841);
nor U658 (N_658,In_908,In_134);
and U659 (N_659,In_168,In_98);
nor U660 (N_660,In_221,In_56);
xor U661 (N_661,In_481,In_780);
or U662 (N_662,In_807,In_927);
xor U663 (N_663,In_183,In_695);
nand U664 (N_664,In_975,In_585);
nor U665 (N_665,In_956,In_523);
nor U666 (N_666,In_282,In_280);
and U667 (N_667,In_520,In_794);
nand U668 (N_668,In_54,In_169);
nand U669 (N_669,In_844,In_544);
nand U670 (N_670,In_96,In_493);
and U671 (N_671,In_739,In_778);
and U672 (N_672,In_128,In_946);
nor U673 (N_673,In_691,In_412);
xor U674 (N_674,In_723,In_458);
nor U675 (N_675,In_312,In_97);
xor U676 (N_676,In_806,In_923);
xor U677 (N_677,In_485,In_712);
or U678 (N_678,In_325,In_889);
nand U679 (N_679,In_871,In_831);
or U680 (N_680,In_589,In_164);
nor U681 (N_681,In_295,In_221);
and U682 (N_682,In_349,In_470);
xor U683 (N_683,In_805,In_848);
nand U684 (N_684,In_515,In_409);
xor U685 (N_685,In_2,In_491);
xor U686 (N_686,In_943,In_942);
and U687 (N_687,In_702,In_319);
nand U688 (N_688,In_497,In_417);
xor U689 (N_689,In_534,In_84);
and U690 (N_690,In_209,In_784);
and U691 (N_691,In_70,In_638);
nand U692 (N_692,In_63,In_633);
nand U693 (N_693,In_742,In_837);
and U694 (N_694,In_186,In_627);
nor U695 (N_695,In_434,In_468);
or U696 (N_696,In_690,In_219);
xnor U697 (N_697,In_33,In_818);
nor U698 (N_698,In_759,In_541);
nor U699 (N_699,In_346,In_454);
nor U700 (N_700,In_77,In_380);
nor U701 (N_701,In_401,In_842);
xor U702 (N_702,In_877,In_217);
nor U703 (N_703,In_848,In_240);
and U704 (N_704,In_997,In_301);
and U705 (N_705,In_559,In_331);
and U706 (N_706,In_879,In_830);
or U707 (N_707,In_651,In_75);
nand U708 (N_708,In_970,In_147);
nor U709 (N_709,In_154,In_854);
nor U710 (N_710,In_210,In_451);
nor U711 (N_711,In_15,In_636);
or U712 (N_712,In_390,In_911);
xor U713 (N_713,In_557,In_403);
and U714 (N_714,In_306,In_732);
or U715 (N_715,In_10,In_490);
or U716 (N_716,In_876,In_440);
and U717 (N_717,In_287,In_980);
xor U718 (N_718,In_243,In_803);
or U719 (N_719,In_666,In_330);
and U720 (N_720,In_676,In_395);
nor U721 (N_721,In_569,In_158);
xor U722 (N_722,In_893,In_144);
nor U723 (N_723,In_324,In_547);
and U724 (N_724,In_160,In_527);
xor U725 (N_725,In_140,In_846);
or U726 (N_726,In_510,In_771);
xnor U727 (N_727,In_416,In_811);
xnor U728 (N_728,In_155,In_396);
xor U729 (N_729,In_675,In_288);
or U730 (N_730,In_700,In_242);
or U731 (N_731,In_92,In_916);
nand U732 (N_732,In_449,In_660);
and U733 (N_733,In_28,In_83);
xor U734 (N_734,In_266,In_352);
and U735 (N_735,In_766,In_987);
nor U736 (N_736,In_693,In_768);
nand U737 (N_737,In_339,In_811);
xor U738 (N_738,In_626,In_641);
xnor U739 (N_739,In_104,In_513);
xnor U740 (N_740,In_88,In_547);
nor U741 (N_741,In_191,In_638);
nand U742 (N_742,In_602,In_551);
nand U743 (N_743,In_830,In_50);
and U744 (N_744,In_161,In_51);
nand U745 (N_745,In_222,In_412);
xnor U746 (N_746,In_453,In_275);
nand U747 (N_747,In_652,In_941);
and U748 (N_748,In_529,In_382);
xor U749 (N_749,In_720,In_383);
or U750 (N_750,In_632,In_642);
or U751 (N_751,In_674,In_879);
nand U752 (N_752,In_212,In_453);
or U753 (N_753,In_801,In_901);
nor U754 (N_754,In_285,In_914);
and U755 (N_755,In_600,In_262);
nand U756 (N_756,In_803,In_560);
nand U757 (N_757,In_239,In_914);
xor U758 (N_758,In_759,In_395);
and U759 (N_759,In_94,In_540);
xor U760 (N_760,In_588,In_929);
or U761 (N_761,In_361,In_863);
nor U762 (N_762,In_909,In_551);
or U763 (N_763,In_270,In_753);
nand U764 (N_764,In_143,In_29);
nor U765 (N_765,In_929,In_382);
nand U766 (N_766,In_499,In_272);
and U767 (N_767,In_942,In_133);
and U768 (N_768,In_446,In_322);
nor U769 (N_769,In_56,In_513);
and U770 (N_770,In_391,In_363);
and U771 (N_771,In_914,In_901);
nor U772 (N_772,In_710,In_523);
nor U773 (N_773,In_121,In_500);
nand U774 (N_774,In_78,In_398);
nand U775 (N_775,In_472,In_843);
xor U776 (N_776,In_432,In_468);
xnor U777 (N_777,In_191,In_80);
nor U778 (N_778,In_640,In_365);
xor U779 (N_779,In_196,In_122);
nand U780 (N_780,In_498,In_924);
or U781 (N_781,In_459,In_274);
nand U782 (N_782,In_341,In_357);
nor U783 (N_783,In_965,In_617);
nand U784 (N_784,In_393,In_435);
nor U785 (N_785,In_149,In_156);
or U786 (N_786,In_168,In_750);
or U787 (N_787,In_610,In_9);
or U788 (N_788,In_884,In_561);
xnor U789 (N_789,In_617,In_301);
xnor U790 (N_790,In_980,In_647);
or U791 (N_791,In_861,In_24);
xnor U792 (N_792,In_348,In_531);
nor U793 (N_793,In_332,In_552);
or U794 (N_794,In_25,In_751);
nand U795 (N_795,In_94,In_434);
and U796 (N_796,In_990,In_465);
nand U797 (N_797,In_262,In_373);
and U798 (N_798,In_410,In_816);
or U799 (N_799,In_116,In_758);
or U800 (N_800,In_576,In_148);
nand U801 (N_801,In_357,In_503);
nand U802 (N_802,In_135,In_889);
nor U803 (N_803,In_365,In_566);
or U804 (N_804,In_90,In_398);
xor U805 (N_805,In_808,In_682);
or U806 (N_806,In_826,In_741);
and U807 (N_807,In_778,In_288);
or U808 (N_808,In_579,In_667);
and U809 (N_809,In_633,In_991);
nand U810 (N_810,In_116,In_235);
xnor U811 (N_811,In_685,In_265);
xnor U812 (N_812,In_369,In_210);
or U813 (N_813,In_1,In_378);
nand U814 (N_814,In_648,In_35);
nand U815 (N_815,In_533,In_635);
nor U816 (N_816,In_364,In_550);
nand U817 (N_817,In_211,In_749);
nand U818 (N_818,In_596,In_216);
or U819 (N_819,In_884,In_199);
xnor U820 (N_820,In_337,In_57);
or U821 (N_821,In_417,In_773);
or U822 (N_822,In_650,In_224);
and U823 (N_823,In_924,In_156);
nand U824 (N_824,In_254,In_993);
or U825 (N_825,In_763,In_550);
xnor U826 (N_826,In_467,In_449);
nor U827 (N_827,In_715,In_943);
nand U828 (N_828,In_545,In_275);
xor U829 (N_829,In_789,In_217);
xor U830 (N_830,In_434,In_859);
xor U831 (N_831,In_921,In_753);
or U832 (N_832,In_705,In_840);
and U833 (N_833,In_652,In_422);
nand U834 (N_834,In_960,In_789);
or U835 (N_835,In_977,In_706);
nor U836 (N_836,In_873,In_727);
and U837 (N_837,In_530,In_947);
xor U838 (N_838,In_536,In_180);
or U839 (N_839,In_826,In_146);
nand U840 (N_840,In_831,In_717);
nor U841 (N_841,In_963,In_314);
or U842 (N_842,In_770,In_530);
or U843 (N_843,In_442,In_451);
xnor U844 (N_844,In_372,In_248);
xor U845 (N_845,In_974,In_746);
or U846 (N_846,In_667,In_993);
xor U847 (N_847,In_762,In_800);
xor U848 (N_848,In_893,In_299);
and U849 (N_849,In_202,In_33);
or U850 (N_850,In_326,In_862);
or U851 (N_851,In_266,In_222);
nand U852 (N_852,In_735,In_271);
and U853 (N_853,In_874,In_123);
nand U854 (N_854,In_28,In_344);
nor U855 (N_855,In_201,In_219);
xnor U856 (N_856,In_250,In_5);
nor U857 (N_857,In_590,In_422);
and U858 (N_858,In_812,In_628);
nor U859 (N_859,In_188,In_161);
xor U860 (N_860,In_355,In_901);
nor U861 (N_861,In_269,In_576);
or U862 (N_862,In_672,In_788);
xnor U863 (N_863,In_784,In_88);
nor U864 (N_864,In_427,In_961);
or U865 (N_865,In_51,In_270);
or U866 (N_866,In_583,In_833);
and U867 (N_867,In_716,In_27);
and U868 (N_868,In_291,In_824);
and U869 (N_869,In_385,In_625);
nor U870 (N_870,In_65,In_845);
nor U871 (N_871,In_128,In_65);
nor U872 (N_872,In_706,In_114);
and U873 (N_873,In_462,In_612);
nor U874 (N_874,In_500,In_360);
xor U875 (N_875,In_237,In_52);
and U876 (N_876,In_357,In_304);
nand U877 (N_877,In_825,In_819);
and U878 (N_878,In_79,In_57);
nand U879 (N_879,In_490,In_331);
nor U880 (N_880,In_841,In_648);
nand U881 (N_881,In_598,In_784);
and U882 (N_882,In_895,In_801);
or U883 (N_883,In_458,In_623);
or U884 (N_884,In_889,In_422);
xnor U885 (N_885,In_639,In_505);
nand U886 (N_886,In_982,In_112);
and U887 (N_887,In_756,In_118);
and U888 (N_888,In_374,In_719);
and U889 (N_889,In_952,In_36);
and U890 (N_890,In_22,In_538);
xnor U891 (N_891,In_852,In_267);
and U892 (N_892,In_627,In_773);
nand U893 (N_893,In_501,In_135);
nor U894 (N_894,In_906,In_111);
nor U895 (N_895,In_497,In_816);
xnor U896 (N_896,In_692,In_645);
nor U897 (N_897,In_129,In_275);
nand U898 (N_898,In_192,In_118);
nor U899 (N_899,In_978,In_2);
and U900 (N_900,In_314,In_602);
xnor U901 (N_901,In_50,In_388);
nand U902 (N_902,In_938,In_437);
nor U903 (N_903,In_780,In_615);
and U904 (N_904,In_830,In_900);
xnor U905 (N_905,In_796,In_429);
xor U906 (N_906,In_333,In_60);
xor U907 (N_907,In_461,In_235);
xnor U908 (N_908,In_266,In_304);
or U909 (N_909,In_759,In_642);
or U910 (N_910,In_227,In_748);
xor U911 (N_911,In_822,In_483);
and U912 (N_912,In_307,In_272);
nor U913 (N_913,In_526,In_841);
or U914 (N_914,In_341,In_194);
nand U915 (N_915,In_806,In_168);
xnor U916 (N_916,In_429,In_780);
xnor U917 (N_917,In_260,In_437);
nor U918 (N_918,In_855,In_286);
nor U919 (N_919,In_83,In_838);
and U920 (N_920,In_800,In_344);
or U921 (N_921,In_92,In_33);
and U922 (N_922,In_446,In_160);
nor U923 (N_923,In_463,In_222);
xor U924 (N_924,In_748,In_183);
nand U925 (N_925,In_124,In_583);
nor U926 (N_926,In_366,In_21);
and U927 (N_927,In_832,In_77);
xnor U928 (N_928,In_256,In_360);
and U929 (N_929,In_951,In_859);
nor U930 (N_930,In_46,In_108);
nor U931 (N_931,In_465,In_924);
xor U932 (N_932,In_29,In_444);
xor U933 (N_933,In_435,In_230);
nor U934 (N_934,In_590,In_521);
xnor U935 (N_935,In_687,In_792);
or U936 (N_936,In_43,In_956);
nor U937 (N_937,In_838,In_487);
or U938 (N_938,In_325,In_210);
nor U939 (N_939,In_529,In_758);
xnor U940 (N_940,In_433,In_546);
and U941 (N_941,In_474,In_118);
xnor U942 (N_942,In_283,In_639);
or U943 (N_943,In_159,In_599);
nor U944 (N_944,In_571,In_568);
nand U945 (N_945,In_915,In_482);
nor U946 (N_946,In_801,In_849);
or U947 (N_947,In_810,In_734);
or U948 (N_948,In_929,In_5);
or U949 (N_949,In_509,In_525);
and U950 (N_950,In_916,In_419);
or U951 (N_951,In_435,In_379);
or U952 (N_952,In_524,In_12);
xnor U953 (N_953,In_484,In_719);
and U954 (N_954,In_462,In_949);
and U955 (N_955,In_707,In_342);
nand U956 (N_956,In_326,In_229);
nor U957 (N_957,In_465,In_423);
nor U958 (N_958,In_82,In_913);
and U959 (N_959,In_486,In_63);
and U960 (N_960,In_898,In_766);
xnor U961 (N_961,In_507,In_52);
and U962 (N_962,In_821,In_519);
xnor U963 (N_963,In_866,In_772);
xor U964 (N_964,In_43,In_859);
and U965 (N_965,In_126,In_106);
nand U966 (N_966,In_938,In_426);
nand U967 (N_967,In_334,In_110);
nor U968 (N_968,In_5,In_999);
nor U969 (N_969,In_734,In_891);
and U970 (N_970,In_576,In_705);
nor U971 (N_971,In_19,In_495);
nand U972 (N_972,In_222,In_734);
nand U973 (N_973,In_728,In_323);
and U974 (N_974,In_522,In_491);
and U975 (N_975,In_650,In_210);
or U976 (N_976,In_103,In_213);
or U977 (N_977,In_94,In_288);
and U978 (N_978,In_683,In_112);
and U979 (N_979,In_82,In_241);
nor U980 (N_980,In_249,In_690);
nand U981 (N_981,In_733,In_855);
xor U982 (N_982,In_22,In_77);
nand U983 (N_983,In_774,In_282);
and U984 (N_984,In_17,In_243);
nand U985 (N_985,In_368,In_577);
xor U986 (N_986,In_100,In_178);
nand U987 (N_987,In_293,In_543);
or U988 (N_988,In_463,In_521);
nand U989 (N_989,In_612,In_461);
and U990 (N_990,In_185,In_825);
nor U991 (N_991,In_681,In_876);
xnor U992 (N_992,In_563,In_392);
nor U993 (N_993,In_394,In_259);
and U994 (N_994,In_803,In_475);
or U995 (N_995,In_261,In_178);
xor U996 (N_996,In_499,In_136);
nor U997 (N_997,In_795,In_672);
or U998 (N_998,In_273,In_92);
xnor U999 (N_999,In_600,In_559);
nand U1000 (N_1000,In_108,In_804);
or U1001 (N_1001,In_476,In_881);
or U1002 (N_1002,In_288,In_835);
or U1003 (N_1003,In_237,In_627);
and U1004 (N_1004,In_177,In_748);
or U1005 (N_1005,In_460,In_631);
nor U1006 (N_1006,In_376,In_661);
or U1007 (N_1007,In_297,In_549);
nand U1008 (N_1008,In_391,In_251);
nor U1009 (N_1009,In_906,In_400);
or U1010 (N_1010,In_610,In_531);
nor U1011 (N_1011,In_307,In_980);
and U1012 (N_1012,In_503,In_15);
or U1013 (N_1013,In_687,In_131);
or U1014 (N_1014,In_507,In_108);
nor U1015 (N_1015,In_811,In_719);
xnor U1016 (N_1016,In_643,In_36);
or U1017 (N_1017,In_73,In_941);
or U1018 (N_1018,In_345,In_943);
nand U1019 (N_1019,In_620,In_123);
and U1020 (N_1020,In_459,In_456);
or U1021 (N_1021,In_650,In_16);
or U1022 (N_1022,In_764,In_899);
nand U1023 (N_1023,In_475,In_690);
nand U1024 (N_1024,In_753,In_971);
and U1025 (N_1025,In_664,In_400);
nand U1026 (N_1026,In_801,In_401);
nand U1027 (N_1027,In_622,In_86);
or U1028 (N_1028,In_166,In_763);
and U1029 (N_1029,In_102,In_663);
nand U1030 (N_1030,In_612,In_374);
and U1031 (N_1031,In_561,In_137);
nand U1032 (N_1032,In_538,In_122);
xnor U1033 (N_1033,In_816,In_727);
or U1034 (N_1034,In_811,In_995);
and U1035 (N_1035,In_14,In_142);
or U1036 (N_1036,In_323,In_767);
nor U1037 (N_1037,In_903,In_809);
nor U1038 (N_1038,In_867,In_548);
or U1039 (N_1039,In_917,In_821);
nor U1040 (N_1040,In_420,In_590);
nor U1041 (N_1041,In_63,In_804);
xor U1042 (N_1042,In_986,In_210);
xnor U1043 (N_1043,In_743,In_666);
xnor U1044 (N_1044,In_290,In_78);
or U1045 (N_1045,In_796,In_11);
or U1046 (N_1046,In_594,In_402);
or U1047 (N_1047,In_226,In_607);
xor U1048 (N_1048,In_827,In_972);
xor U1049 (N_1049,In_514,In_19);
nand U1050 (N_1050,In_823,In_187);
or U1051 (N_1051,In_920,In_215);
nand U1052 (N_1052,In_301,In_3);
and U1053 (N_1053,In_240,In_117);
or U1054 (N_1054,In_488,In_63);
nor U1055 (N_1055,In_0,In_258);
or U1056 (N_1056,In_206,In_475);
xnor U1057 (N_1057,In_915,In_930);
or U1058 (N_1058,In_472,In_909);
xor U1059 (N_1059,In_709,In_847);
or U1060 (N_1060,In_233,In_729);
and U1061 (N_1061,In_652,In_87);
or U1062 (N_1062,In_216,In_104);
nand U1063 (N_1063,In_184,In_10);
nor U1064 (N_1064,In_825,In_901);
nor U1065 (N_1065,In_243,In_38);
nand U1066 (N_1066,In_444,In_529);
nand U1067 (N_1067,In_291,In_966);
xor U1068 (N_1068,In_89,In_310);
xor U1069 (N_1069,In_175,In_118);
xor U1070 (N_1070,In_79,In_437);
and U1071 (N_1071,In_261,In_185);
nand U1072 (N_1072,In_356,In_718);
nand U1073 (N_1073,In_669,In_746);
and U1074 (N_1074,In_922,In_889);
or U1075 (N_1075,In_941,In_927);
nor U1076 (N_1076,In_678,In_128);
nor U1077 (N_1077,In_508,In_711);
xor U1078 (N_1078,In_725,In_381);
and U1079 (N_1079,In_531,In_723);
and U1080 (N_1080,In_609,In_262);
xor U1081 (N_1081,In_571,In_32);
or U1082 (N_1082,In_800,In_51);
or U1083 (N_1083,In_46,In_775);
nor U1084 (N_1084,In_505,In_297);
or U1085 (N_1085,In_645,In_254);
xor U1086 (N_1086,In_211,In_472);
nand U1087 (N_1087,In_542,In_620);
nand U1088 (N_1088,In_595,In_755);
xnor U1089 (N_1089,In_109,In_832);
nor U1090 (N_1090,In_470,In_736);
or U1091 (N_1091,In_958,In_344);
nand U1092 (N_1092,In_741,In_342);
or U1093 (N_1093,In_751,In_953);
nor U1094 (N_1094,In_509,In_365);
nand U1095 (N_1095,In_498,In_552);
or U1096 (N_1096,In_732,In_731);
xnor U1097 (N_1097,In_337,In_804);
and U1098 (N_1098,In_848,In_273);
or U1099 (N_1099,In_314,In_925);
nor U1100 (N_1100,In_606,In_782);
or U1101 (N_1101,In_393,In_246);
nor U1102 (N_1102,In_211,In_589);
or U1103 (N_1103,In_546,In_227);
xnor U1104 (N_1104,In_755,In_102);
nor U1105 (N_1105,In_96,In_739);
nor U1106 (N_1106,In_188,In_632);
xnor U1107 (N_1107,In_318,In_277);
or U1108 (N_1108,In_642,In_885);
xnor U1109 (N_1109,In_534,In_837);
nor U1110 (N_1110,In_293,In_517);
and U1111 (N_1111,In_677,In_159);
nor U1112 (N_1112,In_669,In_936);
or U1113 (N_1113,In_445,In_722);
and U1114 (N_1114,In_660,In_402);
and U1115 (N_1115,In_483,In_831);
nor U1116 (N_1116,In_703,In_172);
and U1117 (N_1117,In_505,In_711);
nor U1118 (N_1118,In_157,In_634);
or U1119 (N_1119,In_118,In_535);
xor U1120 (N_1120,In_266,In_447);
and U1121 (N_1121,In_750,In_337);
and U1122 (N_1122,In_234,In_116);
or U1123 (N_1123,In_130,In_521);
or U1124 (N_1124,In_194,In_475);
nor U1125 (N_1125,In_464,In_991);
or U1126 (N_1126,In_193,In_211);
or U1127 (N_1127,In_647,In_424);
or U1128 (N_1128,In_792,In_585);
xnor U1129 (N_1129,In_319,In_913);
nand U1130 (N_1130,In_805,In_283);
or U1131 (N_1131,In_264,In_69);
nor U1132 (N_1132,In_297,In_883);
nor U1133 (N_1133,In_805,In_547);
nor U1134 (N_1134,In_257,In_779);
xor U1135 (N_1135,In_16,In_386);
nor U1136 (N_1136,In_743,In_760);
nor U1137 (N_1137,In_507,In_621);
nor U1138 (N_1138,In_966,In_876);
nor U1139 (N_1139,In_230,In_266);
xnor U1140 (N_1140,In_570,In_834);
and U1141 (N_1141,In_406,In_300);
xor U1142 (N_1142,In_441,In_15);
or U1143 (N_1143,In_537,In_675);
nor U1144 (N_1144,In_383,In_429);
xor U1145 (N_1145,In_82,In_663);
and U1146 (N_1146,In_971,In_155);
xnor U1147 (N_1147,In_6,In_580);
and U1148 (N_1148,In_201,In_861);
nor U1149 (N_1149,In_187,In_169);
nor U1150 (N_1150,In_127,In_230);
xor U1151 (N_1151,In_452,In_348);
xnor U1152 (N_1152,In_45,In_89);
or U1153 (N_1153,In_391,In_810);
or U1154 (N_1154,In_812,In_25);
and U1155 (N_1155,In_289,In_377);
and U1156 (N_1156,In_558,In_703);
and U1157 (N_1157,In_293,In_696);
xor U1158 (N_1158,In_292,In_948);
nor U1159 (N_1159,In_931,In_155);
or U1160 (N_1160,In_555,In_779);
nand U1161 (N_1161,In_378,In_372);
and U1162 (N_1162,In_464,In_962);
nand U1163 (N_1163,In_358,In_685);
or U1164 (N_1164,In_357,In_604);
xnor U1165 (N_1165,In_398,In_94);
nor U1166 (N_1166,In_273,In_202);
and U1167 (N_1167,In_588,In_894);
xor U1168 (N_1168,In_215,In_100);
nor U1169 (N_1169,In_431,In_289);
nor U1170 (N_1170,In_140,In_266);
nor U1171 (N_1171,In_662,In_457);
nand U1172 (N_1172,In_415,In_539);
xnor U1173 (N_1173,In_536,In_669);
or U1174 (N_1174,In_124,In_140);
or U1175 (N_1175,In_487,In_64);
and U1176 (N_1176,In_971,In_257);
nand U1177 (N_1177,In_814,In_670);
nor U1178 (N_1178,In_380,In_974);
and U1179 (N_1179,In_793,In_384);
nor U1180 (N_1180,In_953,In_192);
xnor U1181 (N_1181,In_75,In_721);
xor U1182 (N_1182,In_366,In_368);
or U1183 (N_1183,In_286,In_509);
or U1184 (N_1184,In_407,In_750);
nand U1185 (N_1185,In_605,In_189);
nor U1186 (N_1186,In_802,In_590);
or U1187 (N_1187,In_177,In_999);
or U1188 (N_1188,In_896,In_323);
xnor U1189 (N_1189,In_465,In_331);
xor U1190 (N_1190,In_945,In_882);
xnor U1191 (N_1191,In_316,In_606);
nand U1192 (N_1192,In_492,In_283);
and U1193 (N_1193,In_87,In_191);
nand U1194 (N_1194,In_881,In_412);
nor U1195 (N_1195,In_826,In_317);
nor U1196 (N_1196,In_850,In_747);
or U1197 (N_1197,In_276,In_349);
and U1198 (N_1198,In_869,In_373);
or U1199 (N_1199,In_520,In_602);
xnor U1200 (N_1200,In_679,In_77);
xor U1201 (N_1201,In_641,In_471);
xor U1202 (N_1202,In_492,In_932);
xnor U1203 (N_1203,In_30,In_176);
and U1204 (N_1204,In_965,In_152);
nand U1205 (N_1205,In_772,In_355);
or U1206 (N_1206,In_872,In_325);
nor U1207 (N_1207,In_916,In_710);
nand U1208 (N_1208,In_30,In_865);
xnor U1209 (N_1209,In_805,In_998);
nand U1210 (N_1210,In_67,In_18);
or U1211 (N_1211,In_765,In_143);
or U1212 (N_1212,In_985,In_720);
nand U1213 (N_1213,In_412,In_58);
or U1214 (N_1214,In_582,In_852);
and U1215 (N_1215,In_462,In_965);
or U1216 (N_1216,In_522,In_300);
or U1217 (N_1217,In_537,In_930);
or U1218 (N_1218,In_470,In_276);
xor U1219 (N_1219,In_361,In_909);
nor U1220 (N_1220,In_217,In_441);
nor U1221 (N_1221,In_557,In_63);
xor U1222 (N_1222,In_698,In_877);
and U1223 (N_1223,In_857,In_54);
nor U1224 (N_1224,In_697,In_419);
nor U1225 (N_1225,In_506,In_347);
and U1226 (N_1226,In_561,In_316);
nor U1227 (N_1227,In_666,In_459);
or U1228 (N_1228,In_570,In_930);
nand U1229 (N_1229,In_949,In_123);
nor U1230 (N_1230,In_395,In_486);
xnor U1231 (N_1231,In_554,In_46);
nor U1232 (N_1232,In_877,In_440);
nor U1233 (N_1233,In_194,In_910);
and U1234 (N_1234,In_98,In_124);
nand U1235 (N_1235,In_142,In_158);
nor U1236 (N_1236,In_392,In_302);
or U1237 (N_1237,In_265,In_299);
xor U1238 (N_1238,In_11,In_932);
nand U1239 (N_1239,In_606,In_758);
or U1240 (N_1240,In_255,In_827);
and U1241 (N_1241,In_703,In_454);
xor U1242 (N_1242,In_926,In_82);
nor U1243 (N_1243,In_738,In_380);
xor U1244 (N_1244,In_888,In_308);
and U1245 (N_1245,In_222,In_220);
nand U1246 (N_1246,In_19,In_286);
xnor U1247 (N_1247,In_351,In_239);
or U1248 (N_1248,In_971,In_377);
or U1249 (N_1249,In_766,In_109);
xnor U1250 (N_1250,In_429,In_99);
and U1251 (N_1251,In_618,In_392);
xor U1252 (N_1252,In_705,In_644);
xnor U1253 (N_1253,In_666,In_66);
xnor U1254 (N_1254,In_925,In_842);
and U1255 (N_1255,In_761,In_556);
xor U1256 (N_1256,In_575,In_190);
xnor U1257 (N_1257,In_481,In_834);
or U1258 (N_1258,In_82,In_705);
xor U1259 (N_1259,In_352,In_703);
or U1260 (N_1260,In_732,In_396);
nor U1261 (N_1261,In_313,In_420);
and U1262 (N_1262,In_931,In_198);
and U1263 (N_1263,In_746,In_148);
or U1264 (N_1264,In_484,In_730);
and U1265 (N_1265,In_188,In_739);
and U1266 (N_1266,In_780,In_364);
nand U1267 (N_1267,In_504,In_809);
nor U1268 (N_1268,In_423,In_104);
or U1269 (N_1269,In_959,In_932);
xnor U1270 (N_1270,In_890,In_735);
xor U1271 (N_1271,In_998,In_423);
xor U1272 (N_1272,In_963,In_212);
xnor U1273 (N_1273,In_964,In_676);
and U1274 (N_1274,In_705,In_209);
xnor U1275 (N_1275,In_245,In_707);
xnor U1276 (N_1276,In_434,In_549);
and U1277 (N_1277,In_476,In_40);
and U1278 (N_1278,In_669,In_340);
or U1279 (N_1279,In_647,In_957);
xor U1280 (N_1280,In_626,In_818);
nand U1281 (N_1281,In_702,In_465);
xnor U1282 (N_1282,In_553,In_667);
and U1283 (N_1283,In_522,In_0);
and U1284 (N_1284,In_712,In_705);
and U1285 (N_1285,In_877,In_868);
or U1286 (N_1286,In_102,In_403);
or U1287 (N_1287,In_712,In_838);
nor U1288 (N_1288,In_942,In_886);
xor U1289 (N_1289,In_871,In_217);
nand U1290 (N_1290,In_4,In_901);
and U1291 (N_1291,In_482,In_307);
nand U1292 (N_1292,In_722,In_535);
nand U1293 (N_1293,In_921,In_819);
xnor U1294 (N_1294,In_458,In_441);
nor U1295 (N_1295,In_259,In_187);
nor U1296 (N_1296,In_101,In_836);
nand U1297 (N_1297,In_234,In_903);
nand U1298 (N_1298,In_617,In_975);
or U1299 (N_1299,In_366,In_946);
or U1300 (N_1300,In_51,In_564);
or U1301 (N_1301,In_564,In_512);
or U1302 (N_1302,In_756,In_449);
nand U1303 (N_1303,In_574,In_634);
and U1304 (N_1304,In_998,In_397);
nor U1305 (N_1305,In_530,In_407);
or U1306 (N_1306,In_346,In_906);
and U1307 (N_1307,In_816,In_4);
nor U1308 (N_1308,In_493,In_489);
or U1309 (N_1309,In_862,In_718);
or U1310 (N_1310,In_770,In_389);
nand U1311 (N_1311,In_310,In_83);
xor U1312 (N_1312,In_693,In_806);
or U1313 (N_1313,In_600,In_471);
and U1314 (N_1314,In_48,In_931);
nor U1315 (N_1315,In_579,In_7);
xnor U1316 (N_1316,In_387,In_901);
xnor U1317 (N_1317,In_838,In_586);
and U1318 (N_1318,In_235,In_771);
xnor U1319 (N_1319,In_689,In_480);
nor U1320 (N_1320,In_89,In_736);
xor U1321 (N_1321,In_854,In_290);
nand U1322 (N_1322,In_802,In_857);
and U1323 (N_1323,In_883,In_927);
nand U1324 (N_1324,In_224,In_271);
and U1325 (N_1325,In_872,In_43);
xnor U1326 (N_1326,In_375,In_779);
or U1327 (N_1327,In_930,In_666);
nor U1328 (N_1328,In_758,In_561);
or U1329 (N_1329,In_800,In_875);
nand U1330 (N_1330,In_971,In_863);
nor U1331 (N_1331,In_59,In_892);
and U1332 (N_1332,In_182,In_941);
or U1333 (N_1333,In_226,In_989);
xor U1334 (N_1334,In_330,In_966);
nor U1335 (N_1335,In_806,In_902);
or U1336 (N_1336,In_643,In_161);
nor U1337 (N_1337,In_825,In_566);
nor U1338 (N_1338,In_480,In_928);
nor U1339 (N_1339,In_467,In_398);
nor U1340 (N_1340,In_84,In_121);
or U1341 (N_1341,In_563,In_558);
and U1342 (N_1342,In_653,In_806);
and U1343 (N_1343,In_589,In_471);
nand U1344 (N_1344,In_434,In_621);
nand U1345 (N_1345,In_867,In_995);
nand U1346 (N_1346,In_556,In_580);
xor U1347 (N_1347,In_94,In_7);
or U1348 (N_1348,In_230,In_917);
xor U1349 (N_1349,In_83,In_55);
or U1350 (N_1350,In_507,In_711);
or U1351 (N_1351,In_796,In_376);
or U1352 (N_1352,In_955,In_573);
nor U1353 (N_1353,In_472,In_384);
or U1354 (N_1354,In_868,In_753);
nor U1355 (N_1355,In_688,In_187);
nand U1356 (N_1356,In_683,In_161);
xor U1357 (N_1357,In_422,In_648);
nand U1358 (N_1358,In_828,In_845);
nor U1359 (N_1359,In_490,In_273);
or U1360 (N_1360,In_763,In_288);
xnor U1361 (N_1361,In_619,In_455);
nand U1362 (N_1362,In_386,In_257);
nor U1363 (N_1363,In_675,In_756);
nand U1364 (N_1364,In_210,In_924);
nor U1365 (N_1365,In_93,In_427);
nor U1366 (N_1366,In_61,In_266);
xor U1367 (N_1367,In_552,In_577);
nor U1368 (N_1368,In_385,In_808);
nor U1369 (N_1369,In_382,In_80);
and U1370 (N_1370,In_20,In_298);
and U1371 (N_1371,In_764,In_825);
nand U1372 (N_1372,In_172,In_474);
nand U1373 (N_1373,In_729,In_63);
xnor U1374 (N_1374,In_965,In_460);
and U1375 (N_1375,In_555,In_803);
and U1376 (N_1376,In_525,In_688);
nand U1377 (N_1377,In_152,In_601);
nand U1378 (N_1378,In_10,In_582);
xor U1379 (N_1379,In_72,In_703);
nand U1380 (N_1380,In_610,In_446);
nand U1381 (N_1381,In_565,In_647);
or U1382 (N_1382,In_376,In_358);
or U1383 (N_1383,In_407,In_800);
or U1384 (N_1384,In_997,In_4);
nand U1385 (N_1385,In_973,In_941);
xor U1386 (N_1386,In_608,In_681);
and U1387 (N_1387,In_204,In_73);
and U1388 (N_1388,In_658,In_533);
nand U1389 (N_1389,In_309,In_367);
nand U1390 (N_1390,In_915,In_151);
and U1391 (N_1391,In_971,In_855);
or U1392 (N_1392,In_392,In_120);
and U1393 (N_1393,In_163,In_881);
or U1394 (N_1394,In_918,In_320);
and U1395 (N_1395,In_316,In_860);
or U1396 (N_1396,In_616,In_302);
nand U1397 (N_1397,In_683,In_724);
xnor U1398 (N_1398,In_999,In_595);
nor U1399 (N_1399,In_819,In_155);
xor U1400 (N_1400,In_409,In_610);
and U1401 (N_1401,In_213,In_513);
nor U1402 (N_1402,In_927,In_27);
nor U1403 (N_1403,In_917,In_133);
or U1404 (N_1404,In_407,In_780);
nand U1405 (N_1405,In_150,In_973);
nand U1406 (N_1406,In_354,In_494);
xnor U1407 (N_1407,In_711,In_843);
or U1408 (N_1408,In_0,In_356);
nand U1409 (N_1409,In_953,In_823);
or U1410 (N_1410,In_607,In_719);
xnor U1411 (N_1411,In_585,In_233);
or U1412 (N_1412,In_791,In_433);
or U1413 (N_1413,In_719,In_186);
nor U1414 (N_1414,In_846,In_703);
and U1415 (N_1415,In_553,In_545);
and U1416 (N_1416,In_231,In_268);
xor U1417 (N_1417,In_360,In_764);
and U1418 (N_1418,In_645,In_349);
nor U1419 (N_1419,In_940,In_605);
or U1420 (N_1420,In_468,In_649);
or U1421 (N_1421,In_984,In_262);
nand U1422 (N_1422,In_317,In_278);
xor U1423 (N_1423,In_441,In_917);
nor U1424 (N_1424,In_38,In_890);
or U1425 (N_1425,In_214,In_964);
and U1426 (N_1426,In_134,In_3);
nor U1427 (N_1427,In_398,In_681);
nand U1428 (N_1428,In_55,In_586);
nand U1429 (N_1429,In_772,In_120);
nor U1430 (N_1430,In_887,In_311);
nor U1431 (N_1431,In_541,In_679);
or U1432 (N_1432,In_147,In_609);
or U1433 (N_1433,In_427,In_431);
nand U1434 (N_1434,In_650,In_966);
or U1435 (N_1435,In_726,In_464);
nor U1436 (N_1436,In_37,In_962);
nor U1437 (N_1437,In_809,In_33);
and U1438 (N_1438,In_926,In_301);
and U1439 (N_1439,In_230,In_757);
or U1440 (N_1440,In_44,In_768);
and U1441 (N_1441,In_704,In_876);
nand U1442 (N_1442,In_992,In_775);
xnor U1443 (N_1443,In_894,In_698);
nor U1444 (N_1444,In_709,In_543);
and U1445 (N_1445,In_831,In_300);
nor U1446 (N_1446,In_852,In_666);
or U1447 (N_1447,In_777,In_174);
xor U1448 (N_1448,In_788,In_983);
nand U1449 (N_1449,In_619,In_420);
xor U1450 (N_1450,In_996,In_444);
or U1451 (N_1451,In_241,In_929);
xor U1452 (N_1452,In_126,In_139);
nor U1453 (N_1453,In_98,In_494);
nand U1454 (N_1454,In_367,In_627);
nand U1455 (N_1455,In_168,In_675);
nand U1456 (N_1456,In_302,In_443);
nand U1457 (N_1457,In_1,In_176);
or U1458 (N_1458,In_620,In_156);
xnor U1459 (N_1459,In_878,In_776);
and U1460 (N_1460,In_186,In_681);
or U1461 (N_1461,In_2,In_661);
nor U1462 (N_1462,In_372,In_276);
or U1463 (N_1463,In_513,In_164);
or U1464 (N_1464,In_272,In_429);
xnor U1465 (N_1465,In_415,In_676);
nand U1466 (N_1466,In_514,In_613);
or U1467 (N_1467,In_553,In_973);
nand U1468 (N_1468,In_284,In_802);
xor U1469 (N_1469,In_919,In_271);
nand U1470 (N_1470,In_368,In_224);
nor U1471 (N_1471,In_678,In_727);
xnor U1472 (N_1472,In_501,In_452);
nor U1473 (N_1473,In_158,In_369);
and U1474 (N_1474,In_894,In_842);
nand U1475 (N_1475,In_59,In_409);
or U1476 (N_1476,In_87,In_671);
and U1477 (N_1477,In_240,In_782);
or U1478 (N_1478,In_398,In_993);
nand U1479 (N_1479,In_789,In_779);
or U1480 (N_1480,In_381,In_512);
xor U1481 (N_1481,In_702,In_463);
xor U1482 (N_1482,In_752,In_374);
or U1483 (N_1483,In_361,In_643);
xnor U1484 (N_1484,In_82,In_747);
or U1485 (N_1485,In_540,In_245);
and U1486 (N_1486,In_761,In_668);
xnor U1487 (N_1487,In_789,In_927);
nor U1488 (N_1488,In_603,In_353);
xor U1489 (N_1489,In_650,In_847);
xnor U1490 (N_1490,In_340,In_874);
nand U1491 (N_1491,In_58,In_970);
nor U1492 (N_1492,In_475,In_626);
or U1493 (N_1493,In_867,In_17);
nor U1494 (N_1494,In_456,In_683);
xnor U1495 (N_1495,In_895,In_916);
nand U1496 (N_1496,In_197,In_506);
or U1497 (N_1497,In_990,In_883);
xor U1498 (N_1498,In_821,In_343);
xor U1499 (N_1499,In_944,In_941);
xor U1500 (N_1500,In_220,In_357);
and U1501 (N_1501,In_557,In_597);
nand U1502 (N_1502,In_638,In_455);
nand U1503 (N_1503,In_411,In_199);
and U1504 (N_1504,In_517,In_368);
nand U1505 (N_1505,In_787,In_798);
nand U1506 (N_1506,In_767,In_682);
and U1507 (N_1507,In_449,In_589);
nand U1508 (N_1508,In_265,In_619);
nor U1509 (N_1509,In_106,In_356);
and U1510 (N_1510,In_875,In_480);
and U1511 (N_1511,In_940,In_131);
and U1512 (N_1512,In_815,In_211);
nand U1513 (N_1513,In_64,In_531);
nand U1514 (N_1514,In_665,In_661);
and U1515 (N_1515,In_480,In_150);
or U1516 (N_1516,In_214,In_746);
or U1517 (N_1517,In_168,In_730);
xnor U1518 (N_1518,In_442,In_626);
nor U1519 (N_1519,In_408,In_686);
xnor U1520 (N_1520,In_786,In_360);
and U1521 (N_1521,In_216,In_781);
or U1522 (N_1522,In_854,In_270);
nand U1523 (N_1523,In_654,In_964);
and U1524 (N_1524,In_965,In_845);
and U1525 (N_1525,In_64,In_615);
or U1526 (N_1526,In_626,In_610);
xnor U1527 (N_1527,In_652,In_950);
and U1528 (N_1528,In_66,In_351);
xor U1529 (N_1529,In_354,In_440);
nor U1530 (N_1530,In_697,In_572);
nor U1531 (N_1531,In_463,In_756);
nand U1532 (N_1532,In_136,In_83);
nand U1533 (N_1533,In_791,In_508);
nor U1534 (N_1534,In_714,In_450);
nand U1535 (N_1535,In_531,In_698);
xor U1536 (N_1536,In_230,In_673);
nor U1537 (N_1537,In_715,In_824);
nand U1538 (N_1538,In_407,In_633);
nor U1539 (N_1539,In_721,In_344);
nand U1540 (N_1540,In_519,In_968);
nor U1541 (N_1541,In_402,In_257);
nand U1542 (N_1542,In_524,In_945);
nand U1543 (N_1543,In_50,In_280);
xor U1544 (N_1544,In_803,In_824);
and U1545 (N_1545,In_208,In_690);
nand U1546 (N_1546,In_295,In_514);
nand U1547 (N_1547,In_512,In_959);
and U1548 (N_1548,In_441,In_1);
nand U1549 (N_1549,In_82,In_695);
or U1550 (N_1550,In_246,In_69);
xor U1551 (N_1551,In_709,In_892);
or U1552 (N_1552,In_676,In_660);
nor U1553 (N_1553,In_321,In_397);
nor U1554 (N_1554,In_533,In_245);
xnor U1555 (N_1555,In_935,In_163);
xnor U1556 (N_1556,In_874,In_392);
nand U1557 (N_1557,In_778,In_351);
xor U1558 (N_1558,In_970,In_948);
nand U1559 (N_1559,In_751,In_528);
nand U1560 (N_1560,In_10,In_289);
xnor U1561 (N_1561,In_391,In_538);
or U1562 (N_1562,In_773,In_907);
or U1563 (N_1563,In_516,In_74);
nand U1564 (N_1564,In_245,In_76);
xor U1565 (N_1565,In_839,In_51);
or U1566 (N_1566,In_823,In_404);
or U1567 (N_1567,In_822,In_360);
nand U1568 (N_1568,In_495,In_241);
xor U1569 (N_1569,In_809,In_607);
and U1570 (N_1570,In_896,In_219);
nor U1571 (N_1571,In_834,In_591);
nand U1572 (N_1572,In_69,In_11);
nand U1573 (N_1573,In_884,In_121);
xnor U1574 (N_1574,In_384,In_737);
or U1575 (N_1575,In_139,In_674);
nor U1576 (N_1576,In_692,In_589);
xnor U1577 (N_1577,In_78,In_282);
and U1578 (N_1578,In_432,In_610);
xor U1579 (N_1579,In_569,In_651);
nand U1580 (N_1580,In_532,In_761);
and U1581 (N_1581,In_28,In_701);
and U1582 (N_1582,In_442,In_636);
or U1583 (N_1583,In_135,In_564);
xnor U1584 (N_1584,In_159,In_491);
xor U1585 (N_1585,In_100,In_884);
nand U1586 (N_1586,In_960,In_688);
and U1587 (N_1587,In_696,In_41);
and U1588 (N_1588,In_532,In_902);
or U1589 (N_1589,In_705,In_324);
nor U1590 (N_1590,In_746,In_717);
and U1591 (N_1591,In_362,In_980);
and U1592 (N_1592,In_459,In_474);
xnor U1593 (N_1593,In_163,In_160);
and U1594 (N_1594,In_775,In_569);
nand U1595 (N_1595,In_175,In_394);
and U1596 (N_1596,In_277,In_449);
nor U1597 (N_1597,In_164,In_432);
or U1598 (N_1598,In_346,In_868);
and U1599 (N_1599,In_299,In_379);
nor U1600 (N_1600,In_643,In_788);
or U1601 (N_1601,In_735,In_83);
nand U1602 (N_1602,In_634,In_368);
nand U1603 (N_1603,In_435,In_487);
xor U1604 (N_1604,In_885,In_704);
xor U1605 (N_1605,In_80,In_499);
nor U1606 (N_1606,In_941,In_221);
or U1607 (N_1607,In_550,In_559);
or U1608 (N_1608,In_291,In_564);
nand U1609 (N_1609,In_560,In_184);
and U1610 (N_1610,In_516,In_601);
or U1611 (N_1611,In_256,In_129);
and U1612 (N_1612,In_624,In_40);
and U1613 (N_1613,In_968,In_473);
nor U1614 (N_1614,In_67,In_376);
nand U1615 (N_1615,In_117,In_510);
nor U1616 (N_1616,In_903,In_210);
and U1617 (N_1617,In_460,In_423);
or U1618 (N_1618,In_678,In_997);
nand U1619 (N_1619,In_988,In_740);
or U1620 (N_1620,In_390,In_902);
nand U1621 (N_1621,In_548,In_417);
nor U1622 (N_1622,In_482,In_64);
and U1623 (N_1623,In_315,In_831);
and U1624 (N_1624,In_475,In_155);
xor U1625 (N_1625,In_479,In_78);
xor U1626 (N_1626,In_450,In_98);
or U1627 (N_1627,In_135,In_537);
nand U1628 (N_1628,In_91,In_462);
nand U1629 (N_1629,In_182,In_200);
or U1630 (N_1630,In_137,In_575);
and U1631 (N_1631,In_732,In_102);
nor U1632 (N_1632,In_511,In_51);
nand U1633 (N_1633,In_8,In_56);
nand U1634 (N_1634,In_129,In_777);
nor U1635 (N_1635,In_210,In_401);
nor U1636 (N_1636,In_983,In_624);
and U1637 (N_1637,In_932,In_494);
xor U1638 (N_1638,In_786,In_561);
nand U1639 (N_1639,In_69,In_687);
xnor U1640 (N_1640,In_710,In_69);
or U1641 (N_1641,In_314,In_207);
or U1642 (N_1642,In_525,In_470);
nor U1643 (N_1643,In_721,In_210);
nor U1644 (N_1644,In_770,In_652);
and U1645 (N_1645,In_475,In_823);
xnor U1646 (N_1646,In_735,In_66);
and U1647 (N_1647,In_162,In_443);
nand U1648 (N_1648,In_380,In_583);
nor U1649 (N_1649,In_253,In_280);
nand U1650 (N_1650,In_9,In_551);
xnor U1651 (N_1651,In_751,In_638);
nand U1652 (N_1652,In_725,In_623);
nor U1653 (N_1653,In_930,In_458);
nor U1654 (N_1654,In_324,In_172);
xnor U1655 (N_1655,In_59,In_256);
and U1656 (N_1656,In_568,In_900);
nand U1657 (N_1657,In_375,In_141);
nand U1658 (N_1658,In_421,In_369);
nor U1659 (N_1659,In_102,In_600);
nor U1660 (N_1660,In_532,In_132);
nor U1661 (N_1661,In_134,In_523);
nand U1662 (N_1662,In_752,In_646);
or U1663 (N_1663,In_535,In_500);
nand U1664 (N_1664,In_56,In_668);
or U1665 (N_1665,In_159,In_655);
nand U1666 (N_1666,In_338,In_948);
nand U1667 (N_1667,In_926,In_475);
or U1668 (N_1668,In_93,In_367);
and U1669 (N_1669,In_692,In_743);
nor U1670 (N_1670,In_637,In_276);
and U1671 (N_1671,In_916,In_291);
nand U1672 (N_1672,In_927,In_313);
nor U1673 (N_1673,In_162,In_786);
xnor U1674 (N_1674,In_198,In_734);
nor U1675 (N_1675,In_18,In_651);
and U1676 (N_1676,In_246,In_877);
xor U1677 (N_1677,In_778,In_692);
and U1678 (N_1678,In_668,In_855);
or U1679 (N_1679,In_5,In_459);
or U1680 (N_1680,In_444,In_438);
xnor U1681 (N_1681,In_591,In_347);
nand U1682 (N_1682,In_217,In_193);
and U1683 (N_1683,In_457,In_284);
nand U1684 (N_1684,In_70,In_613);
and U1685 (N_1685,In_360,In_133);
nor U1686 (N_1686,In_69,In_832);
xnor U1687 (N_1687,In_360,In_285);
and U1688 (N_1688,In_38,In_240);
nor U1689 (N_1689,In_983,In_66);
nor U1690 (N_1690,In_681,In_630);
or U1691 (N_1691,In_966,In_345);
nor U1692 (N_1692,In_378,In_956);
or U1693 (N_1693,In_736,In_837);
xor U1694 (N_1694,In_702,In_942);
xor U1695 (N_1695,In_158,In_172);
xor U1696 (N_1696,In_220,In_317);
xnor U1697 (N_1697,In_333,In_217);
and U1698 (N_1698,In_684,In_477);
nor U1699 (N_1699,In_349,In_379);
and U1700 (N_1700,In_349,In_157);
nor U1701 (N_1701,In_233,In_116);
nand U1702 (N_1702,In_328,In_598);
nor U1703 (N_1703,In_592,In_480);
and U1704 (N_1704,In_79,In_322);
or U1705 (N_1705,In_506,In_41);
and U1706 (N_1706,In_999,In_124);
nand U1707 (N_1707,In_892,In_451);
and U1708 (N_1708,In_980,In_666);
or U1709 (N_1709,In_162,In_446);
and U1710 (N_1710,In_19,In_526);
xnor U1711 (N_1711,In_388,In_239);
xnor U1712 (N_1712,In_7,In_724);
and U1713 (N_1713,In_854,In_544);
or U1714 (N_1714,In_857,In_25);
and U1715 (N_1715,In_13,In_376);
xnor U1716 (N_1716,In_914,In_704);
nand U1717 (N_1717,In_507,In_303);
nor U1718 (N_1718,In_212,In_285);
xor U1719 (N_1719,In_524,In_917);
xnor U1720 (N_1720,In_17,In_416);
or U1721 (N_1721,In_124,In_912);
or U1722 (N_1722,In_784,In_867);
nor U1723 (N_1723,In_94,In_111);
xnor U1724 (N_1724,In_384,In_374);
xor U1725 (N_1725,In_473,In_721);
or U1726 (N_1726,In_406,In_798);
and U1727 (N_1727,In_512,In_944);
xnor U1728 (N_1728,In_304,In_216);
and U1729 (N_1729,In_538,In_792);
nor U1730 (N_1730,In_722,In_20);
nand U1731 (N_1731,In_603,In_919);
xor U1732 (N_1732,In_966,In_901);
or U1733 (N_1733,In_737,In_352);
or U1734 (N_1734,In_654,In_425);
or U1735 (N_1735,In_811,In_364);
and U1736 (N_1736,In_60,In_276);
or U1737 (N_1737,In_397,In_268);
nand U1738 (N_1738,In_984,In_531);
or U1739 (N_1739,In_817,In_630);
or U1740 (N_1740,In_289,In_378);
or U1741 (N_1741,In_824,In_258);
xor U1742 (N_1742,In_766,In_313);
nor U1743 (N_1743,In_368,In_444);
xnor U1744 (N_1744,In_900,In_318);
nor U1745 (N_1745,In_737,In_584);
and U1746 (N_1746,In_625,In_776);
nor U1747 (N_1747,In_580,In_535);
and U1748 (N_1748,In_971,In_567);
nand U1749 (N_1749,In_704,In_960);
nand U1750 (N_1750,In_622,In_313);
nand U1751 (N_1751,In_728,In_446);
or U1752 (N_1752,In_384,In_91);
or U1753 (N_1753,In_991,In_527);
xnor U1754 (N_1754,In_240,In_42);
and U1755 (N_1755,In_378,In_722);
xor U1756 (N_1756,In_460,In_544);
nand U1757 (N_1757,In_843,In_754);
nor U1758 (N_1758,In_437,In_115);
xor U1759 (N_1759,In_496,In_873);
and U1760 (N_1760,In_821,In_817);
nand U1761 (N_1761,In_148,In_484);
xnor U1762 (N_1762,In_692,In_780);
and U1763 (N_1763,In_632,In_680);
or U1764 (N_1764,In_176,In_470);
or U1765 (N_1765,In_548,In_116);
nand U1766 (N_1766,In_762,In_632);
nor U1767 (N_1767,In_960,In_730);
nor U1768 (N_1768,In_113,In_349);
and U1769 (N_1769,In_87,In_566);
nand U1770 (N_1770,In_923,In_27);
nor U1771 (N_1771,In_191,In_724);
nor U1772 (N_1772,In_198,In_53);
or U1773 (N_1773,In_391,In_20);
and U1774 (N_1774,In_846,In_498);
nand U1775 (N_1775,In_104,In_852);
or U1776 (N_1776,In_287,In_999);
nand U1777 (N_1777,In_205,In_579);
nor U1778 (N_1778,In_262,In_946);
nand U1779 (N_1779,In_268,In_386);
or U1780 (N_1780,In_848,In_280);
nand U1781 (N_1781,In_595,In_792);
xor U1782 (N_1782,In_118,In_280);
and U1783 (N_1783,In_916,In_947);
xor U1784 (N_1784,In_72,In_583);
nand U1785 (N_1785,In_446,In_854);
or U1786 (N_1786,In_981,In_553);
xnor U1787 (N_1787,In_525,In_555);
nor U1788 (N_1788,In_754,In_991);
or U1789 (N_1789,In_564,In_255);
nor U1790 (N_1790,In_430,In_973);
xnor U1791 (N_1791,In_830,In_623);
and U1792 (N_1792,In_960,In_506);
or U1793 (N_1793,In_633,In_238);
or U1794 (N_1794,In_662,In_999);
xnor U1795 (N_1795,In_58,In_553);
nand U1796 (N_1796,In_22,In_689);
and U1797 (N_1797,In_248,In_876);
nand U1798 (N_1798,In_81,In_292);
nand U1799 (N_1799,In_427,In_962);
and U1800 (N_1800,In_181,In_517);
xnor U1801 (N_1801,In_738,In_638);
or U1802 (N_1802,In_130,In_68);
nor U1803 (N_1803,In_945,In_406);
nand U1804 (N_1804,In_796,In_187);
nand U1805 (N_1805,In_306,In_223);
and U1806 (N_1806,In_625,In_371);
and U1807 (N_1807,In_685,In_606);
xor U1808 (N_1808,In_172,In_480);
or U1809 (N_1809,In_516,In_962);
nand U1810 (N_1810,In_124,In_858);
and U1811 (N_1811,In_68,In_73);
and U1812 (N_1812,In_866,In_688);
nor U1813 (N_1813,In_447,In_805);
nand U1814 (N_1814,In_30,In_845);
or U1815 (N_1815,In_137,In_174);
nand U1816 (N_1816,In_938,In_378);
nand U1817 (N_1817,In_172,In_76);
nor U1818 (N_1818,In_167,In_263);
xor U1819 (N_1819,In_136,In_826);
xor U1820 (N_1820,In_840,In_150);
xnor U1821 (N_1821,In_163,In_602);
and U1822 (N_1822,In_440,In_660);
or U1823 (N_1823,In_95,In_199);
nor U1824 (N_1824,In_176,In_181);
nor U1825 (N_1825,In_847,In_128);
xor U1826 (N_1826,In_55,In_963);
nand U1827 (N_1827,In_375,In_550);
nor U1828 (N_1828,In_530,In_171);
nand U1829 (N_1829,In_343,In_739);
and U1830 (N_1830,In_442,In_251);
nor U1831 (N_1831,In_820,In_2);
or U1832 (N_1832,In_260,In_810);
xnor U1833 (N_1833,In_6,In_28);
nand U1834 (N_1834,In_695,In_461);
and U1835 (N_1835,In_835,In_684);
nor U1836 (N_1836,In_95,In_966);
xnor U1837 (N_1837,In_454,In_473);
nor U1838 (N_1838,In_427,In_613);
nand U1839 (N_1839,In_411,In_494);
or U1840 (N_1840,In_321,In_731);
xor U1841 (N_1841,In_900,In_320);
and U1842 (N_1842,In_48,In_798);
nor U1843 (N_1843,In_32,In_784);
and U1844 (N_1844,In_442,In_301);
or U1845 (N_1845,In_929,In_106);
nand U1846 (N_1846,In_356,In_973);
nor U1847 (N_1847,In_994,In_193);
and U1848 (N_1848,In_680,In_851);
nor U1849 (N_1849,In_392,In_544);
nand U1850 (N_1850,In_745,In_272);
xnor U1851 (N_1851,In_683,In_336);
and U1852 (N_1852,In_708,In_189);
nand U1853 (N_1853,In_330,In_474);
xor U1854 (N_1854,In_62,In_617);
nand U1855 (N_1855,In_927,In_742);
nand U1856 (N_1856,In_137,In_38);
and U1857 (N_1857,In_681,In_227);
nand U1858 (N_1858,In_43,In_156);
or U1859 (N_1859,In_52,In_912);
xnor U1860 (N_1860,In_809,In_211);
and U1861 (N_1861,In_149,In_658);
nor U1862 (N_1862,In_290,In_352);
or U1863 (N_1863,In_833,In_170);
and U1864 (N_1864,In_751,In_722);
or U1865 (N_1865,In_330,In_509);
nor U1866 (N_1866,In_987,In_648);
or U1867 (N_1867,In_469,In_254);
xor U1868 (N_1868,In_617,In_906);
xor U1869 (N_1869,In_939,In_837);
and U1870 (N_1870,In_999,In_869);
nor U1871 (N_1871,In_100,In_440);
xnor U1872 (N_1872,In_410,In_675);
nor U1873 (N_1873,In_433,In_679);
nand U1874 (N_1874,In_196,In_663);
or U1875 (N_1875,In_943,In_408);
or U1876 (N_1876,In_527,In_712);
nor U1877 (N_1877,In_886,In_902);
nand U1878 (N_1878,In_786,In_977);
or U1879 (N_1879,In_939,In_895);
xor U1880 (N_1880,In_197,In_940);
nor U1881 (N_1881,In_925,In_441);
xor U1882 (N_1882,In_57,In_534);
nand U1883 (N_1883,In_334,In_658);
or U1884 (N_1884,In_807,In_14);
nand U1885 (N_1885,In_536,In_243);
or U1886 (N_1886,In_400,In_111);
xnor U1887 (N_1887,In_585,In_892);
or U1888 (N_1888,In_894,In_70);
or U1889 (N_1889,In_691,In_712);
and U1890 (N_1890,In_193,In_934);
and U1891 (N_1891,In_447,In_858);
and U1892 (N_1892,In_259,In_86);
nor U1893 (N_1893,In_984,In_115);
and U1894 (N_1894,In_741,In_68);
xnor U1895 (N_1895,In_593,In_281);
xor U1896 (N_1896,In_141,In_307);
and U1897 (N_1897,In_226,In_13);
xor U1898 (N_1898,In_137,In_345);
nand U1899 (N_1899,In_462,In_22);
or U1900 (N_1900,In_733,In_931);
nor U1901 (N_1901,In_901,In_307);
xor U1902 (N_1902,In_652,In_846);
nand U1903 (N_1903,In_551,In_333);
and U1904 (N_1904,In_632,In_492);
xnor U1905 (N_1905,In_555,In_895);
or U1906 (N_1906,In_472,In_948);
nor U1907 (N_1907,In_641,In_570);
or U1908 (N_1908,In_942,In_972);
and U1909 (N_1909,In_619,In_362);
xnor U1910 (N_1910,In_327,In_959);
or U1911 (N_1911,In_16,In_916);
and U1912 (N_1912,In_110,In_657);
and U1913 (N_1913,In_423,In_482);
nor U1914 (N_1914,In_718,In_469);
nor U1915 (N_1915,In_633,In_939);
xor U1916 (N_1916,In_919,In_184);
nor U1917 (N_1917,In_372,In_286);
nand U1918 (N_1918,In_74,In_504);
nor U1919 (N_1919,In_152,In_723);
and U1920 (N_1920,In_840,In_752);
xnor U1921 (N_1921,In_667,In_919);
and U1922 (N_1922,In_337,In_627);
nand U1923 (N_1923,In_320,In_83);
nand U1924 (N_1924,In_680,In_724);
nand U1925 (N_1925,In_587,In_25);
nor U1926 (N_1926,In_155,In_451);
nor U1927 (N_1927,In_138,In_824);
or U1928 (N_1928,In_985,In_209);
and U1929 (N_1929,In_453,In_443);
xnor U1930 (N_1930,In_196,In_873);
or U1931 (N_1931,In_191,In_572);
xor U1932 (N_1932,In_175,In_354);
nand U1933 (N_1933,In_590,In_575);
nand U1934 (N_1934,In_386,In_86);
and U1935 (N_1935,In_769,In_312);
xor U1936 (N_1936,In_200,In_509);
nand U1937 (N_1937,In_73,In_226);
nor U1938 (N_1938,In_475,In_465);
xor U1939 (N_1939,In_562,In_505);
or U1940 (N_1940,In_950,In_437);
nor U1941 (N_1941,In_785,In_731);
and U1942 (N_1942,In_717,In_136);
nand U1943 (N_1943,In_957,In_522);
and U1944 (N_1944,In_984,In_51);
nand U1945 (N_1945,In_236,In_820);
and U1946 (N_1946,In_600,In_222);
nor U1947 (N_1947,In_24,In_161);
or U1948 (N_1948,In_418,In_864);
xor U1949 (N_1949,In_655,In_122);
xnor U1950 (N_1950,In_224,In_516);
nor U1951 (N_1951,In_426,In_369);
and U1952 (N_1952,In_588,In_231);
xor U1953 (N_1953,In_706,In_561);
or U1954 (N_1954,In_352,In_631);
or U1955 (N_1955,In_379,In_461);
and U1956 (N_1956,In_5,In_304);
xnor U1957 (N_1957,In_415,In_773);
nand U1958 (N_1958,In_235,In_729);
nand U1959 (N_1959,In_412,In_138);
nor U1960 (N_1960,In_951,In_217);
and U1961 (N_1961,In_592,In_339);
xor U1962 (N_1962,In_22,In_487);
nand U1963 (N_1963,In_391,In_333);
xnor U1964 (N_1964,In_535,In_625);
xnor U1965 (N_1965,In_71,In_813);
and U1966 (N_1966,In_565,In_304);
nand U1967 (N_1967,In_483,In_116);
nand U1968 (N_1968,In_692,In_928);
nor U1969 (N_1969,In_701,In_488);
or U1970 (N_1970,In_120,In_584);
nand U1971 (N_1971,In_239,In_947);
xor U1972 (N_1972,In_433,In_123);
nor U1973 (N_1973,In_377,In_28);
and U1974 (N_1974,In_672,In_180);
and U1975 (N_1975,In_13,In_648);
xnor U1976 (N_1976,In_162,In_800);
nor U1977 (N_1977,In_680,In_622);
or U1978 (N_1978,In_828,In_228);
xnor U1979 (N_1979,In_756,In_575);
or U1980 (N_1980,In_34,In_594);
nand U1981 (N_1981,In_803,In_408);
xnor U1982 (N_1982,In_45,In_917);
or U1983 (N_1983,In_420,In_706);
xor U1984 (N_1984,In_125,In_143);
xor U1985 (N_1985,In_579,In_886);
and U1986 (N_1986,In_626,In_9);
nand U1987 (N_1987,In_967,In_199);
or U1988 (N_1988,In_190,In_607);
nand U1989 (N_1989,In_803,In_27);
and U1990 (N_1990,In_67,In_383);
xnor U1991 (N_1991,In_36,In_203);
and U1992 (N_1992,In_868,In_648);
nor U1993 (N_1993,In_520,In_910);
and U1994 (N_1994,In_966,In_952);
and U1995 (N_1995,In_804,In_3);
or U1996 (N_1996,In_985,In_139);
nand U1997 (N_1997,In_183,In_407);
xnor U1998 (N_1998,In_61,In_708);
nor U1999 (N_1999,In_829,In_360);
nand U2000 (N_2000,In_602,In_6);
nor U2001 (N_2001,In_640,In_719);
or U2002 (N_2002,In_419,In_763);
nor U2003 (N_2003,In_203,In_419);
nor U2004 (N_2004,In_523,In_522);
nand U2005 (N_2005,In_765,In_664);
or U2006 (N_2006,In_383,In_763);
nand U2007 (N_2007,In_999,In_534);
nand U2008 (N_2008,In_79,In_353);
nand U2009 (N_2009,In_178,In_516);
xnor U2010 (N_2010,In_860,In_294);
xnor U2011 (N_2011,In_365,In_54);
nand U2012 (N_2012,In_789,In_268);
nand U2013 (N_2013,In_62,In_602);
nor U2014 (N_2014,In_869,In_759);
nor U2015 (N_2015,In_256,In_281);
or U2016 (N_2016,In_58,In_221);
nand U2017 (N_2017,In_15,In_443);
nand U2018 (N_2018,In_693,In_139);
nor U2019 (N_2019,In_933,In_157);
nand U2020 (N_2020,In_738,In_578);
or U2021 (N_2021,In_456,In_441);
nor U2022 (N_2022,In_398,In_519);
xnor U2023 (N_2023,In_252,In_998);
nor U2024 (N_2024,In_113,In_243);
and U2025 (N_2025,In_717,In_766);
nor U2026 (N_2026,In_445,In_497);
nand U2027 (N_2027,In_489,In_149);
nor U2028 (N_2028,In_525,In_17);
xnor U2029 (N_2029,In_57,In_742);
and U2030 (N_2030,In_477,In_552);
nand U2031 (N_2031,In_961,In_548);
or U2032 (N_2032,In_556,In_462);
nand U2033 (N_2033,In_966,In_46);
nor U2034 (N_2034,In_997,In_503);
and U2035 (N_2035,In_707,In_61);
nand U2036 (N_2036,In_640,In_820);
nand U2037 (N_2037,In_118,In_781);
nor U2038 (N_2038,In_592,In_768);
xor U2039 (N_2039,In_555,In_646);
or U2040 (N_2040,In_908,In_909);
and U2041 (N_2041,In_402,In_771);
nor U2042 (N_2042,In_948,In_146);
or U2043 (N_2043,In_259,In_729);
and U2044 (N_2044,In_798,In_280);
nand U2045 (N_2045,In_755,In_888);
or U2046 (N_2046,In_652,In_113);
or U2047 (N_2047,In_9,In_501);
nand U2048 (N_2048,In_386,In_489);
and U2049 (N_2049,In_144,In_963);
or U2050 (N_2050,In_241,In_704);
xor U2051 (N_2051,In_727,In_73);
nor U2052 (N_2052,In_338,In_353);
and U2053 (N_2053,In_318,In_218);
or U2054 (N_2054,In_447,In_892);
nand U2055 (N_2055,In_120,In_707);
or U2056 (N_2056,In_349,In_14);
xnor U2057 (N_2057,In_90,In_764);
nand U2058 (N_2058,In_44,In_690);
or U2059 (N_2059,In_272,In_394);
nand U2060 (N_2060,In_401,In_939);
nor U2061 (N_2061,In_205,In_161);
or U2062 (N_2062,In_19,In_778);
nor U2063 (N_2063,In_60,In_129);
or U2064 (N_2064,In_197,In_86);
and U2065 (N_2065,In_394,In_879);
or U2066 (N_2066,In_858,In_889);
or U2067 (N_2067,In_325,In_479);
and U2068 (N_2068,In_123,In_325);
nand U2069 (N_2069,In_275,In_250);
nor U2070 (N_2070,In_787,In_320);
or U2071 (N_2071,In_765,In_689);
and U2072 (N_2072,In_469,In_273);
nor U2073 (N_2073,In_45,In_291);
nor U2074 (N_2074,In_603,In_328);
or U2075 (N_2075,In_546,In_735);
or U2076 (N_2076,In_173,In_620);
or U2077 (N_2077,In_289,In_629);
nand U2078 (N_2078,In_879,In_740);
xnor U2079 (N_2079,In_397,In_754);
or U2080 (N_2080,In_263,In_269);
nor U2081 (N_2081,In_443,In_759);
nor U2082 (N_2082,In_251,In_533);
nand U2083 (N_2083,In_756,In_797);
and U2084 (N_2084,In_204,In_130);
nand U2085 (N_2085,In_577,In_805);
and U2086 (N_2086,In_957,In_967);
xnor U2087 (N_2087,In_739,In_746);
and U2088 (N_2088,In_49,In_90);
or U2089 (N_2089,In_609,In_863);
xnor U2090 (N_2090,In_882,In_528);
or U2091 (N_2091,In_538,In_836);
nand U2092 (N_2092,In_263,In_606);
nand U2093 (N_2093,In_120,In_863);
and U2094 (N_2094,In_84,In_592);
xor U2095 (N_2095,In_105,In_979);
or U2096 (N_2096,In_543,In_568);
and U2097 (N_2097,In_411,In_861);
or U2098 (N_2098,In_86,In_193);
and U2099 (N_2099,In_394,In_569);
and U2100 (N_2100,In_645,In_564);
nand U2101 (N_2101,In_594,In_437);
nand U2102 (N_2102,In_938,In_699);
nor U2103 (N_2103,In_89,In_646);
nand U2104 (N_2104,In_138,In_75);
or U2105 (N_2105,In_533,In_133);
nand U2106 (N_2106,In_334,In_363);
nor U2107 (N_2107,In_987,In_967);
and U2108 (N_2108,In_227,In_542);
and U2109 (N_2109,In_142,In_85);
nor U2110 (N_2110,In_122,In_296);
nand U2111 (N_2111,In_68,In_39);
and U2112 (N_2112,In_468,In_16);
xor U2113 (N_2113,In_351,In_381);
xor U2114 (N_2114,In_267,In_245);
and U2115 (N_2115,In_933,In_348);
nand U2116 (N_2116,In_793,In_941);
and U2117 (N_2117,In_678,In_265);
nor U2118 (N_2118,In_331,In_949);
or U2119 (N_2119,In_789,In_650);
nand U2120 (N_2120,In_540,In_417);
or U2121 (N_2121,In_152,In_186);
nand U2122 (N_2122,In_133,In_775);
nor U2123 (N_2123,In_95,In_904);
nand U2124 (N_2124,In_868,In_423);
and U2125 (N_2125,In_310,In_962);
nor U2126 (N_2126,In_99,In_722);
nand U2127 (N_2127,In_837,In_280);
nand U2128 (N_2128,In_156,In_3);
nor U2129 (N_2129,In_474,In_80);
xnor U2130 (N_2130,In_913,In_176);
nor U2131 (N_2131,In_222,In_122);
nor U2132 (N_2132,In_746,In_384);
nor U2133 (N_2133,In_586,In_600);
nor U2134 (N_2134,In_31,In_772);
nand U2135 (N_2135,In_294,In_34);
nand U2136 (N_2136,In_632,In_719);
or U2137 (N_2137,In_466,In_817);
or U2138 (N_2138,In_876,In_587);
and U2139 (N_2139,In_90,In_923);
nand U2140 (N_2140,In_341,In_122);
xnor U2141 (N_2141,In_445,In_481);
xor U2142 (N_2142,In_876,In_660);
nor U2143 (N_2143,In_459,In_151);
nor U2144 (N_2144,In_946,In_461);
nor U2145 (N_2145,In_926,In_705);
xnor U2146 (N_2146,In_951,In_364);
or U2147 (N_2147,In_723,In_33);
xor U2148 (N_2148,In_191,In_309);
nand U2149 (N_2149,In_821,In_165);
nand U2150 (N_2150,In_202,In_401);
nand U2151 (N_2151,In_115,In_213);
or U2152 (N_2152,In_298,In_500);
nand U2153 (N_2153,In_884,In_54);
nor U2154 (N_2154,In_482,In_812);
xor U2155 (N_2155,In_332,In_892);
xor U2156 (N_2156,In_765,In_714);
nand U2157 (N_2157,In_914,In_618);
xor U2158 (N_2158,In_220,In_20);
xor U2159 (N_2159,In_817,In_233);
nor U2160 (N_2160,In_601,In_462);
nor U2161 (N_2161,In_383,In_933);
or U2162 (N_2162,In_785,In_265);
nand U2163 (N_2163,In_359,In_89);
and U2164 (N_2164,In_812,In_837);
or U2165 (N_2165,In_370,In_580);
and U2166 (N_2166,In_871,In_250);
or U2167 (N_2167,In_958,In_497);
xor U2168 (N_2168,In_124,In_337);
nor U2169 (N_2169,In_647,In_152);
nand U2170 (N_2170,In_42,In_894);
or U2171 (N_2171,In_372,In_687);
nand U2172 (N_2172,In_684,In_460);
xor U2173 (N_2173,In_49,In_862);
xor U2174 (N_2174,In_964,In_679);
or U2175 (N_2175,In_663,In_905);
nor U2176 (N_2176,In_27,In_325);
and U2177 (N_2177,In_616,In_369);
nor U2178 (N_2178,In_566,In_1);
xnor U2179 (N_2179,In_143,In_139);
and U2180 (N_2180,In_630,In_927);
nor U2181 (N_2181,In_199,In_740);
nor U2182 (N_2182,In_512,In_613);
nand U2183 (N_2183,In_954,In_489);
nor U2184 (N_2184,In_416,In_83);
xor U2185 (N_2185,In_516,In_665);
and U2186 (N_2186,In_652,In_532);
nor U2187 (N_2187,In_220,In_262);
or U2188 (N_2188,In_514,In_593);
nor U2189 (N_2189,In_877,In_482);
xor U2190 (N_2190,In_439,In_205);
nand U2191 (N_2191,In_615,In_429);
nor U2192 (N_2192,In_750,In_173);
nand U2193 (N_2193,In_907,In_375);
nand U2194 (N_2194,In_37,In_617);
nor U2195 (N_2195,In_837,In_789);
nand U2196 (N_2196,In_309,In_874);
and U2197 (N_2197,In_227,In_208);
xor U2198 (N_2198,In_799,In_647);
and U2199 (N_2199,In_572,In_566);
nand U2200 (N_2200,In_981,In_756);
nand U2201 (N_2201,In_897,In_844);
nor U2202 (N_2202,In_7,In_464);
nand U2203 (N_2203,In_28,In_660);
and U2204 (N_2204,In_227,In_32);
nand U2205 (N_2205,In_903,In_143);
nor U2206 (N_2206,In_27,In_824);
or U2207 (N_2207,In_879,In_385);
nor U2208 (N_2208,In_880,In_338);
or U2209 (N_2209,In_827,In_978);
xnor U2210 (N_2210,In_206,In_56);
xnor U2211 (N_2211,In_7,In_767);
xor U2212 (N_2212,In_691,In_227);
xnor U2213 (N_2213,In_829,In_894);
or U2214 (N_2214,In_110,In_471);
nand U2215 (N_2215,In_999,In_277);
or U2216 (N_2216,In_443,In_101);
nor U2217 (N_2217,In_559,In_353);
and U2218 (N_2218,In_875,In_258);
and U2219 (N_2219,In_534,In_532);
nand U2220 (N_2220,In_333,In_565);
and U2221 (N_2221,In_263,In_61);
and U2222 (N_2222,In_445,In_599);
nand U2223 (N_2223,In_349,In_445);
xnor U2224 (N_2224,In_908,In_325);
and U2225 (N_2225,In_453,In_268);
nand U2226 (N_2226,In_763,In_528);
nand U2227 (N_2227,In_795,In_282);
xnor U2228 (N_2228,In_971,In_840);
nand U2229 (N_2229,In_385,In_101);
nand U2230 (N_2230,In_288,In_595);
nand U2231 (N_2231,In_771,In_875);
nor U2232 (N_2232,In_420,In_714);
and U2233 (N_2233,In_256,In_642);
xnor U2234 (N_2234,In_403,In_813);
nor U2235 (N_2235,In_701,In_443);
xnor U2236 (N_2236,In_930,In_83);
nor U2237 (N_2237,In_122,In_191);
nand U2238 (N_2238,In_382,In_613);
nor U2239 (N_2239,In_556,In_958);
and U2240 (N_2240,In_77,In_214);
and U2241 (N_2241,In_126,In_489);
nor U2242 (N_2242,In_76,In_7);
xor U2243 (N_2243,In_448,In_243);
nor U2244 (N_2244,In_655,In_547);
nor U2245 (N_2245,In_11,In_559);
and U2246 (N_2246,In_116,In_384);
nor U2247 (N_2247,In_582,In_961);
or U2248 (N_2248,In_334,In_892);
xor U2249 (N_2249,In_279,In_250);
and U2250 (N_2250,In_641,In_863);
and U2251 (N_2251,In_272,In_365);
nor U2252 (N_2252,In_223,In_535);
nand U2253 (N_2253,In_356,In_964);
nand U2254 (N_2254,In_546,In_24);
xor U2255 (N_2255,In_2,In_980);
nor U2256 (N_2256,In_535,In_4);
nor U2257 (N_2257,In_894,In_775);
xnor U2258 (N_2258,In_545,In_926);
nor U2259 (N_2259,In_737,In_248);
and U2260 (N_2260,In_864,In_991);
and U2261 (N_2261,In_521,In_755);
or U2262 (N_2262,In_625,In_624);
xnor U2263 (N_2263,In_4,In_62);
nor U2264 (N_2264,In_672,In_639);
or U2265 (N_2265,In_854,In_597);
nand U2266 (N_2266,In_784,In_64);
or U2267 (N_2267,In_992,In_816);
and U2268 (N_2268,In_500,In_163);
xnor U2269 (N_2269,In_963,In_832);
and U2270 (N_2270,In_516,In_504);
nor U2271 (N_2271,In_37,In_370);
nor U2272 (N_2272,In_365,In_347);
or U2273 (N_2273,In_382,In_878);
nor U2274 (N_2274,In_807,In_767);
nor U2275 (N_2275,In_165,In_666);
nand U2276 (N_2276,In_885,In_124);
or U2277 (N_2277,In_910,In_753);
or U2278 (N_2278,In_518,In_845);
and U2279 (N_2279,In_918,In_115);
nand U2280 (N_2280,In_264,In_716);
nand U2281 (N_2281,In_208,In_435);
and U2282 (N_2282,In_837,In_499);
xor U2283 (N_2283,In_788,In_449);
or U2284 (N_2284,In_753,In_560);
nand U2285 (N_2285,In_395,In_849);
nand U2286 (N_2286,In_188,In_436);
nand U2287 (N_2287,In_148,In_852);
nand U2288 (N_2288,In_288,In_347);
nor U2289 (N_2289,In_132,In_751);
nor U2290 (N_2290,In_434,In_87);
or U2291 (N_2291,In_589,In_81);
and U2292 (N_2292,In_95,In_83);
and U2293 (N_2293,In_430,In_631);
or U2294 (N_2294,In_357,In_366);
or U2295 (N_2295,In_752,In_326);
xor U2296 (N_2296,In_881,In_255);
xor U2297 (N_2297,In_931,In_716);
or U2298 (N_2298,In_34,In_310);
nor U2299 (N_2299,In_267,In_413);
nand U2300 (N_2300,In_865,In_510);
nor U2301 (N_2301,In_151,In_276);
or U2302 (N_2302,In_330,In_205);
xnor U2303 (N_2303,In_107,In_329);
nor U2304 (N_2304,In_189,In_842);
nand U2305 (N_2305,In_680,In_22);
or U2306 (N_2306,In_61,In_225);
nor U2307 (N_2307,In_997,In_323);
nor U2308 (N_2308,In_368,In_124);
nor U2309 (N_2309,In_93,In_828);
nand U2310 (N_2310,In_38,In_940);
or U2311 (N_2311,In_397,In_865);
nor U2312 (N_2312,In_533,In_321);
nor U2313 (N_2313,In_314,In_904);
nor U2314 (N_2314,In_774,In_900);
and U2315 (N_2315,In_5,In_202);
xor U2316 (N_2316,In_181,In_302);
nor U2317 (N_2317,In_597,In_386);
or U2318 (N_2318,In_663,In_123);
nand U2319 (N_2319,In_234,In_628);
or U2320 (N_2320,In_677,In_84);
and U2321 (N_2321,In_899,In_635);
and U2322 (N_2322,In_958,In_396);
nor U2323 (N_2323,In_363,In_472);
or U2324 (N_2324,In_953,In_277);
or U2325 (N_2325,In_449,In_959);
and U2326 (N_2326,In_584,In_748);
nor U2327 (N_2327,In_683,In_439);
or U2328 (N_2328,In_878,In_318);
or U2329 (N_2329,In_233,In_394);
xor U2330 (N_2330,In_882,In_656);
xnor U2331 (N_2331,In_446,In_234);
xor U2332 (N_2332,In_256,In_611);
nand U2333 (N_2333,In_971,In_749);
nand U2334 (N_2334,In_641,In_446);
nand U2335 (N_2335,In_508,In_709);
or U2336 (N_2336,In_207,In_8);
or U2337 (N_2337,In_760,In_39);
nor U2338 (N_2338,In_985,In_505);
or U2339 (N_2339,In_595,In_257);
and U2340 (N_2340,In_717,In_690);
and U2341 (N_2341,In_421,In_961);
nand U2342 (N_2342,In_575,In_303);
and U2343 (N_2343,In_97,In_648);
nor U2344 (N_2344,In_304,In_642);
and U2345 (N_2345,In_511,In_520);
xor U2346 (N_2346,In_741,In_736);
and U2347 (N_2347,In_570,In_241);
nor U2348 (N_2348,In_852,In_611);
xnor U2349 (N_2349,In_95,In_861);
nor U2350 (N_2350,In_142,In_993);
and U2351 (N_2351,In_334,In_821);
nand U2352 (N_2352,In_32,In_106);
xor U2353 (N_2353,In_169,In_621);
and U2354 (N_2354,In_911,In_752);
and U2355 (N_2355,In_142,In_804);
and U2356 (N_2356,In_565,In_818);
nor U2357 (N_2357,In_918,In_507);
and U2358 (N_2358,In_49,In_207);
and U2359 (N_2359,In_783,In_663);
nand U2360 (N_2360,In_814,In_897);
nand U2361 (N_2361,In_827,In_520);
or U2362 (N_2362,In_78,In_390);
xnor U2363 (N_2363,In_371,In_707);
xnor U2364 (N_2364,In_489,In_996);
or U2365 (N_2365,In_247,In_817);
nor U2366 (N_2366,In_711,In_189);
nand U2367 (N_2367,In_241,In_610);
or U2368 (N_2368,In_586,In_493);
nand U2369 (N_2369,In_299,In_335);
or U2370 (N_2370,In_778,In_250);
xor U2371 (N_2371,In_517,In_950);
xnor U2372 (N_2372,In_740,In_219);
xor U2373 (N_2373,In_188,In_817);
xnor U2374 (N_2374,In_384,In_219);
nor U2375 (N_2375,In_836,In_482);
xor U2376 (N_2376,In_669,In_895);
or U2377 (N_2377,In_879,In_856);
nor U2378 (N_2378,In_581,In_507);
xor U2379 (N_2379,In_689,In_620);
nand U2380 (N_2380,In_28,In_554);
or U2381 (N_2381,In_65,In_663);
or U2382 (N_2382,In_97,In_523);
nand U2383 (N_2383,In_613,In_489);
nand U2384 (N_2384,In_389,In_249);
and U2385 (N_2385,In_119,In_330);
nor U2386 (N_2386,In_60,In_207);
or U2387 (N_2387,In_649,In_24);
xnor U2388 (N_2388,In_212,In_845);
nand U2389 (N_2389,In_104,In_357);
nand U2390 (N_2390,In_901,In_280);
or U2391 (N_2391,In_749,In_149);
or U2392 (N_2392,In_353,In_714);
or U2393 (N_2393,In_617,In_217);
nor U2394 (N_2394,In_568,In_744);
nor U2395 (N_2395,In_30,In_745);
or U2396 (N_2396,In_597,In_833);
nor U2397 (N_2397,In_770,In_267);
nand U2398 (N_2398,In_403,In_891);
nor U2399 (N_2399,In_484,In_563);
xnor U2400 (N_2400,In_648,In_15);
nand U2401 (N_2401,In_771,In_408);
or U2402 (N_2402,In_684,In_40);
xor U2403 (N_2403,In_237,In_317);
and U2404 (N_2404,In_856,In_464);
and U2405 (N_2405,In_472,In_910);
nor U2406 (N_2406,In_258,In_891);
xnor U2407 (N_2407,In_861,In_584);
and U2408 (N_2408,In_443,In_149);
nor U2409 (N_2409,In_161,In_428);
xor U2410 (N_2410,In_351,In_681);
xor U2411 (N_2411,In_181,In_265);
and U2412 (N_2412,In_687,In_373);
nand U2413 (N_2413,In_65,In_591);
nor U2414 (N_2414,In_797,In_422);
nand U2415 (N_2415,In_74,In_894);
nand U2416 (N_2416,In_156,In_956);
nand U2417 (N_2417,In_642,In_460);
nor U2418 (N_2418,In_291,In_29);
nand U2419 (N_2419,In_36,In_902);
nor U2420 (N_2420,In_840,In_146);
and U2421 (N_2421,In_593,In_435);
nor U2422 (N_2422,In_766,In_500);
nor U2423 (N_2423,In_101,In_604);
or U2424 (N_2424,In_602,In_37);
nor U2425 (N_2425,In_559,In_47);
and U2426 (N_2426,In_870,In_666);
nor U2427 (N_2427,In_850,In_449);
nor U2428 (N_2428,In_577,In_230);
nand U2429 (N_2429,In_999,In_995);
xor U2430 (N_2430,In_312,In_622);
or U2431 (N_2431,In_898,In_755);
and U2432 (N_2432,In_351,In_37);
or U2433 (N_2433,In_984,In_934);
and U2434 (N_2434,In_409,In_815);
xnor U2435 (N_2435,In_52,In_707);
xor U2436 (N_2436,In_420,In_201);
nand U2437 (N_2437,In_52,In_316);
nand U2438 (N_2438,In_96,In_836);
and U2439 (N_2439,In_116,In_177);
nor U2440 (N_2440,In_568,In_391);
or U2441 (N_2441,In_712,In_651);
nor U2442 (N_2442,In_982,In_140);
and U2443 (N_2443,In_674,In_661);
xor U2444 (N_2444,In_229,In_171);
nand U2445 (N_2445,In_774,In_4);
nand U2446 (N_2446,In_780,In_957);
nand U2447 (N_2447,In_656,In_828);
or U2448 (N_2448,In_659,In_416);
xnor U2449 (N_2449,In_446,In_36);
nand U2450 (N_2450,In_350,In_691);
nand U2451 (N_2451,In_994,In_477);
nand U2452 (N_2452,In_315,In_162);
or U2453 (N_2453,In_121,In_784);
nand U2454 (N_2454,In_548,In_60);
xnor U2455 (N_2455,In_674,In_979);
or U2456 (N_2456,In_617,In_195);
or U2457 (N_2457,In_777,In_270);
and U2458 (N_2458,In_904,In_566);
and U2459 (N_2459,In_745,In_149);
nor U2460 (N_2460,In_75,In_169);
and U2461 (N_2461,In_854,In_345);
and U2462 (N_2462,In_64,In_217);
nor U2463 (N_2463,In_951,In_262);
nor U2464 (N_2464,In_260,In_531);
xor U2465 (N_2465,In_670,In_252);
or U2466 (N_2466,In_901,In_55);
and U2467 (N_2467,In_811,In_806);
nand U2468 (N_2468,In_17,In_824);
nand U2469 (N_2469,In_610,In_386);
and U2470 (N_2470,In_501,In_370);
nor U2471 (N_2471,In_282,In_601);
nand U2472 (N_2472,In_371,In_894);
and U2473 (N_2473,In_642,In_101);
xor U2474 (N_2474,In_348,In_645);
and U2475 (N_2475,In_534,In_739);
xnor U2476 (N_2476,In_18,In_613);
or U2477 (N_2477,In_317,In_769);
nand U2478 (N_2478,In_806,In_912);
or U2479 (N_2479,In_80,In_372);
nand U2480 (N_2480,In_292,In_139);
or U2481 (N_2481,In_766,In_331);
nor U2482 (N_2482,In_797,In_933);
and U2483 (N_2483,In_6,In_669);
nor U2484 (N_2484,In_792,In_228);
or U2485 (N_2485,In_540,In_922);
nor U2486 (N_2486,In_4,In_753);
nand U2487 (N_2487,In_320,In_486);
nand U2488 (N_2488,In_915,In_407);
nand U2489 (N_2489,In_936,In_693);
nand U2490 (N_2490,In_226,In_71);
nor U2491 (N_2491,In_721,In_678);
nand U2492 (N_2492,In_627,In_986);
and U2493 (N_2493,In_281,In_621);
xnor U2494 (N_2494,In_529,In_154);
xor U2495 (N_2495,In_318,In_351);
nor U2496 (N_2496,In_352,In_295);
nand U2497 (N_2497,In_87,In_134);
nor U2498 (N_2498,In_479,In_186);
or U2499 (N_2499,In_23,In_264);
or U2500 (N_2500,N_1303,N_920);
nor U2501 (N_2501,N_873,N_2017);
nor U2502 (N_2502,N_1390,N_859);
and U2503 (N_2503,N_1228,N_977);
nor U2504 (N_2504,N_1644,N_1423);
xnor U2505 (N_2505,N_1200,N_2224);
and U2506 (N_2506,N_563,N_1655);
nor U2507 (N_2507,N_1460,N_955);
nor U2508 (N_2508,N_1272,N_291);
xnor U2509 (N_2509,N_659,N_2437);
and U2510 (N_2510,N_2070,N_858);
nor U2511 (N_2511,N_588,N_2374);
xnor U2512 (N_2512,N_205,N_2357);
or U2513 (N_2513,N_182,N_978);
nand U2514 (N_2514,N_1977,N_1727);
and U2515 (N_2515,N_2207,N_965);
nand U2516 (N_2516,N_1140,N_2032);
nor U2517 (N_2517,N_1610,N_729);
xor U2518 (N_2518,N_465,N_1542);
xor U2519 (N_2519,N_1535,N_2185);
nand U2520 (N_2520,N_913,N_386);
nand U2521 (N_2521,N_470,N_673);
and U2522 (N_2522,N_1818,N_1601);
nor U2523 (N_2523,N_878,N_1674);
xor U2524 (N_2524,N_1860,N_2058);
xor U2525 (N_2525,N_2305,N_2129);
nor U2526 (N_2526,N_1420,N_199);
and U2527 (N_2527,N_382,N_807);
and U2528 (N_2528,N_2469,N_1507);
xor U2529 (N_2529,N_277,N_1821);
nor U2530 (N_2530,N_2268,N_1903);
nor U2531 (N_2531,N_1236,N_1964);
nand U2532 (N_2532,N_294,N_50);
nor U2533 (N_2533,N_356,N_2132);
xnor U2534 (N_2534,N_2333,N_2218);
and U2535 (N_2535,N_2149,N_1855);
nand U2536 (N_2536,N_1467,N_610);
xor U2537 (N_2537,N_379,N_552);
or U2538 (N_2538,N_1654,N_394);
or U2539 (N_2539,N_942,N_1558);
nand U2540 (N_2540,N_1804,N_887);
xnor U2541 (N_2541,N_572,N_2148);
nand U2542 (N_2542,N_266,N_240);
nand U2543 (N_2543,N_90,N_246);
and U2544 (N_2544,N_970,N_593);
xor U2545 (N_2545,N_498,N_1809);
nand U2546 (N_2546,N_2192,N_2281);
nand U2547 (N_2547,N_502,N_698);
and U2548 (N_2548,N_1697,N_148);
or U2549 (N_2549,N_249,N_1884);
xor U2550 (N_2550,N_1552,N_1788);
nand U2551 (N_2551,N_1623,N_1770);
and U2552 (N_2552,N_587,N_554);
or U2553 (N_2553,N_2030,N_104);
and U2554 (N_2554,N_2461,N_928);
and U2555 (N_2555,N_1650,N_1624);
xnor U2556 (N_2556,N_1800,N_1871);
nand U2557 (N_2557,N_337,N_2433);
nor U2558 (N_2558,N_11,N_540);
and U2559 (N_2559,N_1919,N_334);
nor U2560 (N_2560,N_722,N_1497);
nor U2561 (N_2561,N_1757,N_418);
nand U2562 (N_2562,N_58,N_2340);
and U2563 (N_2563,N_1725,N_1033);
and U2564 (N_2564,N_2042,N_1211);
or U2565 (N_2565,N_2183,N_15);
nand U2566 (N_2566,N_527,N_385);
or U2567 (N_2567,N_1438,N_1444);
nand U2568 (N_2568,N_931,N_2242);
nor U2569 (N_2569,N_835,N_1119);
or U2570 (N_2570,N_1811,N_2353);
nand U2571 (N_2571,N_57,N_2270);
nand U2572 (N_2572,N_72,N_757);
and U2573 (N_2573,N_2152,N_391);
xnor U2574 (N_2574,N_143,N_1575);
and U2575 (N_2575,N_414,N_1027);
and U2576 (N_2576,N_1353,N_1431);
or U2577 (N_2577,N_128,N_98);
or U2578 (N_2578,N_1791,N_1408);
nand U2579 (N_2579,N_656,N_717);
nand U2580 (N_2580,N_2015,N_864);
or U2581 (N_2581,N_1087,N_1908);
xor U2582 (N_2582,N_426,N_944);
and U2583 (N_2583,N_2468,N_902);
or U2584 (N_2584,N_522,N_579);
nand U2585 (N_2585,N_2170,N_2458);
or U2586 (N_2586,N_1392,N_1916);
nor U2587 (N_2587,N_2171,N_1837);
xor U2588 (N_2588,N_506,N_2179);
nor U2589 (N_2589,N_1581,N_144);
xor U2590 (N_2590,N_983,N_383);
xnor U2591 (N_2591,N_1726,N_145);
xor U2592 (N_2592,N_1984,N_2254);
nor U2593 (N_2593,N_1443,N_2089);
nor U2594 (N_2594,N_734,N_1068);
nor U2595 (N_2595,N_333,N_1812);
or U2596 (N_2596,N_1611,N_1936);
or U2597 (N_2597,N_1694,N_126);
nor U2598 (N_2598,N_1894,N_218);
or U2599 (N_2599,N_2232,N_400);
nor U2600 (N_2600,N_1371,N_708);
nor U2601 (N_2601,N_574,N_2229);
or U2602 (N_2602,N_2079,N_643);
and U2603 (N_2603,N_2298,N_832);
or U2604 (N_2604,N_863,N_845);
nand U2605 (N_2605,N_1273,N_2448);
nand U2606 (N_2606,N_367,N_2198);
nor U2607 (N_2607,N_677,N_1844);
nor U2608 (N_2608,N_855,N_164);
or U2609 (N_2609,N_2429,N_323);
nand U2610 (N_2610,N_1415,N_131);
nand U2611 (N_2611,N_2431,N_2425);
and U2612 (N_2612,N_231,N_2273);
and U2613 (N_2613,N_699,N_1014);
or U2614 (N_2614,N_1579,N_730);
nor U2615 (N_2615,N_915,N_953);
xor U2616 (N_2616,N_89,N_380);
nand U2617 (N_2617,N_2105,N_653);
xnor U2618 (N_2618,N_193,N_260);
nor U2619 (N_2619,N_397,N_860);
nor U2620 (N_2620,N_1637,N_2013);
or U2621 (N_2621,N_1279,N_2368);
xor U2622 (N_2622,N_740,N_471);
nand U2623 (N_2623,N_19,N_1970);
nor U2624 (N_2624,N_828,N_1025);
nor U2625 (N_2625,N_2278,N_1959);
xor U2626 (N_2626,N_631,N_2409);
or U2627 (N_2627,N_2059,N_176);
and U2628 (N_2628,N_2205,N_529);
nand U2629 (N_2629,N_2110,N_620);
nor U2630 (N_2630,N_2190,N_20);
nand U2631 (N_2631,N_1618,N_91);
xor U2632 (N_2632,N_51,N_1638);
nand U2633 (N_2633,N_1801,N_2440);
and U2634 (N_2634,N_839,N_165);
xnor U2635 (N_2635,N_1024,N_1474);
and U2636 (N_2636,N_1396,N_1834);
xnor U2637 (N_2637,N_1950,N_768);
or U2638 (N_2638,N_48,N_453);
or U2639 (N_2639,N_1101,N_2057);
xor U2640 (N_2640,N_2483,N_2066);
xnor U2641 (N_2641,N_2209,N_1670);
xnor U2642 (N_2642,N_1966,N_84);
and U2643 (N_2643,N_1583,N_519);
and U2644 (N_2644,N_1123,N_2403);
nand U2645 (N_2645,N_1196,N_213);
or U2646 (N_2646,N_2260,N_350);
xor U2647 (N_2647,N_1516,N_1180);
nor U2648 (N_2648,N_2494,N_151);
nand U2649 (N_2649,N_1931,N_1873);
xnor U2650 (N_2650,N_1243,N_1993);
and U2651 (N_2651,N_329,N_767);
nand U2652 (N_2652,N_2166,N_1354);
or U2653 (N_2653,N_1785,N_1244);
nor U2654 (N_2654,N_1240,N_2343);
xnor U2655 (N_2655,N_949,N_384);
and U2656 (N_2656,N_1949,N_810);
and U2657 (N_2657,N_2300,N_799);
nand U2658 (N_2658,N_1849,N_1178);
nor U2659 (N_2659,N_1326,N_428);
nand U2660 (N_2660,N_1040,N_2028);
nand U2661 (N_2661,N_1707,N_1224);
nand U2662 (N_2662,N_880,N_306);
nor U2663 (N_2663,N_448,N_1736);
xnor U2664 (N_2664,N_1247,N_756);
or U2665 (N_2665,N_71,N_1487);
xor U2666 (N_2666,N_338,N_626);
and U2667 (N_2667,N_1179,N_843);
or U2668 (N_2668,N_1400,N_2316);
xnor U2669 (N_2669,N_897,N_821);
or U2670 (N_2670,N_1759,N_963);
nand U2671 (N_2671,N_1473,N_2401);
nand U2672 (N_2672,N_1632,N_2350);
nor U2673 (N_2673,N_2354,N_1495);
or U2674 (N_2674,N_504,N_476);
and U2675 (N_2675,N_302,N_362);
and U2676 (N_2676,N_622,N_561);
and U2677 (N_2677,N_1532,N_1898);
xor U2678 (N_2678,N_455,N_1716);
xor U2679 (N_2679,N_43,N_836);
xor U2680 (N_2680,N_2314,N_748);
nand U2681 (N_2681,N_1518,N_1216);
nor U2682 (N_2682,N_893,N_633);
nand U2683 (N_2683,N_2308,N_937);
xor U2684 (N_2684,N_2499,N_848);
nor U2685 (N_2685,N_2049,N_1389);
xnor U2686 (N_2686,N_444,N_2085);
xor U2687 (N_2687,N_2294,N_876);
and U2688 (N_2688,N_1671,N_736);
and U2689 (N_2689,N_230,N_1163);
nand U2690 (N_2690,N_117,N_1207);
nor U2691 (N_2691,N_2258,N_2012);
nor U2692 (N_2692,N_896,N_619);
and U2693 (N_2693,N_744,N_1066);
nor U2694 (N_2694,N_2169,N_478);
and U2695 (N_2695,N_1692,N_1345);
nor U2696 (N_2696,N_2027,N_2492);
and U2697 (N_2697,N_1475,N_1797);
or U2698 (N_2698,N_263,N_241);
nand U2699 (N_2699,N_1194,N_2051);
xor U2700 (N_2700,N_1472,N_1159);
xor U2701 (N_2701,N_1700,N_1234);
and U2702 (N_2702,N_582,N_1749);
or U2703 (N_2703,N_420,N_1626);
or U2704 (N_2704,N_1410,N_275);
nor U2705 (N_2705,N_1897,N_1939);
nor U2706 (N_2706,N_403,N_1793);
nor U2707 (N_2707,N_239,N_505);
nor U2708 (N_2708,N_889,N_1242);
xor U2709 (N_2709,N_2193,N_492);
and U2710 (N_2710,N_763,N_1065);
nor U2711 (N_2711,N_641,N_18);
nand U2712 (N_2712,N_512,N_974);
or U2713 (N_2713,N_2150,N_150);
xor U2714 (N_2714,N_1300,N_1827);
nand U2715 (N_2715,N_2119,N_1015);
nor U2716 (N_2716,N_1582,N_2269);
nor U2717 (N_2717,N_1085,N_1649);
nor U2718 (N_2718,N_2102,N_1803);
nand U2719 (N_2719,N_1419,N_207);
xnor U2720 (N_2720,N_1730,N_1237);
nor U2721 (N_2721,N_564,N_1538);
xor U2722 (N_2722,N_2050,N_840);
and U2723 (N_2723,N_1492,N_305);
nor U2724 (N_2724,N_2126,N_1447);
nand U2725 (N_2725,N_2370,N_228);
nand U2726 (N_2726,N_483,N_583);
and U2727 (N_2727,N_1110,N_288);
nand U2728 (N_2728,N_1543,N_589);
and U2729 (N_2729,N_1695,N_1795);
or U2730 (N_2730,N_2053,N_724);
nand U2731 (N_2731,N_2462,N_2178);
xnor U2732 (N_2732,N_1886,N_1879);
or U2733 (N_2733,N_1245,N_2317);
or U2734 (N_2734,N_2140,N_1957);
xor U2735 (N_2735,N_851,N_621);
or U2736 (N_2736,N_2093,N_1851);
and U2737 (N_2737,N_2362,N_419);
nor U2738 (N_2738,N_1591,N_2231);
and U2739 (N_2739,N_867,N_211);
nand U2740 (N_2740,N_1344,N_2011);
nor U2741 (N_2741,N_2134,N_1045);
or U2742 (N_2742,N_1561,N_908);
and U2743 (N_2743,N_1878,N_1848);
nor U2744 (N_2744,N_2167,N_2211);
nand U2745 (N_2745,N_1266,N_1121);
or U2746 (N_2746,N_1790,N_1126);
or U2747 (N_2747,N_1625,N_2306);
and U2748 (N_2748,N_737,N_1038);
xor U2749 (N_2749,N_1867,N_718);
nand U2750 (N_2750,N_2020,N_2124);
xor U2751 (N_2751,N_136,N_2388);
nor U2752 (N_2752,N_1041,N_1062);
and U2753 (N_2753,N_1019,N_1604);
and U2754 (N_2754,N_2476,N_2275);
nand U2755 (N_2755,N_2098,N_547);
xnor U2756 (N_2756,N_1328,N_856);
xnor U2757 (N_2757,N_2355,N_1668);
nor U2758 (N_2758,N_751,N_542);
nor U2759 (N_2759,N_106,N_1092);
nand U2760 (N_2760,N_689,N_1464);
or U2761 (N_2761,N_494,N_186);
and U2762 (N_2762,N_210,N_1728);
nand U2763 (N_2763,N_66,N_468);
nand U2764 (N_2764,N_2453,N_1646);
or U2765 (N_2765,N_2094,N_109);
xnor U2766 (N_2766,N_1359,N_709);
or U2767 (N_2767,N_1678,N_61);
xor U2768 (N_2768,N_2128,N_99);
nand U2769 (N_2769,N_1521,N_776);
nand U2770 (N_2770,N_413,N_2136);
or U2771 (N_2771,N_1437,N_2029);
xor U2772 (N_2772,N_1208,N_158);
nand U2773 (N_2773,N_1160,N_25);
and U2774 (N_2774,N_1098,N_1029);
or U2775 (N_2775,N_269,N_849);
xor U2776 (N_2776,N_120,N_954);
nand U2777 (N_2777,N_1007,N_2288);
nor U2778 (N_2778,N_1004,N_888);
xnor U2779 (N_2779,N_987,N_87);
nand U2780 (N_2780,N_1767,N_988);
nand U2781 (N_2781,N_687,N_611);
or U2782 (N_2782,N_951,N_1687);
nand U2783 (N_2783,N_1454,N_1167);
xnor U2784 (N_2784,N_67,N_1985);
and U2785 (N_2785,N_2221,N_2376);
and U2786 (N_2786,N_69,N_254);
nand U2787 (N_2787,N_2424,N_735);
or U2788 (N_2788,N_1992,N_1373);
or U2789 (N_2789,N_674,N_999);
or U2790 (N_2790,N_1968,N_499);
or U2791 (N_2791,N_2324,N_119);
or U2792 (N_2792,N_2485,N_947);
xor U2793 (N_2793,N_1336,N_1325);
nor U2794 (N_2794,N_2396,N_267);
nor U2795 (N_2795,N_2498,N_573);
and U2796 (N_2796,N_1841,N_1926);
nor U2797 (N_2797,N_1717,N_1084);
or U2798 (N_2798,N_819,N_1991);
xnor U2799 (N_2799,N_1370,N_392);
nor U2800 (N_2800,N_232,N_919);
nand U2801 (N_2801,N_10,N_1763);
xnor U2802 (N_2802,N_1613,N_154);
and U2803 (N_2803,N_943,N_1348);
nor U2804 (N_2804,N_909,N_615);
or U2805 (N_2805,N_1289,N_927);
or U2806 (N_2806,N_1217,N_1599);
xnor U2807 (N_2807,N_319,N_1258);
and U2808 (N_2808,N_1455,N_1560);
and U2809 (N_2809,N_256,N_600);
and U2810 (N_2810,N_175,N_2226);
nand U2811 (N_2811,N_1924,N_793);
xor U2812 (N_2812,N_1608,N_1302);
nand U2813 (N_2813,N_27,N_679);
and U2814 (N_2814,N_1755,N_2491);
nor U2815 (N_2815,N_2095,N_1127);
and U2816 (N_2816,N_1284,N_2031);
or U2817 (N_2817,N_95,N_261);
nand U2818 (N_2818,N_1122,N_576);
nand U2819 (N_2819,N_423,N_1680);
and U2820 (N_2820,N_477,N_544);
xor U2821 (N_2821,N_777,N_301);
nand U2822 (N_2822,N_311,N_1622);
nor U2823 (N_2823,N_1439,N_2386);
or U2824 (N_2824,N_628,N_597);
or U2825 (N_2825,N_882,N_224);
and U2826 (N_2826,N_2202,N_1783);
xor U2827 (N_2827,N_2172,N_1973);
nand U2828 (N_2828,N_1295,N_1323);
nor U2829 (N_2829,N_2115,N_2361);
nand U2830 (N_2830,N_866,N_1733);
and U2831 (N_2831,N_2087,N_1810);
or U2832 (N_2832,N_486,N_2452);
and U2833 (N_2833,N_1135,N_969);
xor U2834 (N_2834,N_1746,N_1833);
nor U2835 (N_2835,N_1206,N_725);
and U2836 (N_2836,N_688,N_749);
and U2837 (N_2837,N_1564,N_49);
xnor U2838 (N_2838,N_1338,N_1340);
and U2839 (N_2839,N_2236,N_596);
xnor U2840 (N_2840,N_775,N_904);
nor U2841 (N_2841,N_1164,N_1221);
or U2842 (N_2842,N_437,N_1524);
xor U2843 (N_2843,N_1527,N_1088);
nand U2844 (N_2844,N_1866,N_1256);
nor U2845 (N_2845,N_1453,N_1861);
nor U2846 (N_2846,N_1904,N_2381);
and U2847 (N_2847,N_1001,N_676);
nor U2848 (N_2848,N_1271,N_8);
or U2849 (N_2849,N_1037,N_1401);
or U2850 (N_2850,N_416,N_809);
or U2851 (N_2851,N_2342,N_2266);
or U2852 (N_2852,N_903,N_1108);
and U2853 (N_2853,N_2043,N_1506);
nand U2854 (N_2854,N_571,N_2402);
nor U2855 (N_2855,N_962,N_222);
or U2856 (N_2856,N_1635,N_1259);
and U2857 (N_2857,N_862,N_1570);
nand U2858 (N_2858,N_1719,N_912);
xnor U2859 (N_2859,N_443,N_1696);
xnor U2860 (N_2860,N_1580,N_2328);
nor U2861 (N_2861,N_399,N_1852);
xor U2862 (N_2862,N_1100,N_31);
xnor U2863 (N_2863,N_515,N_525);
nor U2864 (N_2864,N_1523,N_2397);
xnor U2865 (N_2865,N_1836,N_94);
and U2866 (N_2866,N_2197,N_883);
or U2867 (N_2867,N_1238,N_9);
xor U2868 (N_2868,N_295,N_1718);
nand U2869 (N_2869,N_351,N_1927);
xnor U2870 (N_2870,N_1141,N_1483);
nor U2871 (N_2871,N_1077,N_939);
nand U2872 (N_2872,N_753,N_1805);
nand U2873 (N_2873,N_741,N_1778);
nor U2874 (N_2874,N_1036,N_2142);
xnor U2875 (N_2875,N_1307,N_607);
or U2876 (N_2876,N_490,N_1079);
or U2877 (N_2877,N_332,N_467);
nor U2878 (N_2878,N_989,N_818);
or U2879 (N_2879,N_853,N_39);
and U2880 (N_2880,N_2117,N_183);
nor U2881 (N_2881,N_1055,N_1563);
or U2882 (N_2882,N_702,N_340);
nand U2883 (N_2883,N_773,N_901);
xnor U2884 (N_2884,N_1227,N_435);
nor U2885 (N_2885,N_1776,N_2088);
and U2886 (N_2886,N_541,N_1682);
or U2887 (N_2887,N_2372,N_162);
nor U2888 (N_2888,N_92,N_1704);
xor U2889 (N_2889,N_1023,N_389);
nand U2890 (N_2890,N_303,N_1118);
nor U2891 (N_2891,N_1422,N_405);
or U2892 (N_2892,N_513,N_891);
or U2893 (N_2893,N_1548,N_2123);
nand U2894 (N_2894,N_1052,N_2336);
nand U2895 (N_2895,N_1509,N_997);
xnor U2896 (N_2896,N_2456,N_2139);
or U2897 (N_2897,N_1616,N_545);
or U2898 (N_2898,N_1779,N_1907);
nand U2899 (N_2899,N_1910,N_2442);
and U2900 (N_2900,N_2297,N_1424);
nor U2901 (N_2901,N_1864,N_1076);
nand U2902 (N_2902,N_2276,N_584);
nand U2903 (N_2903,N_1488,N_1299);
nor U2904 (N_2904,N_2349,N_1691);
and U2905 (N_2905,N_1290,N_1598);
nand U2906 (N_2906,N_1421,N_1089);
and U2907 (N_2907,N_1010,N_52);
xor U2908 (N_2908,N_1462,N_2201);
xnor U2909 (N_2909,N_2359,N_1030);
or U2910 (N_2910,N_1539,N_296);
and U2911 (N_2911,N_868,N_1577);
nand U2912 (N_2912,N_123,N_1265);
or U2913 (N_2913,N_2038,N_1060);
xor U2914 (N_2914,N_1944,N_349);
nand U2915 (N_2915,N_2364,N_1899);
nand U2916 (N_2916,N_663,N_658);
xor U2917 (N_2917,N_238,N_761);
nor U2918 (N_2918,N_2428,N_320);
and U2919 (N_2919,N_1741,N_21);
nor U2920 (N_2920,N_874,N_1330);
and U2921 (N_2921,N_1293,N_2147);
nor U2922 (N_2922,N_262,N_2472);
nor U2923 (N_2923,N_861,N_787);
or U2924 (N_2924,N_137,N_1380);
and U2925 (N_2925,N_1490,N_35);
nand U2926 (N_2926,N_961,N_2156);
and U2927 (N_2927,N_216,N_2225);
nand U2928 (N_2928,N_546,N_2182);
xor U2929 (N_2929,N_197,N_2259);
nand U2930 (N_2930,N_1578,N_2175);
and U2931 (N_2931,N_2451,N_187);
or U2932 (N_2932,N_754,N_2250);
and U2933 (N_2933,N_1209,N_184);
nand U2934 (N_2934,N_614,N_2321);
nand U2935 (N_2935,N_1989,N_669);
xnor U2936 (N_2936,N_929,N_782);
or U2937 (N_2937,N_2125,N_1133);
nor U2938 (N_2938,N_1193,N_80);
nand U2939 (N_2939,N_2358,N_2052);
nor U2940 (N_2940,N_412,N_2318);
xnor U2941 (N_2941,N_2293,N_952);
xor U2942 (N_2942,N_376,N_1006);
nand U2943 (N_2943,N_457,N_2417);
or U2944 (N_2944,N_1854,N_759);
nand U2945 (N_2945,N_1659,N_335);
or U2946 (N_2946,N_2161,N_233);
and U2947 (N_2947,N_2375,N_2296);
nor U2948 (N_2948,N_64,N_2113);
nor U2949 (N_2949,N_466,N_347);
nand U2950 (N_2950,N_834,N_325);
and U2951 (N_2951,N_852,N_1471);
nor U2952 (N_2952,N_683,N_1195);
or U2953 (N_2953,N_341,N_857);
and U2954 (N_2954,N_1870,N_1189);
nor U2955 (N_2955,N_1892,N_1983);
xnor U2956 (N_2956,N_705,N_2035);
nand U2957 (N_2957,N_364,N_1187);
and U2958 (N_2958,N_2426,N_916);
nand U2959 (N_2959,N_1929,N_114);
or U2960 (N_2960,N_2217,N_134);
nor U2961 (N_2961,N_113,N_712);
or U2962 (N_2962,N_950,N_2463);
nor U2963 (N_2963,N_439,N_1436);
xor U2964 (N_2964,N_1175,N_691);
xor U2965 (N_2965,N_992,N_2120);
nor U2966 (N_2966,N_2307,N_697);
or U2967 (N_2967,N_1830,N_1994);
xor U2968 (N_2968,N_2007,N_149);
nor U2969 (N_2969,N_838,N_1642);
and U2970 (N_2970,N_1843,N_996);
nor U2971 (N_2971,N_219,N_1349);
or U2972 (N_2972,N_1152,N_47);
or U2973 (N_2973,N_1574,N_1105);
nor U2974 (N_2974,N_2008,N_2338);
nor U2975 (N_2975,N_1090,N_1061);
and U2976 (N_2976,N_2144,N_1170);
and U2977 (N_2977,N_141,N_36);
xnor U2978 (N_2978,N_2072,N_1314);
nor U2979 (N_2979,N_122,N_1522);
and U2980 (N_2980,N_1925,N_1965);
xnor U2981 (N_2981,N_1607,N_427);
nand U2982 (N_2982,N_2344,N_817);
nor U2983 (N_2983,N_46,N_1813);
and U2984 (N_2984,N_704,N_501);
nor U2985 (N_2985,N_1751,N_206);
or U2986 (N_2986,N_1405,N_533);
and U2987 (N_2987,N_1322,N_2116);
nor U2988 (N_2988,N_1762,N_1394);
or U2989 (N_2989,N_764,N_2191);
nor U2990 (N_2990,N_161,N_1683);
nor U2991 (N_2991,N_1009,N_398);
nand U2992 (N_2992,N_214,N_474);
xnor U2993 (N_2993,N_2018,N_191);
nor U2994 (N_2994,N_2138,N_243);
and U2995 (N_2995,N_45,N_558);
nand U2996 (N_2996,N_1967,N_1657);
xor U2997 (N_2997,N_450,N_2497);
nand U2998 (N_2998,N_2228,N_1080);
and U2999 (N_2999,N_1496,N_1186);
and U3000 (N_3000,N_1070,N_1633);
nand U3001 (N_3001,N_2060,N_1890);
nand U3002 (N_3002,N_694,N_1241);
or U3003 (N_3003,N_1546,N_2003);
or U3004 (N_3004,N_1139,N_177);
and U3005 (N_3005,N_1734,N_1278);
nand U3006 (N_3006,N_1434,N_1287);
nor U3007 (N_3007,N_2223,N_1433);
and U3008 (N_3008,N_1450,N_844);
and U3009 (N_3009,N_985,N_153);
xor U3010 (N_3010,N_1945,N_378);
xor U3011 (N_3011,N_2495,N_181);
or U3012 (N_3012,N_1183,N_2097);
nor U3013 (N_3013,N_720,N_1645);
and U3014 (N_3014,N_2212,N_454);
and U3015 (N_3015,N_1951,N_1856);
xnor U3016 (N_3016,N_2131,N_1395);
xor U3017 (N_3017,N_346,N_1463);
nor U3018 (N_3018,N_1489,N_813);
and U3019 (N_3019,N_2026,N_2473);
or U3020 (N_3020,N_2257,N_1885);
or U3021 (N_3021,N_2249,N_445);
xor U3022 (N_3022,N_1586,N_565);
nor U3023 (N_3023,N_514,N_1641);
nand U3024 (N_3024,N_1947,N_2313);
and U3025 (N_3025,N_2157,N_1268);
or U3026 (N_3026,N_1219,N_671);
and U3027 (N_3027,N_100,N_1210);
nand U3028 (N_3028,N_1491,N_1865);
nor U3029 (N_3029,N_200,N_1103);
xnor U3030 (N_3030,N_1376,N_2077);
xor U3031 (N_3031,N_1430,N_2399);
xnor U3032 (N_3032,N_2036,N_1305);
xor U3033 (N_3033,N_2290,N_850);
or U3034 (N_3034,N_1587,N_518);
nand U3035 (N_3035,N_1915,N_451);
or U3036 (N_3036,N_1282,N_854);
nand U3037 (N_3037,N_1296,N_1043);
nor U3038 (N_3038,N_1976,N_2413);
nor U3039 (N_3039,N_278,N_758);
nor U3040 (N_3040,N_159,N_982);
or U3041 (N_3041,N_1231,N_1102);
nor U3042 (N_3042,N_133,N_2391);
nand U3043 (N_3043,N_1677,N_1137);
or U3044 (N_3044,N_609,N_811);
nand U3045 (N_3045,N_1585,N_252);
nand U3046 (N_3046,N_1112,N_1789);
and U3047 (N_3047,N_310,N_825);
and U3048 (N_3048,N_2222,N_1708);
nor U3049 (N_3049,N_1162,N_2325);
or U3050 (N_3050,N_695,N_1409);
xnor U3051 (N_3051,N_1858,N_1955);
nand U3052 (N_3052,N_2286,N_523);
xnor U3053 (N_3053,N_1201,N_23);
nor U3054 (N_3054,N_473,N_2380);
xnor U3055 (N_3055,N_2378,N_907);
xor U3056 (N_3056,N_1690,N_1952);
nand U3057 (N_3057,N_1566,N_60);
or U3058 (N_3058,N_110,N_2041);
or U3059 (N_3059,N_1269,N_1545);
and U3060 (N_3060,N_2369,N_623);
xnor U3061 (N_3061,N_1018,N_2046);
or U3062 (N_3062,N_336,N_1005);
or U3063 (N_3063,N_2311,N_1998);
or U3064 (N_3064,N_1044,N_2454);
xor U3065 (N_3065,N_270,N_1958);
xnor U3066 (N_3066,N_531,N_1845);
xor U3067 (N_3067,N_1107,N_1154);
nor U3068 (N_3068,N_488,N_682);
and U3069 (N_3069,N_1887,N_1619);
or U3070 (N_3070,N_739,N_1872);
nand U3071 (N_3071,N_2345,N_1740);
xnor U3072 (N_3072,N_1600,N_1132);
nor U3073 (N_3073,N_1835,N_2083);
or U3074 (N_3074,N_1752,N_559);
and U3075 (N_3075,N_1341,N_1435);
and U3076 (N_3076,N_430,N_2208);
nand U3077 (N_3077,N_265,N_2214);
and U3078 (N_3078,N_1699,N_1372);
xnor U3079 (N_3079,N_460,N_693);
nand U3080 (N_3080,N_959,N_1920);
or U3081 (N_3081,N_1316,N_1263);
xnor U3082 (N_3082,N_2080,N_316);
xnor U3083 (N_3083,N_1343,N_2466);
nand U3084 (N_3084,N_1306,N_792);
xnor U3085 (N_3085,N_2406,N_824);
and U3086 (N_3086,N_2267,N_2383);
or U3087 (N_3087,N_847,N_1771);
xnor U3088 (N_3088,N_662,N_2235);
and U3089 (N_3089,N_290,N_2371);
nand U3090 (N_3090,N_1722,N_2351);
nor U3091 (N_3091,N_872,N_801);
nand U3092 (N_3092,N_804,N_1351);
or U3093 (N_3093,N_2347,N_1525);
or U3094 (N_3094,N_2247,N_1321);
xor U3095 (N_3095,N_1481,N_1653);
nand U3096 (N_3096,N_2216,N_1003);
and U3097 (N_3097,N_304,N_733);
nor U3098 (N_3098,N_577,N_2244);
or U3099 (N_3099,N_814,N_1064);
xor U3100 (N_3100,N_1145,N_1177);
or U3101 (N_3101,N_387,N_2496);
nand U3102 (N_3102,N_1629,N_791);
and U3103 (N_3103,N_1337,N_1597);
or U3104 (N_3104,N_1375,N_1962);
nor U3105 (N_3105,N_1254,N_1053);
nand U3106 (N_3106,N_1280,N_971);
xor U3107 (N_3107,N_833,N_2151);
nand U3108 (N_3108,N_2410,N_1468);
nand U3109 (N_3109,N_766,N_1979);
or U3110 (N_3110,N_1486,N_1312);
xnor U3111 (N_3111,N_1011,N_1091);
nor U3112 (N_3112,N_299,N_2470);
or U3113 (N_3113,N_2477,N_409);
or U3114 (N_3114,N_1963,N_932);
or U3115 (N_3115,N_264,N_592);
nand U3116 (N_3116,N_156,N_672);
xnor U3117 (N_3117,N_1643,N_1393);
nor U3118 (N_3118,N_223,N_1173);
and U3119 (N_3119,N_2330,N_298);
nor U3120 (N_3120,N_1125,N_1658);
nor U3121 (N_3121,N_1477,N_1880);
nor U3122 (N_3122,N_2040,N_638);
or U3123 (N_3123,N_1526,N_1933);
nor U3124 (N_3124,N_1875,N_1559);
and U3125 (N_3125,N_481,N_1502);
nor U3126 (N_3126,N_993,N_745);
and U3127 (N_3127,N_1595,N_1493);
nor U3128 (N_3128,N_2240,N_1550);
and U3129 (N_3129,N_2280,N_447);
nand U3130 (N_3130,N_976,N_648);
nand U3131 (N_3131,N_956,N_2455);
nand U3132 (N_3132,N_1381,N_2465);
and U3133 (N_3133,N_991,N_1647);
and U3134 (N_3134,N_152,N_142);
and U3135 (N_3135,N_1515,N_1829);
or U3136 (N_3136,N_2251,N_1192);
nor U3137 (N_3137,N_1428,N_2100);
nand U3138 (N_3138,N_972,N_2420);
nand U3139 (N_3139,N_2173,N_632);
and U3140 (N_3140,N_1981,N_1331);
xor U3141 (N_3141,N_2174,N_2238);
or U3142 (N_3142,N_2432,N_1660);
xor U3143 (N_3143,N_284,N_1510);
nand U3144 (N_3144,N_2023,N_118);
nand U3145 (N_3145,N_1075,N_646);
nand U3146 (N_3146,N_2055,N_1176);
xnor U3147 (N_3147,N_1735,N_778);
or U3148 (N_3148,N_1511,N_536);
and U3149 (N_3149,N_1083,N_924);
nand U3150 (N_3150,N_820,N_1383);
xnor U3151 (N_3151,N_1684,N_1067);
nor U3152 (N_3152,N_710,N_359);
nor U3153 (N_3153,N_1008,N_493);
and U3154 (N_3154,N_1048,N_968);
nand U3155 (N_3155,N_530,N_1275);
nand U3156 (N_3156,N_922,N_1798);
or U3157 (N_3157,N_1335,N_464);
and U3158 (N_3158,N_1213,N_1799);
nor U3159 (N_3159,N_185,N_283);
nand U3160 (N_3160,N_1760,N_348);
nand U3161 (N_3161,N_1461,N_1203);
nand U3162 (N_3162,N_229,N_1034);
or U3163 (N_3163,N_1665,N_550);
xor U3164 (N_3164,N_2210,N_603);
and U3165 (N_3165,N_508,N_1562);
nor U3166 (N_3166,N_147,N_2418);
nand U3167 (N_3167,N_2075,N_1745);
xor U3168 (N_3168,N_225,N_1026);
xnor U3169 (N_3169,N_1784,N_259);
nor U3170 (N_3170,N_2444,N_1534);
nor U3171 (N_3171,N_2000,N_1768);
xnor U3172 (N_3172,N_2480,N_1839);
nor U3173 (N_3173,N_369,N_2438);
and U3174 (N_3174,N_1151,N_2227);
nor U3175 (N_3175,N_1960,N_1500);
or U3176 (N_3176,N_1425,N_377);
and U3177 (N_3177,N_534,N_83);
nand U3178 (N_3178,N_1120,N_1136);
and U3179 (N_3179,N_2081,N_914);
nor U3180 (N_3180,N_2421,N_1820);
and U3181 (N_3181,N_666,N_429);
nor U3182 (N_3182,N_1109,N_96);
nor U3183 (N_3183,N_82,N_321);
and U3184 (N_3184,N_2385,N_203);
nor U3185 (N_3185,N_1448,N_375);
nor U3186 (N_3186,N_608,N_170);
xnor U3187 (N_3187,N_570,N_800);
nor U3188 (N_3188,N_1451,N_798);
or U3189 (N_3189,N_981,N_101);
nand U3190 (N_3190,N_2194,N_1418);
xor U3191 (N_3191,N_2246,N_556);
nor U3192 (N_3192,N_2319,N_507);
xnor U3193 (N_3193,N_1503,N_879);
nand U3194 (N_3194,N_635,N_685);
xor U3195 (N_3195,N_2203,N_1403);
xnor U3196 (N_3196,N_1986,N_485);
xnor U3197 (N_3197,N_1666,N_1743);
nor U3198 (N_3198,N_116,N_877);
nor U3199 (N_3199,N_1166,N_1603);
and U3200 (N_3200,N_2,N_55);
nor U3201 (N_3201,N_1368,N_1721);
xor U3202 (N_3202,N_711,N_2450);
nor U3203 (N_3203,N_1458,N_179);
nand U3204 (N_3204,N_2487,N_282);
nand U3205 (N_3205,N_841,N_2379);
nand U3206 (N_3206,N_2245,N_130);
or U3207 (N_3207,N_509,N_2004);
nor U3208 (N_3208,N_2002,N_16);
or U3209 (N_3209,N_815,N_1630);
xnor U3210 (N_3210,N_934,N_1764);
or U3211 (N_3211,N_253,N_469);
or U3212 (N_3212,N_1168,N_1877);
xnor U3213 (N_3213,N_1485,N_462);
nand U3214 (N_3214,N_1384,N_242);
or U3215 (N_3215,N_892,N_1606);
nor U3216 (N_3216,N_634,N_204);
xor U3217 (N_3217,N_651,N_1703);
or U3218 (N_3218,N_2241,N_2389);
xnor U3219 (N_3219,N_1071,N_1197);
xor U3220 (N_3220,N_746,N_1054);
nor U3221 (N_3221,N_1652,N_1895);
and U3222 (N_3222,N_1753,N_2436);
xor U3223 (N_3223,N_268,N_1099);
nand U3224 (N_3224,N_1361,N_1917);
and U3225 (N_3225,N_1000,N_293);
nand U3226 (N_3226,N_491,N_1286);
or U3227 (N_3227,N_410,N_1602);
xnor U3228 (N_3228,N_647,N_1441);
nand U3229 (N_3229,N_1215,N_1253);
nor U3230 (N_3230,N_62,N_372);
nand U3231 (N_3231,N_7,N_495);
and U3232 (N_3232,N_979,N_381);
and U3233 (N_3233,N_797,N_318);
or U3234 (N_3234,N_2490,N_2215);
nor U3235 (N_3235,N_108,N_1367);
nand U3236 (N_3236,N_1932,N_459);
xnor U3237 (N_3237,N_2111,N_2107);
nand U3238 (N_3238,N_613,N_984);
xnor U3239 (N_3239,N_1554,N_2320);
or U3240 (N_3240,N_1149,N_1853);
nor U3241 (N_3241,N_1457,N_41);
and U3242 (N_3242,N_1342,N_328);
xor U3243 (N_3243,N_743,N_1360);
and U3244 (N_3244,N_63,N_762);
nand U3245 (N_3245,N_30,N_1831);
xor U3246 (N_3246,N_107,N_366);
or U3247 (N_3247,N_681,N_723);
or U3248 (N_3248,N_480,N_135);
nand U3249 (N_3249,N_2363,N_3);
nor U3250 (N_3250,N_911,N_1593);
or U3251 (N_3251,N_1131,N_317);
xnor U3252 (N_3252,N_926,N_1146);
or U3253 (N_3253,N_1569,N_706);
xor U3254 (N_3254,N_1116,N_2384);
nor U3255 (N_3255,N_1772,N_2356);
and U3256 (N_3256,N_1081,N_627);
xnor U3257 (N_3257,N_2071,N_1937);
xor U3258 (N_3258,N_2118,N_1826);
or U3259 (N_3259,N_772,N_449);
xnor U3260 (N_3260,N_788,N_2186);
and U3261 (N_3261,N_590,N_2309);
or U3262 (N_3262,N_780,N_605);
xor U3263 (N_3263,N_14,N_2048);
nand U3264 (N_3264,N_1365,N_339);
xnor U3265 (N_3265,N_322,N_728);
nor U3266 (N_3266,N_816,N_1334);
or U3267 (N_3267,N_1594,N_1673);
and U3268 (N_3268,N_2292,N_1445);
and U3269 (N_3269,N_1233,N_1928);
or U3270 (N_3270,N_1188,N_180);
and U3271 (N_3271,N_2272,N_2263);
nand U3272 (N_3272,N_2181,N_1530);
xor U3273 (N_3273,N_831,N_1051);
xnor U3274 (N_3274,N_980,N_2122);
or U3275 (N_3275,N_1313,N_2127);
or U3276 (N_3276,N_2078,N_1513);
nand U3277 (N_3277,N_1786,N_1298);
nor U3278 (N_3278,N_1816,N_1547);
xor U3279 (N_3279,N_1283,N_560);
and U3280 (N_3280,N_822,N_221);
or U3281 (N_3281,N_692,N_1059);
and U3282 (N_3282,N_355,N_2339);
nand U3283 (N_3283,N_2006,N_2160);
xnor U3284 (N_3284,N_172,N_779);
and U3285 (N_3285,N_2063,N_388);
nor U3286 (N_3286,N_1627,N_923);
or U3287 (N_3287,N_17,N_40);
or U3288 (N_3288,N_649,N_1782);
and U3289 (N_3289,N_1229,N_2009);
and U3290 (N_3290,N_869,N_2415);
or U3291 (N_3291,N_169,N_553);
nand U3292 (N_3292,N_675,N_1369);
xnor U3293 (N_3293,N_2408,N_1883);
xnor U3294 (N_3294,N_535,N_1505);
or U3295 (N_3295,N_140,N_1288);
xor U3296 (N_3296,N_1881,N_500);
nor U3297 (N_3297,N_360,N_188);
and U3298 (N_3298,N_1769,N_1840);
nor U3299 (N_3299,N_2303,N_503);
nor U3300 (N_3300,N_111,N_1386);
nand U3301 (N_3301,N_945,N_313);
or U3302 (N_3302,N_38,N_1427);
nand U3303 (N_3303,N_1249,N_1311);
xnor U3304 (N_3304,N_769,N_411);
nor U3305 (N_3305,N_701,N_703);
nand U3306 (N_3306,N_2239,N_1459);
nand U3307 (N_3307,N_124,N_1218);
nand U3308 (N_3308,N_1732,N_604);
xor U3309 (N_3309,N_1551,N_2061);
or U3310 (N_3310,N_2289,N_2423);
and U3311 (N_3311,N_1688,N_2481);
or U3312 (N_3312,N_826,N_2084);
and U3313 (N_3313,N_102,N_1182);
or U3314 (N_3314,N_900,N_2199);
nor U3315 (N_3315,N_781,N_279);
nor U3316 (N_3316,N_581,N_1094);
xnor U3317 (N_3317,N_1185,N_524);
nor U3318 (N_3318,N_1097,N_1794);
nor U3319 (N_3319,N_967,N_2206);
xnor U3320 (N_3320,N_1114,N_1556);
and U3321 (N_3321,N_1571,N_1918);
or U3322 (N_3322,N_1723,N_285);
or U3323 (N_3323,N_1397,N_1022);
or U3324 (N_3324,N_2395,N_202);
nand U3325 (N_3325,N_1285,N_4);
or U3326 (N_3326,N_1096,N_155);
and U3327 (N_3327,N_715,N_2039);
and U3328 (N_3328,N_2065,N_794);
nand U3329 (N_3329,N_1590,N_2103);
xnor U3330 (N_3330,N_1806,N_1824);
or U3331 (N_3331,N_1796,N_732);
xor U3332 (N_3332,N_1358,N_112);
nor U3333 (N_3333,N_1264,N_2114);
or U3334 (N_3334,N_2133,N_1662);
or U3335 (N_3335,N_309,N_1702);
and U3336 (N_3336,N_998,N_727);
xnor U3337 (N_3337,N_2054,N_1147);
nor U3338 (N_3338,N_1225,N_1357);
nand U3339 (N_3339,N_1969,N_1775);
nand U3340 (N_3340,N_1220,N_194);
xor U3341 (N_3341,N_2219,N_2412);
nor U3342 (N_3342,N_236,N_2255);
nand U3343 (N_3343,N_73,N_208);
or U3344 (N_3344,N_404,N_244);
and U3345 (N_3345,N_1501,N_215);
xor U3346 (N_3346,N_1446,N_1914);
xnor U3347 (N_3347,N_2411,N_1150);
nor U3348 (N_3348,N_935,N_74);
or U3349 (N_3349,N_664,N_837);
xnor U3350 (N_3350,N_127,N_1540);
nor U3351 (N_3351,N_938,N_2334);
xnor U3352 (N_3352,N_1555,N_1214);
or U3353 (N_3353,N_1308,N_789);
and U3354 (N_3354,N_132,N_568);
or U3355 (N_3355,N_660,N_1270);
nor U3356 (N_3356,N_407,N_1617);
and U3357 (N_3357,N_1900,N_1063);
and U3358 (N_3358,N_484,N_1656);
nor U3359 (N_3359,N_1943,N_752);
nor U3360 (N_3360,N_446,N_1822);
nand U3361 (N_3361,N_1350,N_1706);
xnor U3362 (N_3362,N_257,N_1329);
or U3363 (N_3363,N_1808,N_463);
nand U3364 (N_3364,N_1484,N_948);
or U3365 (N_3365,N_1480,N_2291);
nor U3366 (N_3366,N_1553,N_167);
xnor U3367 (N_3367,N_713,N_1346);
nand U3368 (N_3368,N_70,N_2112);
and U3369 (N_3369,N_1319,N_1961);
and U3370 (N_3370,N_1198,N_549);
nand U3371 (N_3371,N_1859,N_870);
and U3372 (N_3372,N_1995,N_595);
or U3373 (N_3373,N_871,N_1385);
nor U3374 (N_3374,N_933,N_1508);
or U3375 (N_3375,N_612,N_1882);
and U3376 (N_3376,N_452,N_2101);
nor U3377 (N_3377,N_958,N_2387);
xor U3378 (N_3378,N_138,N_1028);
nand U3379 (N_3379,N_905,N_1017);
xnor U3380 (N_3380,N_1921,N_28);
or U3381 (N_3381,N_567,N_2445);
nand U3382 (N_3382,N_1407,N_654);
nor U3383 (N_3383,N_2443,N_1807);
and U3384 (N_3384,N_1681,N_1544);
xor U3385 (N_3385,N_1251,N_1148);
xor U3386 (N_3386,N_1095,N_755);
and U3387 (N_3387,N_1378,N_2146);
nor U3388 (N_3388,N_2154,N_1387);
nand U3389 (N_3389,N_1324,N_1246);
xnor U3390 (N_3390,N_1648,N_2302);
nand U3391 (N_3391,N_1056,N_2163);
nor U3392 (N_3392,N_2196,N_2233);
and U3393 (N_3393,N_575,N_2188);
nor U3394 (N_3394,N_1988,N_1568);
or U3395 (N_3395,N_657,N_1614);
xor U3396 (N_3396,N_2062,N_1404);
xnor U3397 (N_3397,N_1332,N_220);
xnor U3398 (N_3398,N_1181,N_1398);
nor U3399 (N_3399,N_76,N_1874);
or U3400 (N_3400,N_1169,N_1035);
nor U3401 (N_3401,N_2400,N_1588);
nor U3402 (N_3402,N_32,N_1698);
nand U3403 (N_3403,N_2047,N_1787);
nand U3404 (N_3404,N_2248,N_1823);
xnor U3405 (N_3405,N_406,N_684);
or U3406 (N_3406,N_1115,N_1987);
or U3407 (N_3407,N_1971,N_750);
or U3408 (N_3408,N_1124,N_13);
nand U3409 (N_3409,N_129,N_2033);
or U3410 (N_3410,N_248,N_2315);
or U3411 (N_3411,N_1399,N_785);
or U3412 (N_3412,N_1724,N_1499);
and U3413 (N_3413,N_716,N_1664);
nor U3414 (N_3414,N_2180,N_370);
nand U3415 (N_3415,N_636,N_910);
and U3416 (N_3416,N_461,N_1631);
or U3417 (N_3417,N_1469,N_1172);
nand U3418 (N_3418,N_1202,N_2200);
nor U3419 (N_3419,N_363,N_12);
or U3420 (N_3420,N_731,N_280);
and U3421 (N_3421,N_539,N_1713);
xnor U3422 (N_3422,N_1301,N_1274);
or U3423 (N_3423,N_103,N_805);
or U3424 (N_3424,N_1046,N_2014);
nor U3425 (N_3425,N_59,N_707);
and U3426 (N_3426,N_827,N_24);
and U3427 (N_3427,N_986,N_1996);
xnor U3428 (N_3428,N_2265,N_440);
nor U3429 (N_3429,N_606,N_2045);
nand U3430 (N_3430,N_2021,N_829);
nand U3431 (N_3431,N_1031,N_1498);
and U3432 (N_3432,N_1541,N_2332);
nor U3433 (N_3433,N_217,N_1413);
nand U3434 (N_3434,N_806,N_994);
and U3435 (N_3435,N_2439,N_1909);
xnor U3436 (N_3436,N_670,N_936);
nand U3437 (N_3437,N_315,N_198);
and U3438 (N_3438,N_1990,N_1974);
nor U3439 (N_3439,N_2165,N_289);
or U3440 (N_3440,N_357,N_415);
and U3441 (N_3441,N_1317,N_1382);
xnor U3442 (N_3442,N_1640,N_212);
nand U3443 (N_3443,N_925,N_422);
xor U3444 (N_3444,N_390,N_1828);
xnor U3445 (N_3445,N_930,N_2405);
nor U3446 (N_3446,N_1134,N_2213);
nor U3447 (N_3447,N_1737,N_408);
xor U3448 (N_3448,N_234,N_526);
xnor U3449 (N_3449,N_2108,N_1528);
nor U3450 (N_3450,N_1117,N_1520);
xor U3451 (N_3451,N_2204,N_2069);
or U3452 (N_3452,N_2310,N_1257);
nor U3453 (N_3453,N_1838,N_1414);
or U3454 (N_3454,N_2274,N_1032);
nor U3455 (N_3455,N_1689,N_1923);
nand U3456 (N_3456,N_2312,N_1589);
and U3457 (N_3457,N_2482,N_396);
or U3458 (N_3458,N_1412,N_1466);
and U3459 (N_3459,N_274,N_2484);
or U3460 (N_3460,N_1261,N_1869);
xnor U3461 (N_3461,N_2143,N_1802);
xnor U3462 (N_3462,N_510,N_2091);
xnor U3463 (N_3463,N_650,N_1073);
or U3464 (N_3464,N_1315,N_585);
nand U3465 (N_3465,N_425,N_326);
nor U3466 (N_3466,N_1567,N_796);
nor U3467 (N_3467,N_1930,N_1165);
and U3468 (N_3468,N_2010,N_1106);
nor U3469 (N_3469,N_1158,N_2073);
xor U3470 (N_3470,N_1938,N_616);
nor U3471 (N_3471,N_1780,N_417);
nand U3472 (N_3472,N_1153,N_201);
nor U3473 (N_3473,N_86,N_54);
xnor U3474 (N_3474,N_1842,N_1104);
nand U3475 (N_3475,N_747,N_1239);
and U3476 (N_3476,N_1975,N_1078);
nand U3477 (N_3477,N_686,N_1142);
nor U3478 (N_3478,N_173,N_2285);
nor U3479 (N_3479,N_431,N_1531);
and U3480 (N_3480,N_823,N_1922);
and U3481 (N_3481,N_1402,N_2434);
xnor U3482 (N_3482,N_2422,N_245);
or U3483 (N_3483,N_1049,N_1519);
and U3484 (N_3484,N_1157,N_2390);
nor U3485 (N_3485,N_195,N_436);
nor U3486 (N_3486,N_680,N_1191);
and U3487 (N_3487,N_286,N_85);
or U3488 (N_3488,N_1934,N_795);
or U3489 (N_3489,N_5,N_2479);
nor U3490 (N_3490,N_2329,N_2252);
xnor U3491 (N_3491,N_1281,N_1529);
xor U3492 (N_3492,N_1199,N_1190);
nand U3493 (N_3493,N_361,N_2407);
xnor U3494 (N_3494,N_2168,N_964);
or U3495 (N_3495,N_2279,N_1710);
nand U3496 (N_3496,N_292,N_1250);
xor U3497 (N_3497,N_401,N_358);
or U3498 (N_3498,N_1130,N_1896);
or U3499 (N_3499,N_1002,N_1074);
xor U3500 (N_3500,N_516,N_1156);
nor U3501 (N_3501,N_655,N_1714);
nand U3502 (N_3502,N_973,N_1817);
nand U3503 (N_3503,N_1476,N_2435);
nor U3504 (N_3504,N_77,N_2237);
or U3505 (N_3505,N_324,N_497);
nor U3506 (N_3506,N_1391,N_1517);
or U3507 (N_3507,N_1748,N_1935);
or U3508 (N_3508,N_639,N_2176);
and U3509 (N_3509,N_1956,N_2365);
xor U3510 (N_3510,N_1576,N_786);
nor U3511 (N_3511,N_1047,N_1);
nand U3512 (N_3512,N_2446,N_738);
or U3513 (N_3513,N_2327,N_1758);
xor U3514 (N_3514,N_2243,N_2360);
nand U3515 (N_3515,N_1742,N_1411);
and U3516 (N_3516,N_1470,N_433);
xnor U3517 (N_3517,N_1504,N_1712);
xor U3518 (N_3518,N_1388,N_591);
nand U3519 (N_3519,N_2074,N_2441);
xor U3520 (N_3520,N_1711,N_2271);
nor U3521 (N_3521,N_157,N_966);
or U3522 (N_3522,N_1686,N_2090);
nor U3523 (N_3523,N_1374,N_2137);
nor U3524 (N_3524,N_479,N_93);
or U3525 (N_3525,N_1537,N_1536);
and U3526 (N_3526,N_1230,N_2352);
or U3527 (N_3527,N_881,N_678);
nand U3528 (N_3528,N_192,N_2471);
or U3529 (N_3529,N_189,N_511);
and U3530 (N_3530,N_594,N_226);
and U3531 (N_3531,N_2299,N_1478);
xor U3532 (N_3532,N_957,N_2382);
nand U3533 (N_3533,N_1262,N_2393);
or U3534 (N_3534,N_168,N_617);
nor U3535 (N_3535,N_146,N_2001);
or U3536 (N_3536,N_1174,N_42);
and U3537 (N_3537,N_941,N_1761);
or U3538 (N_3538,N_354,N_487);
xor U3539 (N_3539,N_1557,N_517);
nor U3540 (N_3540,N_2234,N_6);
xor U3541 (N_3541,N_1940,N_2474);
xor U3542 (N_3542,N_783,N_1953);
or U3543 (N_3543,N_2005,N_139);
nand U3544 (N_3544,N_726,N_34);
or U3545 (N_3545,N_630,N_1889);
or U3546 (N_3546,N_1972,N_770);
xor U3547 (N_3547,N_1573,N_1549);
and U3548 (N_3548,N_2022,N_441);
xnor U3549 (N_3549,N_1416,N_2092);
and U3550 (N_3550,N_1913,N_171);
and U3551 (N_3551,N_1277,N_373);
nand U3552 (N_3552,N_368,N_1333);
or U3553 (N_3553,N_1267,N_1356);
xor U3554 (N_3554,N_331,N_68);
nand U3555 (N_3555,N_300,N_190);
nand U3556 (N_3556,N_2493,N_1715);
nor U3557 (N_3557,N_906,N_1143);
nor U3558 (N_3558,N_2025,N_1161);
nor U3559 (N_3559,N_1584,N_2295);
and U3560 (N_3560,N_774,N_314);
and U3561 (N_3561,N_812,N_719);
and U3562 (N_3562,N_115,N_2323);
nor U3563 (N_3563,N_2398,N_2044);
nand U3564 (N_3564,N_1309,N_1363);
and U3565 (N_3565,N_2457,N_760);
and U3566 (N_3566,N_22,N_365);
and U3567 (N_3567,N_637,N_1494);
or U3568 (N_3568,N_601,N_1815);
and U3569 (N_3569,N_1766,N_1072);
and U3570 (N_3570,N_1204,N_1868);
or U3571 (N_3571,N_166,N_1223);
nand U3572 (N_3572,N_1747,N_352);
nand U3573 (N_3573,N_2109,N_1129);
or U3574 (N_3574,N_2427,N_1620);
nand U3575 (N_3575,N_1086,N_1327);
or U3576 (N_3576,N_2130,N_1184);
or U3577 (N_3577,N_424,N_421);
and U3578 (N_3578,N_438,N_1609);
nand U3579 (N_3579,N_2460,N_121);
and U3580 (N_3580,N_1876,N_1893);
and U3581 (N_3581,N_1948,N_1113);
nand U3582 (N_3582,N_33,N_1781);
nand U3583 (N_3583,N_281,N_1533);
nor U3584 (N_3584,N_1906,N_432);
or U3585 (N_3585,N_1013,N_2341);
nand U3586 (N_3586,N_784,N_2331);
or U3587 (N_3587,N_1744,N_661);
xor U3588 (N_3588,N_1406,N_2135);
nand U3589 (N_3589,N_629,N_548);
xnor U3590 (N_3590,N_2373,N_308);
nand U3591 (N_3591,N_2394,N_2253);
or U3592 (N_3592,N_258,N_1364);
nor U3593 (N_3593,N_652,N_1417);
and U3594 (N_3594,N_2145,N_975);
xor U3595 (N_3595,N_898,N_88);
or U3596 (N_3596,N_1738,N_1226);
and U3597 (N_3597,N_393,N_586);
nand U3598 (N_3598,N_842,N_1615);
nand U3599 (N_3599,N_580,N_1825);
and U3600 (N_3600,N_2024,N_1941);
and U3601 (N_3601,N_2404,N_53);
or U3602 (N_3602,N_771,N_1720);
xnor U3603 (N_3603,N_625,N_2034);
nand U3604 (N_3604,N_434,N_555);
xor U3605 (N_3605,N_2348,N_899);
nor U3606 (N_3606,N_489,N_765);
nor U3607 (N_3607,N_2282,N_2121);
or U3608 (N_3608,N_44,N_1636);
xnor U3609 (N_3609,N_1362,N_803);
nor U3610 (N_3610,N_960,N_343);
nand U3611 (N_3611,N_330,N_1729);
nor U3612 (N_3612,N_1693,N_37);
nand U3613 (N_3613,N_482,N_374);
or U3614 (N_3614,N_29,N_624);
or U3615 (N_3615,N_2326,N_2367);
and U3616 (N_3616,N_125,N_2283);
or U3617 (N_3617,N_830,N_790);
nor U3618 (N_3618,N_237,N_2067);
nor U3619 (N_3619,N_2064,N_1846);
xnor U3620 (N_3620,N_1291,N_1621);
nand U3621 (N_3621,N_1069,N_1320);
and U3622 (N_3622,N_1661,N_1057);
or U3623 (N_3623,N_2304,N_1138);
xor U3624 (N_3624,N_297,N_344);
or U3625 (N_3625,N_566,N_642);
xnor U3626 (N_3626,N_1294,N_2153);
and U3627 (N_3627,N_2287,N_1111);
nor U3628 (N_3628,N_1980,N_2082);
nand U3629 (N_3629,N_2164,N_1012);
or U3630 (N_3630,N_2346,N_287);
or U3631 (N_3631,N_1452,N_1304);
and U3632 (N_3632,N_342,N_345);
nand U3633 (N_3633,N_721,N_1756);
and U3634 (N_3634,N_1978,N_1093);
or U3635 (N_3635,N_2155,N_1679);
nor U3636 (N_3636,N_2419,N_640);
and U3637 (N_3637,N_402,N_1792);
nand U3638 (N_3638,N_714,N_1205);
nand U3639 (N_3639,N_2464,N_1318);
nor U3640 (N_3640,N_1847,N_618);
nor U3641 (N_3641,N_1082,N_865);
nor U3642 (N_3642,N_808,N_1612);
and U3643 (N_3643,N_2099,N_1155);
xnor U3644 (N_3644,N_668,N_1905);
and U3645 (N_3645,N_496,N_1819);
or U3646 (N_3646,N_81,N_2335);
or U3647 (N_3647,N_2264,N_312);
nand U3648 (N_3648,N_2261,N_2220);
or U3649 (N_3649,N_2414,N_1297);
nor U3650 (N_3650,N_1777,N_1709);
nor U3651 (N_3651,N_2177,N_1999);
and U3652 (N_3652,N_667,N_1891);
xnor U3653 (N_3653,N_475,N_921);
nor U3654 (N_3654,N_272,N_2366);
nand U3655 (N_3655,N_1366,N_1514);
nor U3656 (N_3656,N_2016,N_2184);
nor U3657 (N_3657,N_1651,N_1667);
and U3658 (N_3658,N_990,N_442);
xnor U3659 (N_3659,N_472,N_2162);
nor U3660 (N_3660,N_247,N_690);
nand U3661 (N_3661,N_1750,N_1669);
nand U3662 (N_3662,N_1911,N_1252);
nor U3663 (N_3663,N_1912,N_1260);
or U3664 (N_3664,N_2019,N_1512);
nand U3665 (N_3665,N_537,N_56);
nor U3666 (N_3666,N_1377,N_2467);
nor U3667 (N_3667,N_1276,N_2284);
nand U3668 (N_3668,N_1946,N_2056);
and U3669 (N_3669,N_1235,N_602);
nand U3670 (N_3670,N_995,N_1255);
nor U3671 (N_3671,N_160,N_105);
or U3672 (N_3672,N_2488,N_2337);
nand U3673 (N_3673,N_1050,N_1739);
xor U3674 (N_3674,N_875,N_1144);
nor U3675 (N_3675,N_2096,N_1954);
or U3676 (N_3676,N_1672,N_276);
nor U3677 (N_3677,N_327,N_235);
xnor U3678 (N_3678,N_371,N_1596);
and U3679 (N_3679,N_65,N_551);
or U3680 (N_3680,N_1171,N_1676);
xnor U3681 (N_3681,N_1773,N_2449);
nor U3682 (N_3682,N_1765,N_97);
and U3683 (N_3683,N_1572,N_1456);
or U3684 (N_3684,N_1982,N_1347);
or U3685 (N_3685,N_2301,N_1942);
xnor U3686 (N_3686,N_2392,N_2277);
or U3687 (N_3687,N_1016,N_2377);
nand U3688 (N_3688,N_1701,N_1042);
nor U3689 (N_3689,N_1814,N_1663);
nand U3690 (N_3690,N_886,N_1429);
xor U3691 (N_3691,N_894,N_696);
nor U3692 (N_3692,N_895,N_353);
xnor U3693 (N_3693,N_2104,N_543);
or U3694 (N_3694,N_528,N_1432);
or U3695 (N_3695,N_1605,N_645);
nor U3696 (N_3696,N_1379,N_1021);
or U3697 (N_3697,N_2489,N_196);
nor U3698 (N_3698,N_1675,N_700);
nand U3699 (N_3699,N_1902,N_2262);
or U3700 (N_3700,N_1774,N_250);
nor U3701 (N_3701,N_644,N_665);
xor U3702 (N_3702,N_2416,N_1997);
nor U3703 (N_3703,N_2459,N_2447);
nor U3704 (N_3704,N_1440,N_520);
or U3705 (N_3705,N_532,N_458);
xnor U3706 (N_3706,N_599,N_163);
nand U3707 (N_3707,N_1339,N_940);
xnor U3708 (N_3708,N_209,N_78);
and U3709 (N_3709,N_2141,N_562);
and U3710 (N_3710,N_1212,N_1639);
or U3711 (N_3711,N_917,N_890);
or U3712 (N_3712,N_2068,N_1222);
nor U3713 (N_3713,N_1634,N_557);
or U3714 (N_3714,N_2086,N_1355);
nand U3715 (N_3715,N_1731,N_1020);
or U3716 (N_3716,N_271,N_26);
nor U3717 (N_3717,N_946,N_598);
or U3718 (N_3718,N_456,N_918);
nand U3719 (N_3719,N_569,N_1832);
and U3720 (N_3720,N_2037,N_1850);
nand U3721 (N_3721,N_273,N_174);
nor U3722 (N_3722,N_538,N_1754);
nor U3723 (N_3723,N_1592,N_1628);
nor U3724 (N_3724,N_1058,N_1232);
nor U3725 (N_3725,N_742,N_1901);
or U3726 (N_3726,N_307,N_846);
and U3727 (N_3727,N_1310,N_1888);
xnor U3728 (N_3728,N_2195,N_2486);
or U3729 (N_3729,N_255,N_521);
or U3730 (N_3730,N_884,N_2322);
nand U3731 (N_3731,N_1685,N_802);
xnor U3732 (N_3732,N_1426,N_1482);
nand U3733 (N_3733,N_1705,N_1248);
nor U3734 (N_3734,N_227,N_2430);
nand U3735 (N_3735,N_1479,N_578);
nor U3736 (N_3736,N_1449,N_1862);
nor U3737 (N_3737,N_1352,N_0);
and U3738 (N_3738,N_178,N_395);
nor U3739 (N_3739,N_2478,N_1292);
or U3740 (N_3740,N_2159,N_2230);
xor U3741 (N_3741,N_2475,N_1442);
nand U3742 (N_3742,N_1565,N_2106);
xor U3743 (N_3743,N_1039,N_1857);
nor U3744 (N_3744,N_251,N_2256);
or U3745 (N_3745,N_885,N_2076);
nand U3746 (N_3746,N_2158,N_2189);
xor U3747 (N_3747,N_79,N_1863);
xnor U3748 (N_3748,N_2187,N_75);
xnor U3749 (N_3749,N_1465,N_1128);
nor U3750 (N_3750,N_10,N_2028);
or U3751 (N_3751,N_1709,N_10);
xor U3752 (N_3752,N_943,N_304);
and U3753 (N_3753,N_986,N_191);
nor U3754 (N_3754,N_754,N_1928);
and U3755 (N_3755,N_1538,N_752);
or U3756 (N_3756,N_2262,N_1730);
nand U3757 (N_3757,N_1911,N_1011);
and U3758 (N_3758,N_2273,N_682);
nor U3759 (N_3759,N_2030,N_215);
or U3760 (N_3760,N_730,N_110);
and U3761 (N_3761,N_1538,N_66);
nor U3762 (N_3762,N_2135,N_2134);
nand U3763 (N_3763,N_2096,N_1851);
and U3764 (N_3764,N_1531,N_2411);
nor U3765 (N_3765,N_2008,N_571);
nor U3766 (N_3766,N_585,N_2376);
or U3767 (N_3767,N_1175,N_2409);
xor U3768 (N_3768,N_1123,N_95);
xor U3769 (N_3769,N_2384,N_53);
and U3770 (N_3770,N_1652,N_676);
nand U3771 (N_3771,N_913,N_1122);
or U3772 (N_3772,N_2235,N_510);
nor U3773 (N_3773,N_175,N_2446);
and U3774 (N_3774,N_1231,N_2188);
nand U3775 (N_3775,N_1269,N_1724);
nand U3776 (N_3776,N_199,N_810);
or U3777 (N_3777,N_382,N_2023);
xor U3778 (N_3778,N_184,N_282);
xor U3779 (N_3779,N_1044,N_2473);
or U3780 (N_3780,N_937,N_240);
nand U3781 (N_3781,N_2393,N_1788);
xor U3782 (N_3782,N_195,N_2109);
or U3783 (N_3783,N_380,N_2476);
nand U3784 (N_3784,N_761,N_1245);
nor U3785 (N_3785,N_1148,N_1907);
and U3786 (N_3786,N_270,N_138);
and U3787 (N_3787,N_648,N_768);
nor U3788 (N_3788,N_2077,N_1296);
nor U3789 (N_3789,N_1062,N_40);
or U3790 (N_3790,N_793,N_539);
or U3791 (N_3791,N_0,N_1879);
and U3792 (N_3792,N_80,N_1362);
and U3793 (N_3793,N_1259,N_35);
or U3794 (N_3794,N_621,N_1808);
nand U3795 (N_3795,N_1543,N_1613);
xor U3796 (N_3796,N_483,N_1293);
xnor U3797 (N_3797,N_718,N_282);
nand U3798 (N_3798,N_1528,N_1341);
nor U3799 (N_3799,N_1148,N_2417);
xnor U3800 (N_3800,N_715,N_2114);
nor U3801 (N_3801,N_1614,N_452);
nor U3802 (N_3802,N_1216,N_173);
and U3803 (N_3803,N_1385,N_1199);
and U3804 (N_3804,N_2346,N_207);
and U3805 (N_3805,N_46,N_2211);
xor U3806 (N_3806,N_2047,N_1869);
nor U3807 (N_3807,N_2343,N_213);
and U3808 (N_3808,N_1972,N_1390);
and U3809 (N_3809,N_2056,N_915);
xnor U3810 (N_3810,N_2295,N_326);
or U3811 (N_3811,N_1794,N_2228);
nand U3812 (N_3812,N_850,N_1912);
nor U3813 (N_3813,N_640,N_412);
and U3814 (N_3814,N_604,N_2407);
nand U3815 (N_3815,N_2059,N_1253);
nand U3816 (N_3816,N_667,N_1460);
and U3817 (N_3817,N_1859,N_1690);
nor U3818 (N_3818,N_312,N_1019);
nand U3819 (N_3819,N_1515,N_1863);
nand U3820 (N_3820,N_1891,N_2407);
and U3821 (N_3821,N_2445,N_2164);
xor U3822 (N_3822,N_97,N_149);
nor U3823 (N_3823,N_1816,N_898);
or U3824 (N_3824,N_2363,N_1003);
nand U3825 (N_3825,N_1744,N_1846);
nor U3826 (N_3826,N_333,N_65);
or U3827 (N_3827,N_1336,N_933);
nand U3828 (N_3828,N_2495,N_495);
nor U3829 (N_3829,N_1310,N_2011);
nand U3830 (N_3830,N_526,N_1924);
nand U3831 (N_3831,N_828,N_725);
or U3832 (N_3832,N_351,N_217);
nand U3833 (N_3833,N_1435,N_208);
nand U3834 (N_3834,N_1502,N_1109);
or U3835 (N_3835,N_1461,N_107);
xnor U3836 (N_3836,N_39,N_1081);
or U3837 (N_3837,N_2409,N_101);
nand U3838 (N_3838,N_2099,N_476);
nor U3839 (N_3839,N_2412,N_1202);
nand U3840 (N_3840,N_1264,N_1255);
and U3841 (N_3841,N_647,N_485);
nand U3842 (N_3842,N_139,N_1623);
nand U3843 (N_3843,N_117,N_1075);
and U3844 (N_3844,N_1315,N_2470);
or U3845 (N_3845,N_2331,N_387);
xnor U3846 (N_3846,N_1017,N_1119);
or U3847 (N_3847,N_979,N_2040);
or U3848 (N_3848,N_2478,N_815);
and U3849 (N_3849,N_2273,N_1277);
or U3850 (N_3850,N_1064,N_1391);
nor U3851 (N_3851,N_1463,N_1113);
or U3852 (N_3852,N_1859,N_2444);
nand U3853 (N_3853,N_1615,N_2017);
nand U3854 (N_3854,N_1268,N_1122);
or U3855 (N_3855,N_2001,N_131);
xnor U3856 (N_3856,N_598,N_762);
xnor U3857 (N_3857,N_1377,N_2183);
xor U3858 (N_3858,N_158,N_2001);
and U3859 (N_3859,N_1631,N_1590);
xnor U3860 (N_3860,N_262,N_1927);
nor U3861 (N_3861,N_2112,N_1858);
xnor U3862 (N_3862,N_1584,N_1214);
xor U3863 (N_3863,N_1673,N_189);
nor U3864 (N_3864,N_2212,N_225);
xor U3865 (N_3865,N_1714,N_735);
nor U3866 (N_3866,N_1814,N_1309);
nand U3867 (N_3867,N_1935,N_515);
nor U3868 (N_3868,N_671,N_1711);
nand U3869 (N_3869,N_473,N_2358);
nor U3870 (N_3870,N_1735,N_893);
nor U3871 (N_3871,N_661,N_2084);
nor U3872 (N_3872,N_1080,N_228);
or U3873 (N_3873,N_2395,N_1748);
and U3874 (N_3874,N_2161,N_309);
nand U3875 (N_3875,N_2382,N_1103);
xor U3876 (N_3876,N_821,N_1743);
and U3877 (N_3877,N_294,N_1062);
xor U3878 (N_3878,N_1197,N_2210);
and U3879 (N_3879,N_1486,N_636);
or U3880 (N_3880,N_312,N_1448);
or U3881 (N_3881,N_283,N_180);
xnor U3882 (N_3882,N_584,N_91);
or U3883 (N_3883,N_556,N_2045);
and U3884 (N_3884,N_551,N_442);
nor U3885 (N_3885,N_113,N_2337);
xnor U3886 (N_3886,N_1251,N_1452);
nand U3887 (N_3887,N_1702,N_383);
nor U3888 (N_3888,N_1154,N_1748);
and U3889 (N_3889,N_155,N_1976);
or U3890 (N_3890,N_1767,N_2067);
and U3891 (N_3891,N_1506,N_2433);
and U3892 (N_3892,N_202,N_534);
nor U3893 (N_3893,N_2304,N_1411);
and U3894 (N_3894,N_2131,N_2249);
and U3895 (N_3895,N_531,N_754);
nor U3896 (N_3896,N_1839,N_1673);
or U3897 (N_3897,N_1571,N_2263);
xnor U3898 (N_3898,N_444,N_876);
xor U3899 (N_3899,N_983,N_1676);
or U3900 (N_3900,N_2473,N_1017);
xor U3901 (N_3901,N_434,N_936);
or U3902 (N_3902,N_524,N_882);
and U3903 (N_3903,N_2138,N_785);
nand U3904 (N_3904,N_2385,N_1959);
or U3905 (N_3905,N_562,N_1108);
xnor U3906 (N_3906,N_1422,N_1622);
nand U3907 (N_3907,N_1647,N_97);
nor U3908 (N_3908,N_1234,N_3);
nor U3909 (N_3909,N_18,N_1322);
nor U3910 (N_3910,N_356,N_2200);
nor U3911 (N_3911,N_2003,N_70);
nor U3912 (N_3912,N_2387,N_800);
or U3913 (N_3913,N_2373,N_1661);
nor U3914 (N_3914,N_955,N_2051);
nand U3915 (N_3915,N_2498,N_1619);
or U3916 (N_3916,N_1742,N_2024);
nand U3917 (N_3917,N_2442,N_824);
nor U3918 (N_3918,N_1225,N_568);
and U3919 (N_3919,N_2311,N_1875);
nor U3920 (N_3920,N_432,N_2458);
or U3921 (N_3921,N_1210,N_849);
nand U3922 (N_3922,N_1105,N_755);
xnor U3923 (N_3923,N_2308,N_658);
nor U3924 (N_3924,N_1159,N_1663);
and U3925 (N_3925,N_1513,N_749);
nand U3926 (N_3926,N_1420,N_1827);
xor U3927 (N_3927,N_2007,N_1806);
or U3928 (N_3928,N_1769,N_1003);
nor U3929 (N_3929,N_1936,N_1524);
nor U3930 (N_3930,N_194,N_2377);
nor U3931 (N_3931,N_693,N_1654);
nand U3932 (N_3932,N_508,N_2134);
or U3933 (N_3933,N_2370,N_10);
or U3934 (N_3934,N_1202,N_1985);
or U3935 (N_3935,N_1183,N_1735);
nor U3936 (N_3936,N_411,N_2081);
nand U3937 (N_3937,N_1747,N_543);
nor U3938 (N_3938,N_2068,N_1879);
nor U3939 (N_3939,N_942,N_1093);
nand U3940 (N_3940,N_613,N_80);
nor U3941 (N_3941,N_909,N_955);
or U3942 (N_3942,N_2455,N_1373);
nor U3943 (N_3943,N_1989,N_250);
nand U3944 (N_3944,N_2091,N_1365);
or U3945 (N_3945,N_2129,N_659);
nand U3946 (N_3946,N_2138,N_2223);
nor U3947 (N_3947,N_1281,N_195);
or U3948 (N_3948,N_2283,N_342);
or U3949 (N_3949,N_1105,N_252);
xnor U3950 (N_3950,N_773,N_1443);
xnor U3951 (N_3951,N_1501,N_1508);
nor U3952 (N_3952,N_2475,N_658);
or U3953 (N_3953,N_394,N_359);
nand U3954 (N_3954,N_756,N_1175);
xor U3955 (N_3955,N_1619,N_873);
xor U3956 (N_3956,N_53,N_2057);
xnor U3957 (N_3957,N_573,N_176);
and U3958 (N_3958,N_2165,N_2383);
xor U3959 (N_3959,N_2251,N_1571);
nor U3960 (N_3960,N_155,N_2424);
or U3961 (N_3961,N_816,N_432);
and U3962 (N_3962,N_477,N_1544);
nor U3963 (N_3963,N_815,N_258);
nor U3964 (N_3964,N_884,N_437);
and U3965 (N_3965,N_1277,N_2075);
nand U3966 (N_3966,N_494,N_1695);
and U3967 (N_3967,N_1680,N_741);
or U3968 (N_3968,N_729,N_1233);
xor U3969 (N_3969,N_1032,N_994);
xnor U3970 (N_3970,N_292,N_490);
and U3971 (N_3971,N_2381,N_630);
and U3972 (N_3972,N_663,N_1092);
or U3973 (N_3973,N_1426,N_990);
or U3974 (N_3974,N_1183,N_2016);
or U3975 (N_3975,N_1511,N_676);
xor U3976 (N_3976,N_1324,N_152);
nor U3977 (N_3977,N_1584,N_1233);
nor U3978 (N_3978,N_596,N_1369);
xor U3979 (N_3979,N_2452,N_56);
or U3980 (N_3980,N_1289,N_115);
nor U3981 (N_3981,N_2176,N_1983);
xnor U3982 (N_3982,N_345,N_1458);
and U3983 (N_3983,N_767,N_1749);
xnor U3984 (N_3984,N_1483,N_1939);
nand U3985 (N_3985,N_368,N_2376);
nand U3986 (N_3986,N_2235,N_1752);
and U3987 (N_3987,N_617,N_2328);
or U3988 (N_3988,N_1317,N_1633);
nor U3989 (N_3989,N_2311,N_2422);
or U3990 (N_3990,N_259,N_2384);
nand U3991 (N_3991,N_1260,N_148);
nor U3992 (N_3992,N_1773,N_1275);
nand U3993 (N_3993,N_2213,N_2317);
nor U3994 (N_3994,N_1916,N_29);
xnor U3995 (N_3995,N_1274,N_342);
and U3996 (N_3996,N_1827,N_1220);
or U3997 (N_3997,N_1053,N_295);
or U3998 (N_3998,N_408,N_1695);
or U3999 (N_3999,N_1543,N_1988);
or U4000 (N_4000,N_474,N_428);
and U4001 (N_4001,N_168,N_1933);
nand U4002 (N_4002,N_2177,N_2317);
and U4003 (N_4003,N_1545,N_418);
nand U4004 (N_4004,N_1063,N_984);
nor U4005 (N_4005,N_1422,N_839);
and U4006 (N_4006,N_1228,N_70);
nor U4007 (N_4007,N_1168,N_871);
nand U4008 (N_4008,N_1595,N_2390);
or U4009 (N_4009,N_4,N_799);
or U4010 (N_4010,N_1836,N_2141);
nor U4011 (N_4011,N_2297,N_914);
nor U4012 (N_4012,N_2026,N_669);
or U4013 (N_4013,N_1990,N_1544);
nor U4014 (N_4014,N_2179,N_417);
nand U4015 (N_4015,N_1268,N_1286);
nor U4016 (N_4016,N_731,N_2380);
nor U4017 (N_4017,N_907,N_2462);
and U4018 (N_4018,N_1675,N_1962);
or U4019 (N_4019,N_525,N_967);
and U4020 (N_4020,N_1506,N_194);
nor U4021 (N_4021,N_1465,N_1727);
or U4022 (N_4022,N_1426,N_527);
xor U4023 (N_4023,N_261,N_1101);
or U4024 (N_4024,N_537,N_1015);
nand U4025 (N_4025,N_1006,N_1961);
xnor U4026 (N_4026,N_1439,N_2413);
and U4027 (N_4027,N_2313,N_150);
xor U4028 (N_4028,N_2443,N_104);
or U4029 (N_4029,N_1391,N_1518);
xor U4030 (N_4030,N_2293,N_32);
nor U4031 (N_4031,N_101,N_1167);
nor U4032 (N_4032,N_1966,N_2082);
nor U4033 (N_4033,N_1443,N_669);
nor U4034 (N_4034,N_1,N_254);
and U4035 (N_4035,N_1916,N_1515);
nand U4036 (N_4036,N_2407,N_263);
nor U4037 (N_4037,N_2298,N_1799);
or U4038 (N_4038,N_569,N_702);
nand U4039 (N_4039,N_2288,N_1766);
nand U4040 (N_4040,N_796,N_1686);
or U4041 (N_4041,N_1743,N_696);
and U4042 (N_4042,N_959,N_1832);
and U4043 (N_4043,N_2491,N_2418);
nand U4044 (N_4044,N_2308,N_1573);
nand U4045 (N_4045,N_35,N_1046);
or U4046 (N_4046,N_1024,N_2304);
nand U4047 (N_4047,N_1559,N_807);
or U4048 (N_4048,N_2193,N_1060);
nand U4049 (N_4049,N_455,N_2081);
or U4050 (N_4050,N_2076,N_1714);
and U4051 (N_4051,N_1669,N_1821);
and U4052 (N_4052,N_963,N_1384);
or U4053 (N_4053,N_700,N_864);
nand U4054 (N_4054,N_789,N_836);
or U4055 (N_4055,N_1018,N_2109);
and U4056 (N_4056,N_1171,N_2249);
nor U4057 (N_4057,N_1696,N_1236);
xor U4058 (N_4058,N_1422,N_842);
and U4059 (N_4059,N_845,N_933);
nor U4060 (N_4060,N_1905,N_937);
nand U4061 (N_4061,N_2347,N_833);
xor U4062 (N_4062,N_1072,N_2294);
nand U4063 (N_4063,N_1491,N_1804);
or U4064 (N_4064,N_1524,N_689);
nor U4065 (N_4065,N_1380,N_1275);
and U4066 (N_4066,N_1537,N_1398);
xnor U4067 (N_4067,N_2190,N_1122);
nor U4068 (N_4068,N_2377,N_1886);
xnor U4069 (N_4069,N_1513,N_115);
or U4070 (N_4070,N_1925,N_1181);
xnor U4071 (N_4071,N_95,N_2326);
nand U4072 (N_4072,N_938,N_1777);
or U4073 (N_4073,N_2053,N_953);
and U4074 (N_4074,N_2366,N_169);
xor U4075 (N_4075,N_479,N_602);
and U4076 (N_4076,N_1507,N_1971);
or U4077 (N_4077,N_1227,N_2206);
or U4078 (N_4078,N_536,N_1730);
xnor U4079 (N_4079,N_1945,N_1319);
or U4080 (N_4080,N_961,N_1570);
or U4081 (N_4081,N_566,N_329);
xor U4082 (N_4082,N_842,N_653);
and U4083 (N_4083,N_2387,N_2341);
or U4084 (N_4084,N_1312,N_1473);
nand U4085 (N_4085,N_1360,N_866);
or U4086 (N_4086,N_1494,N_1190);
nand U4087 (N_4087,N_674,N_2141);
or U4088 (N_4088,N_279,N_1358);
or U4089 (N_4089,N_1174,N_1630);
xor U4090 (N_4090,N_2292,N_2117);
xor U4091 (N_4091,N_2138,N_1883);
or U4092 (N_4092,N_1609,N_1608);
xnor U4093 (N_4093,N_2148,N_146);
xor U4094 (N_4094,N_1652,N_1781);
xor U4095 (N_4095,N_2110,N_1185);
and U4096 (N_4096,N_291,N_1043);
nor U4097 (N_4097,N_330,N_1941);
xnor U4098 (N_4098,N_308,N_2413);
or U4099 (N_4099,N_2334,N_99);
xnor U4100 (N_4100,N_1908,N_745);
and U4101 (N_4101,N_1693,N_176);
xnor U4102 (N_4102,N_1508,N_432);
and U4103 (N_4103,N_1542,N_836);
nand U4104 (N_4104,N_2211,N_1541);
nand U4105 (N_4105,N_272,N_669);
nand U4106 (N_4106,N_700,N_546);
xnor U4107 (N_4107,N_1787,N_1135);
xor U4108 (N_4108,N_410,N_82);
xor U4109 (N_4109,N_832,N_853);
or U4110 (N_4110,N_2042,N_1042);
nor U4111 (N_4111,N_570,N_1095);
nand U4112 (N_4112,N_521,N_1496);
xor U4113 (N_4113,N_2127,N_30);
nand U4114 (N_4114,N_947,N_2257);
nor U4115 (N_4115,N_787,N_2409);
nor U4116 (N_4116,N_1698,N_192);
or U4117 (N_4117,N_626,N_1490);
nand U4118 (N_4118,N_2270,N_944);
and U4119 (N_4119,N_1682,N_1668);
and U4120 (N_4120,N_2080,N_52);
and U4121 (N_4121,N_2347,N_852);
and U4122 (N_4122,N_2003,N_2060);
nand U4123 (N_4123,N_1570,N_1529);
nand U4124 (N_4124,N_2043,N_1648);
xnor U4125 (N_4125,N_1458,N_377);
and U4126 (N_4126,N_1870,N_689);
xnor U4127 (N_4127,N_1558,N_1031);
nor U4128 (N_4128,N_708,N_2377);
xnor U4129 (N_4129,N_641,N_393);
and U4130 (N_4130,N_776,N_1135);
and U4131 (N_4131,N_441,N_333);
and U4132 (N_4132,N_249,N_558);
xnor U4133 (N_4133,N_906,N_755);
or U4134 (N_4134,N_2338,N_1088);
nand U4135 (N_4135,N_1007,N_2018);
nand U4136 (N_4136,N_400,N_1867);
nor U4137 (N_4137,N_2277,N_1252);
xnor U4138 (N_4138,N_2181,N_1563);
or U4139 (N_4139,N_2237,N_369);
xnor U4140 (N_4140,N_555,N_2159);
or U4141 (N_4141,N_1149,N_144);
and U4142 (N_4142,N_2203,N_531);
nand U4143 (N_4143,N_1374,N_570);
or U4144 (N_4144,N_1012,N_1625);
nor U4145 (N_4145,N_8,N_1048);
and U4146 (N_4146,N_2126,N_1617);
xor U4147 (N_4147,N_1356,N_688);
xor U4148 (N_4148,N_989,N_2351);
or U4149 (N_4149,N_1501,N_1701);
or U4150 (N_4150,N_2351,N_1670);
xor U4151 (N_4151,N_1207,N_893);
nor U4152 (N_4152,N_392,N_893);
xor U4153 (N_4153,N_1552,N_1122);
nand U4154 (N_4154,N_1657,N_1415);
nand U4155 (N_4155,N_1411,N_1891);
or U4156 (N_4156,N_666,N_1738);
and U4157 (N_4157,N_2048,N_2343);
xor U4158 (N_4158,N_669,N_1752);
nor U4159 (N_4159,N_960,N_2098);
nor U4160 (N_4160,N_579,N_1715);
xnor U4161 (N_4161,N_2034,N_535);
nand U4162 (N_4162,N_1963,N_1065);
or U4163 (N_4163,N_2229,N_1933);
or U4164 (N_4164,N_234,N_1168);
and U4165 (N_4165,N_1407,N_794);
xor U4166 (N_4166,N_506,N_337);
or U4167 (N_4167,N_2202,N_571);
and U4168 (N_4168,N_898,N_959);
and U4169 (N_4169,N_1047,N_147);
nor U4170 (N_4170,N_898,N_1352);
and U4171 (N_4171,N_2343,N_2145);
or U4172 (N_4172,N_1836,N_594);
and U4173 (N_4173,N_2360,N_486);
xnor U4174 (N_4174,N_918,N_1596);
and U4175 (N_4175,N_1776,N_744);
xor U4176 (N_4176,N_2322,N_1965);
nand U4177 (N_4177,N_1518,N_2364);
and U4178 (N_4178,N_444,N_402);
and U4179 (N_4179,N_292,N_1874);
nor U4180 (N_4180,N_972,N_470);
or U4181 (N_4181,N_1981,N_1036);
nor U4182 (N_4182,N_1483,N_2431);
nand U4183 (N_4183,N_1898,N_115);
xnor U4184 (N_4184,N_913,N_2389);
and U4185 (N_4185,N_1929,N_2442);
nor U4186 (N_4186,N_805,N_882);
or U4187 (N_4187,N_1311,N_1711);
nor U4188 (N_4188,N_1237,N_1112);
and U4189 (N_4189,N_743,N_2463);
or U4190 (N_4190,N_328,N_2181);
nand U4191 (N_4191,N_2258,N_2134);
xnor U4192 (N_4192,N_119,N_240);
nor U4193 (N_4193,N_1480,N_958);
nor U4194 (N_4194,N_1655,N_1922);
xnor U4195 (N_4195,N_2293,N_2176);
or U4196 (N_4196,N_786,N_710);
and U4197 (N_4197,N_2364,N_1366);
or U4198 (N_4198,N_1332,N_2216);
and U4199 (N_4199,N_1598,N_328);
nor U4200 (N_4200,N_2056,N_2095);
or U4201 (N_4201,N_1326,N_489);
xnor U4202 (N_4202,N_1869,N_19);
and U4203 (N_4203,N_1039,N_863);
xor U4204 (N_4204,N_946,N_778);
or U4205 (N_4205,N_1950,N_1792);
xnor U4206 (N_4206,N_830,N_883);
nand U4207 (N_4207,N_1155,N_649);
or U4208 (N_4208,N_1647,N_1079);
nand U4209 (N_4209,N_2379,N_1002);
and U4210 (N_4210,N_2098,N_1928);
xnor U4211 (N_4211,N_2449,N_443);
or U4212 (N_4212,N_214,N_2382);
or U4213 (N_4213,N_714,N_995);
nor U4214 (N_4214,N_97,N_814);
xnor U4215 (N_4215,N_1277,N_515);
and U4216 (N_4216,N_1446,N_2310);
nand U4217 (N_4217,N_1493,N_1898);
or U4218 (N_4218,N_1749,N_2184);
or U4219 (N_4219,N_1232,N_2299);
and U4220 (N_4220,N_251,N_443);
and U4221 (N_4221,N_812,N_305);
xnor U4222 (N_4222,N_2452,N_49);
or U4223 (N_4223,N_358,N_1600);
nand U4224 (N_4224,N_2217,N_2070);
or U4225 (N_4225,N_1921,N_1608);
xor U4226 (N_4226,N_421,N_1315);
or U4227 (N_4227,N_700,N_1739);
nand U4228 (N_4228,N_604,N_351);
xnor U4229 (N_4229,N_472,N_178);
or U4230 (N_4230,N_678,N_1588);
and U4231 (N_4231,N_1930,N_1833);
xnor U4232 (N_4232,N_1824,N_1265);
and U4233 (N_4233,N_1805,N_335);
xor U4234 (N_4234,N_373,N_2120);
nand U4235 (N_4235,N_1842,N_2292);
nor U4236 (N_4236,N_1541,N_2021);
or U4237 (N_4237,N_1593,N_1179);
nand U4238 (N_4238,N_804,N_1058);
and U4239 (N_4239,N_627,N_2447);
nand U4240 (N_4240,N_594,N_1537);
and U4241 (N_4241,N_1553,N_468);
or U4242 (N_4242,N_360,N_1208);
nand U4243 (N_4243,N_569,N_428);
nor U4244 (N_4244,N_2423,N_263);
nor U4245 (N_4245,N_1679,N_211);
or U4246 (N_4246,N_1573,N_2202);
and U4247 (N_4247,N_2122,N_551);
xnor U4248 (N_4248,N_1287,N_459);
or U4249 (N_4249,N_2463,N_1961);
nand U4250 (N_4250,N_2410,N_190);
or U4251 (N_4251,N_1794,N_1850);
and U4252 (N_4252,N_1731,N_1254);
and U4253 (N_4253,N_2273,N_1763);
or U4254 (N_4254,N_114,N_1722);
or U4255 (N_4255,N_1326,N_1702);
xor U4256 (N_4256,N_516,N_157);
or U4257 (N_4257,N_376,N_1988);
and U4258 (N_4258,N_1601,N_1921);
nor U4259 (N_4259,N_702,N_1460);
xnor U4260 (N_4260,N_2154,N_2029);
or U4261 (N_4261,N_717,N_1427);
nand U4262 (N_4262,N_2200,N_2052);
nor U4263 (N_4263,N_488,N_621);
nor U4264 (N_4264,N_1754,N_841);
xnor U4265 (N_4265,N_528,N_2369);
nand U4266 (N_4266,N_2474,N_874);
and U4267 (N_4267,N_2428,N_1859);
nor U4268 (N_4268,N_2136,N_533);
and U4269 (N_4269,N_1547,N_420);
or U4270 (N_4270,N_2347,N_2140);
xnor U4271 (N_4271,N_1946,N_1810);
nor U4272 (N_4272,N_1200,N_133);
nor U4273 (N_4273,N_1781,N_877);
nor U4274 (N_4274,N_616,N_1323);
and U4275 (N_4275,N_213,N_597);
nand U4276 (N_4276,N_243,N_2445);
and U4277 (N_4277,N_2222,N_2480);
or U4278 (N_4278,N_2227,N_1997);
and U4279 (N_4279,N_457,N_188);
nand U4280 (N_4280,N_1864,N_2220);
or U4281 (N_4281,N_2078,N_1922);
xnor U4282 (N_4282,N_2008,N_2290);
or U4283 (N_4283,N_2488,N_669);
nand U4284 (N_4284,N_1984,N_1588);
or U4285 (N_4285,N_2080,N_637);
xor U4286 (N_4286,N_803,N_330);
xnor U4287 (N_4287,N_1597,N_447);
or U4288 (N_4288,N_191,N_1532);
nand U4289 (N_4289,N_704,N_560);
xor U4290 (N_4290,N_355,N_1578);
xor U4291 (N_4291,N_2263,N_360);
or U4292 (N_4292,N_251,N_2072);
or U4293 (N_4293,N_1138,N_138);
xnor U4294 (N_4294,N_768,N_206);
nand U4295 (N_4295,N_2387,N_1994);
nor U4296 (N_4296,N_1019,N_212);
nand U4297 (N_4297,N_5,N_1563);
or U4298 (N_4298,N_1187,N_2160);
and U4299 (N_4299,N_1897,N_1619);
nand U4300 (N_4300,N_353,N_2051);
xnor U4301 (N_4301,N_1623,N_1355);
xor U4302 (N_4302,N_1158,N_1880);
and U4303 (N_4303,N_2450,N_1222);
and U4304 (N_4304,N_1402,N_1512);
and U4305 (N_4305,N_1299,N_132);
nand U4306 (N_4306,N_1650,N_1662);
xor U4307 (N_4307,N_372,N_2317);
and U4308 (N_4308,N_1860,N_1297);
nand U4309 (N_4309,N_1303,N_403);
or U4310 (N_4310,N_327,N_1993);
or U4311 (N_4311,N_533,N_474);
nor U4312 (N_4312,N_848,N_105);
or U4313 (N_4313,N_954,N_1223);
and U4314 (N_4314,N_47,N_233);
xor U4315 (N_4315,N_2071,N_2008);
nor U4316 (N_4316,N_608,N_704);
and U4317 (N_4317,N_573,N_1389);
nor U4318 (N_4318,N_2434,N_375);
nor U4319 (N_4319,N_2059,N_483);
nor U4320 (N_4320,N_1405,N_465);
and U4321 (N_4321,N_1786,N_842);
nor U4322 (N_4322,N_1065,N_2097);
and U4323 (N_4323,N_1508,N_862);
nor U4324 (N_4324,N_1788,N_830);
xnor U4325 (N_4325,N_2312,N_630);
or U4326 (N_4326,N_566,N_1224);
nand U4327 (N_4327,N_2131,N_1187);
or U4328 (N_4328,N_1010,N_1173);
xnor U4329 (N_4329,N_1153,N_1477);
xnor U4330 (N_4330,N_865,N_1167);
and U4331 (N_4331,N_2048,N_341);
nand U4332 (N_4332,N_1212,N_1647);
nand U4333 (N_4333,N_89,N_1340);
and U4334 (N_4334,N_340,N_1450);
or U4335 (N_4335,N_1637,N_1894);
and U4336 (N_4336,N_1819,N_2002);
xor U4337 (N_4337,N_764,N_926);
or U4338 (N_4338,N_2415,N_2141);
nand U4339 (N_4339,N_434,N_2142);
xnor U4340 (N_4340,N_1226,N_1770);
and U4341 (N_4341,N_2481,N_646);
xor U4342 (N_4342,N_807,N_2106);
nand U4343 (N_4343,N_1502,N_1675);
nor U4344 (N_4344,N_1887,N_1634);
nand U4345 (N_4345,N_1917,N_1245);
xor U4346 (N_4346,N_585,N_178);
xnor U4347 (N_4347,N_1105,N_674);
nor U4348 (N_4348,N_1666,N_2308);
nand U4349 (N_4349,N_2217,N_457);
xor U4350 (N_4350,N_739,N_363);
nor U4351 (N_4351,N_1257,N_1739);
xor U4352 (N_4352,N_802,N_509);
or U4353 (N_4353,N_61,N_1898);
and U4354 (N_4354,N_1832,N_157);
nor U4355 (N_4355,N_2172,N_2438);
nand U4356 (N_4356,N_2051,N_283);
or U4357 (N_4357,N_1900,N_1276);
nor U4358 (N_4358,N_184,N_2344);
nor U4359 (N_4359,N_1235,N_1332);
and U4360 (N_4360,N_1740,N_327);
xor U4361 (N_4361,N_1680,N_2163);
xnor U4362 (N_4362,N_387,N_1672);
xor U4363 (N_4363,N_2243,N_1725);
nand U4364 (N_4364,N_1365,N_1054);
and U4365 (N_4365,N_1980,N_2420);
nor U4366 (N_4366,N_2078,N_1284);
nand U4367 (N_4367,N_1591,N_282);
nand U4368 (N_4368,N_90,N_1130);
and U4369 (N_4369,N_491,N_2413);
xnor U4370 (N_4370,N_1397,N_1589);
xor U4371 (N_4371,N_186,N_1424);
nor U4372 (N_4372,N_2344,N_1235);
or U4373 (N_4373,N_2460,N_1234);
nor U4374 (N_4374,N_944,N_2003);
or U4375 (N_4375,N_1494,N_1135);
or U4376 (N_4376,N_1968,N_913);
nand U4377 (N_4377,N_701,N_1288);
and U4378 (N_4378,N_94,N_2165);
xor U4379 (N_4379,N_484,N_240);
and U4380 (N_4380,N_1330,N_809);
xnor U4381 (N_4381,N_693,N_772);
nor U4382 (N_4382,N_2175,N_822);
or U4383 (N_4383,N_120,N_63);
and U4384 (N_4384,N_1990,N_450);
nand U4385 (N_4385,N_270,N_199);
xnor U4386 (N_4386,N_1115,N_111);
nand U4387 (N_4387,N_1296,N_921);
xor U4388 (N_4388,N_573,N_1010);
or U4389 (N_4389,N_1156,N_339);
xor U4390 (N_4390,N_1471,N_974);
nor U4391 (N_4391,N_2220,N_338);
nand U4392 (N_4392,N_2080,N_1922);
or U4393 (N_4393,N_178,N_1430);
and U4394 (N_4394,N_1616,N_1300);
and U4395 (N_4395,N_2465,N_1164);
nor U4396 (N_4396,N_668,N_2475);
xnor U4397 (N_4397,N_1995,N_2086);
xor U4398 (N_4398,N_1671,N_211);
xnor U4399 (N_4399,N_109,N_2313);
and U4400 (N_4400,N_939,N_704);
xnor U4401 (N_4401,N_965,N_449);
nor U4402 (N_4402,N_31,N_1384);
or U4403 (N_4403,N_2351,N_124);
or U4404 (N_4404,N_2374,N_1280);
and U4405 (N_4405,N_1034,N_1269);
nor U4406 (N_4406,N_688,N_549);
or U4407 (N_4407,N_2120,N_1872);
or U4408 (N_4408,N_2120,N_1664);
nor U4409 (N_4409,N_1477,N_974);
nand U4410 (N_4410,N_1191,N_1928);
nor U4411 (N_4411,N_269,N_1473);
nand U4412 (N_4412,N_462,N_2045);
or U4413 (N_4413,N_314,N_206);
or U4414 (N_4414,N_1847,N_2174);
xor U4415 (N_4415,N_2483,N_1964);
xor U4416 (N_4416,N_741,N_36);
or U4417 (N_4417,N_1478,N_27);
nor U4418 (N_4418,N_1619,N_781);
or U4419 (N_4419,N_120,N_707);
or U4420 (N_4420,N_309,N_2217);
nor U4421 (N_4421,N_1248,N_1569);
and U4422 (N_4422,N_1117,N_2132);
and U4423 (N_4423,N_166,N_1810);
or U4424 (N_4424,N_1775,N_45);
and U4425 (N_4425,N_1294,N_106);
and U4426 (N_4426,N_199,N_2116);
nor U4427 (N_4427,N_2395,N_464);
nor U4428 (N_4428,N_1379,N_1150);
nand U4429 (N_4429,N_2058,N_2093);
xor U4430 (N_4430,N_307,N_854);
and U4431 (N_4431,N_1558,N_113);
xnor U4432 (N_4432,N_945,N_576);
or U4433 (N_4433,N_2381,N_1743);
nand U4434 (N_4434,N_236,N_1192);
xnor U4435 (N_4435,N_2088,N_2273);
and U4436 (N_4436,N_966,N_1791);
nand U4437 (N_4437,N_1124,N_2326);
xnor U4438 (N_4438,N_59,N_600);
nor U4439 (N_4439,N_2433,N_69);
xnor U4440 (N_4440,N_1172,N_972);
xor U4441 (N_4441,N_1353,N_538);
and U4442 (N_4442,N_2033,N_1985);
and U4443 (N_4443,N_2055,N_299);
nor U4444 (N_4444,N_694,N_1966);
nand U4445 (N_4445,N_1758,N_1710);
and U4446 (N_4446,N_1664,N_474);
and U4447 (N_4447,N_2196,N_406);
xor U4448 (N_4448,N_1556,N_1391);
or U4449 (N_4449,N_1597,N_173);
xor U4450 (N_4450,N_1807,N_602);
xor U4451 (N_4451,N_34,N_3);
or U4452 (N_4452,N_1393,N_183);
and U4453 (N_4453,N_364,N_536);
nand U4454 (N_4454,N_1202,N_292);
nor U4455 (N_4455,N_720,N_671);
and U4456 (N_4456,N_1931,N_2488);
nor U4457 (N_4457,N_2314,N_1247);
xor U4458 (N_4458,N_2022,N_398);
and U4459 (N_4459,N_305,N_1203);
nand U4460 (N_4460,N_710,N_2117);
nor U4461 (N_4461,N_1791,N_882);
nor U4462 (N_4462,N_2392,N_1143);
nand U4463 (N_4463,N_536,N_1003);
and U4464 (N_4464,N_1362,N_797);
and U4465 (N_4465,N_1716,N_1344);
xor U4466 (N_4466,N_620,N_2084);
and U4467 (N_4467,N_1628,N_2359);
or U4468 (N_4468,N_1416,N_1916);
and U4469 (N_4469,N_2130,N_1656);
and U4470 (N_4470,N_2125,N_646);
nor U4471 (N_4471,N_133,N_1910);
xnor U4472 (N_4472,N_2216,N_1579);
nor U4473 (N_4473,N_546,N_1725);
or U4474 (N_4474,N_1190,N_1161);
nand U4475 (N_4475,N_1574,N_634);
nor U4476 (N_4476,N_1104,N_179);
and U4477 (N_4477,N_64,N_2461);
and U4478 (N_4478,N_1345,N_683);
and U4479 (N_4479,N_2091,N_1120);
xnor U4480 (N_4480,N_2300,N_538);
and U4481 (N_4481,N_1155,N_2177);
nand U4482 (N_4482,N_1915,N_2411);
nor U4483 (N_4483,N_43,N_2316);
nand U4484 (N_4484,N_1772,N_2277);
nand U4485 (N_4485,N_2118,N_975);
or U4486 (N_4486,N_1099,N_2155);
nand U4487 (N_4487,N_656,N_1590);
nor U4488 (N_4488,N_1559,N_994);
xnor U4489 (N_4489,N_2071,N_1275);
and U4490 (N_4490,N_314,N_277);
nand U4491 (N_4491,N_166,N_1684);
nor U4492 (N_4492,N_1233,N_1468);
xor U4493 (N_4493,N_2445,N_164);
nand U4494 (N_4494,N_577,N_179);
and U4495 (N_4495,N_2245,N_459);
nor U4496 (N_4496,N_302,N_1191);
xor U4497 (N_4497,N_223,N_997);
or U4498 (N_4498,N_886,N_1357);
nand U4499 (N_4499,N_1679,N_1798);
nand U4500 (N_4500,N_1426,N_1744);
nor U4501 (N_4501,N_379,N_1698);
and U4502 (N_4502,N_1321,N_738);
nand U4503 (N_4503,N_1930,N_2110);
or U4504 (N_4504,N_677,N_753);
or U4505 (N_4505,N_690,N_1233);
xnor U4506 (N_4506,N_115,N_1242);
and U4507 (N_4507,N_166,N_802);
nor U4508 (N_4508,N_966,N_974);
nand U4509 (N_4509,N_1587,N_590);
nand U4510 (N_4510,N_2253,N_668);
and U4511 (N_4511,N_1137,N_2412);
or U4512 (N_4512,N_2222,N_323);
and U4513 (N_4513,N_678,N_1715);
nand U4514 (N_4514,N_338,N_506);
nor U4515 (N_4515,N_1876,N_980);
xnor U4516 (N_4516,N_1260,N_241);
or U4517 (N_4517,N_2132,N_2119);
nand U4518 (N_4518,N_60,N_1372);
and U4519 (N_4519,N_1476,N_1058);
nand U4520 (N_4520,N_1657,N_2476);
or U4521 (N_4521,N_729,N_2452);
or U4522 (N_4522,N_2408,N_1748);
xnor U4523 (N_4523,N_331,N_1548);
nor U4524 (N_4524,N_1819,N_2446);
or U4525 (N_4525,N_1469,N_1788);
nand U4526 (N_4526,N_1407,N_1533);
or U4527 (N_4527,N_286,N_1474);
and U4528 (N_4528,N_928,N_71);
or U4529 (N_4529,N_178,N_2251);
nand U4530 (N_4530,N_2378,N_2431);
nand U4531 (N_4531,N_397,N_48);
or U4532 (N_4532,N_401,N_1878);
nand U4533 (N_4533,N_273,N_1967);
xnor U4534 (N_4534,N_2462,N_358);
or U4535 (N_4535,N_2299,N_729);
nor U4536 (N_4536,N_1715,N_1622);
nand U4537 (N_4537,N_676,N_737);
nor U4538 (N_4538,N_1936,N_714);
nand U4539 (N_4539,N_778,N_2466);
xor U4540 (N_4540,N_1589,N_1160);
xor U4541 (N_4541,N_777,N_2122);
and U4542 (N_4542,N_1342,N_1469);
nand U4543 (N_4543,N_631,N_307);
nand U4544 (N_4544,N_2154,N_2045);
or U4545 (N_4545,N_1845,N_784);
and U4546 (N_4546,N_15,N_2166);
nand U4547 (N_4547,N_594,N_642);
nand U4548 (N_4548,N_1164,N_1836);
and U4549 (N_4549,N_2161,N_1839);
and U4550 (N_4550,N_1997,N_2361);
xor U4551 (N_4551,N_2363,N_544);
xnor U4552 (N_4552,N_1016,N_1564);
nand U4553 (N_4553,N_59,N_1858);
and U4554 (N_4554,N_377,N_795);
nor U4555 (N_4555,N_93,N_251);
xnor U4556 (N_4556,N_2490,N_1975);
or U4557 (N_4557,N_1171,N_73);
and U4558 (N_4558,N_708,N_2084);
and U4559 (N_4559,N_1011,N_182);
or U4560 (N_4560,N_1872,N_1477);
xnor U4561 (N_4561,N_2466,N_2114);
and U4562 (N_4562,N_426,N_1675);
nand U4563 (N_4563,N_723,N_125);
nor U4564 (N_4564,N_521,N_1516);
and U4565 (N_4565,N_259,N_1317);
xnor U4566 (N_4566,N_1132,N_448);
nor U4567 (N_4567,N_1930,N_1946);
or U4568 (N_4568,N_2436,N_1232);
or U4569 (N_4569,N_1790,N_128);
or U4570 (N_4570,N_1886,N_421);
and U4571 (N_4571,N_1851,N_1048);
nand U4572 (N_4572,N_604,N_938);
nor U4573 (N_4573,N_1336,N_2376);
nand U4574 (N_4574,N_889,N_1342);
xnor U4575 (N_4575,N_2014,N_1688);
nor U4576 (N_4576,N_1416,N_784);
or U4577 (N_4577,N_2289,N_503);
nand U4578 (N_4578,N_1358,N_1587);
nor U4579 (N_4579,N_1654,N_165);
xor U4580 (N_4580,N_2268,N_267);
nor U4581 (N_4581,N_1156,N_318);
xnor U4582 (N_4582,N_152,N_718);
or U4583 (N_4583,N_965,N_620);
nand U4584 (N_4584,N_1079,N_542);
and U4585 (N_4585,N_1780,N_982);
or U4586 (N_4586,N_434,N_2244);
and U4587 (N_4587,N_883,N_1288);
nor U4588 (N_4588,N_401,N_133);
nor U4589 (N_4589,N_1462,N_2039);
xnor U4590 (N_4590,N_768,N_708);
or U4591 (N_4591,N_50,N_731);
or U4592 (N_4592,N_456,N_2369);
and U4593 (N_4593,N_1084,N_239);
or U4594 (N_4594,N_1942,N_1395);
or U4595 (N_4595,N_1169,N_1595);
xor U4596 (N_4596,N_602,N_2023);
or U4597 (N_4597,N_183,N_781);
and U4598 (N_4598,N_1819,N_2137);
nand U4599 (N_4599,N_2475,N_813);
nor U4600 (N_4600,N_29,N_606);
nor U4601 (N_4601,N_321,N_2132);
xor U4602 (N_4602,N_1158,N_700);
or U4603 (N_4603,N_1772,N_2348);
or U4604 (N_4604,N_2072,N_1460);
or U4605 (N_4605,N_1124,N_1490);
xnor U4606 (N_4606,N_1280,N_1197);
and U4607 (N_4607,N_545,N_41);
xnor U4608 (N_4608,N_2204,N_1334);
nand U4609 (N_4609,N_306,N_2056);
nor U4610 (N_4610,N_173,N_529);
and U4611 (N_4611,N_1229,N_553);
nor U4612 (N_4612,N_1569,N_442);
xor U4613 (N_4613,N_1889,N_696);
or U4614 (N_4614,N_143,N_321);
nor U4615 (N_4615,N_2205,N_256);
nor U4616 (N_4616,N_1025,N_1326);
nor U4617 (N_4617,N_11,N_1646);
and U4618 (N_4618,N_299,N_761);
or U4619 (N_4619,N_2182,N_1344);
or U4620 (N_4620,N_2284,N_278);
nor U4621 (N_4621,N_1547,N_1937);
nor U4622 (N_4622,N_210,N_1946);
xor U4623 (N_4623,N_925,N_500);
or U4624 (N_4624,N_2203,N_1077);
or U4625 (N_4625,N_539,N_1555);
nand U4626 (N_4626,N_2240,N_398);
or U4627 (N_4627,N_2406,N_1291);
nor U4628 (N_4628,N_1512,N_1180);
or U4629 (N_4629,N_2351,N_1392);
nand U4630 (N_4630,N_1412,N_1509);
or U4631 (N_4631,N_7,N_2421);
nor U4632 (N_4632,N_1431,N_1382);
xor U4633 (N_4633,N_213,N_690);
nand U4634 (N_4634,N_286,N_2151);
and U4635 (N_4635,N_907,N_1463);
nand U4636 (N_4636,N_123,N_887);
and U4637 (N_4637,N_637,N_2084);
and U4638 (N_4638,N_1070,N_1769);
nand U4639 (N_4639,N_88,N_2412);
nand U4640 (N_4640,N_61,N_2144);
or U4641 (N_4641,N_1920,N_608);
and U4642 (N_4642,N_1551,N_267);
nand U4643 (N_4643,N_1696,N_1373);
nand U4644 (N_4644,N_618,N_2296);
xor U4645 (N_4645,N_1388,N_929);
and U4646 (N_4646,N_450,N_2419);
nor U4647 (N_4647,N_821,N_2457);
and U4648 (N_4648,N_822,N_1859);
nand U4649 (N_4649,N_961,N_2055);
nand U4650 (N_4650,N_191,N_1099);
and U4651 (N_4651,N_1772,N_1488);
nand U4652 (N_4652,N_870,N_2240);
xor U4653 (N_4653,N_900,N_275);
or U4654 (N_4654,N_148,N_2251);
or U4655 (N_4655,N_1803,N_337);
or U4656 (N_4656,N_2093,N_1406);
and U4657 (N_4657,N_906,N_823);
or U4658 (N_4658,N_2235,N_2391);
or U4659 (N_4659,N_1018,N_2076);
nand U4660 (N_4660,N_819,N_2297);
or U4661 (N_4661,N_196,N_545);
nor U4662 (N_4662,N_2060,N_2145);
or U4663 (N_4663,N_2231,N_1793);
xor U4664 (N_4664,N_1500,N_1131);
xor U4665 (N_4665,N_2163,N_2318);
nand U4666 (N_4666,N_873,N_672);
and U4667 (N_4667,N_1923,N_2323);
nor U4668 (N_4668,N_994,N_1860);
xor U4669 (N_4669,N_1724,N_494);
xnor U4670 (N_4670,N_2456,N_1016);
and U4671 (N_4671,N_2149,N_1151);
nor U4672 (N_4672,N_2122,N_16);
and U4673 (N_4673,N_1405,N_951);
xnor U4674 (N_4674,N_1365,N_1863);
or U4675 (N_4675,N_2222,N_2099);
or U4676 (N_4676,N_2206,N_2185);
xnor U4677 (N_4677,N_2348,N_1665);
and U4678 (N_4678,N_2178,N_2151);
nor U4679 (N_4679,N_870,N_2410);
or U4680 (N_4680,N_1417,N_1961);
xor U4681 (N_4681,N_955,N_2418);
or U4682 (N_4682,N_1301,N_2354);
nand U4683 (N_4683,N_564,N_883);
or U4684 (N_4684,N_393,N_1069);
and U4685 (N_4685,N_2022,N_1090);
and U4686 (N_4686,N_1281,N_284);
nand U4687 (N_4687,N_2497,N_2246);
nand U4688 (N_4688,N_432,N_484);
and U4689 (N_4689,N_1286,N_2099);
and U4690 (N_4690,N_1384,N_151);
nand U4691 (N_4691,N_1379,N_505);
or U4692 (N_4692,N_678,N_17);
or U4693 (N_4693,N_513,N_600);
or U4694 (N_4694,N_1258,N_171);
nor U4695 (N_4695,N_806,N_1270);
or U4696 (N_4696,N_1427,N_1897);
xnor U4697 (N_4697,N_1637,N_2121);
nor U4698 (N_4698,N_1354,N_830);
xor U4699 (N_4699,N_564,N_1269);
nand U4700 (N_4700,N_828,N_2354);
xnor U4701 (N_4701,N_2177,N_241);
and U4702 (N_4702,N_89,N_1985);
or U4703 (N_4703,N_1086,N_969);
and U4704 (N_4704,N_1268,N_794);
nand U4705 (N_4705,N_2412,N_1291);
nand U4706 (N_4706,N_2459,N_1930);
xnor U4707 (N_4707,N_1507,N_1346);
nor U4708 (N_4708,N_1921,N_581);
or U4709 (N_4709,N_1175,N_1713);
and U4710 (N_4710,N_612,N_1604);
xnor U4711 (N_4711,N_2265,N_971);
or U4712 (N_4712,N_2242,N_384);
or U4713 (N_4713,N_1765,N_1188);
xnor U4714 (N_4714,N_110,N_354);
nand U4715 (N_4715,N_1858,N_2272);
nor U4716 (N_4716,N_2176,N_1141);
and U4717 (N_4717,N_969,N_1038);
xnor U4718 (N_4718,N_456,N_1810);
nor U4719 (N_4719,N_1776,N_1193);
and U4720 (N_4720,N_173,N_456);
or U4721 (N_4721,N_255,N_1859);
nor U4722 (N_4722,N_1727,N_1429);
nor U4723 (N_4723,N_1606,N_1243);
and U4724 (N_4724,N_824,N_2382);
and U4725 (N_4725,N_1283,N_2070);
and U4726 (N_4726,N_338,N_194);
or U4727 (N_4727,N_2126,N_2331);
or U4728 (N_4728,N_1411,N_1553);
nor U4729 (N_4729,N_2320,N_1793);
xor U4730 (N_4730,N_315,N_195);
or U4731 (N_4731,N_1911,N_429);
xor U4732 (N_4732,N_2237,N_1111);
or U4733 (N_4733,N_1578,N_1503);
and U4734 (N_4734,N_144,N_882);
nor U4735 (N_4735,N_947,N_2072);
nor U4736 (N_4736,N_2048,N_2463);
or U4737 (N_4737,N_1452,N_54);
nor U4738 (N_4738,N_1624,N_1305);
and U4739 (N_4739,N_632,N_1742);
xor U4740 (N_4740,N_711,N_1438);
nor U4741 (N_4741,N_1730,N_1148);
nand U4742 (N_4742,N_399,N_2011);
or U4743 (N_4743,N_658,N_692);
and U4744 (N_4744,N_1536,N_1326);
and U4745 (N_4745,N_52,N_2068);
and U4746 (N_4746,N_335,N_1636);
or U4747 (N_4747,N_775,N_259);
xnor U4748 (N_4748,N_1132,N_1717);
nand U4749 (N_4749,N_118,N_2152);
xnor U4750 (N_4750,N_51,N_368);
and U4751 (N_4751,N_137,N_2188);
nor U4752 (N_4752,N_2120,N_2000);
xnor U4753 (N_4753,N_604,N_984);
nand U4754 (N_4754,N_2114,N_912);
nand U4755 (N_4755,N_746,N_731);
and U4756 (N_4756,N_787,N_1922);
or U4757 (N_4757,N_2272,N_454);
xor U4758 (N_4758,N_1016,N_1347);
or U4759 (N_4759,N_1911,N_2007);
nor U4760 (N_4760,N_1157,N_826);
or U4761 (N_4761,N_2189,N_2156);
and U4762 (N_4762,N_1446,N_1771);
xor U4763 (N_4763,N_209,N_750);
and U4764 (N_4764,N_1755,N_1356);
or U4765 (N_4765,N_488,N_392);
or U4766 (N_4766,N_276,N_1940);
xor U4767 (N_4767,N_315,N_1277);
and U4768 (N_4768,N_2264,N_952);
xor U4769 (N_4769,N_2247,N_887);
xor U4770 (N_4770,N_2224,N_1701);
or U4771 (N_4771,N_1230,N_1198);
xor U4772 (N_4772,N_308,N_1342);
and U4773 (N_4773,N_1797,N_1295);
xor U4774 (N_4774,N_851,N_1782);
nor U4775 (N_4775,N_1166,N_1872);
nand U4776 (N_4776,N_1635,N_2325);
or U4777 (N_4777,N_2365,N_1839);
and U4778 (N_4778,N_2200,N_1698);
nand U4779 (N_4779,N_826,N_2149);
xnor U4780 (N_4780,N_1270,N_1132);
or U4781 (N_4781,N_1158,N_1900);
xnor U4782 (N_4782,N_195,N_2212);
nor U4783 (N_4783,N_1192,N_388);
nor U4784 (N_4784,N_1955,N_602);
and U4785 (N_4785,N_1449,N_678);
and U4786 (N_4786,N_1696,N_1099);
nand U4787 (N_4787,N_2118,N_1536);
nor U4788 (N_4788,N_876,N_559);
nor U4789 (N_4789,N_1041,N_1097);
nand U4790 (N_4790,N_280,N_461);
or U4791 (N_4791,N_2489,N_2158);
and U4792 (N_4792,N_1887,N_1055);
nor U4793 (N_4793,N_1460,N_2292);
nand U4794 (N_4794,N_2027,N_2332);
or U4795 (N_4795,N_1843,N_71);
or U4796 (N_4796,N_319,N_102);
and U4797 (N_4797,N_544,N_792);
nor U4798 (N_4798,N_729,N_1631);
and U4799 (N_4799,N_2215,N_741);
xnor U4800 (N_4800,N_751,N_1371);
nand U4801 (N_4801,N_1700,N_2065);
and U4802 (N_4802,N_2398,N_1719);
and U4803 (N_4803,N_1820,N_2010);
nor U4804 (N_4804,N_1862,N_853);
nand U4805 (N_4805,N_538,N_236);
xnor U4806 (N_4806,N_149,N_1013);
nand U4807 (N_4807,N_265,N_824);
or U4808 (N_4808,N_740,N_1355);
or U4809 (N_4809,N_317,N_2301);
xor U4810 (N_4810,N_1773,N_1210);
xor U4811 (N_4811,N_1309,N_1483);
xor U4812 (N_4812,N_320,N_1334);
and U4813 (N_4813,N_2013,N_892);
xnor U4814 (N_4814,N_1450,N_1366);
or U4815 (N_4815,N_1049,N_230);
or U4816 (N_4816,N_1225,N_165);
and U4817 (N_4817,N_36,N_1695);
nor U4818 (N_4818,N_2105,N_783);
xor U4819 (N_4819,N_804,N_1970);
and U4820 (N_4820,N_1706,N_137);
xnor U4821 (N_4821,N_1656,N_1439);
or U4822 (N_4822,N_1719,N_777);
nand U4823 (N_4823,N_516,N_766);
nand U4824 (N_4824,N_545,N_1131);
nand U4825 (N_4825,N_1107,N_406);
or U4826 (N_4826,N_988,N_1603);
xor U4827 (N_4827,N_1836,N_508);
nor U4828 (N_4828,N_1187,N_2460);
or U4829 (N_4829,N_1378,N_774);
or U4830 (N_4830,N_352,N_171);
nor U4831 (N_4831,N_4,N_1999);
or U4832 (N_4832,N_2014,N_1735);
or U4833 (N_4833,N_1798,N_1973);
nand U4834 (N_4834,N_817,N_2343);
and U4835 (N_4835,N_1248,N_865);
and U4836 (N_4836,N_1739,N_40);
nor U4837 (N_4837,N_1230,N_1563);
and U4838 (N_4838,N_1740,N_2296);
nor U4839 (N_4839,N_1203,N_1264);
xor U4840 (N_4840,N_1604,N_1092);
xor U4841 (N_4841,N_1602,N_1542);
and U4842 (N_4842,N_913,N_1725);
xnor U4843 (N_4843,N_1573,N_2371);
or U4844 (N_4844,N_384,N_1854);
nand U4845 (N_4845,N_1564,N_1679);
and U4846 (N_4846,N_2028,N_493);
and U4847 (N_4847,N_2477,N_1182);
nand U4848 (N_4848,N_794,N_1257);
nand U4849 (N_4849,N_972,N_40);
and U4850 (N_4850,N_883,N_1633);
nand U4851 (N_4851,N_1764,N_1841);
nor U4852 (N_4852,N_1015,N_1319);
xor U4853 (N_4853,N_2475,N_1914);
or U4854 (N_4854,N_1318,N_2097);
xnor U4855 (N_4855,N_1237,N_2193);
or U4856 (N_4856,N_164,N_631);
nor U4857 (N_4857,N_548,N_2498);
or U4858 (N_4858,N_834,N_490);
xor U4859 (N_4859,N_2353,N_2369);
or U4860 (N_4860,N_2122,N_1136);
or U4861 (N_4861,N_766,N_2043);
xnor U4862 (N_4862,N_1631,N_1452);
nor U4863 (N_4863,N_2031,N_137);
xnor U4864 (N_4864,N_360,N_633);
nand U4865 (N_4865,N_744,N_945);
or U4866 (N_4866,N_1660,N_2283);
nand U4867 (N_4867,N_955,N_153);
nor U4868 (N_4868,N_402,N_1207);
and U4869 (N_4869,N_1932,N_198);
or U4870 (N_4870,N_314,N_2417);
or U4871 (N_4871,N_80,N_1384);
nor U4872 (N_4872,N_287,N_1314);
xor U4873 (N_4873,N_1342,N_832);
and U4874 (N_4874,N_2141,N_1209);
nand U4875 (N_4875,N_1665,N_2050);
or U4876 (N_4876,N_469,N_2332);
and U4877 (N_4877,N_1571,N_1319);
nand U4878 (N_4878,N_633,N_2169);
and U4879 (N_4879,N_1121,N_2355);
xnor U4880 (N_4880,N_2049,N_537);
xor U4881 (N_4881,N_919,N_2108);
xnor U4882 (N_4882,N_1880,N_539);
nor U4883 (N_4883,N_1613,N_1742);
and U4884 (N_4884,N_627,N_1141);
or U4885 (N_4885,N_440,N_1940);
nor U4886 (N_4886,N_2167,N_621);
xor U4887 (N_4887,N_576,N_1902);
xnor U4888 (N_4888,N_2321,N_1262);
and U4889 (N_4889,N_2277,N_220);
nor U4890 (N_4890,N_1050,N_2036);
and U4891 (N_4891,N_303,N_565);
xnor U4892 (N_4892,N_890,N_982);
xnor U4893 (N_4893,N_1520,N_2013);
or U4894 (N_4894,N_2457,N_49);
nand U4895 (N_4895,N_1567,N_169);
or U4896 (N_4896,N_1591,N_1356);
nor U4897 (N_4897,N_2099,N_2318);
and U4898 (N_4898,N_1365,N_2056);
nand U4899 (N_4899,N_1900,N_2068);
nor U4900 (N_4900,N_2453,N_974);
nor U4901 (N_4901,N_2316,N_1559);
nor U4902 (N_4902,N_204,N_2034);
nand U4903 (N_4903,N_2132,N_633);
nor U4904 (N_4904,N_2482,N_2045);
xnor U4905 (N_4905,N_2155,N_2392);
nor U4906 (N_4906,N_46,N_1910);
xnor U4907 (N_4907,N_743,N_803);
nor U4908 (N_4908,N_374,N_801);
xnor U4909 (N_4909,N_1772,N_328);
nand U4910 (N_4910,N_734,N_1664);
and U4911 (N_4911,N_1427,N_1582);
xnor U4912 (N_4912,N_2041,N_307);
or U4913 (N_4913,N_2149,N_921);
nand U4914 (N_4914,N_1463,N_1352);
nand U4915 (N_4915,N_771,N_2003);
nand U4916 (N_4916,N_1774,N_2188);
xnor U4917 (N_4917,N_1914,N_1964);
xor U4918 (N_4918,N_1055,N_546);
nand U4919 (N_4919,N_130,N_320);
nand U4920 (N_4920,N_1351,N_1626);
xnor U4921 (N_4921,N_1801,N_907);
xnor U4922 (N_4922,N_626,N_2217);
and U4923 (N_4923,N_858,N_2278);
or U4924 (N_4924,N_398,N_1002);
nor U4925 (N_4925,N_2217,N_136);
and U4926 (N_4926,N_1005,N_848);
nor U4927 (N_4927,N_256,N_1710);
xor U4928 (N_4928,N_1966,N_101);
xor U4929 (N_4929,N_475,N_2178);
nor U4930 (N_4930,N_1030,N_5);
and U4931 (N_4931,N_1836,N_428);
nor U4932 (N_4932,N_879,N_2283);
xnor U4933 (N_4933,N_1791,N_1269);
nor U4934 (N_4934,N_1805,N_1271);
or U4935 (N_4935,N_1480,N_695);
or U4936 (N_4936,N_2157,N_866);
or U4937 (N_4937,N_2370,N_1532);
nor U4938 (N_4938,N_1612,N_2348);
and U4939 (N_4939,N_516,N_736);
xor U4940 (N_4940,N_2451,N_1024);
and U4941 (N_4941,N_174,N_808);
xnor U4942 (N_4942,N_1385,N_2064);
xnor U4943 (N_4943,N_1873,N_2386);
or U4944 (N_4944,N_1397,N_1468);
or U4945 (N_4945,N_2226,N_2285);
or U4946 (N_4946,N_2400,N_1729);
nor U4947 (N_4947,N_275,N_601);
xor U4948 (N_4948,N_2396,N_356);
xnor U4949 (N_4949,N_295,N_1195);
nand U4950 (N_4950,N_2282,N_2461);
nor U4951 (N_4951,N_1306,N_599);
and U4952 (N_4952,N_360,N_68);
xnor U4953 (N_4953,N_2069,N_2472);
nor U4954 (N_4954,N_2360,N_747);
and U4955 (N_4955,N_1669,N_1330);
xnor U4956 (N_4956,N_1826,N_1460);
and U4957 (N_4957,N_2457,N_2478);
xnor U4958 (N_4958,N_679,N_1660);
or U4959 (N_4959,N_2172,N_2341);
nand U4960 (N_4960,N_393,N_291);
nand U4961 (N_4961,N_1605,N_1161);
xnor U4962 (N_4962,N_13,N_830);
and U4963 (N_4963,N_331,N_119);
and U4964 (N_4964,N_649,N_2396);
or U4965 (N_4965,N_338,N_1619);
xor U4966 (N_4966,N_1276,N_280);
nor U4967 (N_4967,N_1397,N_86);
nor U4968 (N_4968,N_2487,N_2219);
nand U4969 (N_4969,N_182,N_2417);
or U4970 (N_4970,N_43,N_901);
nor U4971 (N_4971,N_609,N_681);
nand U4972 (N_4972,N_2331,N_16);
nand U4973 (N_4973,N_419,N_865);
nand U4974 (N_4974,N_1588,N_1991);
and U4975 (N_4975,N_1007,N_826);
and U4976 (N_4976,N_1047,N_1698);
nor U4977 (N_4977,N_305,N_2472);
xnor U4978 (N_4978,N_1937,N_1534);
xnor U4979 (N_4979,N_2182,N_666);
xnor U4980 (N_4980,N_2128,N_1574);
or U4981 (N_4981,N_1587,N_278);
nor U4982 (N_4982,N_1604,N_1602);
xor U4983 (N_4983,N_2101,N_283);
nand U4984 (N_4984,N_1818,N_1538);
or U4985 (N_4985,N_2050,N_1729);
or U4986 (N_4986,N_915,N_1793);
nand U4987 (N_4987,N_1486,N_127);
and U4988 (N_4988,N_1761,N_1290);
nor U4989 (N_4989,N_1640,N_1175);
and U4990 (N_4990,N_1505,N_2002);
nor U4991 (N_4991,N_2067,N_2269);
and U4992 (N_4992,N_1341,N_1196);
nand U4993 (N_4993,N_1508,N_1038);
and U4994 (N_4994,N_319,N_57);
xor U4995 (N_4995,N_744,N_1304);
nand U4996 (N_4996,N_186,N_1712);
xnor U4997 (N_4997,N_2170,N_1155);
and U4998 (N_4998,N_2346,N_146);
nand U4999 (N_4999,N_1372,N_2269);
or U5000 (N_5000,N_3476,N_2825);
and U5001 (N_5001,N_4328,N_2822);
xor U5002 (N_5002,N_4016,N_4914);
and U5003 (N_5003,N_3864,N_4055);
xor U5004 (N_5004,N_3865,N_4299);
and U5005 (N_5005,N_2760,N_4641);
or U5006 (N_5006,N_3946,N_3034);
and U5007 (N_5007,N_2886,N_2968);
nand U5008 (N_5008,N_3736,N_4755);
and U5009 (N_5009,N_2965,N_2980);
xor U5010 (N_5010,N_4876,N_4414);
xor U5011 (N_5011,N_4428,N_4570);
or U5012 (N_5012,N_3772,N_4271);
nand U5013 (N_5013,N_4024,N_4788);
xnor U5014 (N_5014,N_4488,N_4495);
xor U5015 (N_5015,N_3113,N_4880);
nand U5016 (N_5016,N_4511,N_4619);
or U5017 (N_5017,N_2568,N_2748);
nor U5018 (N_5018,N_4600,N_3211);
nor U5019 (N_5019,N_4628,N_4468);
xor U5020 (N_5020,N_3453,N_3685);
xor U5021 (N_5021,N_3284,N_4996);
or U5022 (N_5022,N_2949,N_4941);
or U5023 (N_5023,N_3237,N_3831);
or U5024 (N_5024,N_3123,N_3018);
or U5025 (N_5025,N_4999,N_3812);
xnor U5026 (N_5026,N_4070,N_2946);
and U5027 (N_5027,N_4168,N_4404);
nand U5028 (N_5028,N_4951,N_3760);
and U5029 (N_5029,N_4122,N_2974);
or U5030 (N_5030,N_4547,N_4329);
or U5031 (N_5031,N_4860,N_4543);
nand U5032 (N_5032,N_3862,N_4808);
nor U5033 (N_5033,N_4871,N_4903);
nand U5034 (N_5034,N_4804,N_3385);
nand U5035 (N_5035,N_4593,N_2837);
nand U5036 (N_5036,N_3935,N_3548);
nand U5037 (N_5037,N_3912,N_3182);
or U5038 (N_5038,N_2923,N_4051);
nand U5039 (N_5039,N_3855,N_4998);
or U5040 (N_5040,N_3972,N_3206);
xor U5041 (N_5041,N_3923,N_4451);
xor U5042 (N_5042,N_3636,N_4418);
xnor U5043 (N_5043,N_2653,N_4062);
or U5044 (N_5044,N_3360,N_2792);
nor U5045 (N_5045,N_3531,N_4481);
xnor U5046 (N_5046,N_3981,N_3014);
nand U5047 (N_5047,N_3857,N_4585);
xnor U5048 (N_5048,N_3756,N_2868);
and U5049 (N_5049,N_2830,N_4144);
xnor U5050 (N_5050,N_4370,N_4194);
and U5051 (N_5051,N_4198,N_4268);
and U5052 (N_5052,N_3042,N_3767);
nand U5053 (N_5053,N_4534,N_2671);
or U5054 (N_5054,N_3418,N_3401);
nand U5055 (N_5055,N_4360,N_2800);
nand U5056 (N_5056,N_4665,N_4560);
xnor U5057 (N_5057,N_4548,N_3980);
nand U5058 (N_5058,N_4963,N_4792);
nand U5059 (N_5059,N_3136,N_2855);
nand U5060 (N_5060,N_2715,N_3882);
xnor U5061 (N_5061,N_3201,N_3277);
nor U5062 (N_5062,N_3352,N_3754);
and U5063 (N_5063,N_3390,N_4470);
xnor U5064 (N_5064,N_4234,N_3996);
and U5065 (N_5065,N_3902,N_3883);
and U5066 (N_5066,N_4777,N_3260);
nand U5067 (N_5067,N_3431,N_3116);
or U5068 (N_5068,N_3101,N_3905);
or U5069 (N_5069,N_3396,N_4659);
and U5070 (N_5070,N_3122,N_4475);
and U5071 (N_5071,N_2544,N_4503);
or U5072 (N_5072,N_3255,N_3643);
nand U5073 (N_5073,N_4724,N_4126);
and U5074 (N_5074,N_4710,N_2744);
xor U5075 (N_5075,N_3055,N_3843);
or U5076 (N_5076,N_4306,N_2700);
xor U5077 (N_5077,N_3199,N_4806);
and U5078 (N_5078,N_2746,N_4293);
nand U5079 (N_5079,N_4921,N_4900);
or U5080 (N_5080,N_4345,N_2719);
and U5081 (N_5081,N_4629,N_2766);
xor U5082 (N_5082,N_3022,N_4893);
and U5083 (N_5083,N_3547,N_2801);
nand U5084 (N_5084,N_3373,N_3381);
nor U5085 (N_5085,N_4915,N_3465);
and U5086 (N_5086,N_3387,N_4330);
xor U5087 (N_5087,N_3421,N_4945);
and U5088 (N_5088,N_2948,N_3545);
nand U5089 (N_5089,N_2687,N_3698);
or U5090 (N_5090,N_2935,N_4797);
or U5091 (N_5091,N_3577,N_3721);
or U5092 (N_5092,N_2768,N_2915);
or U5093 (N_5093,N_3499,N_3152);
xnor U5094 (N_5094,N_2682,N_4142);
or U5095 (N_5095,N_3927,N_4182);
xor U5096 (N_5096,N_4979,N_3572);
or U5097 (N_5097,N_4850,N_2651);
and U5098 (N_5098,N_2625,N_3750);
and U5099 (N_5099,N_3737,N_2922);
xnor U5100 (N_5100,N_3100,N_4054);
nor U5101 (N_5101,N_2545,N_2689);
nor U5102 (N_5102,N_3319,N_4048);
and U5103 (N_5103,N_3312,N_4013);
nor U5104 (N_5104,N_3674,N_4852);
xnor U5105 (N_5105,N_2897,N_3522);
xor U5106 (N_5106,N_4913,N_2758);
nand U5107 (N_5107,N_3082,N_3880);
nor U5108 (N_5108,N_4376,N_4721);
and U5109 (N_5109,N_2884,N_2628);
xor U5110 (N_5110,N_2989,N_3976);
nor U5111 (N_5111,N_2503,N_4321);
xnor U5112 (N_5112,N_3099,N_2951);
nand U5113 (N_5113,N_2741,N_3484);
nor U5114 (N_5114,N_4416,N_3823);
nor U5115 (N_5115,N_2600,N_3096);
or U5116 (N_5116,N_4137,N_4214);
or U5117 (N_5117,N_2961,N_3509);
or U5118 (N_5118,N_3542,N_2918);
or U5119 (N_5119,N_4978,N_3949);
and U5120 (N_5120,N_4249,N_4188);
xnor U5121 (N_5121,N_2505,N_4577);
or U5122 (N_5122,N_3305,N_3748);
xor U5123 (N_5123,N_3094,N_4744);
and U5124 (N_5124,N_3384,N_2848);
or U5125 (N_5125,N_4036,N_4459);
nor U5126 (N_5126,N_4356,N_4892);
nand U5127 (N_5127,N_2888,N_2597);
and U5128 (N_5128,N_3322,N_4292);
nor U5129 (N_5129,N_2854,N_3723);
and U5130 (N_5130,N_3826,N_3303);
xnor U5131 (N_5131,N_2693,N_2970);
nor U5132 (N_5132,N_3253,N_2941);
nand U5133 (N_5133,N_4564,N_3730);
nor U5134 (N_5134,N_2732,N_4566);
nor U5135 (N_5135,N_2815,N_2634);
and U5136 (N_5136,N_3372,N_4680);
nor U5137 (N_5137,N_2838,N_4441);
xor U5138 (N_5138,N_3064,N_4103);
nand U5139 (N_5139,N_4639,N_2718);
xnor U5140 (N_5140,N_4906,N_3406);
nor U5141 (N_5141,N_2958,N_3498);
xor U5142 (N_5142,N_3874,N_4601);
xnor U5143 (N_5143,N_3435,N_3899);
and U5144 (N_5144,N_4264,N_4474);
nor U5145 (N_5145,N_4857,N_4709);
nor U5146 (N_5146,N_3759,N_2692);
nor U5147 (N_5147,N_2893,N_2878);
xnor U5148 (N_5148,N_3818,N_4507);
nor U5149 (N_5149,N_4056,N_3457);
or U5150 (N_5150,N_3516,N_4023);
nor U5151 (N_5151,N_2602,N_3671);
xor U5152 (N_5152,N_2564,N_2519);
or U5153 (N_5153,N_4040,N_3445);
nor U5154 (N_5154,N_4325,N_3139);
nor U5155 (N_5155,N_4358,N_4510);
nand U5156 (N_5156,N_2812,N_4853);
or U5157 (N_5157,N_2660,N_3588);
or U5158 (N_5158,N_2799,N_3463);
xor U5159 (N_5159,N_2985,N_2947);
and U5160 (N_5160,N_2779,N_3174);
nor U5161 (N_5161,N_3187,N_4782);
nand U5162 (N_5162,N_4487,N_3991);
or U5163 (N_5163,N_2934,N_3359);
or U5164 (N_5164,N_3716,N_4196);
and U5165 (N_5165,N_4947,N_3106);
nand U5166 (N_5166,N_3087,N_3472);
nand U5167 (N_5167,N_2930,N_2726);
or U5168 (N_5168,N_2806,N_3554);
and U5169 (N_5169,N_4695,N_4009);
xor U5170 (N_5170,N_4938,N_4750);
xnor U5171 (N_5171,N_3567,N_3241);
xor U5172 (N_5172,N_2510,N_2684);
or U5173 (N_5173,N_3274,N_4020);
xnor U5174 (N_5174,N_3138,N_2705);
xor U5175 (N_5175,N_4789,N_3568);
or U5176 (N_5176,N_2709,N_3778);
or U5177 (N_5177,N_4387,N_2533);
nor U5178 (N_5178,N_2680,N_4435);
nor U5179 (N_5179,N_4827,N_3316);
nor U5180 (N_5180,N_3180,N_3937);
and U5181 (N_5181,N_3611,N_4883);
xnor U5182 (N_5182,N_3849,N_2767);
and U5183 (N_5183,N_2857,N_4956);
nand U5184 (N_5184,N_3487,N_4855);
or U5185 (N_5185,N_4377,N_4044);
or U5186 (N_5186,N_4663,N_2944);
nand U5187 (N_5187,N_4170,N_4443);
nand U5188 (N_5188,N_4650,N_3782);
nand U5189 (N_5189,N_2502,N_3466);
and U5190 (N_5190,N_4412,N_3659);
or U5191 (N_5191,N_3986,N_4865);
or U5192 (N_5192,N_3550,N_4727);
and U5193 (N_5193,N_3813,N_3291);
nand U5194 (N_5194,N_3668,N_4616);
nor U5195 (N_5195,N_3622,N_4497);
nand U5196 (N_5196,N_2557,N_3785);
or U5197 (N_5197,N_4201,N_3173);
and U5198 (N_5198,N_4357,N_4537);
nand U5199 (N_5199,N_2647,N_3944);
nor U5200 (N_5200,N_3814,N_3332);
or U5201 (N_5201,N_4074,N_4960);
xor U5202 (N_5202,N_2525,N_3389);
xor U5203 (N_5203,N_2882,N_4241);
and U5204 (N_5204,N_4192,N_4694);
nand U5205 (N_5205,N_4713,N_3467);
and U5206 (N_5206,N_2515,N_3692);
nand U5207 (N_5207,N_2637,N_4397);
xor U5208 (N_5208,N_2865,N_2781);
nand U5209 (N_5209,N_3158,N_4807);
xor U5210 (N_5210,N_3596,N_3225);
xor U5211 (N_5211,N_3459,N_3348);
nor U5212 (N_5212,N_4714,N_4720);
nand U5213 (N_5213,N_3115,N_3337);
xor U5214 (N_5214,N_4994,N_3829);
and U5215 (N_5215,N_2819,N_3661);
and U5216 (N_5216,N_3680,N_4244);
and U5217 (N_5217,N_3176,N_2743);
xnor U5218 (N_5218,N_4820,N_3534);
or U5219 (N_5219,N_2939,N_4542);
nand U5220 (N_5220,N_3085,N_4532);
nand U5221 (N_5221,N_4668,N_4526);
or U5222 (N_5222,N_2887,N_2959);
nor U5223 (N_5223,N_4688,N_4590);
and U5224 (N_5224,N_4562,N_3266);
nor U5225 (N_5225,N_3217,N_3514);
nor U5226 (N_5226,N_3575,N_4780);
nor U5227 (N_5227,N_4551,N_3504);
nand U5228 (N_5228,N_4219,N_4627);
xnor U5229 (N_5229,N_2501,N_3931);
nand U5230 (N_5230,N_3335,N_4167);
and U5231 (N_5231,N_2728,N_3691);
nand U5232 (N_5232,N_4540,N_3677);
or U5233 (N_5233,N_4402,N_4283);
nand U5234 (N_5234,N_3458,N_2754);
and U5235 (N_5235,N_4734,N_3704);
nor U5236 (N_5236,N_3121,N_2713);
or U5237 (N_5237,N_4227,N_3062);
or U5238 (N_5238,N_4613,N_3833);
nand U5239 (N_5239,N_4810,N_4809);
nor U5240 (N_5240,N_3179,N_4552);
xnor U5241 (N_5241,N_4770,N_2658);
or U5242 (N_5242,N_2573,N_3289);
nand U5243 (N_5243,N_2723,N_2864);
and U5244 (N_5244,N_3285,N_3197);
nor U5245 (N_5245,N_4834,N_3888);
nor U5246 (N_5246,N_4350,N_4116);
and U5247 (N_5247,N_4823,N_4848);
or U5248 (N_5248,N_3369,N_4480);
nand U5249 (N_5249,N_4812,N_4513);
xor U5250 (N_5250,N_4598,N_3979);
and U5251 (N_5251,N_4197,N_3362);
or U5252 (N_5252,N_3758,N_4027);
and U5253 (N_5253,N_4046,N_4189);
or U5254 (N_5254,N_2504,N_3343);
or U5255 (N_5255,N_3656,N_2563);
and U5256 (N_5256,N_4677,N_2701);
and U5257 (N_5257,N_3092,N_3330);
and U5258 (N_5258,N_3552,N_3793);
or U5259 (N_5259,N_4015,N_3393);
nand U5260 (N_5260,N_2691,N_4611);
nand U5261 (N_5261,N_2546,N_4242);
or U5262 (N_5262,N_4922,N_4839);
nor U5263 (N_5263,N_2642,N_3690);
or U5264 (N_5264,N_2813,N_2810);
xnor U5265 (N_5265,N_3137,N_3212);
nor U5266 (N_5266,N_3189,N_3500);
xnor U5267 (N_5267,N_3746,N_4614);
nand U5268 (N_5268,N_2761,N_4444);
and U5269 (N_5269,N_4583,N_3461);
nor U5270 (N_5270,N_4644,N_4530);
nand U5271 (N_5271,N_3129,N_3612);
nand U5272 (N_5272,N_3973,N_3825);
xnor U5273 (N_5273,N_4692,N_2873);
nor U5274 (N_5274,N_3910,N_4401);
or U5275 (N_5275,N_4636,N_3642);
nand U5276 (N_5276,N_2871,N_3664);
nor U5277 (N_5277,N_4842,N_3008);
nand U5278 (N_5278,N_2727,N_3625);
or U5279 (N_5279,N_4516,N_3755);
and U5280 (N_5280,N_2526,N_4712);
and U5281 (N_5281,N_4791,N_3815);
nand U5282 (N_5282,N_4943,N_3998);
or U5283 (N_5283,N_3598,N_3836);
or U5284 (N_5284,N_4104,N_4708);
nor U5285 (N_5285,N_3037,N_4178);
or U5286 (N_5286,N_3341,N_3365);
xnor U5287 (N_5287,N_3492,N_4952);
or U5288 (N_5288,N_4990,N_4388);
and U5289 (N_5289,N_4722,N_3148);
nand U5290 (N_5290,N_3870,N_2737);
or U5291 (N_5291,N_3164,N_3320);
or U5292 (N_5292,N_2553,N_3741);
nor U5293 (N_5293,N_3151,N_2736);
and U5294 (N_5294,N_2818,N_4146);
nand U5295 (N_5295,N_2548,N_4685);
nand U5296 (N_5296,N_4141,N_2665);
nor U5297 (N_5297,N_2704,N_2789);
or U5298 (N_5298,N_3735,N_2956);
nor U5299 (N_5299,N_3270,N_2747);
and U5300 (N_5300,N_3951,N_2824);
xor U5301 (N_5301,N_4608,N_3503);
and U5302 (N_5302,N_3809,N_2678);
nor U5303 (N_5303,N_3493,N_4424);
or U5304 (N_5304,N_3226,N_3419);
nor U5305 (N_5305,N_4520,N_4371);
and U5306 (N_5306,N_3326,N_3455);
and U5307 (N_5307,N_3407,N_4037);
and U5308 (N_5308,N_3056,N_3799);
or U5309 (N_5309,N_3725,N_3228);
xor U5310 (N_5310,N_2994,N_4676);
nor U5311 (N_5311,N_3501,N_2880);
nor U5312 (N_5312,N_2931,N_4875);
nor U5313 (N_5313,N_2925,N_3904);
and U5314 (N_5314,N_3454,N_4819);
and U5315 (N_5315,N_4798,N_4961);
and U5316 (N_5316,N_3159,N_3940);
or U5317 (N_5317,N_4786,N_3714);
nand U5318 (N_5318,N_2604,N_4429);
xor U5319 (N_5319,N_4908,N_3846);
nor U5320 (N_5320,N_4517,N_3962);
nand U5321 (N_5321,N_3700,N_4896);
xnor U5322 (N_5322,N_3302,N_3281);
nor U5323 (N_5323,N_3824,N_2753);
and U5324 (N_5324,N_4224,N_2850);
nand U5325 (N_5325,N_4320,N_4014);
xor U5326 (N_5326,N_2797,N_4212);
and U5327 (N_5327,N_4684,N_2697);
and U5328 (N_5328,N_3112,N_3631);
or U5329 (N_5329,N_2927,N_2567);
nand U5330 (N_5330,N_4413,N_4136);
nor U5331 (N_5331,N_4012,N_2677);
or U5332 (N_5332,N_2733,N_2518);
nand U5333 (N_5333,N_3426,N_4887);
nand U5334 (N_5334,N_4851,N_3248);
nand U5335 (N_5335,N_3520,N_4302);
nand U5336 (N_5336,N_4891,N_3403);
xnor U5337 (N_5337,N_3834,N_3822);
and U5338 (N_5338,N_3306,N_3386);
or U5339 (N_5339,N_3188,N_3283);
or U5340 (N_5340,N_3796,N_3294);
xor U5341 (N_5341,N_4061,N_4717);
and U5342 (N_5342,N_4149,N_4374);
nor U5343 (N_5343,N_3525,N_4831);
nand U5344 (N_5344,N_3967,N_4634);
nand U5345 (N_5345,N_4442,N_4001);
nand U5346 (N_5346,N_2769,N_2626);
and U5347 (N_5347,N_3804,N_3939);
or U5348 (N_5348,N_2648,N_3328);
or U5349 (N_5349,N_4822,N_2993);
or U5350 (N_5350,N_4399,N_4307);
or U5351 (N_5351,N_4483,N_4460);
or U5352 (N_5352,N_4607,N_2863);
or U5353 (N_5353,N_4729,N_3429);
nor U5354 (N_5354,N_4512,N_3909);
nand U5355 (N_5355,N_3926,N_2776);
nand U5356 (N_5356,N_4623,N_3959);
and U5357 (N_5357,N_3911,N_4467);
nor U5358 (N_5358,N_3676,N_4899);
nor U5359 (N_5359,N_3314,N_3470);
and U5360 (N_5360,N_4210,N_3339);
and U5361 (N_5361,N_2621,N_4052);
nor U5362 (N_5362,N_3021,N_2829);
and U5363 (N_5363,N_3143,N_3924);
or U5364 (N_5364,N_4995,N_4417);
or U5365 (N_5365,N_3524,N_3762);
and U5366 (N_5366,N_4369,N_4058);
and U5367 (N_5367,N_4987,N_4165);
xor U5368 (N_5368,N_3325,N_3028);
nand U5369 (N_5369,N_2845,N_2729);
nand U5370 (N_5370,N_2963,N_4965);
xnor U5371 (N_5371,N_3618,N_4326);
nor U5372 (N_5372,N_4725,N_3006);
nand U5373 (N_5373,N_3821,N_3383);
xor U5374 (N_5374,N_3859,N_3259);
or U5375 (N_5375,N_3208,N_2631);
or U5376 (N_5376,N_2770,N_3066);
xnor U5377 (N_5377,N_4675,N_4110);
nand U5378 (N_5378,N_3102,N_4486);
and U5379 (N_5379,N_4410,N_3440);
or U5380 (N_5380,N_3263,N_3791);
and U5381 (N_5381,N_4762,N_2773);
xnor U5382 (N_5382,N_4859,N_4661);
nand U5383 (N_5383,N_3518,N_2530);
nor U5384 (N_5384,N_2656,N_2655);
nor U5385 (N_5385,N_2904,N_2675);
and U5386 (N_5386,N_4038,N_4231);
and U5387 (N_5387,N_2992,N_4132);
nand U5388 (N_5388,N_4186,N_3915);
and U5389 (N_5389,N_2551,N_4733);
xor U5390 (N_5390,N_2839,N_4929);
nor U5391 (N_5391,N_4728,N_4449);
nor U5392 (N_5392,N_3350,N_4069);
nand U5393 (N_5393,N_3728,N_4396);
nor U5394 (N_5394,N_3715,N_3293);
xor U5395 (N_5395,N_4790,N_3132);
or U5396 (N_5396,N_2669,N_3246);
nand U5397 (N_5397,N_3264,N_4544);
nand U5398 (N_5398,N_2540,N_4643);
xor U5399 (N_5399,N_4075,N_3433);
and U5400 (N_5400,N_2535,N_4801);
and U5401 (N_5401,N_3287,N_3884);
xor U5402 (N_5402,N_2952,N_4313);
xnor U5403 (N_5403,N_4150,N_2981);
xor U5404 (N_5404,N_3209,N_3649);
nand U5405 (N_5405,N_3792,N_4584);
and U5406 (N_5406,N_4211,N_3726);
or U5407 (N_5407,N_4354,N_4653);
nor U5408 (N_5408,N_2929,N_4436);
and U5409 (N_5409,N_4868,N_3269);
and U5410 (N_5410,N_4456,N_4026);
nand U5411 (N_5411,N_2513,N_2617);
nor U5412 (N_5412,N_3779,N_3686);
xnor U5413 (N_5413,N_4766,N_3017);
nand U5414 (N_5414,N_4079,N_3523);
nor U5415 (N_5415,N_4019,N_2907);
and U5416 (N_5416,N_4458,N_3342);
nor U5417 (N_5417,N_2875,N_3219);
or U5418 (N_5418,N_3171,N_3934);
xor U5419 (N_5419,N_3626,N_4886);
or U5420 (N_5420,N_4706,N_4563);
nor U5421 (N_5421,N_2596,N_2780);
and U5422 (N_5422,N_4230,N_4083);
nor U5423 (N_5423,N_3950,N_3125);
xnor U5424 (N_5424,N_4390,N_4322);
and U5425 (N_5425,N_3679,N_2764);
nor U5426 (N_5426,N_4002,N_3640);
and U5427 (N_5427,N_2580,N_3414);
xor U5428 (N_5428,N_3149,N_3346);
nand U5429 (N_5429,N_3057,N_4776);
and U5430 (N_5430,N_3364,N_3054);
or U5431 (N_5431,N_4151,N_4287);
xor U5432 (N_5432,N_3634,N_3007);
xnor U5433 (N_5433,N_4498,N_4305);
or U5434 (N_5434,N_4976,N_4679);
nor U5435 (N_5435,N_4939,N_3560);
nand U5436 (N_5436,N_4279,N_2514);
nor U5437 (N_5437,N_4318,N_3135);
and U5438 (N_5438,N_3072,N_3184);
and U5439 (N_5439,N_3192,N_3168);
and U5440 (N_5440,N_3616,N_2919);
nor U5441 (N_5441,N_4647,N_3105);
xnor U5442 (N_5442,N_4101,N_4919);
or U5443 (N_5443,N_2576,N_2823);
xor U5444 (N_5444,N_3628,N_2673);
nor U5445 (N_5445,N_2716,N_3720);
xor U5446 (N_5446,N_3408,N_2650);
nand U5447 (N_5447,N_3084,N_4814);
xor U5448 (N_5448,N_3621,N_3783);
nor U5449 (N_5449,N_3078,N_3696);
nor U5450 (N_5450,N_3239,N_2885);
or U5451 (N_5451,N_3947,N_2969);
or U5452 (N_5452,N_4164,N_3593);
nor U5453 (N_5453,N_4113,N_4588);
and U5454 (N_5454,N_2740,N_3710);
and U5455 (N_5455,N_4252,N_4558);
and U5456 (N_5456,N_4100,N_3852);
xnor U5457 (N_5457,N_4832,N_4159);
nor U5458 (N_5458,N_3941,N_2645);
or U5459 (N_5459,N_3437,N_3620);
xnor U5460 (N_5460,N_2905,N_3722);
and U5461 (N_5461,N_4378,N_4139);
nand U5462 (N_5462,N_3035,N_2938);
or U5463 (N_5463,N_4373,N_3965);
nor U5464 (N_5464,N_3029,N_2566);
xor U5465 (N_5465,N_3839,N_3086);
nor U5466 (N_5466,N_4796,N_3617);
or U5467 (N_5467,N_4902,N_4191);
nand U5468 (N_5468,N_3624,N_2734);
nor U5469 (N_5469,N_3126,N_3060);
nor U5470 (N_5470,N_2924,N_4225);
or U5471 (N_5471,N_2835,N_3541);
and U5472 (N_5472,N_2572,N_3356);
nor U5473 (N_5473,N_3321,N_4403);
and U5474 (N_5474,N_3860,N_3955);
nand U5475 (N_5475,N_4254,N_3740);
or U5476 (N_5476,N_4572,N_3845);
and U5477 (N_5477,N_3181,N_4437);
and U5478 (N_5478,N_3673,N_2509);
xor U5479 (N_5479,N_2846,N_4716);
xor U5480 (N_5480,N_3891,N_2703);
and U5481 (N_5481,N_4195,N_3262);
nor U5482 (N_5482,N_3204,N_4145);
nand U5483 (N_5483,N_3930,N_4821);
nor U5484 (N_5484,N_3288,N_4962);
xnor U5485 (N_5485,N_3872,N_2570);
nor U5486 (N_5486,N_4581,N_4660);
xnor U5487 (N_5487,N_4783,N_3890);
xor U5488 (N_5488,N_2569,N_4747);
or U5489 (N_5489,N_2794,N_3297);
nor U5490 (N_5490,N_2785,N_4285);
nand U5491 (N_5491,N_4257,N_3816);
nor U5492 (N_5492,N_4208,N_3918);
nand U5493 (N_5493,N_2817,N_3919);
nor U5494 (N_5494,N_4731,N_4624);
or U5495 (N_5495,N_3300,N_3573);
nor U5496 (N_5496,N_3819,N_4907);
xor U5497 (N_5497,N_4625,N_4657);
and U5498 (N_5498,N_4238,N_3960);
nand U5499 (N_5499,N_3788,N_2611);
xnor U5500 (N_5500,N_4297,N_3011);
and U5501 (N_5501,N_3744,N_2851);
nand U5502 (N_5502,N_4379,N_3046);
and U5503 (N_5503,N_4872,N_4011);
nand U5504 (N_5504,N_3838,N_3650);
or U5505 (N_5505,N_2649,N_3336);
and U5506 (N_5506,N_3252,N_4270);
and U5507 (N_5507,N_3652,N_3662);
and U5508 (N_5508,N_4940,N_3963);
nor U5509 (N_5509,N_3751,N_3895);
xor U5510 (N_5510,N_3988,N_2756);
and U5511 (N_5511,N_4153,N_4580);
nand U5512 (N_5512,N_3693,N_4741);
xor U5513 (N_5513,N_3585,N_4689);
or U5514 (N_5514,N_4539,N_3448);
or U5515 (N_5515,N_3601,N_3805);
or U5516 (N_5516,N_2898,N_3667);
xnor U5517 (N_5517,N_4446,N_3913);
xnor U5518 (N_5518,N_2771,N_2735);
and U5519 (N_5519,N_3608,N_4993);
and U5520 (N_5520,N_2894,N_4096);
or U5521 (N_5521,N_3376,N_2809);
nor U5522 (N_5522,N_2652,N_3229);
xnor U5523 (N_5523,N_2892,N_3800);
xor U5524 (N_5524,N_3000,N_4989);
and U5525 (N_5525,N_4799,N_2654);
or U5526 (N_5526,N_4043,N_4846);
or U5527 (N_5527,N_4398,N_4099);
nand U5528 (N_5528,N_3127,N_3432);
nor U5529 (N_5529,N_3977,N_4553);
xnor U5530 (N_5530,N_3982,N_3706);
nor U5531 (N_5531,N_3663,N_3247);
or U5532 (N_5532,N_4466,N_4311);
nand U5533 (N_5533,N_3511,N_3222);
or U5534 (N_5534,N_3361,N_4226);
nand U5535 (N_5535,N_3957,N_3790);
and U5536 (N_5536,N_4473,N_3658);
xnor U5537 (N_5537,N_3752,N_4578);
or U5538 (N_5538,N_2738,N_2869);
and U5539 (N_5539,N_2696,N_4795);
nor U5540 (N_5540,N_4349,N_4147);
or U5541 (N_5541,N_2788,N_4221);
xnor U5542 (N_5542,N_3602,N_4818);
nor U5543 (N_5543,N_4158,N_3185);
xor U5544 (N_5544,N_3489,N_4282);
nand U5545 (N_5545,N_4484,N_4702);
nand U5546 (N_5546,N_4970,N_3669);
nor U5547 (N_5547,N_3155,N_3952);
nor U5548 (N_5548,N_2856,N_4426);
and U5549 (N_5549,N_3561,N_3162);
nor U5550 (N_5550,N_4064,N_3956);
nor U5551 (N_5551,N_3743,N_4529);
and U5552 (N_5552,N_4575,N_4152);
nand U5553 (N_5553,N_3896,N_4276);
and U5554 (N_5554,N_4973,N_3327);
nand U5555 (N_5555,N_4612,N_3052);
and U5556 (N_5556,N_3394,N_3687);
xnor U5557 (N_5557,N_3851,N_3290);
nand U5558 (N_5558,N_2711,N_2836);
xnor U5559 (N_5559,N_2590,N_2555);
xor U5560 (N_5560,N_4845,N_2558);
nor U5561 (N_5561,N_4163,N_4423);
nor U5562 (N_5562,N_4312,N_3077);
and U5563 (N_5563,N_3128,N_3610);
nand U5564 (N_5564,N_2725,N_2791);
nand U5565 (N_5565,N_4667,N_4393);
and U5566 (N_5566,N_3049,N_4097);
and U5567 (N_5567,N_2523,N_4112);
nor U5568 (N_5568,N_4508,N_3916);
and U5569 (N_5569,N_3196,N_4574);
or U5570 (N_5570,N_3413,N_2609);
and U5571 (N_5571,N_4603,N_2639);
xnor U5572 (N_5572,N_3970,N_3528);
nand U5573 (N_5573,N_4405,N_2559);
and U5574 (N_5574,N_4726,N_3070);
or U5575 (N_5575,N_2714,N_4047);
nor U5576 (N_5576,N_3701,N_3216);
nand U5577 (N_5577,N_4206,N_4095);
nand U5578 (N_5578,N_4130,N_4586);
nand U5579 (N_5579,N_3073,N_3537);
nand U5580 (N_5580,N_3292,N_3771);
and U5581 (N_5581,N_3009,N_4815);
and U5582 (N_5582,N_2763,N_4730);
nand U5583 (N_5583,N_3606,N_4160);
nand U5584 (N_5584,N_2972,N_4118);
or U5585 (N_5585,N_3775,N_3538);
xnor U5586 (N_5586,N_4869,N_3648);
nand U5587 (N_5587,N_4582,N_4916);
nor U5588 (N_5588,N_4383,N_2592);
nor U5589 (N_5589,N_4697,N_4187);
or U5590 (N_5590,N_4289,N_4589);
nor U5591 (N_5591,N_3167,N_3075);
or U5592 (N_5592,N_3402,N_4243);
nor U5593 (N_5593,N_4991,N_4157);
and U5594 (N_5594,N_4005,N_4309);
nand U5595 (N_5595,N_4324,N_3665);
nor U5596 (N_5596,N_4758,N_4533);
xnor U5597 (N_5597,N_3678,N_3278);
xnor U5598 (N_5598,N_4088,N_3144);
and U5599 (N_5599,N_4406,N_3854);
xor U5600 (N_5600,N_3481,N_2537);
or U5601 (N_5601,N_4874,N_2640);
and U5602 (N_5602,N_3850,N_4602);
nor U5603 (N_5603,N_4936,N_4928);
nor U5604 (N_5604,N_4072,N_3731);
and U5605 (N_5605,N_2786,N_2895);
or U5606 (N_5606,N_3773,N_4561);
and U5607 (N_5607,N_3043,N_3681);
or U5608 (N_5608,N_3200,N_2762);
nand U5609 (N_5609,N_2908,N_3841);
xor U5610 (N_5610,N_3301,N_2534);
nor U5611 (N_5611,N_3430,N_4658);
nand U5612 (N_5612,N_3856,N_3984);
xor U5613 (N_5613,N_3579,N_3604);
or U5614 (N_5614,N_2914,N_3145);
and U5615 (N_5615,N_4250,N_3848);
nor U5616 (N_5616,N_4670,N_3502);
nor U5617 (N_5617,N_2973,N_4773);
or U5618 (N_5618,N_3830,N_3382);
and U5619 (N_5619,N_4425,N_3817);
nand U5620 (N_5620,N_3040,N_4485);
and U5621 (N_5621,N_3994,N_3641);
nor U5622 (N_5622,N_4955,N_3623);
nor U5623 (N_5623,N_4997,N_3140);
nor U5624 (N_5624,N_4966,N_3220);
nand U5625 (N_5625,N_4177,N_3033);
or U5626 (N_5626,N_4094,N_3030);
and U5627 (N_5627,N_3985,N_2577);
and U5628 (N_5628,N_4108,N_4964);
nor U5629 (N_5629,N_2943,N_4701);
nor U5630 (N_5630,N_4841,N_2583);
nor U5631 (N_5631,N_3010,N_3273);
xor U5632 (N_5632,N_4439,N_2911);
and U5633 (N_5633,N_4260,N_3398);
and U5634 (N_5634,N_4599,N_2920);
or U5635 (N_5635,N_4518,N_2613);
and U5636 (N_5636,N_3591,N_2793);
and U5637 (N_5637,N_3256,N_2996);
or U5638 (N_5638,N_2912,N_4803);
xor U5639 (N_5639,N_3526,N_3953);
xnor U5640 (N_5640,N_3153,N_4923);
and U5641 (N_5641,N_4696,N_4813);
xor U5642 (N_5642,N_2599,N_2891);
nor U5643 (N_5643,N_4983,N_3280);
and U5644 (N_5644,N_4524,N_3474);
or U5645 (N_5645,N_4904,N_4384);
xor U5646 (N_5646,N_3366,N_3450);
nand U5647 (N_5647,N_4375,N_3802);
nor U5648 (N_5648,N_4353,N_3670);
and U5649 (N_5649,N_3203,N_4986);
nand U5650 (N_5650,N_4032,N_4690);
nand U5651 (N_5651,N_4336,N_4898);
nand U5652 (N_5652,N_4514,N_3999);
and U5653 (N_5653,N_4873,N_4618);
or U5654 (N_5654,N_2903,N_2906);
xor U5655 (N_5655,N_4878,N_4420);
or U5656 (N_5656,N_4434,N_3423);
xnor U5657 (N_5657,N_4262,N_4918);
or U5658 (N_5658,N_4531,N_4610);
nand U5659 (N_5659,N_3657,N_4763);
and U5660 (N_5660,N_2571,N_4751);
or U5661 (N_5661,N_4025,N_4592);
xor U5662 (N_5662,N_3081,N_4840);
nand U5663 (N_5663,N_2594,N_4538);
xnor U5664 (N_5664,N_2870,N_2724);
or U5665 (N_5665,N_4740,N_3235);
nand U5666 (N_5666,N_2636,N_3683);
or U5667 (N_5667,N_4686,N_3798);
xnor U5668 (N_5668,N_4419,N_2842);
and U5669 (N_5669,N_3378,N_4494);
and U5670 (N_5670,N_4018,N_3505);
and U5671 (N_5671,N_4087,N_4748);
xor U5672 (N_5672,N_3416,N_3768);
nor U5673 (N_5673,N_2581,N_2978);
or U5674 (N_5674,N_3130,N_4802);
or U5675 (N_5675,N_4010,N_4671);
or U5676 (N_5676,N_2601,N_4911);
and U5677 (N_5677,N_4265,N_3885);
nor U5678 (N_5678,N_3357,N_4862);
or U5679 (N_5679,N_4339,N_4765);
xor U5680 (N_5680,N_4295,N_3639);
and U5681 (N_5681,N_3495,N_3444);
nor U5682 (N_5682,N_4652,N_3869);
nor U5683 (N_5683,N_2562,N_4501);
nor U5684 (N_5684,N_4746,N_3161);
or U5685 (N_5685,N_3844,N_4674);
nor U5686 (N_5686,N_2765,N_4656);
or U5687 (N_5687,N_4248,N_3257);
or U5688 (N_5688,N_4057,N_4719);
or U5689 (N_5689,N_3299,N_3061);
nand U5690 (N_5690,N_3169,N_3879);
xnor U5691 (N_5691,N_3324,N_2672);
nor U5692 (N_5692,N_4557,N_3150);
or U5693 (N_5693,N_4567,N_3108);
and U5694 (N_5694,N_3801,N_3803);
nand U5695 (N_5695,N_3761,N_4323);
nor U5696 (N_5696,N_3966,N_3992);
nand U5697 (N_5697,N_4981,N_3098);
or U5698 (N_5698,N_4315,N_3218);
xnor U5699 (N_5699,N_4123,N_3589);
nand U5700 (N_5700,N_2790,N_4461);
nand U5701 (N_5701,N_4073,N_3047);
nor U5702 (N_5702,N_2679,N_2745);
nor U5703 (N_5703,N_4368,N_4071);
nand U5704 (N_5704,N_4824,N_3271);
xnor U5705 (N_5705,N_4352,N_4826);
nor U5706 (N_5706,N_4303,N_3363);
and U5707 (N_5707,N_4545,N_3163);
and U5708 (N_5708,N_4760,N_4084);
xor U5709 (N_5709,N_3494,N_3587);
nor U5710 (N_5710,N_4341,N_4199);
nor U5711 (N_5711,N_3317,N_4090);
and U5712 (N_5712,N_4738,N_4666);
or U5713 (N_5713,N_4343,N_4129);
nor U5714 (N_5714,N_3971,N_2782);
nand U5715 (N_5715,N_3739,N_2635);
and U5716 (N_5716,N_4063,N_2722);
nand U5717 (N_5717,N_3842,N_4372);
or U5718 (N_5718,N_3019,N_4228);
nor U5719 (N_5719,N_4867,N_3866);
nand U5720 (N_5720,N_4829,N_4174);
nand U5721 (N_5721,N_4089,N_3551);
xnor U5722 (N_5722,N_4102,N_4263);
nor U5723 (N_5723,N_2730,N_3540);
nand U5724 (N_5724,N_3605,N_3562);
nand U5725 (N_5725,N_3482,N_4346);
nor U5726 (N_5726,N_3840,N_3766);
xor U5727 (N_5727,N_4573,N_3486);
nand U5728 (N_5728,N_3770,N_4218);
nand U5729 (N_5729,N_3404,N_2866);
nand U5730 (N_5730,N_4053,N_2861);
nor U5731 (N_5731,N_4125,N_2517);
xnor U5732 (N_5732,N_3917,N_3308);
or U5733 (N_5733,N_4258,N_3974);
and U5734 (N_5734,N_3776,N_3443);
and U5735 (N_5735,N_4505,N_3797);
or U5736 (N_5736,N_3558,N_2560);
nand U5737 (N_5737,N_4217,N_3377);
and U5738 (N_5738,N_2936,N_2979);
nor U5739 (N_5739,N_4825,N_3711);
xor U5740 (N_5740,N_3039,N_3961);
xor U5741 (N_5741,N_4638,N_3405);
nor U5742 (N_5742,N_4864,N_4651);
or U5743 (N_5743,N_4969,N_4338);
or U5744 (N_5744,N_3227,N_3733);
xor U5745 (N_5745,N_3820,N_4957);
nor U5746 (N_5746,N_4202,N_2500);
nor U5747 (N_5747,N_4098,N_4235);
xor U5748 (N_5748,N_3015,N_4500);
or U5749 (N_5749,N_4462,N_4114);
and U5750 (N_5750,N_3565,N_4984);
xor U5751 (N_5751,N_4067,N_4452);
xor U5752 (N_5752,N_4344,N_3351);
and U5753 (N_5753,N_4579,N_3901);
nor U5754 (N_5754,N_3079,N_4407);
xnor U5755 (N_5755,N_4863,N_4835);
or U5756 (N_5756,N_3422,N_4591);
and U5757 (N_5757,N_3434,N_4890);
nand U5758 (N_5758,N_3861,N_4476);
xor U5759 (N_5759,N_3630,N_3543);
nor U5760 (N_5760,N_4946,N_4972);
and U5761 (N_5761,N_4742,N_4490);
or U5762 (N_5762,N_4756,N_2772);
xnor U5763 (N_5763,N_4715,N_3417);
nand U5764 (N_5764,N_2913,N_3877);
and U5765 (N_5765,N_2550,N_4672);
nor U5766 (N_5766,N_4003,N_2632);
nor U5767 (N_5767,N_3254,N_4982);
nand U5768 (N_5768,N_2967,N_3020);
nor U5769 (N_5769,N_3045,N_2619);
nor U5770 (N_5770,N_3374,N_4361);
or U5771 (N_5771,N_4754,N_2618);
or U5772 (N_5772,N_4917,N_3569);
nor U5773 (N_5773,N_3236,N_4784);
nor U5774 (N_5774,N_4816,N_4365);
nor U5775 (N_5775,N_4595,N_3233);
and U5776 (N_5776,N_2685,N_3051);
and U5777 (N_5777,N_3111,N_3942);
nand U5778 (N_5778,N_2664,N_3392);
nand U5779 (N_5779,N_2928,N_4775);
or U5780 (N_5780,N_4974,N_3993);
or U5781 (N_5781,N_3214,N_3195);
or U5782 (N_5782,N_3240,N_4637);
xor U5783 (N_5783,N_4509,N_4930);
or U5784 (N_5784,N_4000,N_3276);
xnor U5785 (N_5785,N_3038,N_4959);
and U5786 (N_5786,N_3609,N_4183);
and U5787 (N_5787,N_4968,N_3488);
nand U5788 (N_5788,N_4934,N_3876);
nand U5789 (N_5789,N_3738,N_4266);
nor U5790 (N_5790,N_2717,N_4894);
or U5791 (N_5791,N_4337,N_4753);
nor U5792 (N_5792,N_4319,N_3978);
or U5793 (N_5793,N_2593,N_3832);
and U5794 (N_5794,N_3619,N_2623);
nand U5795 (N_5795,N_3323,N_4236);
xor U5796 (N_5796,N_4077,N_2536);
nand U5797 (N_5797,N_2910,N_4185);
or U5798 (N_5798,N_4275,N_2921);
nor U5799 (N_5799,N_3689,N_3638);
xor U5800 (N_5800,N_3091,N_4284);
nor U5801 (N_5801,N_3027,N_3763);
xor U5802 (N_5802,N_4944,N_4392);
or U5803 (N_5803,N_2668,N_3837);
nand U5804 (N_5804,N_4029,N_4596);
xnor U5805 (N_5805,N_3519,N_2516);
or U5806 (N_5806,N_3989,N_3873);
nor U5807 (N_5807,N_4866,N_3666);
and U5808 (N_5808,N_4308,N_3410);
or U5809 (N_5809,N_4794,N_4190);
or U5810 (N_5810,N_3412,N_4173);
nor U5811 (N_5811,N_4800,N_3399);
or U5812 (N_5812,N_2937,N_3059);
nand U5813 (N_5813,N_4897,N_4213);
or U5814 (N_5814,N_3533,N_3090);
or U5815 (N_5815,N_4229,N_4281);
and U5816 (N_5816,N_3210,N_3480);
or U5817 (N_5817,N_3205,N_2707);
and U5818 (N_5818,N_3141,N_3223);
nand U5819 (N_5819,N_2816,N_2977);
and U5820 (N_5820,N_4007,N_3146);
nand U5821 (N_5821,N_4298,N_4937);
or U5822 (N_5822,N_3442,N_3529);
xor U5823 (N_5823,N_4705,N_4764);
xor U5824 (N_5824,N_2807,N_4772);
and U5825 (N_5825,N_4222,N_2607);
and U5826 (N_5826,N_2874,N_3175);
or U5827 (N_5827,N_3329,N_2670);
nand U5828 (N_5828,N_3477,N_3058);
nor U5829 (N_5829,N_2694,N_4215);
xor U5830 (N_5830,N_2616,N_4640);
xor U5831 (N_5831,N_4615,N_3234);
nand U5832 (N_5832,N_4347,N_2739);
xnor U5833 (N_5833,N_3786,N_2630);
or U5834 (N_5834,N_4021,N_4288);
or U5835 (N_5835,N_4774,N_4301);
and U5836 (N_5836,N_3794,N_2561);
xor U5837 (N_5837,N_3958,N_4522);
nor U5838 (N_5838,N_4366,N_3496);
or U5839 (N_5839,N_4761,N_4280);
and U5840 (N_5840,N_4920,N_2757);
nand U5841 (N_5841,N_2954,N_4948);
nor U5842 (N_5842,N_4571,N_4885);
nor U5843 (N_5843,N_2867,N_4035);
nor U5844 (N_5844,N_4992,N_2755);
and U5845 (N_5845,N_3607,N_3041);
or U5846 (N_5846,N_4743,N_3110);
nand U5847 (N_5847,N_4389,N_3464);
and U5848 (N_5848,N_2833,N_2821);
xnor U5849 (N_5849,N_4059,N_3929);
nor U5850 (N_5850,N_3858,N_4438);
nor U5851 (N_5851,N_3244,N_4521);
and U5852 (N_5852,N_2990,N_4617);
nand U5853 (N_5853,N_3370,N_4316);
and U5854 (N_5854,N_4050,N_3478);
nand U5855 (N_5855,N_3093,N_3707);
xor U5856 (N_5856,N_4171,N_4933);
and U5857 (N_5857,N_2841,N_2795);
nand U5858 (N_5858,N_4626,N_4477);
nor U5859 (N_5859,N_4176,N_4335);
or U5860 (N_5860,N_4454,N_3586);
and U5861 (N_5861,N_3764,N_2666);
xor U5862 (N_5862,N_4068,N_3948);
xor U5863 (N_5863,N_3539,N_4359);
or U5864 (N_5864,N_2916,N_3001);
xnor U5865 (N_5865,N_3025,N_4884);
or U5866 (N_5866,N_3938,N_3172);
xnor U5867 (N_5867,N_4447,N_3898);
or U5868 (N_5868,N_4469,N_2749);
and U5869 (N_5869,N_4771,N_4278);
and U5870 (N_5870,N_2787,N_3076);
and U5871 (N_5871,N_3789,N_4749);
xnor U5872 (N_5872,N_4448,N_3215);
nand U5873 (N_5873,N_2995,N_3409);
or U5874 (N_5874,N_3050,N_4042);
or U5875 (N_5875,N_4463,N_2976);
xor U5876 (N_5876,N_4450,N_3635);
xnor U5877 (N_5877,N_3765,N_3827);
and U5878 (N_5878,N_4240,N_3907);
xnor U5879 (N_5879,N_3889,N_3615);
or U5880 (N_5880,N_4367,N_3258);
and U5881 (N_5881,N_4155,N_2917);
nand U5882 (N_5882,N_3688,N_3358);
nor U5883 (N_5883,N_2610,N_3975);
nor U5884 (N_5884,N_4838,N_3795);
xnor U5885 (N_5885,N_4471,N_3900);
or U5886 (N_5886,N_3749,N_3391);
xor U5887 (N_5887,N_2643,N_3987);
xor U5888 (N_5888,N_3990,N_2531);
or U5889 (N_5889,N_3071,N_4683);
or U5890 (N_5890,N_3375,N_4549);
nor U5891 (N_5891,N_4382,N_2860);
or U5892 (N_5892,N_2698,N_4785);
nor U5893 (N_5893,N_4348,N_3004);
nor U5894 (N_5894,N_3475,N_3506);
xor U5895 (N_5895,N_2554,N_3933);
nand U5896 (N_5896,N_3395,N_3333);
xnor U5897 (N_5897,N_4430,N_3983);
nand U5898 (N_5898,N_3564,N_4028);
or U5899 (N_5899,N_4954,N_2622);
nand U5900 (N_5900,N_4034,N_4854);
nor U5901 (N_5901,N_2751,N_3053);
and U5902 (N_5902,N_4080,N_4739);
xnor U5903 (N_5903,N_3109,N_3002);
nand U5904 (N_5904,N_3584,N_3232);
nor U5905 (N_5905,N_3867,N_4380);
xor U5906 (N_5906,N_2901,N_2849);
and U5907 (N_5907,N_3003,N_2775);
and U5908 (N_5908,N_3886,N_2587);
nor U5909 (N_5909,N_4931,N_3718);
nand U5910 (N_5910,N_3581,N_3655);
nand U5911 (N_5911,N_3016,N_4082);
or U5912 (N_5912,N_4482,N_4836);
nor U5913 (N_5913,N_2731,N_3193);
nand U5914 (N_5914,N_4870,N_4277);
nand U5915 (N_5915,N_2527,N_2520);
nand U5916 (N_5916,N_4546,N_4432);
and U5917 (N_5917,N_2549,N_4117);
nor U5918 (N_5918,N_3224,N_4172);
and U5919 (N_5919,N_2629,N_4493);
or U5920 (N_5920,N_3863,N_3313);
nor U5921 (N_5921,N_3732,N_3245);
or U5922 (N_5922,N_2879,N_3614);
nand U5923 (N_5923,N_4386,N_4491);
or U5924 (N_5924,N_4682,N_4039);
and U5925 (N_5925,N_4422,N_3473);
and U5926 (N_5926,N_4778,N_4409);
or U5927 (N_5927,N_3757,N_3157);
and U5928 (N_5928,N_4060,N_3345);
or U5929 (N_5929,N_2584,N_3119);
xnor U5930 (N_5930,N_3647,N_4246);
nand U5931 (N_5931,N_2843,N_2808);
xor U5932 (N_5932,N_4635,N_4455);
nand U5933 (N_5933,N_4958,N_3012);
nand U5934 (N_5934,N_3928,N_3420);
or U5935 (N_5935,N_4092,N_4049);
or U5936 (N_5936,N_3592,N_3191);
nand U5937 (N_5937,N_4924,N_2579);
xnor U5938 (N_5938,N_3069,N_4107);
and U5939 (N_5939,N_3881,N_2686);
nor U5940 (N_5940,N_3811,N_3400);
or U5941 (N_5941,N_2508,N_2695);
and U5942 (N_5942,N_2932,N_4737);
and U5943 (N_5943,N_2661,N_2998);
nor U5944 (N_5944,N_4735,N_2657);
nor U5945 (N_5945,N_4576,N_3460);
and U5946 (N_5946,N_4849,N_4362);
and U5947 (N_5947,N_3921,N_4175);
nand U5948 (N_5948,N_2589,N_2608);
xor U5949 (N_5949,N_3703,N_4895);
nor U5950 (N_5950,N_3508,N_3483);
or U5951 (N_5951,N_2712,N_3513);
or U5952 (N_5952,N_3491,N_4844);
nor U5953 (N_5953,N_4453,N_2811);
nand U5954 (N_5954,N_2582,N_2659);
or U5955 (N_5955,N_4953,N_4355);
nand U5956 (N_5956,N_3745,N_4304);
or U5957 (N_5957,N_2522,N_4223);
and U5958 (N_5958,N_4233,N_3871);
xor U5959 (N_5959,N_4556,N_4594);
nand U5960 (N_5960,N_3705,N_3134);
nand U5961 (N_5961,N_2777,N_2983);
and U5962 (N_5962,N_2612,N_4631);
and U5963 (N_5963,N_3124,N_2552);
xnor U5964 (N_5964,N_3202,N_3747);
nor U5965 (N_5965,N_3644,N_4091);
or U5966 (N_5966,N_3535,N_4912);
xnor U5967 (N_5967,N_3574,N_2784);
or U5968 (N_5968,N_2909,N_3131);
and U5969 (N_5969,N_3456,N_2543);
xor U5970 (N_5970,N_4693,N_4017);
nor U5971 (N_5971,N_2538,N_4078);
xor U5972 (N_5972,N_3194,N_3156);
nor U5973 (N_5973,N_2644,N_3347);
nand U5974 (N_5974,N_3532,N_4408);
and U5975 (N_5975,N_2641,N_3719);
and U5976 (N_5976,N_3708,N_3887);
nand U5977 (N_5977,N_3808,N_3286);
nor U5978 (N_5978,N_3945,N_4209);
nor U5979 (N_5979,N_3954,N_4723);
nor U5980 (N_5980,N_4274,N_3695);
or U5981 (N_5981,N_4273,N_3411);
xnor U5982 (N_5982,N_4622,N_2844);
nand U5983 (N_5983,N_2663,N_4830);
and U5984 (N_5984,N_3694,N_2966);
and U5985 (N_5985,N_3697,N_3868);
xor U5986 (N_5986,N_3684,N_4861);
nand U5987 (N_5987,N_4391,N_3097);
and U5988 (N_5988,N_3925,N_3279);
nand U5989 (N_5989,N_4166,N_2507);
nor U5990 (N_5990,N_2547,N_3063);
and U5991 (N_5991,N_4120,N_3734);
xor U5992 (N_5992,N_3427,N_2662);
nor U5993 (N_5993,N_3425,N_2615);
or U5994 (N_5994,N_2506,N_4156);
nor U5995 (N_5995,N_2902,N_3428);
nand U5996 (N_5996,N_4633,N_4645);
nor U5997 (N_5997,N_3599,N_3653);
xnor U5998 (N_5998,N_3810,N_4843);
xnor U5999 (N_5999,N_4111,N_3438);
and U6000 (N_6000,N_4247,N_4528);
and U6001 (N_6001,N_2847,N_2539);
and U6002 (N_6002,N_3729,N_3997);
and U6003 (N_6003,N_4909,N_3186);
or U6004 (N_6004,N_3590,N_2827);
xnor U6005 (N_6005,N_4269,N_3013);
nor U6006 (N_6006,N_4433,N_4381);
or U6007 (N_6007,N_4008,N_4745);
xnor U6008 (N_6008,N_4879,N_3298);
xnor U6009 (N_6009,N_4143,N_2574);
nor U6010 (N_6010,N_2603,N_3338);
nor U6011 (N_6011,N_2999,N_2896);
or U6012 (N_6012,N_3557,N_4793);
nand U6013 (N_6013,N_2512,N_3583);
nor U6014 (N_6014,N_4207,N_4180);
or U6015 (N_6015,N_3713,N_3777);
xnor U6016 (N_6016,N_3490,N_4033);
and U6017 (N_6017,N_3507,N_2688);
nand U6018 (N_6018,N_4988,N_4504);
xor U6019 (N_6019,N_4587,N_4138);
nand U6020 (N_6020,N_3559,N_4045);
or U6021 (N_6021,N_3892,N_3154);
nor U6022 (N_6022,N_4828,N_3517);
nand U6023 (N_6023,N_3897,N_4457);
and U6024 (N_6024,N_3242,N_2814);
nor U6025 (N_6025,N_3780,N_2598);
nand U6026 (N_6026,N_3295,N_2832);
nand U6027 (N_6027,N_2889,N_2708);
and U6028 (N_6028,N_2804,N_4759);
or U6029 (N_6029,N_4769,N_4779);
or U6030 (N_6030,N_4131,N_3853);
nor U6031 (N_6031,N_3243,N_2955);
xor U6032 (N_6032,N_3580,N_3600);
or U6033 (N_6033,N_4340,N_2962);
and U6034 (N_6034,N_4342,N_3044);
nand U6035 (N_6035,N_3633,N_3282);
and U6036 (N_6036,N_3717,N_4106);
nand U6037 (N_6037,N_4630,N_4314);
or U6038 (N_6038,N_2528,N_3787);
xor U6039 (N_6039,N_4220,N_2834);
nand U6040 (N_6040,N_2840,N_3089);
nand U6041 (N_6041,N_4031,N_3318);
xnor U6042 (N_6042,N_3712,N_3995);
xor U6043 (N_6043,N_4411,N_4066);
and U6044 (N_6044,N_4124,N_4691);
nor U6045 (N_6045,N_3451,N_3578);
xor U6046 (N_6046,N_4465,N_3147);
xor U6047 (N_6047,N_4259,N_4204);
nor U6048 (N_6048,N_3510,N_4237);
or U6049 (N_6049,N_4833,N_2890);
or U6050 (N_6050,N_3651,N_3893);
xnor U6051 (N_6051,N_3452,N_4200);
or U6052 (N_6052,N_3080,N_4317);
or U6053 (N_6053,N_3468,N_4041);
and U6054 (N_6054,N_4148,N_2862);
xor U6055 (N_6055,N_2872,N_3439);
nand U6056 (N_6056,N_3906,N_4888);
xor U6057 (N_6057,N_4006,N_3603);
xor U6058 (N_6058,N_2676,N_2586);
nor U6059 (N_6059,N_4648,N_4506);
nand U6060 (N_6060,N_4882,N_3521);
xor U6061 (N_6061,N_2802,N_2900);
xnor U6062 (N_6062,N_3067,N_4527);
or U6063 (N_6063,N_3627,N_2720);
nor U6064 (N_6064,N_3275,N_3672);
nand U6065 (N_6065,N_3424,N_2828);
or U6066 (N_6066,N_3497,N_3546);
xor U6067 (N_6067,N_4300,N_3355);
xor U6068 (N_6068,N_3367,N_3485);
and U6069 (N_6069,N_3571,N_4093);
nor U6070 (N_6070,N_4400,N_3446);
xor U6071 (N_6071,N_4678,N_3727);
and U6072 (N_6072,N_2826,N_2926);
and U6073 (N_6073,N_2624,N_4267);
nor U6074 (N_6074,N_3943,N_3462);
nor U6075 (N_6075,N_4291,N_2997);
nand U6076 (N_6076,N_2975,N_4757);
and U6077 (N_6077,N_4489,N_3875);
nand U6078 (N_6078,N_2876,N_4004);
nand U6079 (N_6079,N_4105,N_3207);
nor U6080 (N_6080,N_4932,N_2556);
or U6081 (N_6081,N_3702,N_3250);
nand U6082 (N_6082,N_3936,N_3629);
or U6083 (N_6083,N_4030,N_3024);
or U6084 (N_6084,N_4609,N_2859);
xnor U6085 (N_6085,N_3133,N_4332);
or U6086 (N_6086,N_3251,N_2532);
and U6087 (N_6087,N_3088,N_4698);
and U6088 (N_6088,N_3806,N_3527);
xnor U6089 (N_6089,N_3632,N_4334);
or U6090 (N_6090,N_3660,N_2783);
nor U6091 (N_6091,N_2542,N_4927);
nor U6092 (N_6092,N_4128,N_3272);
nand U6093 (N_6093,N_3036,N_3512);
xor U6094 (N_6094,N_3894,N_2933);
xnor U6095 (N_6095,N_4655,N_3032);
and U6096 (N_6096,N_2982,N_4687);
xnor U6097 (N_6097,N_3479,N_4253);
nand U6098 (N_6098,N_4181,N_4421);
nand U6099 (N_6099,N_2759,N_4472);
and U6100 (N_6100,N_2883,N_3556);
xor U6101 (N_6101,N_3165,N_2511);
nand U6102 (N_6102,N_4971,N_3968);
nor U6103 (N_6103,N_4605,N_4977);
or U6104 (N_6104,N_4664,N_3415);
nand U6105 (N_6105,N_4662,N_3114);
nor U6106 (N_6106,N_2881,N_3065);
and U6107 (N_6107,N_4620,N_2591);
or U6108 (N_6108,N_3005,N_3646);
or U6109 (N_6109,N_2899,N_2699);
nor U6110 (N_6110,N_4703,N_4076);
nor U6111 (N_6111,N_4699,N_2942);
nor U6112 (N_6112,N_3969,N_4967);
or U6113 (N_6113,N_4445,N_4536);
nor U6114 (N_6114,N_2853,N_4889);
xor U6115 (N_6115,N_3230,N_3142);
or U6116 (N_6116,N_4554,N_3331);
nand U6117 (N_6117,N_3436,N_3582);
and U6118 (N_6118,N_3530,N_4135);
and U6119 (N_6119,N_3310,N_4555);
nand U6120 (N_6120,N_4119,N_3597);
or U6121 (N_6121,N_4022,N_4781);
and U6122 (N_6122,N_4395,N_3566);
xor U6123 (N_6123,N_3555,N_2831);
nor U6124 (N_6124,N_2960,N_2778);
and U6125 (N_6125,N_3344,N_3221);
or U6126 (N_6126,N_2605,N_4654);
nor U6127 (N_6127,N_4856,N_4711);
xor U6128 (N_6128,N_2541,N_3083);
xnor U6129 (N_6129,N_3576,N_3570);
nor U6130 (N_6130,N_4134,N_3349);
or U6131 (N_6131,N_3682,N_3807);
xor U6132 (N_6132,N_2986,N_4184);
or U6133 (N_6133,N_4394,N_4203);
nor U6134 (N_6134,N_4121,N_2852);
nand U6135 (N_6135,N_4296,N_3515);
nor U6136 (N_6136,N_4154,N_4515);
and U6137 (N_6137,N_4980,N_2646);
nor U6138 (N_6138,N_3654,N_2988);
and U6139 (N_6139,N_3553,N_2752);
xor U6140 (N_6140,N_4479,N_2585);
nor U6141 (N_6141,N_3107,N_3388);
xor U6142 (N_6142,N_3724,N_3920);
nor U6143 (N_6143,N_2950,N_4351);
or U6144 (N_6144,N_3903,N_4926);
nor U6145 (N_6145,N_3190,N_4901);
nor U6146 (N_6146,N_2614,N_3835);
or U6147 (N_6147,N_3847,N_3774);
nor U6148 (N_6148,N_2620,N_3449);
nand U6149 (N_6149,N_4272,N_3048);
nand U6150 (N_6150,N_3675,N_4877);
xnor U6151 (N_6151,N_4569,N_4431);
nand U6152 (N_6152,N_3265,N_3023);
and U6153 (N_6153,N_4905,N_3613);
nor U6154 (N_6154,N_4385,N_3231);
nand U6155 (N_6155,N_3914,N_2750);
nor U6156 (N_6156,N_4881,N_3469);
nor U6157 (N_6157,N_3828,N_4333);
or U6158 (N_6158,N_3637,N_4673);
nand U6159 (N_6159,N_3645,N_4140);
nor U6160 (N_6160,N_4950,N_4239);
and U6161 (N_6161,N_3922,N_3334);
nand U6162 (N_6162,N_3026,N_4942);
and U6163 (N_6163,N_3447,N_4496);
and U6164 (N_6164,N_3117,N_3177);
nor U6165 (N_6165,N_3594,N_3031);
xnor U6166 (N_6166,N_4768,N_4363);
nor U6167 (N_6167,N_4294,N_2606);
nand U6168 (N_6168,N_3340,N_4597);
xnor U6169 (N_6169,N_2721,N_4492);
xor U6170 (N_6170,N_4127,N_3074);
nand U6171 (N_6171,N_2529,N_4732);
or U6172 (N_6172,N_3068,N_4805);
xnor U6173 (N_6173,N_4255,N_4704);
or U6174 (N_6174,N_4837,N_3769);
or U6175 (N_6175,N_4858,N_4193);
nor U6176 (N_6176,N_2798,N_3120);
and U6177 (N_6177,N_4216,N_2706);
xor U6178 (N_6178,N_3441,N_3170);
nand U6179 (N_6179,N_3238,N_3311);
nor U6180 (N_6180,N_4162,N_4261);
nand U6181 (N_6181,N_4718,N_2710);
nor U6182 (N_6182,N_4700,N_2953);
nor U6183 (N_6183,N_2667,N_4310);
xnor U6184 (N_6184,N_4427,N_4681);
and U6185 (N_6185,N_4985,N_3784);
or U6186 (N_6186,N_2627,N_4925);
xnor U6187 (N_6187,N_4179,N_4245);
nand U6188 (N_6188,N_4752,N_2690);
nor U6189 (N_6189,N_4478,N_4935);
and U6190 (N_6190,N_4364,N_4649);
and U6191 (N_6191,N_4621,N_2858);
nor U6192 (N_6192,N_4065,N_4535);
and U6193 (N_6193,N_2683,N_4736);
or U6194 (N_6194,N_2702,N_2805);
xor U6195 (N_6195,N_4256,N_4499);
xnor U6196 (N_6196,N_4109,N_4787);
and U6197 (N_6197,N_3964,N_2638);
nand U6198 (N_6198,N_3354,N_2521);
nand U6199 (N_6199,N_4541,N_2820);
or U6200 (N_6200,N_4642,N_2945);
or U6201 (N_6201,N_3549,N_3118);
xnor U6202 (N_6202,N_3878,N_4811);
xor U6203 (N_6203,N_3379,N_2971);
nor U6204 (N_6204,N_3103,N_3932);
and U6205 (N_6205,N_4646,N_4550);
and U6206 (N_6206,N_2575,N_3268);
nor U6207 (N_6207,N_3249,N_3296);
and U6208 (N_6208,N_2524,N_4085);
nor U6209 (N_6209,N_3213,N_4502);
nor U6210 (N_6210,N_3178,N_4910);
and U6211 (N_6211,N_4949,N_4415);
nor U6212 (N_6212,N_3742,N_3471);
and U6213 (N_6213,N_4707,N_4086);
xnor U6214 (N_6214,N_3095,N_2877);
nor U6215 (N_6215,N_2803,N_3536);
xnor U6216 (N_6216,N_4604,N_3261);
nand U6217 (N_6217,N_3397,N_4606);
and U6218 (N_6218,N_2991,N_4975);
nor U6219 (N_6219,N_4286,N_3563);
and U6220 (N_6220,N_2957,N_2633);
and U6221 (N_6221,N_2595,N_2588);
nor U6222 (N_6222,N_4232,N_4440);
xnor U6223 (N_6223,N_2565,N_2796);
or U6224 (N_6224,N_3166,N_4290);
nand U6225 (N_6225,N_3371,N_3781);
nand U6226 (N_6226,N_3595,N_2578);
and U6227 (N_6227,N_4568,N_4847);
and U6228 (N_6228,N_2940,N_2774);
and U6229 (N_6229,N_4669,N_3307);
xor U6230 (N_6230,N_3709,N_3198);
and U6231 (N_6231,N_2964,N_4632);
nand U6232 (N_6232,N_2987,N_3104);
and U6233 (N_6233,N_4767,N_4331);
xor U6234 (N_6234,N_4523,N_3267);
nor U6235 (N_6235,N_3353,N_3380);
nand U6236 (N_6236,N_3753,N_3699);
or U6237 (N_6237,N_4327,N_4464);
nor U6238 (N_6238,N_3368,N_4559);
and U6239 (N_6239,N_3309,N_4115);
nor U6240 (N_6240,N_4817,N_3183);
nor U6241 (N_6241,N_3544,N_4565);
nand U6242 (N_6242,N_3160,N_2674);
or U6243 (N_6243,N_2984,N_2681);
or U6244 (N_6244,N_4081,N_4161);
nand U6245 (N_6245,N_3304,N_3315);
nor U6246 (N_6246,N_4205,N_4519);
or U6247 (N_6247,N_4169,N_3908);
and U6248 (N_6248,N_2742,N_4525);
nand U6249 (N_6249,N_4133,N_4251);
or U6250 (N_6250,N_3517,N_4590);
and U6251 (N_6251,N_3731,N_4032);
nor U6252 (N_6252,N_2722,N_4891);
nand U6253 (N_6253,N_3052,N_3379);
or U6254 (N_6254,N_2737,N_3964);
nand U6255 (N_6255,N_4792,N_4714);
nand U6256 (N_6256,N_2732,N_4352);
or U6257 (N_6257,N_3028,N_2850);
nand U6258 (N_6258,N_2529,N_3328);
nor U6259 (N_6259,N_4757,N_2618);
and U6260 (N_6260,N_4796,N_3743);
xor U6261 (N_6261,N_3452,N_2781);
xor U6262 (N_6262,N_3433,N_3844);
nand U6263 (N_6263,N_3140,N_3132);
nand U6264 (N_6264,N_3986,N_4869);
or U6265 (N_6265,N_3891,N_2634);
xor U6266 (N_6266,N_3172,N_3127);
and U6267 (N_6267,N_4148,N_3049);
and U6268 (N_6268,N_3647,N_4841);
nand U6269 (N_6269,N_4648,N_2888);
and U6270 (N_6270,N_2509,N_4318);
and U6271 (N_6271,N_2771,N_3946);
and U6272 (N_6272,N_2539,N_4262);
and U6273 (N_6273,N_4198,N_3261);
nor U6274 (N_6274,N_4629,N_4200);
and U6275 (N_6275,N_4198,N_3766);
xor U6276 (N_6276,N_4422,N_4511);
nor U6277 (N_6277,N_4549,N_4124);
nand U6278 (N_6278,N_2880,N_2571);
nand U6279 (N_6279,N_2799,N_3579);
nand U6280 (N_6280,N_3422,N_4053);
and U6281 (N_6281,N_3532,N_3967);
xnor U6282 (N_6282,N_2667,N_4098);
nor U6283 (N_6283,N_4473,N_4953);
nor U6284 (N_6284,N_4283,N_4731);
and U6285 (N_6285,N_3654,N_4290);
nor U6286 (N_6286,N_3236,N_2599);
nand U6287 (N_6287,N_2546,N_4635);
or U6288 (N_6288,N_3637,N_3277);
nor U6289 (N_6289,N_4821,N_4284);
or U6290 (N_6290,N_4917,N_3433);
nand U6291 (N_6291,N_2514,N_3174);
nor U6292 (N_6292,N_3351,N_4843);
or U6293 (N_6293,N_4674,N_2723);
nor U6294 (N_6294,N_4000,N_3890);
nand U6295 (N_6295,N_4680,N_3286);
or U6296 (N_6296,N_2506,N_3807);
or U6297 (N_6297,N_2838,N_4542);
nor U6298 (N_6298,N_4739,N_3012);
and U6299 (N_6299,N_3256,N_4932);
or U6300 (N_6300,N_4929,N_4040);
nand U6301 (N_6301,N_3590,N_2650);
and U6302 (N_6302,N_4770,N_2949);
nor U6303 (N_6303,N_3196,N_4179);
nor U6304 (N_6304,N_3711,N_3241);
or U6305 (N_6305,N_3840,N_4959);
nand U6306 (N_6306,N_3793,N_3403);
and U6307 (N_6307,N_2700,N_2776);
xor U6308 (N_6308,N_3491,N_3752);
nor U6309 (N_6309,N_3790,N_2683);
nor U6310 (N_6310,N_3342,N_4391);
nor U6311 (N_6311,N_3627,N_4273);
and U6312 (N_6312,N_4287,N_4664);
xnor U6313 (N_6313,N_4376,N_2930);
nor U6314 (N_6314,N_4909,N_4170);
nand U6315 (N_6315,N_2613,N_3971);
nand U6316 (N_6316,N_3634,N_3689);
or U6317 (N_6317,N_3844,N_4069);
nor U6318 (N_6318,N_3998,N_4638);
or U6319 (N_6319,N_4954,N_2767);
and U6320 (N_6320,N_3749,N_3508);
nor U6321 (N_6321,N_4980,N_4403);
xnor U6322 (N_6322,N_2879,N_2876);
or U6323 (N_6323,N_3447,N_4524);
or U6324 (N_6324,N_4513,N_2720);
or U6325 (N_6325,N_2610,N_2581);
xor U6326 (N_6326,N_3085,N_4314);
and U6327 (N_6327,N_2958,N_4452);
xnor U6328 (N_6328,N_4231,N_4091);
xor U6329 (N_6329,N_4105,N_3337);
nand U6330 (N_6330,N_2857,N_3825);
nand U6331 (N_6331,N_3358,N_2904);
and U6332 (N_6332,N_4793,N_3267);
nand U6333 (N_6333,N_2982,N_4123);
xnor U6334 (N_6334,N_4129,N_4777);
nor U6335 (N_6335,N_2544,N_4731);
nand U6336 (N_6336,N_2827,N_4565);
nor U6337 (N_6337,N_2960,N_2518);
nand U6338 (N_6338,N_2786,N_3896);
nand U6339 (N_6339,N_4461,N_4902);
or U6340 (N_6340,N_3942,N_2730);
and U6341 (N_6341,N_2528,N_4860);
nand U6342 (N_6342,N_2513,N_2894);
nand U6343 (N_6343,N_4188,N_4820);
or U6344 (N_6344,N_3094,N_3715);
or U6345 (N_6345,N_4707,N_3244);
xor U6346 (N_6346,N_4290,N_3208);
xor U6347 (N_6347,N_3693,N_3783);
nor U6348 (N_6348,N_3915,N_4962);
or U6349 (N_6349,N_4142,N_2878);
or U6350 (N_6350,N_3426,N_4091);
or U6351 (N_6351,N_2738,N_2546);
nand U6352 (N_6352,N_4790,N_3084);
nor U6353 (N_6353,N_4964,N_4958);
or U6354 (N_6354,N_2881,N_4928);
nor U6355 (N_6355,N_3916,N_3905);
and U6356 (N_6356,N_4902,N_3712);
or U6357 (N_6357,N_4528,N_3175);
nor U6358 (N_6358,N_2599,N_3546);
nand U6359 (N_6359,N_3933,N_3239);
nand U6360 (N_6360,N_4116,N_4876);
or U6361 (N_6361,N_3220,N_4133);
or U6362 (N_6362,N_3130,N_3923);
nand U6363 (N_6363,N_4136,N_3834);
or U6364 (N_6364,N_4432,N_4531);
nor U6365 (N_6365,N_4960,N_4641);
nor U6366 (N_6366,N_2550,N_2623);
nand U6367 (N_6367,N_3092,N_2588);
nor U6368 (N_6368,N_4646,N_2832);
nor U6369 (N_6369,N_3297,N_4945);
and U6370 (N_6370,N_4776,N_3082);
and U6371 (N_6371,N_4586,N_4741);
xor U6372 (N_6372,N_3708,N_4049);
nor U6373 (N_6373,N_3318,N_3688);
and U6374 (N_6374,N_2519,N_2990);
nor U6375 (N_6375,N_3469,N_4275);
nand U6376 (N_6376,N_3067,N_4833);
nor U6377 (N_6377,N_4882,N_4758);
xor U6378 (N_6378,N_4625,N_4477);
xor U6379 (N_6379,N_4551,N_3948);
or U6380 (N_6380,N_3656,N_4648);
or U6381 (N_6381,N_3755,N_3746);
or U6382 (N_6382,N_3809,N_4139);
or U6383 (N_6383,N_3950,N_4286);
nor U6384 (N_6384,N_4041,N_3309);
or U6385 (N_6385,N_4313,N_3578);
nor U6386 (N_6386,N_3816,N_2794);
nor U6387 (N_6387,N_3584,N_3714);
and U6388 (N_6388,N_3753,N_4103);
and U6389 (N_6389,N_4212,N_3671);
nor U6390 (N_6390,N_3931,N_3713);
nand U6391 (N_6391,N_3441,N_2781);
or U6392 (N_6392,N_2791,N_4853);
or U6393 (N_6393,N_2982,N_3963);
nor U6394 (N_6394,N_4712,N_3262);
xnor U6395 (N_6395,N_3531,N_4208);
nand U6396 (N_6396,N_3439,N_2723);
or U6397 (N_6397,N_3765,N_4505);
xor U6398 (N_6398,N_3913,N_4816);
nand U6399 (N_6399,N_3813,N_4669);
and U6400 (N_6400,N_3711,N_2537);
xor U6401 (N_6401,N_3161,N_2756);
and U6402 (N_6402,N_4641,N_2532);
xor U6403 (N_6403,N_4997,N_3244);
and U6404 (N_6404,N_4802,N_3205);
xnor U6405 (N_6405,N_4287,N_3633);
nand U6406 (N_6406,N_3231,N_4632);
or U6407 (N_6407,N_4259,N_4409);
or U6408 (N_6408,N_4645,N_3108);
xnor U6409 (N_6409,N_3739,N_2850);
nand U6410 (N_6410,N_2677,N_2967);
xor U6411 (N_6411,N_3745,N_4353);
nand U6412 (N_6412,N_3458,N_3964);
and U6413 (N_6413,N_2625,N_4576);
and U6414 (N_6414,N_4075,N_3262);
nor U6415 (N_6415,N_4881,N_4599);
nor U6416 (N_6416,N_3969,N_3460);
nor U6417 (N_6417,N_4379,N_4458);
or U6418 (N_6418,N_3391,N_2817);
nand U6419 (N_6419,N_2680,N_2884);
nand U6420 (N_6420,N_3984,N_2961);
nor U6421 (N_6421,N_2946,N_3458);
or U6422 (N_6422,N_3127,N_3827);
and U6423 (N_6423,N_4704,N_3565);
and U6424 (N_6424,N_3126,N_4544);
xor U6425 (N_6425,N_3311,N_3723);
nand U6426 (N_6426,N_4086,N_3311);
or U6427 (N_6427,N_3096,N_4106);
nor U6428 (N_6428,N_4090,N_4017);
nand U6429 (N_6429,N_4406,N_4840);
nand U6430 (N_6430,N_4685,N_4617);
xnor U6431 (N_6431,N_4733,N_3127);
nor U6432 (N_6432,N_4138,N_2881);
or U6433 (N_6433,N_4302,N_3010);
or U6434 (N_6434,N_2910,N_4983);
or U6435 (N_6435,N_2522,N_4816);
and U6436 (N_6436,N_4292,N_3879);
and U6437 (N_6437,N_2730,N_4743);
or U6438 (N_6438,N_4380,N_3510);
nor U6439 (N_6439,N_3151,N_4990);
nand U6440 (N_6440,N_3737,N_4183);
xor U6441 (N_6441,N_4177,N_2729);
nor U6442 (N_6442,N_3603,N_3428);
xnor U6443 (N_6443,N_3154,N_2911);
nand U6444 (N_6444,N_2643,N_4850);
xnor U6445 (N_6445,N_3582,N_4710);
or U6446 (N_6446,N_3567,N_3540);
nor U6447 (N_6447,N_2770,N_3496);
nand U6448 (N_6448,N_4032,N_4637);
nand U6449 (N_6449,N_4156,N_4626);
or U6450 (N_6450,N_4200,N_4540);
nand U6451 (N_6451,N_4464,N_2656);
or U6452 (N_6452,N_4368,N_2735);
or U6453 (N_6453,N_4342,N_2582);
xnor U6454 (N_6454,N_4710,N_4742);
nand U6455 (N_6455,N_4879,N_3007);
xor U6456 (N_6456,N_4222,N_4104);
or U6457 (N_6457,N_2779,N_4210);
and U6458 (N_6458,N_4570,N_4030);
xnor U6459 (N_6459,N_3202,N_3570);
nor U6460 (N_6460,N_2516,N_4360);
or U6461 (N_6461,N_3965,N_3247);
and U6462 (N_6462,N_3759,N_3436);
xnor U6463 (N_6463,N_4222,N_4571);
and U6464 (N_6464,N_4924,N_2576);
nor U6465 (N_6465,N_4424,N_3362);
or U6466 (N_6466,N_2587,N_3551);
and U6467 (N_6467,N_2860,N_2796);
xnor U6468 (N_6468,N_3012,N_4456);
and U6469 (N_6469,N_3248,N_4350);
xor U6470 (N_6470,N_4503,N_3193);
xor U6471 (N_6471,N_3302,N_4124);
xnor U6472 (N_6472,N_2709,N_3889);
xnor U6473 (N_6473,N_2540,N_4973);
nand U6474 (N_6474,N_4826,N_4572);
nor U6475 (N_6475,N_2851,N_4717);
nor U6476 (N_6476,N_4904,N_4547);
or U6477 (N_6477,N_3452,N_4940);
nand U6478 (N_6478,N_2847,N_4041);
and U6479 (N_6479,N_2703,N_3348);
or U6480 (N_6480,N_4638,N_3762);
and U6481 (N_6481,N_3289,N_4826);
and U6482 (N_6482,N_3798,N_3696);
xnor U6483 (N_6483,N_3696,N_3660);
and U6484 (N_6484,N_3354,N_2966);
nand U6485 (N_6485,N_4880,N_3067);
nor U6486 (N_6486,N_4924,N_3272);
xor U6487 (N_6487,N_3722,N_2919);
and U6488 (N_6488,N_3740,N_4345);
nand U6489 (N_6489,N_3052,N_3938);
or U6490 (N_6490,N_3981,N_4302);
nor U6491 (N_6491,N_4715,N_2872);
or U6492 (N_6492,N_3584,N_4616);
nand U6493 (N_6493,N_3261,N_3523);
xor U6494 (N_6494,N_4767,N_3806);
xnor U6495 (N_6495,N_4145,N_3516);
xor U6496 (N_6496,N_4252,N_4172);
xnor U6497 (N_6497,N_2511,N_2711);
nor U6498 (N_6498,N_3173,N_4762);
nor U6499 (N_6499,N_3884,N_3845);
nand U6500 (N_6500,N_2963,N_2882);
nand U6501 (N_6501,N_4223,N_4510);
and U6502 (N_6502,N_2604,N_3894);
nor U6503 (N_6503,N_3329,N_3191);
or U6504 (N_6504,N_3665,N_4498);
nand U6505 (N_6505,N_3351,N_4495);
and U6506 (N_6506,N_3880,N_3617);
and U6507 (N_6507,N_2780,N_4815);
xor U6508 (N_6508,N_2914,N_3525);
nand U6509 (N_6509,N_4353,N_4940);
and U6510 (N_6510,N_3108,N_3980);
and U6511 (N_6511,N_2608,N_2564);
nand U6512 (N_6512,N_4416,N_2919);
or U6513 (N_6513,N_3962,N_4080);
nand U6514 (N_6514,N_3810,N_4224);
or U6515 (N_6515,N_4149,N_2618);
and U6516 (N_6516,N_4755,N_3163);
xnor U6517 (N_6517,N_2753,N_2920);
nor U6518 (N_6518,N_2940,N_3255);
xnor U6519 (N_6519,N_4026,N_4164);
nor U6520 (N_6520,N_3020,N_4570);
and U6521 (N_6521,N_2881,N_4087);
and U6522 (N_6522,N_3781,N_3923);
and U6523 (N_6523,N_2629,N_3968);
nand U6524 (N_6524,N_4626,N_3943);
or U6525 (N_6525,N_3701,N_3605);
nor U6526 (N_6526,N_3583,N_3752);
or U6527 (N_6527,N_3308,N_4512);
nand U6528 (N_6528,N_4420,N_4387);
xor U6529 (N_6529,N_3435,N_3820);
and U6530 (N_6530,N_3681,N_4333);
and U6531 (N_6531,N_2929,N_4866);
or U6532 (N_6532,N_4206,N_4848);
xor U6533 (N_6533,N_3443,N_3936);
nor U6534 (N_6534,N_4792,N_3955);
nor U6535 (N_6535,N_4808,N_3732);
nor U6536 (N_6536,N_2730,N_3619);
xnor U6537 (N_6537,N_2911,N_4110);
or U6538 (N_6538,N_2885,N_4147);
or U6539 (N_6539,N_3962,N_3951);
nor U6540 (N_6540,N_3528,N_3901);
nand U6541 (N_6541,N_4721,N_3986);
nand U6542 (N_6542,N_2633,N_4638);
or U6543 (N_6543,N_4410,N_2756);
nor U6544 (N_6544,N_3501,N_4171);
xnor U6545 (N_6545,N_3478,N_2851);
xor U6546 (N_6546,N_4224,N_2965);
and U6547 (N_6547,N_4972,N_3512);
and U6548 (N_6548,N_4067,N_4134);
xor U6549 (N_6549,N_2780,N_2916);
nand U6550 (N_6550,N_3668,N_4682);
xnor U6551 (N_6551,N_4977,N_3486);
or U6552 (N_6552,N_4516,N_4702);
xnor U6553 (N_6553,N_3415,N_4800);
and U6554 (N_6554,N_3908,N_2737);
nor U6555 (N_6555,N_4821,N_3981);
or U6556 (N_6556,N_3623,N_4761);
nand U6557 (N_6557,N_3852,N_3484);
nor U6558 (N_6558,N_3000,N_3660);
nand U6559 (N_6559,N_3429,N_3364);
nand U6560 (N_6560,N_3472,N_3534);
xnor U6561 (N_6561,N_4608,N_4989);
or U6562 (N_6562,N_4090,N_4135);
nand U6563 (N_6563,N_3001,N_3384);
or U6564 (N_6564,N_4599,N_4221);
or U6565 (N_6565,N_4994,N_2510);
xor U6566 (N_6566,N_3909,N_2736);
nand U6567 (N_6567,N_4678,N_2806);
nor U6568 (N_6568,N_3719,N_4957);
and U6569 (N_6569,N_2620,N_3835);
nand U6570 (N_6570,N_4815,N_3390);
xor U6571 (N_6571,N_3557,N_3602);
nand U6572 (N_6572,N_2837,N_2750);
or U6573 (N_6573,N_3093,N_2866);
nor U6574 (N_6574,N_4143,N_2812);
and U6575 (N_6575,N_3898,N_4731);
nand U6576 (N_6576,N_3760,N_2780);
xor U6577 (N_6577,N_4771,N_4369);
or U6578 (N_6578,N_3571,N_3121);
and U6579 (N_6579,N_3840,N_2864);
nor U6580 (N_6580,N_3046,N_3833);
xor U6581 (N_6581,N_4163,N_4317);
nor U6582 (N_6582,N_3138,N_3492);
or U6583 (N_6583,N_3804,N_4510);
nand U6584 (N_6584,N_3443,N_4503);
or U6585 (N_6585,N_4847,N_4815);
xnor U6586 (N_6586,N_3485,N_3417);
or U6587 (N_6587,N_4489,N_3471);
xnor U6588 (N_6588,N_3842,N_3767);
or U6589 (N_6589,N_3372,N_3319);
and U6590 (N_6590,N_4794,N_3112);
or U6591 (N_6591,N_2910,N_2694);
or U6592 (N_6592,N_4569,N_4051);
xor U6593 (N_6593,N_2517,N_4570);
or U6594 (N_6594,N_2721,N_2530);
nand U6595 (N_6595,N_4691,N_4806);
or U6596 (N_6596,N_4706,N_4449);
nor U6597 (N_6597,N_3874,N_3796);
or U6598 (N_6598,N_3291,N_4458);
xor U6599 (N_6599,N_3582,N_2659);
and U6600 (N_6600,N_2715,N_4176);
or U6601 (N_6601,N_4159,N_3921);
and U6602 (N_6602,N_4911,N_2810);
nor U6603 (N_6603,N_2645,N_4634);
or U6604 (N_6604,N_4255,N_4929);
nor U6605 (N_6605,N_3677,N_4269);
nor U6606 (N_6606,N_3321,N_3379);
and U6607 (N_6607,N_3526,N_4745);
or U6608 (N_6608,N_2666,N_4373);
nor U6609 (N_6609,N_3449,N_3844);
or U6610 (N_6610,N_4087,N_4851);
nand U6611 (N_6611,N_3902,N_3789);
xor U6612 (N_6612,N_2781,N_4981);
nand U6613 (N_6613,N_3411,N_4380);
xnor U6614 (N_6614,N_4069,N_3162);
xor U6615 (N_6615,N_2619,N_3951);
nand U6616 (N_6616,N_2505,N_2757);
nand U6617 (N_6617,N_2878,N_4373);
xnor U6618 (N_6618,N_4741,N_4194);
nor U6619 (N_6619,N_2966,N_2666);
and U6620 (N_6620,N_3506,N_3577);
and U6621 (N_6621,N_4547,N_2907);
or U6622 (N_6622,N_4697,N_4904);
or U6623 (N_6623,N_2810,N_3650);
xor U6624 (N_6624,N_4681,N_2829);
xnor U6625 (N_6625,N_2978,N_4731);
nand U6626 (N_6626,N_2996,N_4754);
nor U6627 (N_6627,N_2752,N_2541);
nor U6628 (N_6628,N_3075,N_3040);
nor U6629 (N_6629,N_4662,N_4453);
nand U6630 (N_6630,N_3564,N_3418);
and U6631 (N_6631,N_2662,N_3681);
nor U6632 (N_6632,N_2944,N_3298);
nand U6633 (N_6633,N_2673,N_3909);
and U6634 (N_6634,N_4798,N_4328);
nor U6635 (N_6635,N_4032,N_2952);
nor U6636 (N_6636,N_3607,N_4093);
or U6637 (N_6637,N_4665,N_2962);
nor U6638 (N_6638,N_4198,N_4665);
and U6639 (N_6639,N_3720,N_4315);
nor U6640 (N_6640,N_4603,N_2841);
nand U6641 (N_6641,N_4287,N_3710);
nor U6642 (N_6642,N_3991,N_4284);
and U6643 (N_6643,N_3195,N_3751);
and U6644 (N_6644,N_3120,N_3898);
or U6645 (N_6645,N_3943,N_3935);
nor U6646 (N_6646,N_4272,N_4619);
and U6647 (N_6647,N_4676,N_3385);
and U6648 (N_6648,N_3218,N_3691);
and U6649 (N_6649,N_2891,N_4655);
or U6650 (N_6650,N_3312,N_3729);
nor U6651 (N_6651,N_4811,N_3569);
nand U6652 (N_6652,N_3784,N_4425);
xnor U6653 (N_6653,N_4683,N_4375);
nand U6654 (N_6654,N_4724,N_2710);
and U6655 (N_6655,N_3670,N_3827);
nand U6656 (N_6656,N_2603,N_4138);
nor U6657 (N_6657,N_3372,N_2987);
nor U6658 (N_6658,N_3298,N_4664);
nor U6659 (N_6659,N_3551,N_4231);
nand U6660 (N_6660,N_4312,N_4063);
nor U6661 (N_6661,N_4250,N_4620);
and U6662 (N_6662,N_3018,N_2917);
or U6663 (N_6663,N_4853,N_4119);
and U6664 (N_6664,N_2727,N_4699);
nor U6665 (N_6665,N_4300,N_3123);
nand U6666 (N_6666,N_3237,N_4081);
nor U6667 (N_6667,N_2779,N_4392);
and U6668 (N_6668,N_4317,N_3551);
nor U6669 (N_6669,N_3433,N_2722);
nand U6670 (N_6670,N_4097,N_3670);
xor U6671 (N_6671,N_4891,N_2730);
or U6672 (N_6672,N_4199,N_2690);
nor U6673 (N_6673,N_2506,N_3548);
xor U6674 (N_6674,N_4557,N_3912);
nand U6675 (N_6675,N_2990,N_4616);
nor U6676 (N_6676,N_3585,N_3991);
nor U6677 (N_6677,N_3579,N_4134);
nor U6678 (N_6678,N_3633,N_2841);
nor U6679 (N_6679,N_3200,N_4860);
nor U6680 (N_6680,N_4804,N_4825);
and U6681 (N_6681,N_3973,N_3406);
xor U6682 (N_6682,N_4032,N_4080);
xor U6683 (N_6683,N_4164,N_4653);
or U6684 (N_6684,N_3865,N_3675);
nand U6685 (N_6685,N_2987,N_2771);
xnor U6686 (N_6686,N_4853,N_4762);
nand U6687 (N_6687,N_3320,N_3723);
nor U6688 (N_6688,N_2649,N_3076);
nand U6689 (N_6689,N_4418,N_4536);
and U6690 (N_6690,N_4298,N_3247);
nand U6691 (N_6691,N_4899,N_3151);
nor U6692 (N_6692,N_3789,N_2675);
or U6693 (N_6693,N_4351,N_2959);
and U6694 (N_6694,N_3556,N_3698);
nand U6695 (N_6695,N_4740,N_2704);
and U6696 (N_6696,N_3007,N_4795);
nand U6697 (N_6697,N_4164,N_2501);
nand U6698 (N_6698,N_3461,N_2727);
nand U6699 (N_6699,N_3415,N_2904);
nor U6700 (N_6700,N_2994,N_4859);
nand U6701 (N_6701,N_2714,N_3611);
and U6702 (N_6702,N_3460,N_3614);
nor U6703 (N_6703,N_3139,N_4149);
nand U6704 (N_6704,N_2561,N_2618);
or U6705 (N_6705,N_3296,N_3028);
nand U6706 (N_6706,N_4519,N_4482);
nand U6707 (N_6707,N_2536,N_3126);
and U6708 (N_6708,N_2545,N_4313);
nand U6709 (N_6709,N_3531,N_3102);
or U6710 (N_6710,N_3116,N_3917);
nor U6711 (N_6711,N_4176,N_3221);
nand U6712 (N_6712,N_4493,N_3378);
and U6713 (N_6713,N_3977,N_3435);
and U6714 (N_6714,N_4003,N_3998);
nand U6715 (N_6715,N_3441,N_3098);
or U6716 (N_6716,N_2652,N_4463);
xor U6717 (N_6717,N_4004,N_3790);
or U6718 (N_6718,N_3646,N_4619);
or U6719 (N_6719,N_2641,N_3546);
nor U6720 (N_6720,N_3695,N_3263);
xor U6721 (N_6721,N_4716,N_3831);
xor U6722 (N_6722,N_3141,N_3130);
nor U6723 (N_6723,N_4268,N_4114);
nor U6724 (N_6724,N_4292,N_3775);
nand U6725 (N_6725,N_2630,N_2811);
nand U6726 (N_6726,N_4145,N_4212);
or U6727 (N_6727,N_4725,N_2755);
and U6728 (N_6728,N_4080,N_3037);
nor U6729 (N_6729,N_3109,N_3716);
nor U6730 (N_6730,N_3908,N_2738);
xnor U6731 (N_6731,N_4622,N_4426);
and U6732 (N_6732,N_4880,N_3563);
nand U6733 (N_6733,N_2649,N_3672);
nand U6734 (N_6734,N_4234,N_4243);
nor U6735 (N_6735,N_3629,N_3636);
nand U6736 (N_6736,N_3582,N_4256);
and U6737 (N_6737,N_2505,N_3044);
nor U6738 (N_6738,N_3612,N_4704);
nor U6739 (N_6739,N_2792,N_3133);
nor U6740 (N_6740,N_3690,N_4459);
nand U6741 (N_6741,N_3098,N_4327);
nor U6742 (N_6742,N_3454,N_4665);
nor U6743 (N_6743,N_3114,N_3172);
xnor U6744 (N_6744,N_3983,N_3962);
xor U6745 (N_6745,N_2846,N_4819);
or U6746 (N_6746,N_2690,N_2758);
nand U6747 (N_6747,N_2859,N_4760);
and U6748 (N_6748,N_3236,N_3974);
nor U6749 (N_6749,N_4305,N_2811);
nand U6750 (N_6750,N_4032,N_4582);
or U6751 (N_6751,N_3293,N_3288);
or U6752 (N_6752,N_4893,N_3154);
xnor U6753 (N_6753,N_3824,N_3660);
xor U6754 (N_6754,N_3756,N_3238);
nand U6755 (N_6755,N_3883,N_3313);
and U6756 (N_6756,N_4434,N_4925);
xor U6757 (N_6757,N_4326,N_4134);
or U6758 (N_6758,N_4425,N_3368);
nand U6759 (N_6759,N_3491,N_2747);
xor U6760 (N_6760,N_2934,N_4138);
nor U6761 (N_6761,N_3490,N_2565);
or U6762 (N_6762,N_4314,N_3921);
and U6763 (N_6763,N_2614,N_2738);
and U6764 (N_6764,N_2842,N_3425);
nor U6765 (N_6765,N_3370,N_3458);
nor U6766 (N_6766,N_4199,N_2964);
and U6767 (N_6767,N_3539,N_3248);
xnor U6768 (N_6768,N_3275,N_4222);
xor U6769 (N_6769,N_2537,N_2645);
and U6770 (N_6770,N_3321,N_2981);
nand U6771 (N_6771,N_4460,N_3880);
nor U6772 (N_6772,N_4024,N_3610);
nand U6773 (N_6773,N_2693,N_3618);
or U6774 (N_6774,N_4402,N_3972);
xor U6775 (N_6775,N_4525,N_4922);
or U6776 (N_6776,N_3235,N_2852);
nor U6777 (N_6777,N_2831,N_4543);
nand U6778 (N_6778,N_3549,N_4809);
nor U6779 (N_6779,N_4652,N_3619);
or U6780 (N_6780,N_3879,N_2554);
nor U6781 (N_6781,N_3417,N_4938);
nand U6782 (N_6782,N_3881,N_3234);
xor U6783 (N_6783,N_4672,N_3321);
xor U6784 (N_6784,N_4219,N_3361);
xor U6785 (N_6785,N_4772,N_3323);
and U6786 (N_6786,N_3170,N_3954);
or U6787 (N_6787,N_4995,N_2990);
xnor U6788 (N_6788,N_4247,N_2934);
nor U6789 (N_6789,N_4830,N_4463);
nand U6790 (N_6790,N_2541,N_3318);
nand U6791 (N_6791,N_3986,N_2579);
nor U6792 (N_6792,N_3441,N_2832);
xnor U6793 (N_6793,N_3016,N_4638);
nor U6794 (N_6794,N_4665,N_3113);
nand U6795 (N_6795,N_4108,N_3780);
xor U6796 (N_6796,N_3188,N_2637);
and U6797 (N_6797,N_4114,N_4417);
xnor U6798 (N_6798,N_4569,N_3009);
nand U6799 (N_6799,N_4045,N_4852);
or U6800 (N_6800,N_3295,N_3570);
nor U6801 (N_6801,N_2512,N_3836);
and U6802 (N_6802,N_4481,N_3778);
and U6803 (N_6803,N_3783,N_3211);
xor U6804 (N_6804,N_2633,N_2500);
xnor U6805 (N_6805,N_4154,N_4505);
nor U6806 (N_6806,N_4383,N_2757);
nor U6807 (N_6807,N_2883,N_4735);
nand U6808 (N_6808,N_2755,N_2810);
nor U6809 (N_6809,N_3182,N_3527);
nor U6810 (N_6810,N_4949,N_3337);
nor U6811 (N_6811,N_2774,N_4160);
nand U6812 (N_6812,N_4339,N_4895);
xnor U6813 (N_6813,N_2575,N_4775);
or U6814 (N_6814,N_3719,N_4495);
and U6815 (N_6815,N_4287,N_3751);
xor U6816 (N_6816,N_3928,N_2782);
or U6817 (N_6817,N_3436,N_3587);
and U6818 (N_6818,N_4207,N_3837);
xor U6819 (N_6819,N_3778,N_4240);
xnor U6820 (N_6820,N_3566,N_4411);
or U6821 (N_6821,N_4581,N_3449);
or U6822 (N_6822,N_2956,N_2894);
xnor U6823 (N_6823,N_3036,N_3742);
nor U6824 (N_6824,N_4051,N_3868);
nor U6825 (N_6825,N_4968,N_4497);
nor U6826 (N_6826,N_3398,N_3712);
xor U6827 (N_6827,N_4704,N_4758);
and U6828 (N_6828,N_4524,N_4750);
nor U6829 (N_6829,N_2968,N_4947);
or U6830 (N_6830,N_3098,N_4104);
or U6831 (N_6831,N_4952,N_4567);
and U6832 (N_6832,N_3868,N_2944);
xnor U6833 (N_6833,N_4228,N_2508);
and U6834 (N_6834,N_4729,N_4063);
nand U6835 (N_6835,N_3460,N_3754);
xor U6836 (N_6836,N_2955,N_2857);
nand U6837 (N_6837,N_4818,N_4024);
xor U6838 (N_6838,N_2634,N_3344);
nand U6839 (N_6839,N_4805,N_4172);
nand U6840 (N_6840,N_3283,N_3209);
and U6841 (N_6841,N_4975,N_2769);
and U6842 (N_6842,N_3168,N_4322);
or U6843 (N_6843,N_3906,N_2945);
xor U6844 (N_6844,N_3407,N_4515);
and U6845 (N_6845,N_3846,N_2588);
xor U6846 (N_6846,N_4622,N_3295);
and U6847 (N_6847,N_4138,N_3107);
and U6848 (N_6848,N_4699,N_3157);
nand U6849 (N_6849,N_4569,N_3048);
or U6850 (N_6850,N_3399,N_3641);
nor U6851 (N_6851,N_4420,N_3122);
and U6852 (N_6852,N_3339,N_4385);
and U6853 (N_6853,N_3939,N_4422);
nor U6854 (N_6854,N_3665,N_4579);
or U6855 (N_6855,N_4484,N_4241);
nor U6856 (N_6856,N_3459,N_4112);
or U6857 (N_6857,N_4767,N_4117);
xor U6858 (N_6858,N_3751,N_3821);
nand U6859 (N_6859,N_4048,N_4516);
and U6860 (N_6860,N_3195,N_4292);
xor U6861 (N_6861,N_4308,N_3662);
nand U6862 (N_6862,N_4857,N_3307);
nand U6863 (N_6863,N_4250,N_4636);
xnor U6864 (N_6864,N_3957,N_4104);
nand U6865 (N_6865,N_2525,N_2675);
or U6866 (N_6866,N_3645,N_3649);
nor U6867 (N_6867,N_4340,N_2982);
nor U6868 (N_6868,N_3104,N_3369);
nor U6869 (N_6869,N_3323,N_4978);
or U6870 (N_6870,N_3959,N_3533);
nor U6871 (N_6871,N_4830,N_3235);
xor U6872 (N_6872,N_2820,N_3531);
nand U6873 (N_6873,N_4154,N_4207);
nand U6874 (N_6874,N_2820,N_2770);
nand U6875 (N_6875,N_2855,N_3567);
and U6876 (N_6876,N_4692,N_4313);
and U6877 (N_6877,N_3588,N_4222);
nor U6878 (N_6878,N_3070,N_3201);
and U6879 (N_6879,N_4554,N_4047);
or U6880 (N_6880,N_4239,N_2524);
nand U6881 (N_6881,N_3178,N_4934);
nor U6882 (N_6882,N_4397,N_4907);
nand U6883 (N_6883,N_3729,N_3869);
nor U6884 (N_6884,N_4405,N_3617);
xnor U6885 (N_6885,N_3976,N_2958);
nand U6886 (N_6886,N_3327,N_3519);
nor U6887 (N_6887,N_4283,N_3825);
xor U6888 (N_6888,N_3914,N_4636);
and U6889 (N_6889,N_3195,N_3449);
nand U6890 (N_6890,N_3960,N_3586);
and U6891 (N_6891,N_4820,N_4815);
nor U6892 (N_6892,N_2971,N_2550);
nand U6893 (N_6893,N_4728,N_4587);
nand U6894 (N_6894,N_4325,N_4843);
xnor U6895 (N_6895,N_4445,N_2917);
and U6896 (N_6896,N_3821,N_4181);
or U6897 (N_6897,N_4853,N_2726);
nor U6898 (N_6898,N_2940,N_3465);
nor U6899 (N_6899,N_3277,N_4143);
nor U6900 (N_6900,N_3149,N_4719);
nand U6901 (N_6901,N_3905,N_3067);
nand U6902 (N_6902,N_4429,N_2914);
nor U6903 (N_6903,N_4602,N_2786);
or U6904 (N_6904,N_3315,N_4047);
nor U6905 (N_6905,N_3678,N_3275);
nand U6906 (N_6906,N_3437,N_3945);
nor U6907 (N_6907,N_4756,N_4955);
nand U6908 (N_6908,N_3076,N_3905);
and U6909 (N_6909,N_2520,N_4880);
and U6910 (N_6910,N_2585,N_2885);
xnor U6911 (N_6911,N_4975,N_4296);
or U6912 (N_6912,N_3781,N_4270);
nor U6913 (N_6913,N_4699,N_3421);
nor U6914 (N_6914,N_3383,N_4081);
nand U6915 (N_6915,N_4072,N_3085);
nor U6916 (N_6916,N_4043,N_4664);
or U6917 (N_6917,N_4204,N_2639);
xor U6918 (N_6918,N_2652,N_3340);
xor U6919 (N_6919,N_4583,N_3037);
nor U6920 (N_6920,N_3316,N_3841);
nand U6921 (N_6921,N_4078,N_3203);
nand U6922 (N_6922,N_2906,N_3752);
and U6923 (N_6923,N_4375,N_2625);
or U6924 (N_6924,N_3727,N_3598);
nor U6925 (N_6925,N_3938,N_2726);
nand U6926 (N_6926,N_3981,N_3129);
nand U6927 (N_6927,N_3590,N_2916);
or U6928 (N_6928,N_4187,N_4991);
xnor U6929 (N_6929,N_3045,N_4887);
nor U6930 (N_6930,N_3196,N_4216);
or U6931 (N_6931,N_3357,N_4399);
and U6932 (N_6932,N_4032,N_4549);
and U6933 (N_6933,N_3609,N_4620);
nand U6934 (N_6934,N_4230,N_3326);
nand U6935 (N_6935,N_4289,N_4347);
nor U6936 (N_6936,N_3702,N_4602);
and U6937 (N_6937,N_2632,N_3599);
nand U6938 (N_6938,N_3593,N_4735);
nand U6939 (N_6939,N_3611,N_3267);
nor U6940 (N_6940,N_3138,N_2652);
and U6941 (N_6941,N_4417,N_4186);
or U6942 (N_6942,N_3209,N_4426);
or U6943 (N_6943,N_3589,N_3080);
and U6944 (N_6944,N_4300,N_3346);
nand U6945 (N_6945,N_4760,N_3591);
nor U6946 (N_6946,N_2727,N_3395);
or U6947 (N_6947,N_3274,N_4621);
xor U6948 (N_6948,N_3036,N_3303);
nand U6949 (N_6949,N_2984,N_3351);
nand U6950 (N_6950,N_3410,N_3879);
xor U6951 (N_6951,N_3136,N_3210);
and U6952 (N_6952,N_3627,N_4988);
nor U6953 (N_6953,N_4235,N_4247);
xnor U6954 (N_6954,N_3771,N_3645);
xor U6955 (N_6955,N_3301,N_4512);
xor U6956 (N_6956,N_4026,N_4002);
and U6957 (N_6957,N_3227,N_4667);
nand U6958 (N_6958,N_2933,N_2784);
nand U6959 (N_6959,N_3026,N_3622);
nand U6960 (N_6960,N_4764,N_3982);
or U6961 (N_6961,N_4021,N_3846);
xnor U6962 (N_6962,N_4531,N_2749);
nor U6963 (N_6963,N_4094,N_3943);
nor U6964 (N_6964,N_4410,N_3304);
xnor U6965 (N_6965,N_3931,N_4962);
or U6966 (N_6966,N_4069,N_4368);
xnor U6967 (N_6967,N_3282,N_2788);
and U6968 (N_6968,N_3503,N_4571);
or U6969 (N_6969,N_4790,N_3650);
nor U6970 (N_6970,N_3735,N_4609);
xor U6971 (N_6971,N_4619,N_3030);
or U6972 (N_6972,N_4678,N_4992);
nor U6973 (N_6973,N_2929,N_4894);
and U6974 (N_6974,N_2584,N_4441);
xor U6975 (N_6975,N_4990,N_3209);
xnor U6976 (N_6976,N_3549,N_4627);
and U6977 (N_6977,N_3280,N_4386);
nand U6978 (N_6978,N_3185,N_4427);
or U6979 (N_6979,N_4557,N_4631);
and U6980 (N_6980,N_4730,N_3032);
xnor U6981 (N_6981,N_3780,N_4139);
nor U6982 (N_6982,N_4911,N_4729);
nand U6983 (N_6983,N_2553,N_4788);
xnor U6984 (N_6984,N_3975,N_2963);
and U6985 (N_6985,N_3258,N_3039);
nor U6986 (N_6986,N_3051,N_3703);
nand U6987 (N_6987,N_3375,N_3520);
nor U6988 (N_6988,N_4501,N_2714);
or U6989 (N_6989,N_2788,N_3888);
and U6990 (N_6990,N_4140,N_3260);
nand U6991 (N_6991,N_3841,N_2961);
nor U6992 (N_6992,N_3117,N_3483);
xnor U6993 (N_6993,N_4886,N_3163);
xnor U6994 (N_6994,N_4244,N_3852);
nand U6995 (N_6995,N_4120,N_4476);
nor U6996 (N_6996,N_2890,N_2505);
or U6997 (N_6997,N_4007,N_4639);
nor U6998 (N_6998,N_4163,N_4532);
or U6999 (N_6999,N_4002,N_2565);
or U7000 (N_7000,N_3309,N_2800);
or U7001 (N_7001,N_2788,N_4800);
or U7002 (N_7002,N_3026,N_4306);
nand U7003 (N_7003,N_3653,N_4345);
xor U7004 (N_7004,N_3114,N_4168);
nor U7005 (N_7005,N_3658,N_3133);
or U7006 (N_7006,N_4598,N_4174);
xnor U7007 (N_7007,N_3674,N_2693);
or U7008 (N_7008,N_2665,N_2561);
and U7009 (N_7009,N_2890,N_4750);
or U7010 (N_7010,N_4734,N_4203);
nand U7011 (N_7011,N_4071,N_3928);
nand U7012 (N_7012,N_4814,N_4172);
or U7013 (N_7013,N_4898,N_3933);
or U7014 (N_7014,N_3153,N_4810);
or U7015 (N_7015,N_4631,N_4866);
xor U7016 (N_7016,N_3080,N_3377);
nor U7017 (N_7017,N_3180,N_3659);
nor U7018 (N_7018,N_4250,N_3991);
nor U7019 (N_7019,N_3730,N_4624);
and U7020 (N_7020,N_3726,N_4232);
and U7021 (N_7021,N_4707,N_2907);
nor U7022 (N_7022,N_3911,N_3672);
or U7023 (N_7023,N_3389,N_4638);
or U7024 (N_7024,N_3593,N_4417);
xnor U7025 (N_7025,N_4335,N_3634);
or U7026 (N_7026,N_4688,N_3226);
or U7027 (N_7027,N_4066,N_3342);
xnor U7028 (N_7028,N_2778,N_3114);
xor U7029 (N_7029,N_4043,N_3767);
xnor U7030 (N_7030,N_4333,N_3724);
and U7031 (N_7031,N_3582,N_3987);
nor U7032 (N_7032,N_3221,N_3372);
and U7033 (N_7033,N_2637,N_2942);
xnor U7034 (N_7034,N_3305,N_3208);
or U7035 (N_7035,N_3754,N_2798);
and U7036 (N_7036,N_3102,N_4860);
or U7037 (N_7037,N_3770,N_4951);
nor U7038 (N_7038,N_2657,N_4431);
nand U7039 (N_7039,N_4339,N_2516);
xor U7040 (N_7040,N_3125,N_3342);
nor U7041 (N_7041,N_4081,N_3181);
xnor U7042 (N_7042,N_3532,N_4045);
or U7043 (N_7043,N_2549,N_4465);
or U7044 (N_7044,N_3869,N_4453);
or U7045 (N_7045,N_4818,N_4183);
nor U7046 (N_7046,N_2760,N_4265);
or U7047 (N_7047,N_3643,N_4830);
nor U7048 (N_7048,N_4650,N_3195);
nand U7049 (N_7049,N_4733,N_2790);
nand U7050 (N_7050,N_4586,N_4423);
nor U7051 (N_7051,N_4637,N_3359);
xor U7052 (N_7052,N_2666,N_3195);
nor U7053 (N_7053,N_3506,N_3923);
xnor U7054 (N_7054,N_4380,N_3739);
nand U7055 (N_7055,N_4456,N_3240);
xor U7056 (N_7056,N_2625,N_3850);
or U7057 (N_7057,N_4388,N_4574);
nor U7058 (N_7058,N_4971,N_3821);
and U7059 (N_7059,N_4239,N_3105);
nand U7060 (N_7060,N_4293,N_2519);
nor U7061 (N_7061,N_2515,N_4878);
nand U7062 (N_7062,N_4773,N_4857);
nor U7063 (N_7063,N_2559,N_3938);
xor U7064 (N_7064,N_3871,N_3298);
and U7065 (N_7065,N_2734,N_4566);
nand U7066 (N_7066,N_3949,N_3298);
nor U7067 (N_7067,N_4468,N_3586);
and U7068 (N_7068,N_3649,N_3848);
and U7069 (N_7069,N_2868,N_2730);
nor U7070 (N_7070,N_3514,N_4040);
nor U7071 (N_7071,N_3155,N_2699);
xnor U7072 (N_7072,N_4456,N_3506);
nand U7073 (N_7073,N_2641,N_4852);
or U7074 (N_7074,N_4536,N_3075);
or U7075 (N_7075,N_4533,N_3647);
nand U7076 (N_7076,N_3353,N_3599);
nand U7077 (N_7077,N_4605,N_4368);
nor U7078 (N_7078,N_4328,N_4715);
and U7079 (N_7079,N_3993,N_3780);
xnor U7080 (N_7080,N_3060,N_2524);
nand U7081 (N_7081,N_4305,N_3747);
nor U7082 (N_7082,N_4660,N_4611);
nand U7083 (N_7083,N_3835,N_3236);
or U7084 (N_7084,N_4874,N_3504);
or U7085 (N_7085,N_4750,N_4202);
or U7086 (N_7086,N_2656,N_4965);
or U7087 (N_7087,N_4626,N_4340);
nand U7088 (N_7088,N_3459,N_4386);
or U7089 (N_7089,N_4235,N_4157);
nand U7090 (N_7090,N_3910,N_4523);
and U7091 (N_7091,N_3255,N_4621);
nand U7092 (N_7092,N_3116,N_3440);
nand U7093 (N_7093,N_2943,N_3399);
or U7094 (N_7094,N_2506,N_2521);
nor U7095 (N_7095,N_4437,N_3232);
nor U7096 (N_7096,N_3993,N_4342);
nor U7097 (N_7097,N_3241,N_3356);
nor U7098 (N_7098,N_2505,N_2855);
or U7099 (N_7099,N_4915,N_3110);
and U7100 (N_7100,N_4704,N_3593);
nor U7101 (N_7101,N_3056,N_3303);
nand U7102 (N_7102,N_3316,N_4196);
nand U7103 (N_7103,N_4833,N_3116);
nand U7104 (N_7104,N_3864,N_3423);
or U7105 (N_7105,N_4354,N_2788);
nand U7106 (N_7106,N_3943,N_3876);
and U7107 (N_7107,N_3901,N_4398);
xor U7108 (N_7108,N_4554,N_3229);
xnor U7109 (N_7109,N_4431,N_2817);
nor U7110 (N_7110,N_4969,N_2721);
nor U7111 (N_7111,N_3853,N_3960);
nor U7112 (N_7112,N_4936,N_4692);
nand U7113 (N_7113,N_3255,N_3426);
nor U7114 (N_7114,N_4428,N_4365);
nor U7115 (N_7115,N_3732,N_3320);
xor U7116 (N_7116,N_4466,N_2889);
xor U7117 (N_7117,N_4779,N_3994);
nor U7118 (N_7118,N_4560,N_3225);
nand U7119 (N_7119,N_4279,N_2543);
nand U7120 (N_7120,N_4886,N_3288);
nor U7121 (N_7121,N_3844,N_2816);
xnor U7122 (N_7122,N_3226,N_3585);
nand U7123 (N_7123,N_4907,N_4518);
xor U7124 (N_7124,N_2845,N_4237);
nand U7125 (N_7125,N_4582,N_3216);
nand U7126 (N_7126,N_4413,N_2533);
nand U7127 (N_7127,N_4451,N_3488);
nand U7128 (N_7128,N_3408,N_4249);
nor U7129 (N_7129,N_2768,N_2787);
xnor U7130 (N_7130,N_4274,N_2670);
nor U7131 (N_7131,N_3629,N_3624);
nor U7132 (N_7132,N_3471,N_2668);
xor U7133 (N_7133,N_2793,N_3029);
xnor U7134 (N_7134,N_4268,N_4108);
xor U7135 (N_7135,N_3711,N_2940);
xnor U7136 (N_7136,N_4015,N_4149);
xnor U7137 (N_7137,N_2891,N_3136);
nand U7138 (N_7138,N_4042,N_4192);
or U7139 (N_7139,N_3180,N_4395);
nor U7140 (N_7140,N_3547,N_3045);
nand U7141 (N_7141,N_3024,N_2567);
or U7142 (N_7142,N_3996,N_4947);
xnor U7143 (N_7143,N_4434,N_3994);
or U7144 (N_7144,N_4912,N_3950);
nand U7145 (N_7145,N_3660,N_2875);
xnor U7146 (N_7146,N_4891,N_4167);
nand U7147 (N_7147,N_2854,N_4541);
nor U7148 (N_7148,N_4060,N_4742);
nand U7149 (N_7149,N_3604,N_3017);
nor U7150 (N_7150,N_4634,N_2510);
xnor U7151 (N_7151,N_3253,N_4180);
or U7152 (N_7152,N_4482,N_4198);
nor U7153 (N_7153,N_3292,N_4119);
xnor U7154 (N_7154,N_3927,N_4318);
xnor U7155 (N_7155,N_4283,N_2847);
and U7156 (N_7156,N_4946,N_4054);
nor U7157 (N_7157,N_2712,N_4985);
and U7158 (N_7158,N_4440,N_3134);
nor U7159 (N_7159,N_2802,N_2996);
xor U7160 (N_7160,N_2583,N_4908);
or U7161 (N_7161,N_3702,N_3657);
nand U7162 (N_7162,N_2682,N_2557);
xor U7163 (N_7163,N_3149,N_3988);
and U7164 (N_7164,N_4892,N_2948);
nor U7165 (N_7165,N_3941,N_4719);
nor U7166 (N_7166,N_4419,N_3469);
or U7167 (N_7167,N_4968,N_3983);
or U7168 (N_7168,N_2991,N_2583);
xor U7169 (N_7169,N_4050,N_4440);
xor U7170 (N_7170,N_2665,N_4468);
and U7171 (N_7171,N_2796,N_4948);
or U7172 (N_7172,N_4537,N_4510);
and U7173 (N_7173,N_3490,N_4385);
or U7174 (N_7174,N_3535,N_2618);
or U7175 (N_7175,N_3552,N_2790);
nor U7176 (N_7176,N_4781,N_3774);
xnor U7177 (N_7177,N_3070,N_3153);
or U7178 (N_7178,N_4114,N_3963);
and U7179 (N_7179,N_3930,N_2793);
or U7180 (N_7180,N_3122,N_4398);
nand U7181 (N_7181,N_2566,N_4993);
xor U7182 (N_7182,N_2877,N_3105);
and U7183 (N_7183,N_4110,N_2500);
nor U7184 (N_7184,N_4881,N_3251);
nor U7185 (N_7185,N_3070,N_4176);
nor U7186 (N_7186,N_4588,N_3560);
and U7187 (N_7187,N_3494,N_4528);
nand U7188 (N_7188,N_3581,N_2567);
xor U7189 (N_7189,N_2957,N_2586);
nor U7190 (N_7190,N_3837,N_4293);
and U7191 (N_7191,N_3273,N_4316);
nand U7192 (N_7192,N_3983,N_2747);
nor U7193 (N_7193,N_3741,N_4531);
and U7194 (N_7194,N_4672,N_3680);
nand U7195 (N_7195,N_3296,N_4565);
nand U7196 (N_7196,N_4014,N_4004);
and U7197 (N_7197,N_2712,N_4982);
xor U7198 (N_7198,N_4109,N_4182);
or U7199 (N_7199,N_4107,N_3267);
nand U7200 (N_7200,N_2773,N_4652);
or U7201 (N_7201,N_4837,N_4361);
nand U7202 (N_7202,N_3747,N_3682);
or U7203 (N_7203,N_4169,N_4146);
nand U7204 (N_7204,N_3881,N_3404);
nor U7205 (N_7205,N_3984,N_3326);
nor U7206 (N_7206,N_3581,N_4597);
or U7207 (N_7207,N_4090,N_2771);
nand U7208 (N_7208,N_3868,N_3351);
and U7209 (N_7209,N_4677,N_3416);
nor U7210 (N_7210,N_4551,N_4659);
nand U7211 (N_7211,N_4935,N_3764);
nor U7212 (N_7212,N_3300,N_4850);
or U7213 (N_7213,N_3975,N_4038);
xor U7214 (N_7214,N_2846,N_3697);
nand U7215 (N_7215,N_3654,N_3018);
or U7216 (N_7216,N_4691,N_3198);
and U7217 (N_7217,N_2504,N_2512);
nand U7218 (N_7218,N_4303,N_3652);
nor U7219 (N_7219,N_3148,N_4788);
nor U7220 (N_7220,N_3832,N_3055);
or U7221 (N_7221,N_3312,N_2585);
xnor U7222 (N_7222,N_3542,N_2998);
xor U7223 (N_7223,N_4882,N_4123);
xnor U7224 (N_7224,N_4804,N_4923);
or U7225 (N_7225,N_2798,N_4312);
or U7226 (N_7226,N_4807,N_3088);
nor U7227 (N_7227,N_4606,N_2806);
or U7228 (N_7228,N_4565,N_4957);
xnor U7229 (N_7229,N_3848,N_4918);
xor U7230 (N_7230,N_4410,N_3905);
nor U7231 (N_7231,N_4426,N_3029);
nor U7232 (N_7232,N_4990,N_4498);
and U7233 (N_7233,N_4245,N_3953);
xor U7234 (N_7234,N_4361,N_4277);
nor U7235 (N_7235,N_3792,N_4228);
xnor U7236 (N_7236,N_3303,N_4349);
nand U7237 (N_7237,N_4392,N_3524);
and U7238 (N_7238,N_3722,N_4610);
nor U7239 (N_7239,N_2665,N_3440);
nand U7240 (N_7240,N_4736,N_2668);
nand U7241 (N_7241,N_4754,N_2786);
and U7242 (N_7242,N_2813,N_3243);
nor U7243 (N_7243,N_3278,N_3628);
and U7244 (N_7244,N_4011,N_3023);
nand U7245 (N_7245,N_2576,N_4320);
nand U7246 (N_7246,N_4180,N_3661);
or U7247 (N_7247,N_3220,N_4195);
nand U7248 (N_7248,N_4522,N_2618);
or U7249 (N_7249,N_3523,N_4591);
or U7250 (N_7250,N_2904,N_3985);
nor U7251 (N_7251,N_3546,N_3838);
and U7252 (N_7252,N_4581,N_4650);
and U7253 (N_7253,N_4891,N_3378);
and U7254 (N_7254,N_3864,N_3964);
and U7255 (N_7255,N_4741,N_3959);
or U7256 (N_7256,N_3160,N_3356);
and U7257 (N_7257,N_4861,N_3461);
nor U7258 (N_7258,N_2855,N_2542);
or U7259 (N_7259,N_2858,N_4172);
or U7260 (N_7260,N_4215,N_3476);
nor U7261 (N_7261,N_4089,N_3157);
nor U7262 (N_7262,N_2544,N_3623);
xor U7263 (N_7263,N_2516,N_3831);
nand U7264 (N_7264,N_4609,N_4635);
nor U7265 (N_7265,N_3979,N_3843);
xor U7266 (N_7266,N_2640,N_3113);
nor U7267 (N_7267,N_2638,N_3324);
and U7268 (N_7268,N_4729,N_2909);
nand U7269 (N_7269,N_2656,N_3905);
xnor U7270 (N_7270,N_2549,N_2626);
nand U7271 (N_7271,N_4874,N_3496);
xnor U7272 (N_7272,N_4709,N_2598);
nor U7273 (N_7273,N_2518,N_2568);
xor U7274 (N_7274,N_2841,N_3760);
nand U7275 (N_7275,N_4593,N_2997);
nand U7276 (N_7276,N_4755,N_4914);
nor U7277 (N_7277,N_4794,N_4275);
or U7278 (N_7278,N_3354,N_3227);
nor U7279 (N_7279,N_4454,N_2662);
nand U7280 (N_7280,N_3022,N_4178);
xor U7281 (N_7281,N_4794,N_4723);
or U7282 (N_7282,N_3124,N_3729);
xnor U7283 (N_7283,N_3088,N_3922);
xnor U7284 (N_7284,N_4916,N_4197);
nand U7285 (N_7285,N_3494,N_3625);
nand U7286 (N_7286,N_3425,N_2530);
nand U7287 (N_7287,N_2533,N_3622);
xnor U7288 (N_7288,N_3821,N_3822);
xnor U7289 (N_7289,N_4098,N_4645);
or U7290 (N_7290,N_3300,N_4379);
xor U7291 (N_7291,N_3335,N_3847);
nor U7292 (N_7292,N_2908,N_3959);
or U7293 (N_7293,N_3972,N_4315);
nor U7294 (N_7294,N_3801,N_4983);
or U7295 (N_7295,N_3345,N_3650);
or U7296 (N_7296,N_3552,N_4381);
xnor U7297 (N_7297,N_3681,N_4765);
and U7298 (N_7298,N_3732,N_4439);
xnor U7299 (N_7299,N_4614,N_3221);
nand U7300 (N_7300,N_3656,N_3283);
xnor U7301 (N_7301,N_2700,N_4055);
or U7302 (N_7302,N_2678,N_2530);
and U7303 (N_7303,N_4829,N_2897);
xor U7304 (N_7304,N_2607,N_3655);
and U7305 (N_7305,N_2559,N_3214);
nand U7306 (N_7306,N_2789,N_3287);
nor U7307 (N_7307,N_3529,N_2906);
nor U7308 (N_7308,N_3359,N_4994);
or U7309 (N_7309,N_3647,N_3939);
nand U7310 (N_7310,N_4083,N_2904);
nor U7311 (N_7311,N_3886,N_3231);
nand U7312 (N_7312,N_3788,N_4532);
xnor U7313 (N_7313,N_4828,N_4716);
nand U7314 (N_7314,N_2981,N_2870);
nand U7315 (N_7315,N_4417,N_4906);
nor U7316 (N_7316,N_3916,N_3321);
xor U7317 (N_7317,N_2977,N_3050);
and U7318 (N_7318,N_4640,N_3588);
xnor U7319 (N_7319,N_2982,N_3083);
or U7320 (N_7320,N_3907,N_2919);
or U7321 (N_7321,N_2924,N_3464);
nand U7322 (N_7322,N_3229,N_2958);
xor U7323 (N_7323,N_3273,N_3847);
xnor U7324 (N_7324,N_2513,N_4542);
nand U7325 (N_7325,N_2846,N_3542);
nor U7326 (N_7326,N_3554,N_3851);
nand U7327 (N_7327,N_3585,N_3224);
or U7328 (N_7328,N_4563,N_3187);
nand U7329 (N_7329,N_3905,N_3370);
and U7330 (N_7330,N_2621,N_4778);
or U7331 (N_7331,N_4702,N_3486);
nand U7332 (N_7332,N_4704,N_4100);
nor U7333 (N_7333,N_2890,N_4965);
nand U7334 (N_7334,N_2528,N_2759);
xor U7335 (N_7335,N_4999,N_3805);
xor U7336 (N_7336,N_3185,N_3695);
or U7337 (N_7337,N_4679,N_2641);
nand U7338 (N_7338,N_4654,N_4377);
nand U7339 (N_7339,N_3147,N_3257);
nand U7340 (N_7340,N_4734,N_4900);
nand U7341 (N_7341,N_3698,N_3648);
xnor U7342 (N_7342,N_2730,N_3505);
nand U7343 (N_7343,N_4680,N_4541);
xnor U7344 (N_7344,N_3347,N_3567);
nor U7345 (N_7345,N_2535,N_4361);
xnor U7346 (N_7346,N_4474,N_4160);
xnor U7347 (N_7347,N_3180,N_3412);
and U7348 (N_7348,N_3950,N_4950);
or U7349 (N_7349,N_4575,N_3701);
and U7350 (N_7350,N_4483,N_4156);
or U7351 (N_7351,N_3488,N_3744);
xnor U7352 (N_7352,N_3649,N_3661);
nand U7353 (N_7353,N_3361,N_4563);
or U7354 (N_7354,N_3523,N_4734);
nand U7355 (N_7355,N_4648,N_3151);
or U7356 (N_7356,N_3420,N_2621);
nand U7357 (N_7357,N_3678,N_4697);
or U7358 (N_7358,N_3416,N_4383);
or U7359 (N_7359,N_2652,N_4345);
nand U7360 (N_7360,N_3196,N_4764);
xor U7361 (N_7361,N_4233,N_3465);
nand U7362 (N_7362,N_4858,N_3705);
xor U7363 (N_7363,N_3278,N_4488);
and U7364 (N_7364,N_4066,N_3529);
and U7365 (N_7365,N_3533,N_2925);
nand U7366 (N_7366,N_4848,N_4491);
nand U7367 (N_7367,N_3335,N_4023);
xnor U7368 (N_7368,N_3324,N_4709);
nor U7369 (N_7369,N_4895,N_3030);
nor U7370 (N_7370,N_4204,N_4860);
nor U7371 (N_7371,N_3171,N_3795);
xor U7372 (N_7372,N_3226,N_4268);
or U7373 (N_7373,N_4701,N_4661);
or U7374 (N_7374,N_4382,N_4921);
and U7375 (N_7375,N_3751,N_2979);
nor U7376 (N_7376,N_4984,N_2905);
or U7377 (N_7377,N_3545,N_2939);
xor U7378 (N_7378,N_4314,N_4461);
and U7379 (N_7379,N_4750,N_2822);
xor U7380 (N_7380,N_3486,N_3809);
nor U7381 (N_7381,N_3911,N_4659);
and U7382 (N_7382,N_2958,N_4551);
xor U7383 (N_7383,N_3122,N_3921);
xor U7384 (N_7384,N_3961,N_4019);
nand U7385 (N_7385,N_2766,N_4804);
nand U7386 (N_7386,N_3244,N_3012);
nor U7387 (N_7387,N_3442,N_3572);
nand U7388 (N_7388,N_2805,N_2728);
nand U7389 (N_7389,N_4198,N_4398);
nand U7390 (N_7390,N_3125,N_4871);
or U7391 (N_7391,N_3250,N_3767);
nand U7392 (N_7392,N_4368,N_2586);
nand U7393 (N_7393,N_4063,N_2918);
nor U7394 (N_7394,N_4967,N_4856);
nand U7395 (N_7395,N_2887,N_4681);
xnor U7396 (N_7396,N_4346,N_4177);
nor U7397 (N_7397,N_3338,N_4593);
or U7398 (N_7398,N_3905,N_3467);
nand U7399 (N_7399,N_3860,N_3539);
and U7400 (N_7400,N_3337,N_2898);
and U7401 (N_7401,N_4284,N_3999);
and U7402 (N_7402,N_4786,N_3758);
and U7403 (N_7403,N_3923,N_2693);
nor U7404 (N_7404,N_2927,N_3001);
and U7405 (N_7405,N_3583,N_4700);
or U7406 (N_7406,N_2930,N_2571);
nand U7407 (N_7407,N_4213,N_2678);
xnor U7408 (N_7408,N_2998,N_2987);
and U7409 (N_7409,N_4026,N_2660);
or U7410 (N_7410,N_2605,N_2979);
nor U7411 (N_7411,N_3978,N_2991);
or U7412 (N_7412,N_3391,N_4521);
xnor U7413 (N_7413,N_2588,N_4754);
or U7414 (N_7414,N_2804,N_3432);
nor U7415 (N_7415,N_4371,N_3100);
and U7416 (N_7416,N_4454,N_4528);
and U7417 (N_7417,N_4026,N_4582);
xnor U7418 (N_7418,N_2766,N_4826);
xor U7419 (N_7419,N_2896,N_3446);
nand U7420 (N_7420,N_4743,N_3238);
and U7421 (N_7421,N_2826,N_4586);
nor U7422 (N_7422,N_3496,N_3178);
nor U7423 (N_7423,N_3197,N_4083);
xnor U7424 (N_7424,N_3323,N_4650);
and U7425 (N_7425,N_3722,N_4439);
nor U7426 (N_7426,N_3439,N_2813);
and U7427 (N_7427,N_3546,N_3381);
or U7428 (N_7428,N_2917,N_2849);
or U7429 (N_7429,N_3968,N_2774);
nand U7430 (N_7430,N_2842,N_4468);
nand U7431 (N_7431,N_3232,N_3115);
xor U7432 (N_7432,N_4830,N_3836);
or U7433 (N_7433,N_4407,N_4954);
xnor U7434 (N_7434,N_2849,N_2913);
and U7435 (N_7435,N_3852,N_2578);
xor U7436 (N_7436,N_2615,N_3632);
xnor U7437 (N_7437,N_4126,N_2940);
nand U7438 (N_7438,N_2511,N_3219);
xnor U7439 (N_7439,N_2894,N_3427);
or U7440 (N_7440,N_3922,N_4748);
and U7441 (N_7441,N_3364,N_4973);
xor U7442 (N_7442,N_3935,N_3023);
xor U7443 (N_7443,N_4557,N_4619);
and U7444 (N_7444,N_4847,N_3913);
nand U7445 (N_7445,N_3519,N_3207);
xnor U7446 (N_7446,N_3275,N_2984);
nand U7447 (N_7447,N_2848,N_4326);
nor U7448 (N_7448,N_4283,N_4021);
nor U7449 (N_7449,N_4370,N_3495);
nand U7450 (N_7450,N_3839,N_4002);
nor U7451 (N_7451,N_2706,N_3592);
nand U7452 (N_7452,N_4472,N_4530);
nand U7453 (N_7453,N_4555,N_2748);
and U7454 (N_7454,N_3544,N_3505);
nand U7455 (N_7455,N_4814,N_3830);
nand U7456 (N_7456,N_2557,N_4893);
and U7457 (N_7457,N_3557,N_4475);
nor U7458 (N_7458,N_2872,N_3311);
nand U7459 (N_7459,N_4905,N_4008);
and U7460 (N_7460,N_3870,N_2629);
nand U7461 (N_7461,N_3452,N_4564);
or U7462 (N_7462,N_3083,N_4324);
nor U7463 (N_7463,N_2555,N_4832);
nor U7464 (N_7464,N_3680,N_3856);
nand U7465 (N_7465,N_3573,N_4939);
or U7466 (N_7466,N_3445,N_2543);
or U7467 (N_7467,N_2624,N_4892);
nor U7468 (N_7468,N_4095,N_3702);
nand U7469 (N_7469,N_4432,N_2935);
nor U7470 (N_7470,N_3602,N_3087);
xnor U7471 (N_7471,N_4773,N_4718);
and U7472 (N_7472,N_3066,N_4425);
or U7473 (N_7473,N_4794,N_4263);
or U7474 (N_7474,N_3741,N_3506);
and U7475 (N_7475,N_3210,N_2693);
or U7476 (N_7476,N_4588,N_4630);
nand U7477 (N_7477,N_4768,N_4664);
and U7478 (N_7478,N_4125,N_4515);
nor U7479 (N_7479,N_4579,N_4411);
nor U7480 (N_7480,N_2616,N_3090);
xor U7481 (N_7481,N_3247,N_3643);
xor U7482 (N_7482,N_2566,N_4917);
nor U7483 (N_7483,N_4044,N_3200);
xor U7484 (N_7484,N_4607,N_2877);
nor U7485 (N_7485,N_4957,N_2924);
nand U7486 (N_7486,N_2685,N_3020);
xnor U7487 (N_7487,N_4398,N_4025);
or U7488 (N_7488,N_4249,N_3131);
nor U7489 (N_7489,N_4549,N_4136);
or U7490 (N_7490,N_3883,N_3851);
or U7491 (N_7491,N_3461,N_2720);
and U7492 (N_7492,N_3715,N_2562);
and U7493 (N_7493,N_4050,N_4232);
nand U7494 (N_7494,N_2991,N_3021);
and U7495 (N_7495,N_2853,N_3425);
and U7496 (N_7496,N_4988,N_3208);
xor U7497 (N_7497,N_3373,N_3573);
xnor U7498 (N_7498,N_4705,N_4133);
or U7499 (N_7499,N_4861,N_3882);
nand U7500 (N_7500,N_6823,N_5499);
xor U7501 (N_7501,N_7284,N_5598);
nor U7502 (N_7502,N_6945,N_6999);
xor U7503 (N_7503,N_7375,N_5145);
xnor U7504 (N_7504,N_6644,N_7382);
xnor U7505 (N_7505,N_6726,N_6224);
or U7506 (N_7506,N_7113,N_5975);
or U7507 (N_7507,N_7425,N_5762);
nor U7508 (N_7508,N_5603,N_5847);
nor U7509 (N_7509,N_5819,N_6091);
and U7510 (N_7510,N_6219,N_7434);
or U7511 (N_7511,N_5522,N_6902);
and U7512 (N_7512,N_5963,N_6266);
and U7513 (N_7513,N_6829,N_6756);
nand U7514 (N_7514,N_6708,N_6666);
nand U7515 (N_7515,N_7321,N_7151);
xnor U7516 (N_7516,N_6861,N_6425);
nand U7517 (N_7517,N_6342,N_7359);
xnor U7518 (N_7518,N_7015,N_6865);
or U7519 (N_7519,N_7097,N_6007);
nor U7520 (N_7520,N_5584,N_6156);
or U7521 (N_7521,N_7421,N_5369);
and U7522 (N_7522,N_5310,N_5621);
nor U7523 (N_7523,N_7335,N_5002);
nor U7524 (N_7524,N_7310,N_6080);
or U7525 (N_7525,N_7349,N_5280);
nor U7526 (N_7526,N_5590,N_5570);
nor U7527 (N_7527,N_7183,N_6576);
or U7528 (N_7528,N_5983,N_5639);
nor U7529 (N_7529,N_6888,N_7215);
xnor U7530 (N_7530,N_5944,N_5060);
xnor U7531 (N_7531,N_6974,N_5468);
nand U7532 (N_7532,N_5970,N_7378);
nand U7533 (N_7533,N_5136,N_6258);
or U7534 (N_7534,N_6282,N_5913);
and U7535 (N_7535,N_5801,N_6131);
and U7536 (N_7536,N_6641,N_5740);
and U7537 (N_7537,N_7412,N_6728);
and U7538 (N_7538,N_7338,N_6042);
or U7539 (N_7539,N_6114,N_6142);
and U7540 (N_7540,N_7405,N_6367);
or U7541 (N_7541,N_7307,N_6349);
xnor U7542 (N_7542,N_7363,N_5853);
xnor U7543 (N_7543,N_6578,N_6087);
or U7544 (N_7544,N_6068,N_5936);
or U7545 (N_7545,N_7174,N_5231);
nor U7546 (N_7546,N_6260,N_6281);
nor U7547 (N_7547,N_5770,N_7316);
xnor U7548 (N_7548,N_6365,N_5390);
xor U7549 (N_7549,N_5290,N_6388);
nor U7550 (N_7550,N_5174,N_7201);
nor U7551 (N_7551,N_6181,N_6274);
or U7552 (N_7552,N_7288,N_6261);
nor U7553 (N_7553,N_7271,N_7318);
or U7554 (N_7554,N_7132,N_5079);
nor U7555 (N_7555,N_5443,N_7331);
xor U7556 (N_7556,N_5547,N_6444);
nand U7557 (N_7557,N_5964,N_7374);
nand U7558 (N_7558,N_5643,N_5725);
and U7559 (N_7559,N_7320,N_6504);
nor U7560 (N_7560,N_5305,N_6866);
xor U7561 (N_7561,N_6573,N_5010);
xnor U7562 (N_7562,N_7043,N_7061);
nor U7563 (N_7563,N_6216,N_5015);
xnor U7564 (N_7564,N_5815,N_5967);
xor U7565 (N_7565,N_6556,N_6118);
nand U7566 (N_7566,N_5893,N_6703);
nand U7567 (N_7567,N_7041,N_6712);
or U7568 (N_7568,N_5271,N_7393);
nor U7569 (N_7569,N_7030,N_5228);
xnor U7570 (N_7570,N_6093,N_6437);
nor U7571 (N_7571,N_7347,N_5342);
nand U7572 (N_7572,N_5834,N_6533);
nand U7573 (N_7573,N_5566,N_6662);
and U7574 (N_7574,N_6976,N_6668);
nand U7575 (N_7575,N_5057,N_6429);
nand U7576 (N_7576,N_6110,N_7141);
xor U7577 (N_7577,N_6451,N_5044);
xnor U7578 (N_7578,N_5993,N_6789);
nand U7579 (N_7579,N_6783,N_7031);
and U7580 (N_7580,N_7027,N_6496);
and U7581 (N_7581,N_5950,N_6177);
or U7582 (N_7582,N_6881,N_6936);
xor U7583 (N_7583,N_6409,N_6380);
xor U7584 (N_7584,N_5216,N_7042);
nand U7585 (N_7585,N_6286,N_6507);
nand U7586 (N_7586,N_6162,N_6250);
and U7587 (N_7587,N_5012,N_6815);
or U7588 (N_7588,N_7194,N_7229);
nand U7589 (N_7589,N_7419,N_7235);
nand U7590 (N_7590,N_7009,N_7166);
nor U7591 (N_7591,N_7388,N_6706);
nand U7592 (N_7592,N_5262,N_7472);
xnor U7593 (N_7593,N_7244,N_7251);
or U7594 (N_7594,N_6797,N_6534);
nand U7595 (N_7595,N_6996,N_7119);
nor U7596 (N_7596,N_5772,N_7026);
nand U7597 (N_7597,N_7025,N_7280);
and U7598 (N_7598,N_5450,N_6035);
and U7599 (N_7599,N_5997,N_5160);
and U7600 (N_7600,N_6682,N_5794);
or U7601 (N_7601,N_5065,N_7432);
and U7602 (N_7602,N_7088,N_6824);
and U7603 (N_7603,N_5188,N_7357);
and U7604 (N_7604,N_7051,N_6998);
or U7605 (N_7605,N_6084,N_6964);
nor U7606 (N_7606,N_6227,N_6225);
xor U7607 (N_7607,N_5708,N_6715);
nor U7608 (N_7608,N_6746,N_6923);
and U7609 (N_7609,N_6627,N_5317);
nor U7610 (N_7610,N_7392,N_5719);
nand U7611 (N_7611,N_6940,N_6745);
nand U7612 (N_7612,N_7476,N_7301);
and U7613 (N_7613,N_6434,N_5515);
nand U7614 (N_7614,N_5984,N_6914);
or U7615 (N_7615,N_5977,N_6991);
nor U7616 (N_7616,N_5606,N_5969);
xnor U7617 (N_7617,N_5904,N_5124);
nor U7618 (N_7618,N_6691,N_6594);
xor U7619 (N_7619,N_6036,N_7046);
nor U7620 (N_7620,N_7356,N_6382);
nand U7621 (N_7621,N_7152,N_6220);
and U7622 (N_7622,N_5111,N_6344);
and U7623 (N_7623,N_6055,N_5773);
and U7624 (N_7624,N_7184,N_6678);
and U7625 (N_7625,N_6904,N_7397);
or U7626 (N_7626,N_6000,N_5744);
nor U7627 (N_7627,N_6725,N_6518);
xnor U7628 (N_7628,N_6321,N_5750);
or U7629 (N_7629,N_6102,N_5693);
nand U7630 (N_7630,N_6821,N_5557);
nor U7631 (N_7631,N_7367,N_7283);
or U7632 (N_7632,N_6559,N_6587);
xor U7633 (N_7633,N_7002,N_6639);
nand U7634 (N_7634,N_6734,N_7129);
xor U7635 (N_7635,N_5349,N_5956);
nor U7636 (N_7636,N_5597,N_6681);
and U7637 (N_7637,N_7112,N_6279);
nor U7638 (N_7638,N_5264,N_5144);
and U7639 (N_7639,N_6074,N_7422);
nor U7640 (N_7640,N_5883,N_6383);
and U7641 (N_7641,N_6058,N_6887);
nand U7642 (N_7642,N_5143,N_5743);
xnor U7643 (N_7643,N_5704,N_7096);
xor U7644 (N_7644,N_5223,N_6804);
nand U7645 (N_7645,N_5695,N_6626);
xor U7646 (N_7646,N_5863,N_7438);
nor U7647 (N_7647,N_5745,N_6811);
nor U7648 (N_7648,N_7128,N_5045);
xnor U7649 (N_7649,N_7265,N_7380);
nand U7650 (N_7650,N_5282,N_6060);
nor U7651 (N_7651,N_5101,N_5116);
or U7652 (N_7652,N_6188,N_5351);
or U7653 (N_7653,N_6481,N_6730);
and U7654 (N_7654,N_7457,N_5480);
nor U7655 (N_7655,N_5564,N_5764);
nor U7656 (N_7656,N_5700,N_7262);
nor U7657 (N_7657,N_6401,N_6646);
nand U7658 (N_7658,N_5831,N_5582);
xor U7659 (N_7659,N_5540,N_5358);
or U7660 (N_7660,N_7258,N_5865);
xor U7661 (N_7661,N_6871,N_6189);
nand U7662 (N_7662,N_6950,N_6537);
nor U7663 (N_7663,N_6768,N_5238);
xor U7664 (N_7664,N_5097,N_5998);
and U7665 (N_7665,N_7341,N_6128);
or U7666 (N_7666,N_5510,N_5686);
and U7667 (N_7667,N_6906,N_5475);
or U7668 (N_7668,N_6345,N_5813);
and U7669 (N_7669,N_6347,N_6354);
or U7670 (N_7670,N_6479,N_6612);
xor U7671 (N_7671,N_6795,N_5542);
and U7672 (N_7672,N_6047,N_5359);
and U7673 (N_7673,N_6820,N_6879);
nand U7674 (N_7674,N_5363,N_6530);
and U7675 (N_7675,N_5488,N_5901);
and U7676 (N_7676,N_6148,N_6442);
nor U7677 (N_7677,N_7390,N_6526);
xor U7678 (N_7678,N_6422,N_6930);
nor U7679 (N_7679,N_5086,N_5915);
xnor U7680 (N_7680,N_6929,N_5165);
or U7681 (N_7681,N_7093,N_6366);
and U7682 (N_7682,N_6175,N_5472);
and U7683 (N_7683,N_7358,N_6655);
xnor U7684 (N_7684,N_6222,N_5827);
nor U7685 (N_7685,N_5907,N_6385);
xor U7686 (N_7686,N_6984,N_6294);
nand U7687 (N_7687,N_6669,N_7336);
or U7688 (N_7688,N_6043,N_6315);
xnor U7689 (N_7689,N_7297,N_5183);
nand U7690 (N_7690,N_6732,N_6842);
nand U7691 (N_7691,N_5399,N_6375);
or U7692 (N_7692,N_6452,N_5804);
or U7693 (N_7693,N_5434,N_7077);
and U7694 (N_7694,N_6535,N_5020);
and U7695 (N_7695,N_6436,N_7337);
and U7696 (N_7696,N_5255,N_7238);
or U7697 (N_7697,N_6199,N_5298);
or U7698 (N_7698,N_5133,N_5876);
nand U7699 (N_7699,N_5383,N_5114);
nor U7700 (N_7700,N_7186,N_6474);
or U7701 (N_7701,N_7400,N_5022);
nor U7702 (N_7702,N_6073,N_7342);
or U7703 (N_7703,N_5166,N_6650);
nand U7704 (N_7704,N_7450,N_5529);
nor U7705 (N_7705,N_7123,N_6729);
xnor U7706 (N_7706,N_6816,N_6628);
nand U7707 (N_7707,N_6977,N_5947);
nand U7708 (N_7708,N_5805,N_6283);
and U7709 (N_7709,N_7399,N_7437);
or U7710 (N_7710,N_6997,N_5150);
or U7711 (N_7711,N_5954,N_6982);
nand U7712 (N_7712,N_5852,N_7406);
or U7713 (N_7713,N_7106,N_6277);
nand U7714 (N_7714,N_7228,N_7071);
nand U7715 (N_7715,N_7047,N_7279);
or U7716 (N_7716,N_7188,N_5988);
nand U7717 (N_7717,N_7360,N_7257);
xor U7718 (N_7718,N_5927,N_5215);
xnor U7719 (N_7719,N_7298,N_5089);
xnor U7720 (N_7720,N_5925,N_7154);
nor U7721 (N_7721,N_6499,N_5049);
and U7722 (N_7722,N_7190,N_7192);
xnor U7723 (N_7723,N_7466,N_6711);
nor U7724 (N_7724,N_5170,N_6153);
nand U7725 (N_7725,N_5424,N_6548);
nand U7726 (N_7726,N_6630,N_5072);
and U7727 (N_7727,N_6515,N_5953);
nor U7728 (N_7728,N_6113,N_6104);
xor U7729 (N_7729,N_7082,N_5624);
or U7730 (N_7730,N_5924,N_5830);
or U7731 (N_7731,N_7398,N_7386);
or U7732 (N_7732,N_7091,N_6494);
xnor U7733 (N_7733,N_5674,N_5462);
or U7734 (N_7734,N_6116,N_5670);
or U7735 (N_7735,N_5550,N_7131);
nand U7736 (N_7736,N_5554,N_7126);
and U7737 (N_7737,N_7081,N_7435);
nor U7738 (N_7738,N_5470,N_5800);
xor U7739 (N_7739,N_6608,N_7037);
or U7740 (N_7740,N_7191,N_6405);
xor U7741 (N_7741,N_6079,N_6334);
or U7742 (N_7742,N_5989,N_6268);
and U7743 (N_7743,N_6395,N_7086);
or U7744 (N_7744,N_5483,N_5864);
xor U7745 (N_7745,N_7482,N_7000);
or U7746 (N_7746,N_6280,N_6852);
nand U7747 (N_7747,N_5825,N_6471);
and U7748 (N_7748,N_5287,N_6915);
or U7749 (N_7749,N_5884,N_6891);
nand U7750 (N_7750,N_6198,N_5548);
nand U7751 (N_7751,N_6086,N_6918);
and U7752 (N_7752,N_6632,N_6748);
nand U7753 (N_7753,N_5395,N_6560);
xor U7754 (N_7754,N_5321,N_7087);
nor U7755 (N_7755,N_5220,N_6448);
nand U7756 (N_7756,N_5701,N_6089);
or U7757 (N_7757,N_5581,N_7462);
nor U7758 (N_7758,N_5357,N_7403);
and U7759 (N_7759,N_5236,N_6882);
nor U7760 (N_7760,N_6658,N_7366);
nand U7761 (N_7761,N_5346,N_6317);
nand U7762 (N_7762,N_6617,N_6165);
and U7763 (N_7763,N_7196,N_6392);
nor U7764 (N_7764,N_5610,N_6979);
nand U7765 (N_7765,N_6590,N_7286);
or U7766 (N_7766,N_5257,N_6209);
xnor U7767 (N_7767,N_6406,N_5861);
or U7768 (N_7768,N_6248,N_5664);
or U7769 (N_7769,N_6348,N_5978);
and U7770 (N_7770,N_6327,N_5406);
xor U7771 (N_7771,N_5099,N_5979);
nand U7772 (N_7772,N_5190,N_5688);
nor U7773 (N_7773,N_6989,N_6601);
or U7774 (N_7774,N_6755,N_6004);
or U7775 (N_7775,N_7431,N_5417);
xnor U7776 (N_7776,N_6511,N_6144);
or U7777 (N_7777,N_6012,N_6477);
nor U7778 (N_7778,N_6447,N_7033);
nand U7779 (N_7779,N_6581,N_5103);
nand U7780 (N_7780,N_6886,N_6738);
nor U7781 (N_7781,N_6568,N_5741);
nand U7782 (N_7782,N_7252,N_5172);
xor U7783 (N_7783,N_5648,N_6402);
xor U7784 (N_7784,N_5630,N_5872);
nor U7785 (N_7785,N_7134,N_7311);
and U7786 (N_7786,N_5141,N_5671);
nand U7787 (N_7787,N_7484,N_5836);
nor U7788 (N_7788,N_5625,N_5192);
and U7789 (N_7789,N_6911,N_6202);
xnor U7790 (N_7790,N_5105,N_5793);
xor U7791 (N_7791,N_5712,N_5594);
xor U7792 (N_7792,N_6793,N_6901);
nor U7793 (N_7793,N_7013,N_7084);
nor U7794 (N_7794,N_5660,N_5680);
or U7795 (N_7795,N_5225,N_5713);
nand U7796 (N_7796,N_6832,N_6784);
and U7797 (N_7797,N_7255,N_5528);
or U7798 (N_7798,N_5100,N_5031);
or U7799 (N_7799,N_5339,N_5673);
xor U7800 (N_7800,N_5270,N_6880);
and U7801 (N_7801,N_6358,N_6117);
nor U7802 (N_7802,N_6584,N_7494);
xor U7803 (N_7803,N_5051,N_5251);
and U7804 (N_7804,N_5047,N_5533);
and U7805 (N_7805,N_6521,N_5322);
nor U7806 (N_7806,N_7249,N_6239);
nor U7807 (N_7807,N_7036,N_6384);
nand U7808 (N_7808,N_6446,N_5931);
nand U7809 (N_7809,N_6435,N_5560);
and U7810 (N_7810,N_7195,N_7352);
nor U7811 (N_7811,N_5513,N_6767);
and U7812 (N_7812,N_6551,N_5197);
xor U7813 (N_7813,N_6687,N_6741);
and U7814 (N_7814,N_7424,N_5048);
and U7815 (N_7815,N_5039,N_5909);
nor U7816 (N_7816,N_5024,N_5479);
xnor U7817 (N_7817,N_5593,N_6194);
nor U7818 (N_7818,N_7264,N_7125);
or U7819 (N_7819,N_5285,N_6709);
and U7820 (N_7820,N_7221,N_6701);
nor U7821 (N_7821,N_6067,N_6462);
nand U7822 (N_7822,N_5277,N_7198);
and U7823 (N_7823,N_6120,N_7458);
nand U7824 (N_7824,N_6675,N_6372);
or U7825 (N_7825,N_6747,N_5043);
nand U7826 (N_7826,N_5870,N_6312);
xnor U7827 (N_7827,N_5335,N_7373);
nor U7828 (N_7828,N_7164,N_5849);
and U7829 (N_7829,N_7237,N_5588);
or U7830 (N_7830,N_7068,N_6718);
xnor U7831 (N_7831,N_7109,N_5050);
or U7832 (N_7832,N_5613,N_5033);
and U7833 (N_7833,N_7300,N_5722);
xnor U7834 (N_7834,N_6145,N_5780);
nor U7835 (N_7835,N_6461,N_6762);
or U7836 (N_7836,N_5873,N_6574);
and U7837 (N_7837,N_5921,N_5330);
nand U7838 (N_7838,N_5668,N_7115);
or U7839 (N_7839,N_5908,N_6619);
and U7840 (N_7840,N_5272,N_5627);
xor U7841 (N_7841,N_6799,N_6426);
xor U7842 (N_7842,N_6782,N_6845);
nand U7843 (N_7843,N_7073,N_7491);
nor U7844 (N_7844,N_7079,N_5982);
nand U7845 (N_7845,N_7463,N_7496);
or U7846 (N_7846,N_5019,N_6851);
or U7847 (N_7847,N_5867,N_5640);
and U7848 (N_7848,N_5500,N_6792);
or U7849 (N_7849,N_6735,N_5394);
xnor U7850 (N_7850,N_5961,N_5181);
or U7851 (N_7851,N_5644,N_5677);
nor U7852 (N_7852,N_5182,N_7292);
and U7853 (N_7853,N_6028,N_5672);
nor U7854 (N_7854,N_7023,N_6098);
and U7855 (N_7855,N_5313,N_6583);
or U7856 (N_7856,N_6739,N_6826);
nand U7857 (N_7857,N_6618,N_7350);
and U7858 (N_7858,N_6736,N_5341);
and U7859 (N_7859,N_7022,N_5685);
and U7860 (N_7860,N_5098,N_5037);
or U7861 (N_7861,N_5364,N_5976);
nand U7862 (N_7862,N_6355,N_7459);
nor U7863 (N_7863,N_7245,N_5727);
nor U7864 (N_7864,N_5185,N_5193);
and U7865 (N_7865,N_5345,N_6710);
nor U7866 (N_7866,N_5519,N_6588);
nand U7867 (N_7867,N_5108,N_7075);
nor U7868 (N_7868,N_6847,N_7418);
nand U7869 (N_7869,N_6802,N_7447);
xor U7870 (N_7870,N_5945,N_6063);
nand U7871 (N_7871,N_6167,N_6661);
nand U7872 (N_7872,N_5551,N_5543);
nor U7873 (N_7873,N_6878,N_5854);
and U7874 (N_7874,N_7146,N_7387);
and U7875 (N_7875,N_5615,N_5655);
nand U7876 (N_7876,N_6112,N_6607);
nand U7877 (N_7877,N_6654,N_5076);
xnor U7878 (N_7878,N_6014,N_6256);
and U7879 (N_7879,N_5122,N_6966);
xor U7880 (N_7880,N_7493,N_7239);
xor U7881 (N_7881,N_6753,N_6562);
xnor U7882 (N_7882,N_6941,N_6566);
or U7883 (N_7883,N_7410,N_5308);
nand U7884 (N_7884,N_5401,N_5121);
nand U7885 (N_7885,N_7200,N_5445);
or U7886 (N_7886,N_7001,N_6947);
or U7887 (N_7887,N_6561,N_7404);
or U7888 (N_7888,N_5362,N_7308);
xnor U7889 (N_7889,N_6835,N_7227);
nand U7890 (N_7890,N_6785,N_6252);
and U7891 (N_7891,N_6284,N_5344);
nor U7892 (N_7892,N_5128,N_5159);
and U7893 (N_7893,N_5426,N_6853);
nor U7894 (N_7894,N_5038,N_7060);
xnor U7895 (N_7895,N_6920,N_6656);
and U7896 (N_7896,N_5614,N_5372);
or U7897 (N_7897,N_6430,N_5214);
and U7898 (N_7898,N_6704,N_5213);
nand U7899 (N_7899,N_5546,N_6955);
and U7900 (N_7900,N_7322,N_5527);
or U7901 (N_7901,N_7429,N_7348);
or U7902 (N_7902,N_7460,N_7461);
nor U7903 (N_7903,N_6088,N_7232);
xor U7904 (N_7904,N_7381,N_5903);
or U7905 (N_7905,N_5822,N_5917);
nand U7906 (N_7906,N_6917,N_6555);
xor U7907 (N_7907,N_5061,N_6351);
and U7908 (N_7908,N_7428,N_6257);
nor U7909 (N_7909,N_6700,N_5119);
nor U7910 (N_7910,N_5354,N_6213);
nand U7911 (N_7911,N_7377,N_7291);
nor U7912 (N_7912,N_6772,N_5253);
nor U7913 (N_7913,N_5137,N_6158);
or U7914 (N_7914,N_5843,N_6957);
xor U7915 (N_7915,N_7414,N_6183);
or U7916 (N_7916,N_6176,N_5302);
nand U7917 (N_7917,N_6016,N_6764);
nand U7918 (N_7918,N_6041,N_7481);
xnor U7919 (N_7919,N_6338,N_5348);
or U7920 (N_7920,N_5229,N_6455);
nand U7921 (N_7921,N_6994,N_6803);
nor U7922 (N_7922,N_6039,N_5632);
nand U7923 (N_7923,N_7267,N_7144);
or U7924 (N_7924,N_6263,N_5299);
nor U7925 (N_7925,N_5477,N_6637);
nand U7926 (N_7926,N_5638,N_7278);
and U7927 (N_7927,N_5058,N_6195);
nand U7928 (N_7928,N_5990,N_7171);
nor U7929 (N_7929,N_7140,N_5812);
nor U7930 (N_7930,N_7067,N_6071);
nor U7931 (N_7931,N_5587,N_5735);
xnor U7932 (N_7932,N_7222,N_6961);
or U7933 (N_7933,N_5782,N_6210);
xnor U7934 (N_7934,N_6483,N_6129);
xor U7935 (N_7935,N_5653,N_6987);
or U7936 (N_7936,N_7076,N_7281);
nor U7937 (N_7937,N_6232,N_6983);
or U7938 (N_7938,N_6895,N_6567);
and U7939 (N_7939,N_6407,N_6935);
xor U7940 (N_7940,N_5922,N_6370);
nor U7941 (N_7941,N_6810,N_6275);
or U7942 (N_7942,N_5056,N_5962);
nand U7943 (N_7943,N_5739,N_5748);
nor U7944 (N_7944,N_7230,N_7138);
nand U7945 (N_7945,N_7276,N_7189);
nand U7946 (N_7946,N_5803,N_5142);
nor U7947 (N_7947,N_7103,N_6679);
and U7948 (N_7948,N_5367,N_7483);
or U7949 (N_7949,N_5832,N_5093);
or U7950 (N_7950,N_6775,N_6101);
nor U7951 (N_7951,N_5767,N_5751);
nor U7952 (N_7952,N_6254,N_6652);
and U7953 (N_7953,N_5957,N_5623);
xor U7954 (N_7954,N_6554,N_5579);
or U7955 (N_7955,N_6032,N_6889);
or U7956 (N_7956,N_5720,N_6970);
nor U7957 (N_7957,N_6856,N_5465);
xnor U7958 (N_7958,N_6249,N_6571);
xor U7959 (N_7959,N_5385,N_6648);
and U7960 (N_7960,N_7107,N_6604);
nor U7961 (N_7961,N_5992,N_6026);
nand U7962 (N_7962,N_7116,N_6683);
nand U7963 (N_7963,N_6015,N_7275);
nand U7964 (N_7964,N_6665,N_5571);
or U7965 (N_7965,N_7197,N_6300);
nor U7966 (N_7966,N_7269,N_6070);
nand U7967 (N_7967,N_5402,N_5501);
or U7968 (N_7968,N_5792,N_7490);
nand U7969 (N_7969,N_5366,N_7056);
nand U7970 (N_7970,N_6021,N_5378);
nand U7971 (N_7971,N_7448,N_5059);
nor U7972 (N_7972,N_6285,N_6550);
xor U7973 (N_7973,N_7017,N_5195);
and U7974 (N_7974,N_6475,N_5457);
and U7975 (N_7975,N_5612,N_5572);
nand U7976 (N_7976,N_5416,N_6787);
xnor U7977 (N_7977,N_7181,N_5667);
nor U7978 (N_7978,N_6667,N_6423);
and U7979 (N_7979,N_7379,N_6864);
or U7980 (N_7980,N_6150,N_5286);
nor U7981 (N_7981,N_6528,N_6786);
xnor U7982 (N_7982,N_5736,N_6350);
xor U7983 (N_7983,N_5676,N_6754);
and U7984 (N_7984,N_6305,N_5619);
and U7985 (N_7985,N_5217,N_6536);
nor U7986 (N_7986,N_6427,N_5552);
and U7987 (N_7987,N_6800,N_6883);
and U7988 (N_7988,N_5140,N_5392);
nand U7989 (N_7989,N_5645,N_5030);
nor U7990 (N_7990,N_5490,N_7474);
or U7991 (N_7991,N_5112,N_6522);
and U7992 (N_7992,N_5887,N_6214);
nor U7993 (N_7993,N_5656,N_6868);
nor U7994 (N_7994,N_6932,N_7168);
nand U7995 (N_7995,N_5732,N_7121);
and U7996 (N_7996,N_5910,N_5295);
xor U7997 (N_7997,N_6172,N_6885);
xor U7998 (N_7998,N_7260,N_5897);
nor U7999 (N_7999,N_5332,N_5463);
and U8000 (N_8000,N_6737,N_5697);
xor U8001 (N_8001,N_6519,N_5766);
xnor U8002 (N_8002,N_5934,N_6243);
nand U8003 (N_8003,N_5860,N_6921);
xor U8004 (N_8004,N_5769,N_7040);
and U8005 (N_8005,N_5694,N_7045);
or U8006 (N_8006,N_5177,N_7069);
nand U8007 (N_8007,N_7423,N_6040);
nor U8008 (N_8008,N_5952,N_6833);
nand U8009 (N_8009,N_5629,N_5609);
or U8010 (N_8010,N_5646,N_6009);
nor U8011 (N_8011,N_5946,N_6103);
nand U8012 (N_8012,N_5315,N_5107);
and U8013 (N_8013,N_7206,N_5535);
nor U8014 (N_8014,N_5151,N_5055);
xnor U8015 (N_8015,N_7441,N_6340);
nand U8016 (N_8016,N_5152,N_7035);
or U8017 (N_8017,N_6925,N_7110);
nand U8018 (N_8018,N_7070,N_6971);
nor U8019 (N_8019,N_6001,N_6487);
xor U8020 (N_8020,N_6863,N_6778);
or U8021 (N_8021,N_6398,N_6616);
or U8022 (N_8022,N_6415,N_6251);
nand U8023 (N_8023,N_5336,N_5260);
nor U8024 (N_8024,N_6685,N_6408);
nor U8025 (N_8025,N_5973,N_5244);
and U8026 (N_8026,N_7055,N_6493);
nand U8027 (N_8027,N_5935,N_6020);
xnor U8028 (N_8028,N_6099,N_5484);
nor U8029 (N_8029,N_5338,N_5651);
xor U8030 (N_8030,N_7104,N_5747);
xnor U8031 (N_8031,N_7455,N_5328);
nor U8032 (N_8032,N_6184,N_5888);
nand U8033 (N_8033,N_5200,N_5293);
nand U8034 (N_8034,N_5403,N_5808);
nand U8035 (N_8035,N_7158,N_6206);
or U8036 (N_8036,N_6132,N_6692);
xor U8037 (N_8037,N_5859,N_5691);
xnor U8038 (N_8038,N_6814,N_5898);
or U8039 (N_8039,N_5206,N_5115);
xnor U8040 (N_8040,N_6443,N_5355);
nand U8041 (N_8041,N_6095,N_7178);
and U8042 (N_8042,N_7032,N_5377);
nor U8043 (N_8043,N_5186,N_5340);
and U8044 (N_8044,N_6512,N_5440);
and U8045 (N_8045,N_5237,N_6516);
or U8046 (N_8046,N_6993,N_5666);
xnor U8047 (N_8047,N_5900,N_6038);
nor U8048 (N_8048,N_7346,N_5690);
nand U8049 (N_8049,N_5239,N_5787);
nor U8050 (N_8050,N_6233,N_7114);
and U8051 (N_8051,N_6613,N_5023);
or U8052 (N_8052,N_6322,N_5194);
or U8053 (N_8053,N_5191,N_5297);
nor U8054 (N_8054,N_5309,N_6759);
xnor U8055 (N_8055,N_5514,N_7180);
or U8056 (N_8056,N_5256,N_5835);
nand U8057 (N_8057,N_6255,N_6937);
and U8058 (N_8058,N_5138,N_7306);
nor U8059 (N_8059,N_6975,N_6412);
nor U8060 (N_8060,N_6313,N_7370);
and U8061 (N_8061,N_6111,N_6456);
nand U8062 (N_8062,N_5158,N_5889);
xor U8063 (N_8063,N_7193,N_5459);
and U8064 (N_8064,N_7296,N_6352);
or U8065 (N_8065,N_6288,N_7355);
nor U8066 (N_8066,N_6597,N_7012);
and U8067 (N_8067,N_5706,N_6122);
nand U8068 (N_8068,N_6546,N_6139);
or U8069 (N_8069,N_5289,N_5451);
and U8070 (N_8070,N_5763,N_6359);
or U8071 (N_8071,N_6962,N_6942);
nor U8072 (N_8072,N_5442,N_5784);
and U8073 (N_8073,N_5568,N_6291);
and U8074 (N_8074,N_7065,N_7282);
and U8075 (N_8075,N_7220,N_6677);
nand U8076 (N_8076,N_5932,N_6164);
or U8077 (N_8077,N_6727,N_7157);
nor U8078 (N_8078,N_5189,N_6602);
xor U8079 (N_8079,N_5536,N_5523);
and U8080 (N_8080,N_7340,N_6134);
nand U8081 (N_8081,N_6320,N_7010);
nand U8082 (N_8082,N_6031,N_6819);
and U8083 (N_8083,N_6138,N_7143);
nor U8084 (N_8084,N_7090,N_6264);
xnor U8085 (N_8085,N_5391,N_5840);
xnor U8086 (N_8086,N_5886,N_6485);
nor U8087 (N_8087,N_7345,N_7444);
xor U8088 (N_8088,N_6651,N_5375);
or U8089 (N_8089,N_5261,N_5569);
nor U8090 (N_8090,N_5029,N_6862);
and U8091 (N_8091,N_6107,N_6686);
and U8092 (N_8092,N_6179,N_5125);
xnor U8093 (N_8093,N_5716,N_6017);
xnor U8094 (N_8094,N_7299,N_6170);
nand U8095 (N_8095,N_6822,N_6705);
and U8096 (N_8096,N_5168,N_6369);
xor U8097 (N_8097,N_6598,N_7295);
xnor U8098 (N_8098,N_5951,N_6003);
xnor U8099 (N_8099,N_5016,N_6008);
xnor U8100 (N_8100,N_7159,N_6633);
nand U8101 (N_8101,N_6623,N_5679);
nor U8102 (N_8102,N_5221,N_6149);
or U8103 (N_8103,N_7150,N_7050);
and U8104 (N_8104,N_5288,N_6373);
nand U8105 (N_8105,N_6326,N_5505);
or U8106 (N_8106,N_5202,N_6105);
and U8107 (N_8107,N_7456,N_5127);
nor U8108 (N_8108,N_6094,N_5269);
xnor U8109 (N_8109,N_5862,N_7416);
xnor U8110 (N_8110,N_5242,N_7213);
nor U8111 (N_8111,N_6870,N_5633);
xnor U8112 (N_8112,N_6187,N_5410);
nor U8113 (N_8113,N_5926,N_6716);
or U8114 (N_8114,N_6393,N_6808);
nor U8115 (N_8115,N_6794,N_6827);
nor U8116 (N_8116,N_5393,N_5636);
or U8117 (N_8117,N_5583,N_7179);
and U8118 (N_8118,N_7464,N_6161);
nor U8119 (N_8119,N_6163,N_5368);
xnor U8120 (N_8120,N_5427,N_7253);
nor U8121 (N_8121,N_5585,N_5178);
nor U8122 (N_8122,N_5074,N_5258);
xnor U8123 (N_8123,N_5746,N_6269);
nand U8124 (N_8124,N_5235,N_6159);
and U8125 (N_8125,N_6992,N_7003);
or U8126 (N_8126,N_6674,N_5816);
nor U8127 (N_8127,N_5439,N_6386);
or U8128 (N_8128,N_6464,N_6890);
or U8129 (N_8129,N_6899,N_6525);
or U8130 (N_8130,N_6374,N_5553);
xor U8131 (N_8131,N_5460,N_7368);
xnor U8132 (N_8132,N_6077,N_7383);
nor U8133 (N_8133,N_6877,N_5232);
and U8134 (N_8134,N_6575,N_6939);
nand U8135 (N_8135,N_7409,N_6486);
and U8136 (N_8136,N_6025,N_6377);
xnor U8137 (N_8137,N_6609,N_5974);
xor U8138 (N_8138,N_6603,N_6011);
or U8139 (N_8139,N_7163,N_5503);
xor U8140 (N_8140,N_5826,N_5233);
nand U8141 (N_8141,N_5774,N_5544);
and U8142 (N_8142,N_5005,N_5578);
nand U8143 (N_8143,N_6813,N_5730);
nor U8144 (N_8144,N_6240,N_5064);
and U8145 (N_8145,N_7328,N_6066);
or U8146 (N_8146,N_6642,N_6467);
nand U8147 (N_8147,N_6672,N_5580);
nor U8148 (N_8148,N_5797,N_6173);
and U8149 (N_8149,N_5259,N_7063);
nand U8150 (N_8150,N_6119,N_5066);
nand U8151 (N_8151,N_5491,N_6825);
and U8152 (N_8152,N_5411,N_7334);
or U8153 (N_8153,N_5413,N_7011);
nand U8154 (N_8154,N_5420,N_6052);
xor U8155 (N_8155,N_6247,N_5068);
nand U8156 (N_8156,N_6790,N_6763);
nor U8157 (N_8157,N_5388,N_5760);
and U8158 (N_8158,N_5387,N_5798);
xor U8159 (N_8159,N_6859,N_5398);
xor U8160 (N_8160,N_5123,N_5923);
and U8161 (N_8161,N_5397,N_5234);
or U8162 (N_8162,N_5118,N_6137);
xnor U8163 (N_8163,N_5657,N_6468);
or U8164 (N_8164,N_5948,N_6898);
xnor U8165 (N_8165,N_6565,N_6636);
or U8166 (N_8166,N_7118,N_6053);
and U8167 (N_8167,N_5323,N_6295);
or U8168 (N_8168,N_5595,N_5721);
and U8169 (N_8169,N_5892,N_6152);
and U8170 (N_8170,N_5487,N_6245);
or U8171 (N_8171,N_5911,N_6204);
nand U8172 (N_8172,N_6664,N_6582);
xor U8173 (N_8173,N_7211,N_6126);
and U8174 (N_8174,N_5376,N_5807);
nand U8175 (N_8175,N_7105,N_6972);
and U8176 (N_8176,N_6978,N_6614);
xor U8177 (N_8177,N_5482,N_6469);
and U8178 (N_8178,N_7130,N_5899);
xor U8179 (N_8179,N_6545,N_5596);
and U8180 (N_8180,N_5173,N_6201);
nand U8181 (N_8181,N_6769,N_5882);
nand U8182 (N_8182,N_5203,N_6410);
nor U8183 (N_8183,N_5879,N_7332);
nor U8184 (N_8184,N_5711,N_6506);
xnor U8185 (N_8185,N_5507,N_5283);
and U8186 (N_8186,N_7216,N_6146);
and U8187 (N_8187,N_6178,N_5091);
nor U8188 (N_8188,N_7078,N_5966);
xnor U8189 (N_8189,N_5199,N_5906);
or U8190 (N_8190,N_5069,N_6625);
xor U8191 (N_8191,N_5545,N_6417);
xor U8192 (N_8192,N_5971,N_6585);
and U8193 (N_8193,N_7100,N_6433);
nor U8194 (N_8194,N_6416,N_7108);
nor U8195 (N_8195,N_5318,N_7170);
xnor U8196 (N_8196,N_5224,N_5814);
or U8197 (N_8197,N_6635,N_7391);
and U8198 (N_8198,N_6203,N_6690);
nor U8199 (N_8199,N_6946,N_5296);
and U8200 (N_8200,N_6072,N_5279);
xor U8201 (N_8201,N_5135,N_5777);
nand U8202 (N_8202,N_5404,N_6106);
and U8203 (N_8203,N_6301,N_5541);
and U8204 (N_8204,N_5855,N_6933);
nor U8205 (N_8205,N_6874,N_5486);
or U8206 (N_8206,N_6328,N_7309);
nand U8207 (N_8207,N_5618,N_5508);
and U8208 (N_8208,N_5891,N_6010);
nor U8209 (N_8209,N_6318,N_6547);
nand U8210 (N_8210,N_7016,N_6564);
nor U8211 (N_8211,N_6838,N_6439);
xnor U8212 (N_8212,N_7446,N_7172);
nand U8213 (N_8213,N_5781,N_7389);
and U8214 (N_8214,N_7054,N_6620);
or U8215 (N_8215,N_5496,N_5733);
or U8216 (N_8216,N_5447,N_5084);
and U8217 (N_8217,N_5526,N_7333);
nand U8218 (N_8218,N_6743,N_6419);
nand U8219 (N_8219,N_6463,N_6044);
nor U8220 (N_8220,N_5432,N_5415);
xor U8221 (N_8221,N_7153,N_6325);
or U8222 (N_8222,N_6558,N_7443);
nor U8223 (N_8223,N_6205,N_6289);
xor U8224 (N_8224,N_7289,N_6353);
nor U8225 (N_8225,N_7261,N_5617);
xor U8226 (N_8226,N_6777,N_5267);
nor U8227 (N_8227,N_5169,N_6013);
and U8228 (N_8228,N_5586,N_6341);
xor U8229 (N_8229,N_6723,N_6949);
or U8230 (N_8230,N_6830,N_6660);
xor U8231 (N_8231,N_5300,N_5009);
or U8232 (N_8232,N_5562,N_6160);
and U8233 (N_8233,N_6174,N_5314);
and U8234 (N_8234,N_5075,N_5241);
xor U8235 (N_8235,N_5205,N_5156);
or U8236 (N_8236,N_6593,N_6421);
nand U8237 (N_8237,N_7353,N_7293);
nand U8238 (N_8238,N_5175,N_5090);
nand U8239 (N_8239,N_5555,N_6208);
nand U8240 (N_8240,N_5620,N_5032);
nor U8241 (N_8241,N_6809,N_5775);
and U8242 (N_8242,N_6424,N_7426);
nand U8243 (N_8243,N_6297,N_6046);
nand U8244 (N_8244,N_6758,N_5837);
or U8245 (N_8245,N_6307,N_6900);
nor U8246 (N_8246,N_6907,N_7135);
nand U8247 (N_8247,N_5495,N_6085);
xor U8248 (N_8248,N_6958,N_7384);
or U8249 (N_8249,N_5052,N_7234);
nor U8250 (N_8250,N_5723,N_5675);
nor U8251 (N_8251,N_7465,N_5573);
nand U8252 (N_8252,N_5916,N_5171);
or U8253 (N_8253,N_6869,N_6659);
xnor U8254 (N_8254,N_6302,N_5149);
xnor U8255 (N_8255,N_5851,N_5284);
or U8256 (N_8256,N_5665,N_6460);
nand U8257 (N_8257,N_6151,N_6524);
nand U8258 (N_8258,N_5418,N_5294);
or U8259 (N_8259,N_5972,N_5265);
or U8260 (N_8260,N_5682,N_6125);
xor U8261 (N_8261,N_7470,N_5435);
xnor U8262 (N_8262,N_5006,N_5846);
or U8263 (N_8263,N_5343,N_5078);
or U8264 (N_8264,N_7354,N_5857);
or U8265 (N_8265,N_6143,N_5985);
xnor U8266 (N_8266,N_5602,N_6057);
xnor U8267 (N_8267,N_5478,N_5650);
xnor U8268 (N_8268,N_6244,N_5539);
xnor U8269 (N_8269,N_6123,N_5035);
nor U8270 (N_8270,N_5071,N_5987);
xnor U8271 (N_8271,N_5409,N_7004);
xor U8272 (N_8272,N_5958,N_6371);
xnor U8273 (N_8273,N_6752,N_5866);
nor U8274 (N_8274,N_7019,N_7007);
xnor U8275 (N_8275,N_6963,N_5811);
xor U8276 (N_8276,N_7361,N_5350);
and U8277 (N_8277,N_5408,N_5622);
xor U8278 (N_8278,N_7285,N_7218);
and U8279 (N_8279,N_6140,N_5518);
nand U8280 (N_8280,N_5263,N_6595);
xor U8281 (N_8281,N_6959,N_5412);
nand U8282 (N_8282,N_5929,N_5880);
nand U8283 (N_8283,N_5466,N_6466);
xor U8284 (N_8284,N_6938,N_5511);
xor U8285 (N_8285,N_6470,N_5791);
or U8286 (N_8286,N_6200,N_7136);
or U8287 (N_8287,N_5373,N_5266);
or U8288 (N_8288,N_5806,N_6100);
xnor U8289 (N_8289,N_5247,N_5018);
or U8290 (N_8290,N_7364,N_5890);
and U8291 (N_8291,N_6236,N_6339);
nor U8292 (N_8292,N_5431,N_6896);
and U8293 (N_8293,N_7059,N_7445);
nor U8294 (N_8294,N_5053,N_5429);
xor U8295 (N_8295,N_7236,N_5824);
and U8296 (N_8296,N_6699,N_6894);
xor U8297 (N_8297,N_6520,N_7176);
nand U8298 (N_8298,N_6050,N_5467);
nand U8299 (N_8299,N_5201,N_6024);
or U8300 (N_8300,N_6731,N_5361);
or U8301 (N_8301,N_7451,N_5275);
xor U8302 (N_8302,N_5699,N_5106);
xor U8303 (N_8303,N_7014,N_7165);
nand U8304 (N_8304,N_5353,N_6967);
nor U8305 (N_8305,N_6638,N_6378);
nand U8306 (N_8306,N_6045,N_7243);
nand U8307 (N_8307,N_7371,N_6671);
xor U8308 (N_8308,N_7038,N_7315);
and U8309 (N_8309,N_5311,N_5198);
nor U8310 (N_8310,N_7395,N_6517);
nor U8311 (N_8311,N_6023,N_6127);
nor U8312 (N_8312,N_6653,N_6742);
xor U8313 (N_8313,N_5531,N_7372);
xnor U8314 (N_8314,N_6502,N_5025);
and U8315 (N_8315,N_7270,N_5469);
nor U8316 (N_8316,N_5768,N_6391);
xnor U8317 (N_8317,N_5920,N_5428);
or U8318 (N_8318,N_6510,N_6090);
nand U8319 (N_8319,N_5991,N_7083);
and U8320 (N_8320,N_5524,N_6458);
and U8321 (N_8321,N_5493,N_6924);
nand U8322 (N_8322,N_7240,N_6676);
or U8323 (N_8323,N_5352,N_5601);
nor U8324 (N_8324,N_5131,N_5110);
and U8325 (N_8325,N_6770,N_6606);
or U8326 (N_8326,N_6357,N_7272);
nand U8327 (N_8327,N_7250,N_7497);
or U8328 (N_8328,N_6807,N_7217);
xnor U8329 (N_8329,N_5167,N_7475);
xnor U8330 (N_8330,N_7487,N_6719);
or U8331 (N_8331,N_5687,N_5790);
and U8332 (N_8332,N_6779,N_6440);
nor U8333 (N_8333,N_6673,N_5155);
or U8334 (N_8334,N_5082,N_6875);
and U8335 (N_8335,N_5559,N_7099);
nor U8336 (N_8336,N_6335,N_7287);
and U8337 (N_8337,N_5113,N_6332);
nand U8338 (N_8338,N_5833,N_5386);
nor U8339 (N_8339,N_7223,N_5669);
nor U8340 (N_8340,N_6552,N_5211);
or U8341 (N_8341,N_7024,N_6744);
nor U8342 (N_8342,N_5109,N_5654);
or U8343 (N_8343,N_7098,N_5227);
and U8344 (N_8344,N_6484,N_7127);
nand U8345 (N_8345,N_5092,N_6314);
nor U8346 (N_8346,N_6557,N_5379);
nor U8347 (N_8347,N_5823,N_5405);
and U8348 (N_8348,N_5737,N_7028);
and U8349 (N_8349,N_5534,N_7486);
or U8350 (N_8350,N_7058,N_6362);
and U8351 (N_8351,N_6733,N_5844);
xor U8352 (N_8352,N_6336,N_6828);
or U8353 (N_8353,N_7417,N_5347);
nor U8354 (N_8354,N_6061,N_6969);
and U8355 (N_8355,N_6259,N_5088);
xnor U8356 (N_8356,N_7226,N_5516);
nor U8357 (N_8357,N_5414,N_5877);
nand U8358 (N_8358,N_7385,N_5464);
xor U8359 (N_8359,N_5955,N_7454);
and U8360 (N_8360,N_5129,N_6611);
and U8361 (N_8361,N_6806,N_6580);
and U8362 (N_8362,N_6621,N_7169);
nand U8363 (N_8363,N_5356,N_5252);
xor U8364 (N_8364,N_6954,N_6843);
nand U8365 (N_8365,N_5758,N_7160);
or U8366 (N_8366,N_7402,N_6872);
nand U8367 (N_8367,N_6473,N_6133);
and U8368 (N_8368,N_6333,N_6363);
and U8369 (N_8369,N_6304,N_5698);
nand U8370 (N_8370,N_6501,N_5724);
nand U8371 (N_8371,N_7480,N_5117);
and U8372 (N_8372,N_6505,N_6404);
and U8373 (N_8373,N_6235,N_6185);
and U8374 (N_8374,N_7248,N_7305);
or U8375 (N_8375,N_5783,N_6956);
nand U8376 (N_8376,N_7101,N_6495);
nor U8377 (N_8377,N_6121,N_6513);
nor U8378 (N_8378,N_5635,N_5626);
nor U8379 (N_8379,N_5591,N_5986);
xnor U8380 (N_8380,N_5248,N_6092);
or U8381 (N_8381,N_6361,N_7212);
nand U8382 (N_8382,N_5291,N_5868);
xnor U8383 (N_8383,N_5802,N_7394);
and U8384 (N_8384,N_5759,N_6713);
and U8385 (N_8385,N_5628,N_5726);
and U8386 (N_8386,N_7468,N_6155);
or U8387 (N_8387,N_5446,N_7156);
and U8388 (N_8388,N_7442,N_7449);
or U8389 (N_8389,N_5278,N_6622);
nor U8390 (N_8390,N_5073,N_5785);
nor U8391 (N_8391,N_7415,N_5240);
and U8392 (N_8392,N_5096,N_5734);
or U8393 (N_8393,N_5497,N_5521);
nand U8394 (N_8394,N_6781,N_6801);
nand U8395 (N_8395,N_5574,N_6387);
or U8396 (N_8396,N_5894,N_5874);
nand U8397 (N_8397,N_6995,N_5959);
xor U8398 (N_8398,N_6948,N_5014);
xnor U8399 (N_8399,N_6059,N_5841);
nor U8400 (N_8400,N_6337,N_6476);
nand U8401 (N_8401,N_5757,N_6980);
or U8402 (N_8402,N_5180,N_6207);
nand U8403 (N_8403,N_6276,N_6394);
or U8404 (N_8404,N_7263,N_5753);
or U8405 (N_8405,N_5530,N_5642);
nor U8406 (N_8406,N_6605,N_5083);
or U8407 (N_8407,N_5102,N_6892);
nand U8408 (N_8408,N_6154,N_7325);
nor U8409 (N_8409,N_6817,N_5146);
nor U8410 (N_8410,N_5786,N_6217);
nand U8411 (N_8411,N_6854,N_5692);
nand U8412 (N_8412,N_7396,N_5821);
nor U8413 (N_8413,N_5858,N_6523);
or U8414 (N_8414,N_6909,N_6694);
or U8415 (N_8415,N_6182,N_5163);
xnor U8416 (N_8416,N_5219,N_5875);
and U8417 (N_8417,N_5320,N_5492);
or U8418 (N_8418,N_5881,N_7495);
and U8419 (N_8419,N_6689,N_5274);
nor U8420 (N_8420,N_7277,N_5919);
or U8421 (N_8421,N_5604,N_6850);
nor U8422 (N_8422,N_6542,N_5441);
and U8423 (N_8423,N_5742,N_5077);
and U8424 (N_8424,N_5324,N_7005);
xor U8425 (N_8425,N_6893,N_5631);
nand U8426 (N_8426,N_6919,N_7274);
or U8427 (N_8427,N_6221,N_7327);
nor U8428 (N_8428,N_5563,N_5476);
nor U8429 (N_8429,N_6229,N_6197);
and U8430 (N_8430,N_6048,N_7225);
nor U8431 (N_8431,N_6707,N_6858);
and U8432 (N_8432,N_6457,N_5327);
and U8433 (N_8433,N_6029,N_7207);
and U8434 (N_8434,N_5087,N_5013);
nor U8435 (N_8435,N_5081,N_6498);
xor U8436 (N_8436,N_6065,N_6928);
and U8437 (N_8437,N_5845,N_5996);
or U8438 (N_8438,N_6514,N_6169);
nor U8439 (N_8439,N_5436,N_5382);
or U8440 (N_8440,N_6324,N_5796);
xor U8441 (N_8441,N_6849,N_5485);
nor U8442 (N_8442,N_5506,N_6022);
or U8443 (N_8443,N_6722,N_7317);
and U8444 (N_8444,N_5637,N_6069);
and U8445 (N_8445,N_7095,N_5438);
and U8446 (N_8446,N_6509,N_5702);
and U8447 (N_8447,N_6840,N_6922);
nand U8448 (N_8448,N_6124,N_5714);
nor U8449 (N_8449,N_7066,N_6873);
xnor U8450 (N_8450,N_5828,N_6449);
or U8451 (N_8451,N_5684,N_6532);
and U8452 (N_8452,N_7008,N_5502);
or U8453 (N_8453,N_6631,N_6951);
xnor U8454 (N_8454,N_6246,N_6445);
xor U8455 (N_8455,N_7137,N_6253);
or U8456 (N_8456,N_6290,N_5538);
nor U8457 (N_8457,N_6081,N_6714);
nor U8458 (N_8458,N_7439,N_5134);
and U8459 (N_8459,N_7074,N_7089);
nand U8460 (N_8460,N_5681,N_5810);
xor U8461 (N_8461,N_5230,N_6988);
nand U8462 (N_8462,N_5046,N_7155);
nor U8463 (N_8463,N_5995,N_6490);
xor U8464 (N_8464,N_6953,N_6273);
and U8465 (N_8465,N_5728,N_6702);
or U8466 (N_8466,N_6480,N_7162);
nand U8467 (N_8467,N_5304,N_7351);
xor U8468 (N_8468,N_7427,N_6531);
nor U8469 (N_8469,N_6757,N_6299);
or U8470 (N_8470,N_6791,N_6760);
and U8471 (N_8471,N_7339,N_6459);
nand U8472 (N_8472,N_7362,N_6771);
or U8473 (N_8473,N_7302,N_5576);
nand U8474 (N_8474,N_7498,N_7122);
nand U8475 (N_8475,N_7233,N_5749);
nand U8476 (N_8476,N_6306,N_5011);
nor U8477 (N_8477,N_7478,N_7124);
nor U8478 (N_8478,N_7471,N_5509);
or U8479 (N_8479,N_6952,N_6319);
xor U8480 (N_8480,N_6912,N_5437);
nand U8481 (N_8481,N_6329,N_6724);
xnor U8482 (N_8482,N_6064,N_6538);
xnor U8483 (N_8483,N_6910,N_5207);
xor U8484 (N_8484,N_6343,N_6647);
and U8485 (N_8485,N_6697,N_5641);
or U8486 (N_8486,N_6855,N_5634);
or U8487 (N_8487,N_7241,N_7489);
nand U8488 (N_8488,N_5187,N_5371);
or U8489 (N_8489,N_5292,N_6381);
nand U8490 (N_8490,N_6413,N_5461);
xor U8491 (N_8491,N_6428,N_6400);
nand U8492 (N_8492,N_6166,N_5703);
xnor U8493 (N_8493,N_7256,N_5210);
nand U8494 (N_8494,N_5561,N_6346);
nand U8495 (N_8495,N_6529,N_6643);
nor U8496 (N_8496,N_6267,N_6196);
and U8497 (N_8497,N_7102,N_7473);
nand U8498 (N_8498,N_5455,N_6211);
and U8499 (N_8499,N_6271,N_6926);
nor U8500 (N_8500,N_6130,N_5943);
and U8501 (N_8501,N_7326,N_5471);
nand U8502 (N_8502,N_6818,N_6897);
xor U8503 (N_8503,N_5453,N_5054);
and U8504 (N_8504,N_5494,N_6027);
xor U8505 (N_8505,N_7210,N_6750);
and U8506 (N_8506,N_6193,N_7052);
or U8507 (N_8507,N_6379,N_5161);
and U8508 (N_8508,N_5912,N_5600);
nand U8509 (N_8509,N_5070,N_6773);
nand U8510 (N_8510,N_6287,N_5208);
or U8511 (N_8511,N_6884,N_5652);
or U8512 (N_8512,N_5034,N_7369);
nand U8513 (N_8513,N_5949,N_6293);
or U8514 (N_8514,N_7303,N_5120);
nand U8515 (N_8515,N_6553,N_6798);
and U8516 (N_8516,N_5153,N_7034);
nor U8517 (N_8517,N_5556,N_6688);
nor U8518 (N_8518,N_6857,N_5848);
nor U8519 (N_8519,N_7092,N_5276);
or U8520 (N_8520,N_7177,N_5000);
nand U8521 (N_8521,N_6841,N_6230);
xor U8522 (N_8522,N_6540,N_5312);
xor U8523 (N_8523,N_5778,N_6761);
and U8524 (N_8524,N_7044,N_7214);
or U8525 (N_8525,N_6848,N_5164);
nand U8526 (N_8526,N_6492,N_6489);
nor U8527 (N_8527,N_5334,N_7314);
and U8528 (N_8528,N_7329,N_7202);
nor U8529 (N_8529,N_6805,N_5365);
and U8530 (N_8530,N_6579,N_6860);
nand U8531 (N_8531,N_6774,N_6231);
and U8532 (N_8532,N_5817,N_6765);
or U8533 (N_8533,N_7376,N_5273);
xor U8534 (N_8534,N_5839,N_5820);
nor U8535 (N_8535,N_5914,N_6376);
nand U8536 (N_8536,N_7499,N_5705);
nor U8537 (N_8537,N_6033,N_5063);
or U8538 (N_8538,N_5489,N_6431);
or U8539 (N_8539,N_6108,N_6592);
or U8540 (N_8540,N_5026,N_6018);
nand U8541 (N_8541,N_6136,N_5512);
nor U8542 (N_8542,N_7148,N_6986);
nor U8543 (N_8543,N_6083,N_5930);
or U8544 (N_8544,N_6570,N_6168);
nand U8545 (N_8545,N_7469,N_5968);
and U8546 (N_8546,N_6215,N_6663);
nor U8547 (N_8547,N_7020,N_5939);
nand U8548 (N_8548,N_5755,N_7319);
and U8549 (N_8549,N_6610,N_5938);
xnor U8550 (N_8550,N_6330,N_5829);
nor U8551 (N_8551,N_6563,N_6399);
xor U8552 (N_8552,N_6684,N_6238);
nand U8553 (N_8553,N_7117,N_7167);
nor U8554 (N_8554,N_7323,N_6812);
nand U8555 (N_8555,N_7247,N_6438);
and U8556 (N_8556,N_5196,N_7062);
nand U8557 (N_8557,N_6141,N_5396);
nand U8558 (N_8558,N_5326,N_6019);
and U8559 (N_8559,N_5433,N_5218);
nand U8560 (N_8560,N_5245,N_5659);
nand U8561 (N_8561,N_5422,N_7205);
or U8562 (N_8562,N_5696,N_7203);
nor U8563 (N_8563,N_6640,N_5850);
and U8564 (N_8564,N_6837,N_6212);
and U8565 (N_8565,N_6634,N_6780);
nor U8566 (N_8566,N_5965,N_7209);
nand U8567 (N_8567,N_5080,N_7182);
or U8568 (N_8568,N_7145,N_5856);
nor U8569 (N_8569,N_6944,N_5329);
xor U8570 (N_8570,N_5250,N_6973);
or U8571 (N_8571,N_7294,N_5718);
xnor U8572 (N_8572,N_6157,N_5981);
xnor U8573 (N_8573,N_7477,N_5448);
nor U8574 (N_8574,N_7313,N_6981);
or U8575 (N_8575,N_6397,N_7029);
and U8576 (N_8576,N_5941,N_6482);
or U8577 (N_8577,N_5246,N_5549);
and U8578 (N_8578,N_5809,N_5331);
nand U8579 (N_8579,N_7488,N_6082);
and U8580 (N_8580,N_5567,N_5895);
nor U8581 (N_8581,N_7142,N_5041);
or U8582 (N_8582,N_6549,N_5027);
nand U8583 (N_8583,N_6171,N_5473);
and U8584 (N_8584,N_5607,N_7492);
nor U8585 (N_8585,N_5761,N_5306);
or U8586 (N_8586,N_5788,N_5871);
or U8587 (N_8587,N_5520,N_5337);
xnor U8588 (N_8588,N_7254,N_6599);
xnor U8589 (N_8589,N_6364,N_6272);
xnor U8590 (N_8590,N_5162,N_5611);
and U8591 (N_8591,N_6109,N_5130);
or U8592 (N_8592,N_5902,N_7312);
xor U8593 (N_8593,N_5689,N_6572);
nand U8594 (N_8594,N_5184,N_5148);
and U8595 (N_8595,N_5878,N_5999);
xor U8596 (N_8596,N_7187,N_7304);
xor U8597 (N_8597,N_5204,N_5268);
nor U8598 (N_8598,N_6985,N_5001);
and U8599 (N_8599,N_6135,N_6316);
xnor U8600 (N_8600,N_5423,N_5430);
xor U8601 (N_8601,N_7199,N_5254);
nor U8602 (N_8602,N_5498,N_5709);
nand U8603 (N_8603,N_6766,N_6508);
or U8604 (N_8604,N_7185,N_6242);
nor U8605 (N_8605,N_5176,N_7057);
and U8606 (N_8606,N_5444,N_5717);
and U8607 (N_8607,N_6693,N_6543);
or U8608 (N_8608,N_5738,N_7053);
xnor U8609 (N_8609,N_6749,N_5575);
nand U8610 (N_8610,N_7430,N_6356);
xor U8611 (N_8611,N_6454,N_5249);
and U8612 (N_8612,N_5384,N_7173);
xor U8613 (N_8613,N_6049,N_5942);
xnor U8614 (N_8614,N_5731,N_5017);
nor U8615 (N_8615,N_6943,N_5458);
and U8616 (N_8616,N_7094,N_5004);
nand U8617 (N_8617,N_7413,N_6056);
xnor U8618 (N_8618,N_5333,N_5454);
nor U8619 (N_8619,N_5154,N_5933);
xnor U8620 (N_8620,N_7324,N_7133);
nand U8621 (N_8621,N_6721,N_6418);
and U8622 (N_8622,N_6596,N_7021);
or U8623 (N_8623,N_5400,N_7266);
nand U8624 (N_8624,N_5756,N_6876);
nor U8625 (N_8625,N_5532,N_5647);
or U8626 (N_8626,N_5605,N_5896);
and U8627 (N_8627,N_5715,N_5838);
nor U8628 (N_8628,N_6776,N_5325);
or U8629 (N_8629,N_6308,N_6054);
xnor U8630 (N_8630,N_6541,N_7147);
xnor U8631 (N_8631,N_5008,N_6645);
and U8632 (N_8632,N_6309,N_7111);
nand U8633 (N_8633,N_6839,N_7467);
nand U8634 (N_8634,N_5360,N_5419);
or U8635 (N_8635,N_5885,N_5303);
nand U8636 (N_8636,N_6389,N_6228);
or U8637 (N_8637,N_5678,N_6002);
or U8638 (N_8638,N_6310,N_6180);
nand U8639 (N_8639,N_6934,N_5040);
or U8640 (N_8640,N_7208,N_5608);
xor U8641 (N_8641,N_6186,N_5765);
xor U8642 (N_8642,N_5036,N_5776);
nor U8643 (N_8643,N_5381,N_7330);
nor U8644 (N_8644,N_7290,N_6218);
xor U8645 (N_8645,N_5683,N_5067);
or U8646 (N_8646,N_5301,N_6441);
nor U8647 (N_8647,N_6097,N_6657);
xor U8648 (N_8648,N_6586,N_5937);
nor U8649 (N_8649,N_6298,N_7120);
xor U8650 (N_8650,N_6836,N_6844);
nand U8651 (N_8651,N_6740,N_5104);
nand U8652 (N_8652,N_5085,N_6680);
nand U8653 (N_8653,N_5729,N_6234);
nor U8654 (N_8654,N_6527,N_6788);
and U8655 (N_8655,N_7006,N_5592);
or U8656 (N_8656,N_5710,N_7049);
nor U8657 (N_8657,N_6005,N_6278);
and U8658 (N_8658,N_6096,N_6908);
nor U8659 (N_8659,N_5157,N_5062);
and U8660 (N_8660,N_7344,N_5222);
nor U8661 (N_8661,N_7411,N_5504);
nand U8662 (N_8662,N_6491,N_6696);
or U8663 (N_8663,N_6034,N_5799);
or U8664 (N_8664,N_5028,N_7440);
and U8665 (N_8665,N_5928,N_7064);
nand U8666 (N_8666,N_5179,N_7224);
xnor U8667 (N_8667,N_6396,N_7231);
and U8668 (N_8668,N_5243,N_6037);
nand U8669 (N_8669,N_6265,N_6629);
and U8670 (N_8670,N_6960,N_6488);
and U8671 (N_8671,N_6303,N_5474);
and U8672 (N_8672,N_7436,N_7219);
and U8673 (N_8673,N_5456,N_7408);
xnor U8674 (N_8674,N_6237,N_7161);
xor U8675 (N_8675,N_7149,N_5449);
and U8676 (N_8676,N_6539,N_6905);
xnor U8677 (N_8677,N_6147,N_6292);
nand U8678 (N_8678,N_5869,N_5226);
or U8679 (N_8679,N_7433,N_6751);
or U8680 (N_8680,N_5818,N_5425);
nor U8681 (N_8681,N_5147,N_5599);
or U8682 (N_8682,N_5558,N_6051);
nand U8683 (N_8683,N_5316,N_5212);
and U8684 (N_8684,N_6990,N_5577);
nor U8685 (N_8685,N_6497,N_6296);
nand U8686 (N_8686,N_6450,N_5905);
xor U8687 (N_8687,N_5407,N_7175);
nor U8688 (N_8688,N_5525,N_5940);
nand U8689 (N_8689,N_6323,N_6834);
nor U8690 (N_8690,N_5662,N_6968);
and U8691 (N_8691,N_7246,N_5658);
nand U8692 (N_8692,N_7479,N_6670);
nor U8693 (N_8693,N_5842,N_6368);
xor U8694 (N_8694,N_6115,N_6931);
or U8695 (N_8695,N_6624,N_5481);
or U8696 (N_8696,N_7204,N_6500);
and U8697 (N_8697,N_5565,N_6411);
and U8698 (N_8698,N_7485,N_5918);
or U8699 (N_8699,N_5042,N_5616);
nand U8700 (N_8700,N_5389,N_5209);
and U8701 (N_8701,N_6720,N_5007);
and U8702 (N_8702,N_6717,N_6453);
nand U8703 (N_8703,N_6076,N_7273);
xor U8704 (N_8704,N_7268,N_6262);
xnor U8705 (N_8705,N_6569,N_6577);
nor U8706 (N_8706,N_6030,N_5319);
or U8707 (N_8707,N_5980,N_7048);
nand U8708 (N_8708,N_7085,N_5281);
nor U8709 (N_8709,N_6831,N_6544);
nor U8710 (N_8710,N_6192,N_6796);
or U8711 (N_8711,N_5779,N_6478);
nand U8712 (N_8712,N_5370,N_6075);
nand U8713 (N_8713,N_6615,N_5771);
or U8714 (N_8714,N_7242,N_7139);
nor U8715 (N_8715,N_5021,N_6191);
and U8716 (N_8716,N_6903,N_7407);
or U8717 (N_8717,N_5537,N_5789);
nand U8718 (N_8718,N_6226,N_7080);
nand U8719 (N_8719,N_6403,N_5517);
nor U8720 (N_8720,N_6223,N_5126);
xor U8721 (N_8721,N_5589,N_6270);
nand U8722 (N_8722,N_6591,N_6311);
or U8723 (N_8723,N_6913,N_5663);
nor U8724 (N_8724,N_6698,N_6331);
xnor U8725 (N_8725,N_6360,N_7343);
xnor U8726 (N_8726,N_6846,N_7072);
nand U8727 (N_8727,N_5960,N_5994);
xnor U8728 (N_8728,N_6420,N_6927);
nand U8729 (N_8729,N_6078,N_6465);
and U8730 (N_8730,N_6472,N_5095);
nand U8731 (N_8731,N_5132,N_5421);
and U8732 (N_8732,N_5003,N_5795);
and U8733 (N_8733,N_6414,N_7453);
or U8734 (N_8734,N_5661,N_5754);
xor U8735 (N_8735,N_6589,N_7018);
nor U8736 (N_8736,N_5380,N_6695);
xor U8737 (N_8737,N_7365,N_5307);
and U8738 (N_8738,N_7401,N_7039);
xor U8739 (N_8739,N_5139,N_6867);
xor U8740 (N_8740,N_5452,N_6062);
nor U8741 (N_8741,N_5752,N_6241);
and U8742 (N_8742,N_5707,N_6600);
and U8743 (N_8743,N_6965,N_6503);
nand U8744 (N_8744,N_5649,N_7420);
xnor U8745 (N_8745,N_5374,N_7452);
xnor U8746 (N_8746,N_6006,N_7259);
xor U8747 (N_8747,N_6649,N_6432);
or U8748 (N_8748,N_6190,N_6916);
nor U8749 (N_8749,N_6390,N_5094);
nor U8750 (N_8750,N_7106,N_6588);
nor U8751 (N_8751,N_5747,N_5428);
nand U8752 (N_8752,N_5237,N_6902);
nor U8753 (N_8753,N_5569,N_6683);
xor U8754 (N_8754,N_6289,N_7005);
nor U8755 (N_8755,N_5867,N_6395);
xnor U8756 (N_8756,N_5588,N_5777);
xor U8757 (N_8757,N_7345,N_5214);
xor U8758 (N_8758,N_7380,N_6437);
nor U8759 (N_8759,N_6030,N_5939);
nand U8760 (N_8760,N_5067,N_6946);
and U8761 (N_8761,N_6024,N_5066);
nand U8762 (N_8762,N_5920,N_5739);
or U8763 (N_8763,N_6833,N_5592);
and U8764 (N_8764,N_5593,N_6908);
xor U8765 (N_8765,N_7377,N_7265);
nor U8766 (N_8766,N_7216,N_7482);
or U8767 (N_8767,N_6933,N_6918);
nor U8768 (N_8768,N_5469,N_7119);
xnor U8769 (N_8769,N_5742,N_5584);
xnor U8770 (N_8770,N_6332,N_6930);
nor U8771 (N_8771,N_6220,N_7055);
nand U8772 (N_8772,N_6426,N_5198);
nand U8773 (N_8773,N_6182,N_6375);
and U8774 (N_8774,N_7001,N_6890);
and U8775 (N_8775,N_5512,N_6862);
or U8776 (N_8776,N_5000,N_5514);
nor U8777 (N_8777,N_6882,N_5984);
xor U8778 (N_8778,N_5705,N_7070);
nand U8779 (N_8779,N_5917,N_7044);
and U8780 (N_8780,N_6514,N_5747);
and U8781 (N_8781,N_7460,N_6617);
and U8782 (N_8782,N_6169,N_5300);
xnor U8783 (N_8783,N_6701,N_6712);
nor U8784 (N_8784,N_7167,N_6687);
nand U8785 (N_8785,N_7038,N_6281);
or U8786 (N_8786,N_6131,N_5011);
nand U8787 (N_8787,N_5900,N_5195);
xor U8788 (N_8788,N_6183,N_5371);
nor U8789 (N_8789,N_5188,N_5371);
nand U8790 (N_8790,N_6817,N_7164);
nor U8791 (N_8791,N_5470,N_6465);
or U8792 (N_8792,N_6834,N_7191);
nand U8793 (N_8793,N_5936,N_7405);
xor U8794 (N_8794,N_7064,N_5990);
or U8795 (N_8795,N_7077,N_7371);
nand U8796 (N_8796,N_5078,N_6688);
nor U8797 (N_8797,N_5781,N_6247);
or U8798 (N_8798,N_7047,N_5790);
nor U8799 (N_8799,N_5666,N_5922);
nand U8800 (N_8800,N_5128,N_6512);
nor U8801 (N_8801,N_6326,N_7440);
nor U8802 (N_8802,N_6895,N_5471);
nand U8803 (N_8803,N_5429,N_7212);
and U8804 (N_8804,N_6907,N_7493);
or U8805 (N_8805,N_5128,N_5342);
xnor U8806 (N_8806,N_7329,N_6867);
nor U8807 (N_8807,N_6081,N_5961);
and U8808 (N_8808,N_5877,N_7115);
nand U8809 (N_8809,N_6373,N_5476);
nand U8810 (N_8810,N_7201,N_6296);
xor U8811 (N_8811,N_5628,N_5010);
nand U8812 (N_8812,N_6265,N_5424);
xor U8813 (N_8813,N_6114,N_7250);
and U8814 (N_8814,N_6571,N_6864);
and U8815 (N_8815,N_5998,N_5283);
nor U8816 (N_8816,N_6333,N_6547);
or U8817 (N_8817,N_7080,N_6247);
and U8818 (N_8818,N_5264,N_5853);
or U8819 (N_8819,N_7146,N_6649);
nor U8820 (N_8820,N_5965,N_6664);
or U8821 (N_8821,N_5154,N_5259);
or U8822 (N_8822,N_6774,N_6116);
nor U8823 (N_8823,N_6190,N_6475);
nand U8824 (N_8824,N_6743,N_6310);
nand U8825 (N_8825,N_7075,N_5700);
nand U8826 (N_8826,N_5290,N_7017);
nor U8827 (N_8827,N_6552,N_5744);
or U8828 (N_8828,N_6591,N_5311);
xnor U8829 (N_8829,N_6622,N_5905);
nand U8830 (N_8830,N_6862,N_6678);
xnor U8831 (N_8831,N_7213,N_7088);
or U8832 (N_8832,N_6692,N_7345);
xnor U8833 (N_8833,N_6291,N_5090);
or U8834 (N_8834,N_7453,N_5253);
xor U8835 (N_8835,N_6009,N_5528);
xnor U8836 (N_8836,N_6996,N_5980);
nor U8837 (N_8837,N_7217,N_7162);
xor U8838 (N_8838,N_7201,N_5641);
xnor U8839 (N_8839,N_7200,N_6746);
or U8840 (N_8840,N_6961,N_6937);
and U8841 (N_8841,N_7206,N_6604);
or U8842 (N_8842,N_5091,N_6393);
nor U8843 (N_8843,N_7484,N_7218);
nand U8844 (N_8844,N_5816,N_5727);
nand U8845 (N_8845,N_5195,N_6169);
nor U8846 (N_8846,N_7498,N_5926);
nand U8847 (N_8847,N_7235,N_6232);
nor U8848 (N_8848,N_5468,N_7346);
xor U8849 (N_8849,N_6263,N_7143);
and U8850 (N_8850,N_5019,N_5203);
and U8851 (N_8851,N_6770,N_6003);
xor U8852 (N_8852,N_5012,N_7252);
nand U8853 (N_8853,N_5664,N_5398);
and U8854 (N_8854,N_5649,N_7202);
nand U8855 (N_8855,N_6772,N_6179);
and U8856 (N_8856,N_7379,N_6683);
nor U8857 (N_8857,N_6342,N_6502);
nor U8858 (N_8858,N_5674,N_5763);
nor U8859 (N_8859,N_7162,N_6201);
xor U8860 (N_8860,N_7474,N_7082);
nand U8861 (N_8861,N_6631,N_7197);
xnor U8862 (N_8862,N_6150,N_6606);
or U8863 (N_8863,N_7177,N_7420);
or U8864 (N_8864,N_7101,N_6991);
nand U8865 (N_8865,N_6103,N_6507);
xnor U8866 (N_8866,N_6344,N_6529);
nor U8867 (N_8867,N_5437,N_5295);
or U8868 (N_8868,N_6904,N_5805);
nor U8869 (N_8869,N_6117,N_5737);
xor U8870 (N_8870,N_5452,N_7020);
xnor U8871 (N_8871,N_5889,N_7366);
nor U8872 (N_8872,N_5992,N_6735);
nand U8873 (N_8873,N_6885,N_7057);
nand U8874 (N_8874,N_5643,N_5500);
xor U8875 (N_8875,N_5307,N_6962);
or U8876 (N_8876,N_6688,N_5571);
nor U8877 (N_8877,N_6078,N_6837);
nor U8878 (N_8878,N_5918,N_6336);
nand U8879 (N_8879,N_6440,N_6262);
or U8880 (N_8880,N_5587,N_6190);
nor U8881 (N_8881,N_5141,N_6181);
nor U8882 (N_8882,N_6314,N_6093);
nor U8883 (N_8883,N_7131,N_5682);
nand U8884 (N_8884,N_5945,N_5503);
and U8885 (N_8885,N_6133,N_6608);
or U8886 (N_8886,N_6801,N_7174);
nand U8887 (N_8887,N_5373,N_5383);
xor U8888 (N_8888,N_6846,N_7074);
and U8889 (N_8889,N_7432,N_5681);
and U8890 (N_8890,N_7092,N_7117);
or U8891 (N_8891,N_5861,N_5115);
or U8892 (N_8892,N_6666,N_5615);
nor U8893 (N_8893,N_6605,N_5961);
xor U8894 (N_8894,N_7450,N_7438);
and U8895 (N_8895,N_7156,N_7223);
or U8896 (N_8896,N_6567,N_6216);
or U8897 (N_8897,N_6644,N_6570);
or U8898 (N_8898,N_6531,N_6930);
xor U8899 (N_8899,N_5102,N_6409);
nand U8900 (N_8900,N_5928,N_5894);
nor U8901 (N_8901,N_6005,N_6870);
and U8902 (N_8902,N_5020,N_7204);
nor U8903 (N_8903,N_6390,N_6132);
xor U8904 (N_8904,N_5123,N_5328);
xnor U8905 (N_8905,N_5395,N_5974);
nor U8906 (N_8906,N_6866,N_6114);
or U8907 (N_8907,N_5635,N_6866);
or U8908 (N_8908,N_7340,N_7128);
and U8909 (N_8909,N_7155,N_5340);
or U8910 (N_8910,N_5825,N_6510);
nor U8911 (N_8911,N_6964,N_5797);
nand U8912 (N_8912,N_6634,N_6946);
and U8913 (N_8913,N_5722,N_5591);
or U8914 (N_8914,N_5811,N_7411);
nand U8915 (N_8915,N_5432,N_5396);
nand U8916 (N_8916,N_5455,N_6668);
or U8917 (N_8917,N_5851,N_5561);
nor U8918 (N_8918,N_7215,N_6444);
and U8919 (N_8919,N_5445,N_6447);
xnor U8920 (N_8920,N_5117,N_6620);
xnor U8921 (N_8921,N_5710,N_6397);
or U8922 (N_8922,N_5094,N_5089);
xnor U8923 (N_8923,N_6116,N_7347);
xor U8924 (N_8924,N_6702,N_6309);
and U8925 (N_8925,N_5551,N_6055);
and U8926 (N_8926,N_5771,N_6574);
nand U8927 (N_8927,N_7009,N_7165);
and U8928 (N_8928,N_6671,N_5712);
or U8929 (N_8929,N_5793,N_7081);
xnor U8930 (N_8930,N_6943,N_5352);
nor U8931 (N_8931,N_6765,N_6647);
nor U8932 (N_8932,N_5178,N_5021);
and U8933 (N_8933,N_7457,N_7318);
xor U8934 (N_8934,N_5972,N_5347);
nor U8935 (N_8935,N_6455,N_6489);
or U8936 (N_8936,N_6730,N_6274);
or U8937 (N_8937,N_5812,N_6601);
xnor U8938 (N_8938,N_6229,N_6157);
nor U8939 (N_8939,N_6426,N_6743);
nor U8940 (N_8940,N_6530,N_6168);
xnor U8941 (N_8941,N_5851,N_5332);
nor U8942 (N_8942,N_7066,N_6228);
nor U8943 (N_8943,N_5320,N_7375);
nand U8944 (N_8944,N_6319,N_5991);
xnor U8945 (N_8945,N_5208,N_7375);
xor U8946 (N_8946,N_5233,N_5473);
or U8947 (N_8947,N_7222,N_7313);
nor U8948 (N_8948,N_5274,N_5692);
nor U8949 (N_8949,N_5415,N_6408);
or U8950 (N_8950,N_7048,N_6563);
nand U8951 (N_8951,N_7184,N_5269);
nand U8952 (N_8952,N_7383,N_5025);
xnor U8953 (N_8953,N_6416,N_5082);
nand U8954 (N_8954,N_5010,N_7079);
xor U8955 (N_8955,N_6160,N_7339);
xnor U8956 (N_8956,N_7408,N_6593);
and U8957 (N_8957,N_5631,N_6051);
nor U8958 (N_8958,N_6821,N_5781);
and U8959 (N_8959,N_5040,N_5234);
xor U8960 (N_8960,N_6679,N_7315);
nor U8961 (N_8961,N_7035,N_5070);
nand U8962 (N_8962,N_5938,N_6131);
and U8963 (N_8963,N_5737,N_5409);
nand U8964 (N_8964,N_6478,N_5351);
xnor U8965 (N_8965,N_6901,N_7082);
xor U8966 (N_8966,N_6442,N_6897);
or U8967 (N_8967,N_5222,N_5320);
xnor U8968 (N_8968,N_6628,N_6765);
or U8969 (N_8969,N_6255,N_7193);
or U8970 (N_8970,N_6093,N_6770);
or U8971 (N_8971,N_6008,N_6291);
nor U8972 (N_8972,N_6833,N_6955);
nand U8973 (N_8973,N_5588,N_5643);
and U8974 (N_8974,N_6732,N_5610);
and U8975 (N_8975,N_6901,N_6450);
nor U8976 (N_8976,N_5632,N_6461);
nor U8977 (N_8977,N_6340,N_6273);
nand U8978 (N_8978,N_5989,N_6531);
nor U8979 (N_8979,N_6059,N_5493);
nand U8980 (N_8980,N_7322,N_6652);
nand U8981 (N_8981,N_6627,N_6206);
nand U8982 (N_8982,N_5859,N_6617);
xnor U8983 (N_8983,N_6646,N_5970);
nand U8984 (N_8984,N_5350,N_5858);
xnor U8985 (N_8985,N_6277,N_6859);
and U8986 (N_8986,N_5728,N_7088);
or U8987 (N_8987,N_7213,N_5485);
xor U8988 (N_8988,N_5567,N_6205);
nor U8989 (N_8989,N_7409,N_7312);
and U8990 (N_8990,N_6806,N_6827);
or U8991 (N_8991,N_5540,N_5220);
or U8992 (N_8992,N_5056,N_5444);
or U8993 (N_8993,N_5162,N_6045);
or U8994 (N_8994,N_5835,N_6048);
and U8995 (N_8995,N_5894,N_5381);
or U8996 (N_8996,N_7005,N_5117);
and U8997 (N_8997,N_5684,N_6919);
nor U8998 (N_8998,N_6689,N_6146);
nand U8999 (N_8999,N_5266,N_7167);
nand U9000 (N_9000,N_7426,N_5298);
nor U9001 (N_9001,N_5898,N_5795);
nor U9002 (N_9002,N_6759,N_6804);
nor U9003 (N_9003,N_6085,N_6470);
nand U9004 (N_9004,N_6421,N_7443);
xor U9005 (N_9005,N_5127,N_5121);
xor U9006 (N_9006,N_5734,N_6975);
xnor U9007 (N_9007,N_6259,N_6029);
nand U9008 (N_9008,N_6125,N_7229);
nor U9009 (N_9009,N_6757,N_5889);
or U9010 (N_9010,N_5886,N_6048);
or U9011 (N_9011,N_5166,N_5453);
xor U9012 (N_9012,N_6948,N_5680);
nand U9013 (N_9013,N_5858,N_6315);
xor U9014 (N_9014,N_6816,N_5860);
nand U9015 (N_9015,N_7076,N_6469);
and U9016 (N_9016,N_5397,N_6200);
nor U9017 (N_9017,N_5652,N_6110);
nor U9018 (N_9018,N_7175,N_7049);
xor U9019 (N_9019,N_6456,N_5261);
or U9020 (N_9020,N_5849,N_5162);
or U9021 (N_9021,N_7243,N_5869);
nand U9022 (N_9022,N_6995,N_5622);
nor U9023 (N_9023,N_7241,N_6075);
nand U9024 (N_9024,N_5102,N_7136);
nand U9025 (N_9025,N_6805,N_5411);
or U9026 (N_9026,N_6095,N_7131);
xor U9027 (N_9027,N_6580,N_5893);
and U9028 (N_9028,N_5494,N_5262);
and U9029 (N_9029,N_5514,N_5319);
and U9030 (N_9030,N_6010,N_7192);
or U9031 (N_9031,N_5773,N_5214);
xor U9032 (N_9032,N_7475,N_6745);
and U9033 (N_9033,N_6049,N_7472);
nor U9034 (N_9034,N_5948,N_6105);
nor U9035 (N_9035,N_5287,N_7421);
and U9036 (N_9036,N_5675,N_6218);
nor U9037 (N_9037,N_6764,N_6326);
nand U9038 (N_9038,N_7338,N_6123);
nand U9039 (N_9039,N_5180,N_6691);
nand U9040 (N_9040,N_5150,N_5335);
and U9041 (N_9041,N_6726,N_5881);
nor U9042 (N_9042,N_6669,N_5938);
nand U9043 (N_9043,N_5595,N_5868);
or U9044 (N_9044,N_7466,N_6185);
nor U9045 (N_9045,N_5200,N_7154);
xor U9046 (N_9046,N_6835,N_5549);
xor U9047 (N_9047,N_6146,N_7065);
or U9048 (N_9048,N_6299,N_6955);
or U9049 (N_9049,N_6387,N_6782);
nand U9050 (N_9050,N_6757,N_6501);
nand U9051 (N_9051,N_6152,N_6715);
and U9052 (N_9052,N_7009,N_7057);
nor U9053 (N_9053,N_5347,N_6321);
nand U9054 (N_9054,N_5830,N_7066);
or U9055 (N_9055,N_6875,N_5111);
and U9056 (N_9056,N_6867,N_6635);
xor U9057 (N_9057,N_5303,N_6376);
or U9058 (N_9058,N_6888,N_6836);
and U9059 (N_9059,N_5976,N_7035);
nand U9060 (N_9060,N_5890,N_7078);
xnor U9061 (N_9061,N_5776,N_6597);
or U9062 (N_9062,N_7463,N_6426);
and U9063 (N_9063,N_5771,N_6849);
xnor U9064 (N_9064,N_5839,N_5295);
nand U9065 (N_9065,N_7454,N_6357);
nor U9066 (N_9066,N_6999,N_7231);
xnor U9067 (N_9067,N_5113,N_6691);
and U9068 (N_9068,N_5055,N_6617);
and U9069 (N_9069,N_7028,N_5761);
xor U9070 (N_9070,N_6245,N_6532);
nor U9071 (N_9071,N_6155,N_5132);
xnor U9072 (N_9072,N_5186,N_6476);
nand U9073 (N_9073,N_7013,N_6641);
nand U9074 (N_9074,N_6118,N_6713);
and U9075 (N_9075,N_6894,N_5597);
or U9076 (N_9076,N_6298,N_5468);
and U9077 (N_9077,N_5011,N_7114);
nand U9078 (N_9078,N_7480,N_6696);
nand U9079 (N_9079,N_5058,N_7420);
nand U9080 (N_9080,N_7304,N_5093);
or U9081 (N_9081,N_6785,N_5412);
or U9082 (N_9082,N_6189,N_7083);
nor U9083 (N_9083,N_5826,N_5947);
or U9084 (N_9084,N_6180,N_7235);
nand U9085 (N_9085,N_6419,N_5447);
xnor U9086 (N_9086,N_7069,N_7312);
nand U9087 (N_9087,N_5199,N_6118);
or U9088 (N_9088,N_7359,N_6870);
xnor U9089 (N_9089,N_5608,N_5647);
xnor U9090 (N_9090,N_5380,N_5357);
or U9091 (N_9091,N_6173,N_5555);
nand U9092 (N_9092,N_6526,N_5826);
nand U9093 (N_9093,N_6861,N_6565);
or U9094 (N_9094,N_6164,N_7444);
xnor U9095 (N_9095,N_5842,N_5239);
xor U9096 (N_9096,N_7423,N_7190);
xor U9097 (N_9097,N_5144,N_6525);
and U9098 (N_9098,N_6820,N_5746);
nand U9099 (N_9099,N_5825,N_6564);
nand U9100 (N_9100,N_7213,N_6983);
and U9101 (N_9101,N_5622,N_5614);
nand U9102 (N_9102,N_6122,N_6251);
and U9103 (N_9103,N_5502,N_6105);
nand U9104 (N_9104,N_5656,N_6164);
and U9105 (N_9105,N_6388,N_5997);
nand U9106 (N_9106,N_7492,N_7430);
nor U9107 (N_9107,N_5358,N_6148);
xnor U9108 (N_9108,N_5081,N_5997);
or U9109 (N_9109,N_5434,N_5311);
and U9110 (N_9110,N_5910,N_5973);
nor U9111 (N_9111,N_6806,N_6264);
and U9112 (N_9112,N_5612,N_5659);
xnor U9113 (N_9113,N_5103,N_7076);
and U9114 (N_9114,N_5979,N_7102);
nor U9115 (N_9115,N_7002,N_5683);
nor U9116 (N_9116,N_5515,N_7299);
xnor U9117 (N_9117,N_5319,N_6362);
and U9118 (N_9118,N_5893,N_6092);
nand U9119 (N_9119,N_6283,N_5042);
and U9120 (N_9120,N_5012,N_6964);
nand U9121 (N_9121,N_6174,N_6160);
nor U9122 (N_9122,N_5622,N_5867);
xor U9123 (N_9123,N_5462,N_7229);
or U9124 (N_9124,N_5968,N_7143);
or U9125 (N_9125,N_5078,N_5726);
nand U9126 (N_9126,N_6821,N_5453);
xnor U9127 (N_9127,N_6486,N_7024);
or U9128 (N_9128,N_6477,N_7298);
nor U9129 (N_9129,N_7064,N_7087);
nor U9130 (N_9130,N_6151,N_5428);
xor U9131 (N_9131,N_5237,N_6807);
or U9132 (N_9132,N_5301,N_6804);
xnor U9133 (N_9133,N_7413,N_6744);
nand U9134 (N_9134,N_6771,N_5462);
or U9135 (N_9135,N_7065,N_5931);
nand U9136 (N_9136,N_6821,N_6467);
and U9137 (N_9137,N_5637,N_6422);
nand U9138 (N_9138,N_7427,N_6929);
or U9139 (N_9139,N_6294,N_5709);
nor U9140 (N_9140,N_5295,N_6881);
and U9141 (N_9141,N_7260,N_5972);
and U9142 (N_9142,N_6204,N_6500);
xnor U9143 (N_9143,N_5644,N_5167);
nand U9144 (N_9144,N_6824,N_5974);
or U9145 (N_9145,N_6500,N_5969);
nand U9146 (N_9146,N_5243,N_7469);
and U9147 (N_9147,N_7360,N_6948);
nand U9148 (N_9148,N_5022,N_7219);
or U9149 (N_9149,N_7441,N_5580);
nand U9150 (N_9150,N_6150,N_5211);
and U9151 (N_9151,N_6394,N_6140);
xnor U9152 (N_9152,N_6632,N_7206);
and U9153 (N_9153,N_6742,N_6463);
nand U9154 (N_9154,N_5696,N_5600);
nor U9155 (N_9155,N_6209,N_7310);
nor U9156 (N_9156,N_5823,N_6516);
or U9157 (N_9157,N_7250,N_6571);
or U9158 (N_9158,N_6269,N_7362);
and U9159 (N_9159,N_7019,N_6552);
or U9160 (N_9160,N_6649,N_5364);
or U9161 (N_9161,N_5176,N_5136);
nor U9162 (N_9162,N_5205,N_5453);
xor U9163 (N_9163,N_6351,N_5932);
and U9164 (N_9164,N_6084,N_7388);
or U9165 (N_9165,N_5964,N_6585);
or U9166 (N_9166,N_5083,N_5152);
xor U9167 (N_9167,N_6631,N_5723);
and U9168 (N_9168,N_5803,N_5686);
xnor U9169 (N_9169,N_7104,N_7417);
nor U9170 (N_9170,N_5223,N_5978);
nor U9171 (N_9171,N_7002,N_7023);
nand U9172 (N_9172,N_5202,N_6976);
and U9173 (N_9173,N_7192,N_6323);
xor U9174 (N_9174,N_6832,N_6123);
xor U9175 (N_9175,N_5837,N_6017);
nand U9176 (N_9176,N_5966,N_6406);
nor U9177 (N_9177,N_6859,N_6499);
nand U9178 (N_9178,N_7271,N_6481);
xnor U9179 (N_9179,N_7299,N_5781);
xnor U9180 (N_9180,N_6276,N_7327);
nand U9181 (N_9181,N_7408,N_5854);
and U9182 (N_9182,N_7277,N_6834);
nor U9183 (N_9183,N_7435,N_7279);
xnor U9184 (N_9184,N_7365,N_6102);
or U9185 (N_9185,N_6561,N_7236);
and U9186 (N_9186,N_6229,N_7453);
or U9187 (N_9187,N_5929,N_6542);
or U9188 (N_9188,N_5014,N_6462);
or U9189 (N_9189,N_5318,N_5209);
or U9190 (N_9190,N_6836,N_6277);
or U9191 (N_9191,N_6171,N_5890);
nand U9192 (N_9192,N_5635,N_6659);
xnor U9193 (N_9193,N_5218,N_5593);
or U9194 (N_9194,N_7164,N_5572);
and U9195 (N_9195,N_5524,N_5240);
and U9196 (N_9196,N_6680,N_5399);
and U9197 (N_9197,N_5375,N_6391);
nand U9198 (N_9198,N_5132,N_5589);
or U9199 (N_9199,N_7494,N_5115);
nand U9200 (N_9200,N_5488,N_7341);
xnor U9201 (N_9201,N_7381,N_6391);
xor U9202 (N_9202,N_7408,N_6611);
or U9203 (N_9203,N_5238,N_6158);
xor U9204 (N_9204,N_7157,N_6336);
or U9205 (N_9205,N_5379,N_5530);
xor U9206 (N_9206,N_5678,N_6436);
nor U9207 (N_9207,N_5199,N_6913);
and U9208 (N_9208,N_5398,N_5386);
nand U9209 (N_9209,N_5157,N_5151);
nor U9210 (N_9210,N_6488,N_7170);
nand U9211 (N_9211,N_6997,N_7356);
and U9212 (N_9212,N_6007,N_6902);
nand U9213 (N_9213,N_5786,N_5586);
and U9214 (N_9214,N_6390,N_5815);
nand U9215 (N_9215,N_6343,N_5246);
xor U9216 (N_9216,N_5303,N_6882);
nor U9217 (N_9217,N_5862,N_6283);
and U9218 (N_9218,N_6417,N_5052);
nand U9219 (N_9219,N_5060,N_6409);
nor U9220 (N_9220,N_6483,N_6053);
nor U9221 (N_9221,N_6220,N_5094);
nor U9222 (N_9222,N_5663,N_5145);
nand U9223 (N_9223,N_6462,N_5642);
xor U9224 (N_9224,N_5198,N_7066);
xnor U9225 (N_9225,N_5703,N_6703);
nand U9226 (N_9226,N_6602,N_6279);
or U9227 (N_9227,N_5244,N_5706);
and U9228 (N_9228,N_7321,N_6297);
or U9229 (N_9229,N_6151,N_5600);
nand U9230 (N_9230,N_6238,N_7249);
and U9231 (N_9231,N_5422,N_6866);
nor U9232 (N_9232,N_5938,N_5158);
nor U9233 (N_9233,N_5389,N_5148);
or U9234 (N_9234,N_6112,N_6888);
nor U9235 (N_9235,N_7134,N_7145);
nand U9236 (N_9236,N_7047,N_5665);
or U9237 (N_9237,N_5705,N_5729);
nor U9238 (N_9238,N_6822,N_6172);
nand U9239 (N_9239,N_5966,N_5416);
nand U9240 (N_9240,N_5409,N_5997);
xor U9241 (N_9241,N_6165,N_6504);
nor U9242 (N_9242,N_6696,N_5086);
nand U9243 (N_9243,N_6344,N_7087);
nand U9244 (N_9244,N_7129,N_5370);
nand U9245 (N_9245,N_6998,N_5009);
nand U9246 (N_9246,N_6577,N_6236);
or U9247 (N_9247,N_6471,N_5056);
or U9248 (N_9248,N_5419,N_6125);
or U9249 (N_9249,N_6963,N_6495);
nor U9250 (N_9250,N_7079,N_5174);
and U9251 (N_9251,N_7017,N_5379);
or U9252 (N_9252,N_7384,N_5457);
or U9253 (N_9253,N_6610,N_7278);
nand U9254 (N_9254,N_7068,N_7151);
and U9255 (N_9255,N_5097,N_6258);
xnor U9256 (N_9256,N_5520,N_6480);
xnor U9257 (N_9257,N_5491,N_6380);
xnor U9258 (N_9258,N_6006,N_7288);
nor U9259 (N_9259,N_5349,N_5944);
and U9260 (N_9260,N_7153,N_6099);
or U9261 (N_9261,N_6556,N_5942);
nand U9262 (N_9262,N_6232,N_7061);
nor U9263 (N_9263,N_6245,N_6502);
nand U9264 (N_9264,N_7466,N_5663);
xnor U9265 (N_9265,N_5029,N_5081);
or U9266 (N_9266,N_6517,N_6810);
nand U9267 (N_9267,N_6005,N_7443);
nor U9268 (N_9268,N_6360,N_5695);
nor U9269 (N_9269,N_6792,N_6795);
nor U9270 (N_9270,N_7179,N_5033);
xor U9271 (N_9271,N_6554,N_5825);
xnor U9272 (N_9272,N_7263,N_7042);
xnor U9273 (N_9273,N_5088,N_5560);
xnor U9274 (N_9274,N_7160,N_7075);
and U9275 (N_9275,N_6236,N_6699);
nor U9276 (N_9276,N_7110,N_5694);
xnor U9277 (N_9277,N_7453,N_6242);
nand U9278 (N_9278,N_5133,N_6298);
xor U9279 (N_9279,N_5017,N_5782);
nor U9280 (N_9280,N_7135,N_5452);
xnor U9281 (N_9281,N_7212,N_5087);
xnor U9282 (N_9282,N_6148,N_6653);
xnor U9283 (N_9283,N_6857,N_5252);
nand U9284 (N_9284,N_5849,N_5755);
xnor U9285 (N_9285,N_7031,N_7178);
nor U9286 (N_9286,N_5746,N_5045);
or U9287 (N_9287,N_7100,N_5644);
or U9288 (N_9288,N_7200,N_5966);
xor U9289 (N_9289,N_6888,N_7447);
nor U9290 (N_9290,N_7140,N_5088);
xor U9291 (N_9291,N_5413,N_6297);
nor U9292 (N_9292,N_6624,N_6702);
nand U9293 (N_9293,N_6774,N_5466);
or U9294 (N_9294,N_6700,N_7318);
nor U9295 (N_9295,N_6815,N_5412);
and U9296 (N_9296,N_6049,N_5435);
nand U9297 (N_9297,N_6445,N_7273);
xnor U9298 (N_9298,N_6908,N_7346);
nor U9299 (N_9299,N_5852,N_6675);
and U9300 (N_9300,N_6946,N_5304);
or U9301 (N_9301,N_7090,N_6277);
or U9302 (N_9302,N_6936,N_5499);
nor U9303 (N_9303,N_5877,N_5543);
or U9304 (N_9304,N_5077,N_6825);
and U9305 (N_9305,N_6666,N_7112);
nor U9306 (N_9306,N_6043,N_5534);
and U9307 (N_9307,N_7265,N_7451);
or U9308 (N_9308,N_7177,N_6678);
nor U9309 (N_9309,N_7035,N_6846);
xor U9310 (N_9310,N_6327,N_5158);
nor U9311 (N_9311,N_5531,N_7088);
or U9312 (N_9312,N_7272,N_5073);
and U9313 (N_9313,N_5645,N_7358);
nand U9314 (N_9314,N_6583,N_6584);
nor U9315 (N_9315,N_6485,N_6126);
xnor U9316 (N_9316,N_6999,N_6661);
or U9317 (N_9317,N_6800,N_7196);
nand U9318 (N_9318,N_6176,N_5480);
and U9319 (N_9319,N_5461,N_7207);
nor U9320 (N_9320,N_5269,N_7268);
or U9321 (N_9321,N_6878,N_6348);
or U9322 (N_9322,N_6574,N_5185);
or U9323 (N_9323,N_5486,N_6212);
or U9324 (N_9324,N_7253,N_7211);
xnor U9325 (N_9325,N_5668,N_6154);
and U9326 (N_9326,N_7409,N_5777);
nand U9327 (N_9327,N_6933,N_5239);
nand U9328 (N_9328,N_5793,N_7424);
and U9329 (N_9329,N_5522,N_5734);
or U9330 (N_9330,N_6390,N_5689);
or U9331 (N_9331,N_6817,N_6038);
nor U9332 (N_9332,N_6198,N_6925);
xor U9333 (N_9333,N_5511,N_5653);
nor U9334 (N_9334,N_6196,N_6506);
and U9335 (N_9335,N_7280,N_6616);
and U9336 (N_9336,N_5816,N_7132);
or U9337 (N_9337,N_5992,N_6956);
or U9338 (N_9338,N_6672,N_5671);
or U9339 (N_9339,N_5288,N_5305);
or U9340 (N_9340,N_5134,N_6473);
nor U9341 (N_9341,N_5707,N_5588);
nand U9342 (N_9342,N_7320,N_6566);
and U9343 (N_9343,N_6883,N_6254);
nand U9344 (N_9344,N_5681,N_6971);
nor U9345 (N_9345,N_5793,N_7009);
nor U9346 (N_9346,N_7343,N_7191);
xnor U9347 (N_9347,N_5386,N_7197);
nor U9348 (N_9348,N_6431,N_7051);
and U9349 (N_9349,N_6376,N_6531);
xnor U9350 (N_9350,N_7027,N_6499);
xnor U9351 (N_9351,N_5411,N_5092);
nor U9352 (N_9352,N_6722,N_7420);
nor U9353 (N_9353,N_6294,N_6476);
and U9354 (N_9354,N_5983,N_6088);
nand U9355 (N_9355,N_5108,N_5589);
and U9356 (N_9356,N_5500,N_7169);
nor U9357 (N_9357,N_6727,N_6732);
nand U9358 (N_9358,N_7370,N_6739);
nor U9359 (N_9359,N_6558,N_7240);
nor U9360 (N_9360,N_5729,N_6921);
and U9361 (N_9361,N_7005,N_6316);
xnor U9362 (N_9362,N_7276,N_5719);
and U9363 (N_9363,N_6113,N_5410);
nor U9364 (N_9364,N_5099,N_5909);
nand U9365 (N_9365,N_5858,N_6777);
or U9366 (N_9366,N_7133,N_6774);
and U9367 (N_9367,N_6638,N_6776);
or U9368 (N_9368,N_5111,N_5302);
nor U9369 (N_9369,N_7177,N_7257);
xor U9370 (N_9370,N_5289,N_7032);
xnor U9371 (N_9371,N_5551,N_7437);
nor U9372 (N_9372,N_5709,N_7304);
nand U9373 (N_9373,N_5213,N_7498);
nor U9374 (N_9374,N_6562,N_5332);
nand U9375 (N_9375,N_5753,N_6514);
or U9376 (N_9376,N_7046,N_5212);
xnor U9377 (N_9377,N_6523,N_6926);
xor U9378 (N_9378,N_6946,N_5963);
or U9379 (N_9379,N_5637,N_7006);
or U9380 (N_9380,N_6695,N_7176);
xnor U9381 (N_9381,N_5522,N_6683);
xnor U9382 (N_9382,N_6995,N_5437);
and U9383 (N_9383,N_7074,N_7324);
nor U9384 (N_9384,N_5918,N_7285);
nand U9385 (N_9385,N_6107,N_5597);
or U9386 (N_9386,N_5425,N_6636);
and U9387 (N_9387,N_6194,N_6810);
or U9388 (N_9388,N_6145,N_5270);
xor U9389 (N_9389,N_5124,N_5346);
and U9390 (N_9390,N_5804,N_5022);
or U9391 (N_9391,N_7207,N_6709);
nand U9392 (N_9392,N_6428,N_6680);
xnor U9393 (N_9393,N_6119,N_5692);
and U9394 (N_9394,N_7381,N_5760);
nor U9395 (N_9395,N_6882,N_5967);
xor U9396 (N_9396,N_5186,N_6433);
or U9397 (N_9397,N_6888,N_6754);
and U9398 (N_9398,N_7290,N_5963);
or U9399 (N_9399,N_5753,N_6763);
or U9400 (N_9400,N_7023,N_5685);
xnor U9401 (N_9401,N_5607,N_5815);
and U9402 (N_9402,N_5958,N_6518);
nor U9403 (N_9403,N_6499,N_7401);
nor U9404 (N_9404,N_5351,N_6640);
xnor U9405 (N_9405,N_6681,N_5789);
xnor U9406 (N_9406,N_5310,N_7481);
nor U9407 (N_9407,N_6767,N_6610);
nor U9408 (N_9408,N_5282,N_5794);
nor U9409 (N_9409,N_7392,N_6579);
nand U9410 (N_9410,N_5440,N_6646);
or U9411 (N_9411,N_7025,N_5993);
or U9412 (N_9412,N_6348,N_6072);
nand U9413 (N_9413,N_5394,N_6021);
xor U9414 (N_9414,N_6116,N_5042);
or U9415 (N_9415,N_5578,N_5301);
nand U9416 (N_9416,N_6435,N_6480);
xnor U9417 (N_9417,N_5888,N_6060);
or U9418 (N_9418,N_5017,N_7298);
or U9419 (N_9419,N_6798,N_5013);
or U9420 (N_9420,N_7015,N_7150);
and U9421 (N_9421,N_7219,N_5727);
xnor U9422 (N_9422,N_7398,N_5253);
or U9423 (N_9423,N_6114,N_5448);
xor U9424 (N_9424,N_7370,N_5035);
and U9425 (N_9425,N_6837,N_6219);
nand U9426 (N_9426,N_6851,N_6127);
and U9427 (N_9427,N_5591,N_7112);
nor U9428 (N_9428,N_6711,N_7297);
nor U9429 (N_9429,N_6967,N_5937);
and U9430 (N_9430,N_6566,N_5810);
nand U9431 (N_9431,N_6462,N_6609);
or U9432 (N_9432,N_6041,N_6891);
and U9433 (N_9433,N_7495,N_5909);
nor U9434 (N_9434,N_5380,N_5809);
or U9435 (N_9435,N_7279,N_5375);
and U9436 (N_9436,N_5547,N_6530);
nor U9437 (N_9437,N_5381,N_7040);
nor U9438 (N_9438,N_5018,N_6429);
xor U9439 (N_9439,N_5853,N_6670);
or U9440 (N_9440,N_6594,N_6990);
xor U9441 (N_9441,N_6304,N_6841);
nand U9442 (N_9442,N_6011,N_6321);
xor U9443 (N_9443,N_6782,N_7402);
or U9444 (N_9444,N_5025,N_5646);
and U9445 (N_9445,N_5971,N_5829);
nand U9446 (N_9446,N_5737,N_5629);
or U9447 (N_9447,N_5508,N_6210);
or U9448 (N_9448,N_5789,N_6335);
and U9449 (N_9449,N_7349,N_6381);
or U9450 (N_9450,N_6707,N_7194);
or U9451 (N_9451,N_6864,N_5188);
and U9452 (N_9452,N_6671,N_6667);
or U9453 (N_9453,N_6632,N_6627);
xnor U9454 (N_9454,N_6294,N_5313);
xnor U9455 (N_9455,N_6955,N_5281);
xor U9456 (N_9456,N_5185,N_6106);
nor U9457 (N_9457,N_5150,N_5632);
nand U9458 (N_9458,N_5879,N_6376);
or U9459 (N_9459,N_5869,N_6660);
nor U9460 (N_9460,N_5053,N_5915);
or U9461 (N_9461,N_5048,N_6584);
or U9462 (N_9462,N_7312,N_5081);
xor U9463 (N_9463,N_5027,N_7423);
xnor U9464 (N_9464,N_6373,N_6733);
or U9465 (N_9465,N_6723,N_6860);
or U9466 (N_9466,N_6593,N_7439);
xor U9467 (N_9467,N_6161,N_6568);
or U9468 (N_9468,N_5291,N_6297);
xnor U9469 (N_9469,N_6452,N_5505);
xnor U9470 (N_9470,N_5506,N_5427);
and U9471 (N_9471,N_6199,N_5246);
or U9472 (N_9472,N_6439,N_6627);
nor U9473 (N_9473,N_5989,N_5888);
and U9474 (N_9474,N_5772,N_5145);
xnor U9475 (N_9475,N_6891,N_6308);
or U9476 (N_9476,N_6791,N_5023);
and U9477 (N_9477,N_5856,N_6458);
nand U9478 (N_9478,N_5005,N_5796);
nor U9479 (N_9479,N_6887,N_6384);
nor U9480 (N_9480,N_7098,N_6054);
xor U9481 (N_9481,N_5264,N_6018);
or U9482 (N_9482,N_6401,N_6193);
nand U9483 (N_9483,N_6792,N_7478);
and U9484 (N_9484,N_5628,N_6236);
and U9485 (N_9485,N_7094,N_7342);
xor U9486 (N_9486,N_7226,N_6858);
or U9487 (N_9487,N_6850,N_6436);
or U9488 (N_9488,N_5700,N_5561);
or U9489 (N_9489,N_6593,N_5677);
and U9490 (N_9490,N_6118,N_5143);
and U9491 (N_9491,N_6973,N_5055);
nand U9492 (N_9492,N_6526,N_5094);
or U9493 (N_9493,N_7028,N_5078);
or U9494 (N_9494,N_7093,N_5738);
xor U9495 (N_9495,N_6053,N_6252);
nor U9496 (N_9496,N_6358,N_6498);
nand U9497 (N_9497,N_7399,N_5463);
or U9498 (N_9498,N_6108,N_6472);
or U9499 (N_9499,N_7219,N_6262);
nand U9500 (N_9500,N_5286,N_6527);
xor U9501 (N_9501,N_5313,N_5898);
nor U9502 (N_9502,N_5013,N_5344);
and U9503 (N_9503,N_6616,N_6703);
or U9504 (N_9504,N_6499,N_5148);
nand U9505 (N_9505,N_7119,N_5561);
or U9506 (N_9506,N_5771,N_5589);
nand U9507 (N_9507,N_6479,N_5754);
and U9508 (N_9508,N_7225,N_5065);
and U9509 (N_9509,N_7261,N_6145);
nor U9510 (N_9510,N_5364,N_6215);
nand U9511 (N_9511,N_5966,N_6777);
or U9512 (N_9512,N_6553,N_6099);
xnor U9513 (N_9513,N_5875,N_5506);
or U9514 (N_9514,N_7289,N_6189);
xor U9515 (N_9515,N_7432,N_5613);
nand U9516 (N_9516,N_5932,N_6683);
and U9517 (N_9517,N_7379,N_6564);
and U9518 (N_9518,N_6640,N_5047);
or U9519 (N_9519,N_6908,N_6357);
xor U9520 (N_9520,N_5701,N_5786);
nand U9521 (N_9521,N_5383,N_6308);
xnor U9522 (N_9522,N_7153,N_6209);
nor U9523 (N_9523,N_6142,N_5150);
nor U9524 (N_9524,N_5814,N_5025);
xnor U9525 (N_9525,N_6173,N_6537);
nand U9526 (N_9526,N_5303,N_7420);
nor U9527 (N_9527,N_6391,N_5885);
nor U9528 (N_9528,N_5993,N_5683);
or U9529 (N_9529,N_7033,N_5703);
nor U9530 (N_9530,N_7472,N_7066);
and U9531 (N_9531,N_7212,N_5873);
or U9532 (N_9532,N_5220,N_5199);
or U9533 (N_9533,N_6616,N_7294);
xnor U9534 (N_9534,N_6585,N_5483);
nor U9535 (N_9535,N_6570,N_7297);
xor U9536 (N_9536,N_7021,N_5020);
nor U9537 (N_9537,N_5294,N_7116);
xnor U9538 (N_9538,N_6355,N_6417);
and U9539 (N_9539,N_7246,N_5562);
nor U9540 (N_9540,N_7026,N_5638);
nor U9541 (N_9541,N_6330,N_6701);
nand U9542 (N_9542,N_5459,N_5138);
nor U9543 (N_9543,N_5693,N_5245);
xor U9544 (N_9544,N_6968,N_6963);
or U9545 (N_9545,N_7104,N_6527);
and U9546 (N_9546,N_6823,N_7066);
and U9547 (N_9547,N_5449,N_6143);
nor U9548 (N_9548,N_5198,N_5469);
nor U9549 (N_9549,N_7204,N_7344);
xor U9550 (N_9550,N_5713,N_5262);
or U9551 (N_9551,N_5132,N_7486);
xnor U9552 (N_9552,N_5462,N_7394);
and U9553 (N_9553,N_7107,N_6519);
and U9554 (N_9554,N_6676,N_5021);
xnor U9555 (N_9555,N_7043,N_6252);
nand U9556 (N_9556,N_6579,N_7364);
or U9557 (N_9557,N_5545,N_6346);
xnor U9558 (N_9558,N_5424,N_5994);
nor U9559 (N_9559,N_6228,N_7394);
nand U9560 (N_9560,N_6319,N_7271);
nand U9561 (N_9561,N_7225,N_6125);
and U9562 (N_9562,N_7105,N_7244);
nand U9563 (N_9563,N_6534,N_6212);
nand U9564 (N_9564,N_5233,N_5458);
or U9565 (N_9565,N_5853,N_5367);
xnor U9566 (N_9566,N_5085,N_5123);
or U9567 (N_9567,N_5571,N_5465);
xor U9568 (N_9568,N_6682,N_5255);
and U9569 (N_9569,N_6905,N_6729);
and U9570 (N_9570,N_6422,N_5528);
nand U9571 (N_9571,N_7176,N_5172);
xor U9572 (N_9572,N_6027,N_6762);
xnor U9573 (N_9573,N_6772,N_6471);
xnor U9574 (N_9574,N_6449,N_7388);
nor U9575 (N_9575,N_6807,N_7418);
xor U9576 (N_9576,N_5895,N_7014);
xor U9577 (N_9577,N_5784,N_6768);
or U9578 (N_9578,N_6754,N_6408);
xor U9579 (N_9579,N_6034,N_6770);
nand U9580 (N_9580,N_6867,N_6965);
xnor U9581 (N_9581,N_5887,N_6908);
nor U9582 (N_9582,N_5114,N_5320);
xnor U9583 (N_9583,N_5508,N_6680);
nand U9584 (N_9584,N_6188,N_6031);
and U9585 (N_9585,N_6978,N_5462);
nand U9586 (N_9586,N_6300,N_7055);
and U9587 (N_9587,N_5356,N_6834);
nor U9588 (N_9588,N_6316,N_5850);
nand U9589 (N_9589,N_5928,N_7129);
nand U9590 (N_9590,N_7383,N_5970);
nand U9591 (N_9591,N_6551,N_5369);
nor U9592 (N_9592,N_6054,N_6652);
nor U9593 (N_9593,N_6914,N_6535);
and U9594 (N_9594,N_6368,N_5793);
xor U9595 (N_9595,N_5230,N_6794);
xor U9596 (N_9596,N_6864,N_5833);
and U9597 (N_9597,N_7213,N_7345);
nand U9598 (N_9598,N_5563,N_7030);
xor U9599 (N_9599,N_5058,N_6168);
nor U9600 (N_9600,N_7066,N_7397);
and U9601 (N_9601,N_7202,N_6824);
xor U9602 (N_9602,N_5756,N_5967);
or U9603 (N_9603,N_5559,N_5307);
and U9604 (N_9604,N_6628,N_5871);
nor U9605 (N_9605,N_7150,N_7102);
and U9606 (N_9606,N_5917,N_5250);
nor U9607 (N_9607,N_7279,N_5299);
nand U9608 (N_9608,N_7147,N_5122);
nand U9609 (N_9609,N_7193,N_5793);
and U9610 (N_9610,N_5753,N_5603);
and U9611 (N_9611,N_6204,N_5596);
xnor U9612 (N_9612,N_5295,N_5599);
xnor U9613 (N_9613,N_7192,N_6136);
nor U9614 (N_9614,N_6562,N_6180);
and U9615 (N_9615,N_7441,N_7131);
xnor U9616 (N_9616,N_5008,N_7035);
nor U9617 (N_9617,N_6064,N_6568);
nor U9618 (N_9618,N_5874,N_5944);
and U9619 (N_9619,N_7045,N_7127);
xor U9620 (N_9620,N_7112,N_6066);
or U9621 (N_9621,N_5772,N_7131);
nand U9622 (N_9622,N_5806,N_6463);
xnor U9623 (N_9623,N_5741,N_7279);
nor U9624 (N_9624,N_7130,N_5838);
nor U9625 (N_9625,N_6910,N_5233);
nand U9626 (N_9626,N_6171,N_6969);
nor U9627 (N_9627,N_7399,N_6302);
nor U9628 (N_9628,N_6268,N_7373);
nor U9629 (N_9629,N_5743,N_6877);
nor U9630 (N_9630,N_5031,N_6414);
xnor U9631 (N_9631,N_5949,N_6465);
nor U9632 (N_9632,N_7176,N_5663);
nand U9633 (N_9633,N_5153,N_5781);
nand U9634 (N_9634,N_5036,N_7250);
nor U9635 (N_9635,N_7270,N_6147);
xor U9636 (N_9636,N_5542,N_6090);
nand U9637 (N_9637,N_5378,N_6982);
xor U9638 (N_9638,N_7144,N_6415);
and U9639 (N_9639,N_6209,N_5437);
and U9640 (N_9640,N_5985,N_5055);
and U9641 (N_9641,N_5544,N_5812);
and U9642 (N_9642,N_5963,N_7331);
nand U9643 (N_9643,N_6935,N_7053);
and U9644 (N_9644,N_7229,N_5580);
nand U9645 (N_9645,N_7442,N_6405);
or U9646 (N_9646,N_7132,N_7484);
or U9647 (N_9647,N_5305,N_6682);
or U9648 (N_9648,N_6259,N_5500);
and U9649 (N_9649,N_6546,N_6371);
nand U9650 (N_9650,N_5173,N_5310);
nand U9651 (N_9651,N_5448,N_6471);
xor U9652 (N_9652,N_5816,N_6606);
nand U9653 (N_9653,N_6849,N_6320);
nand U9654 (N_9654,N_5625,N_5027);
or U9655 (N_9655,N_5429,N_6979);
nand U9656 (N_9656,N_6015,N_6681);
or U9657 (N_9657,N_5411,N_7035);
xnor U9658 (N_9658,N_5704,N_7390);
nor U9659 (N_9659,N_5553,N_6316);
xor U9660 (N_9660,N_6865,N_5353);
or U9661 (N_9661,N_5247,N_5861);
nor U9662 (N_9662,N_5915,N_6701);
xor U9663 (N_9663,N_7395,N_7378);
xnor U9664 (N_9664,N_6039,N_5491);
nor U9665 (N_9665,N_6254,N_5734);
or U9666 (N_9666,N_6847,N_6071);
nor U9667 (N_9667,N_7048,N_5765);
and U9668 (N_9668,N_6341,N_6568);
or U9669 (N_9669,N_6114,N_6923);
and U9670 (N_9670,N_7472,N_7304);
nor U9671 (N_9671,N_6436,N_6452);
xnor U9672 (N_9672,N_6495,N_6014);
or U9673 (N_9673,N_5501,N_7038);
or U9674 (N_9674,N_6298,N_6175);
nand U9675 (N_9675,N_7211,N_5540);
and U9676 (N_9676,N_5171,N_5319);
and U9677 (N_9677,N_5982,N_5079);
nor U9678 (N_9678,N_5499,N_7479);
nand U9679 (N_9679,N_7130,N_7105);
nor U9680 (N_9680,N_5500,N_5715);
nand U9681 (N_9681,N_5860,N_6490);
nor U9682 (N_9682,N_5960,N_5350);
nor U9683 (N_9683,N_6188,N_6745);
nor U9684 (N_9684,N_5035,N_6796);
nand U9685 (N_9685,N_6856,N_6328);
and U9686 (N_9686,N_7148,N_7325);
nor U9687 (N_9687,N_5739,N_5962);
nor U9688 (N_9688,N_6784,N_5130);
nand U9689 (N_9689,N_6339,N_5553);
nand U9690 (N_9690,N_5321,N_7041);
nor U9691 (N_9691,N_5321,N_7352);
or U9692 (N_9692,N_6834,N_5639);
nor U9693 (N_9693,N_7227,N_5002);
and U9694 (N_9694,N_7196,N_5492);
or U9695 (N_9695,N_5916,N_6971);
or U9696 (N_9696,N_5669,N_6848);
or U9697 (N_9697,N_5466,N_7089);
and U9698 (N_9698,N_7341,N_5828);
and U9699 (N_9699,N_5406,N_5608);
nand U9700 (N_9700,N_6181,N_5566);
nor U9701 (N_9701,N_5771,N_7255);
nand U9702 (N_9702,N_6216,N_7427);
xor U9703 (N_9703,N_5571,N_6641);
xnor U9704 (N_9704,N_5482,N_6203);
nand U9705 (N_9705,N_6272,N_5109);
xnor U9706 (N_9706,N_5504,N_5907);
and U9707 (N_9707,N_5986,N_6054);
nand U9708 (N_9708,N_6531,N_6390);
nand U9709 (N_9709,N_5885,N_5581);
nand U9710 (N_9710,N_5782,N_7320);
nand U9711 (N_9711,N_5278,N_5353);
nor U9712 (N_9712,N_5317,N_6740);
xor U9713 (N_9713,N_6560,N_7151);
nor U9714 (N_9714,N_5694,N_5692);
and U9715 (N_9715,N_6985,N_5711);
xor U9716 (N_9716,N_5127,N_6941);
nor U9717 (N_9717,N_6652,N_7068);
and U9718 (N_9718,N_5119,N_5725);
nor U9719 (N_9719,N_7161,N_7082);
nor U9720 (N_9720,N_5900,N_6688);
or U9721 (N_9721,N_5910,N_7346);
nand U9722 (N_9722,N_5585,N_7272);
nor U9723 (N_9723,N_6631,N_5247);
nor U9724 (N_9724,N_7367,N_7473);
nand U9725 (N_9725,N_6059,N_7218);
nand U9726 (N_9726,N_5088,N_7061);
nand U9727 (N_9727,N_6963,N_7476);
nand U9728 (N_9728,N_7193,N_6472);
and U9729 (N_9729,N_6915,N_5239);
or U9730 (N_9730,N_5453,N_6482);
nor U9731 (N_9731,N_6239,N_5711);
nand U9732 (N_9732,N_6709,N_5737);
nand U9733 (N_9733,N_6147,N_6006);
or U9734 (N_9734,N_5587,N_7020);
nand U9735 (N_9735,N_5781,N_5497);
nor U9736 (N_9736,N_5216,N_7290);
nand U9737 (N_9737,N_5419,N_6817);
xnor U9738 (N_9738,N_6852,N_5453);
nand U9739 (N_9739,N_5663,N_5160);
or U9740 (N_9740,N_5155,N_6129);
or U9741 (N_9741,N_6067,N_6562);
and U9742 (N_9742,N_7278,N_5646);
nand U9743 (N_9743,N_5004,N_5101);
xor U9744 (N_9744,N_6237,N_5181);
xnor U9745 (N_9745,N_7226,N_7311);
xnor U9746 (N_9746,N_6693,N_5174);
xor U9747 (N_9747,N_6012,N_5009);
and U9748 (N_9748,N_5333,N_6967);
nor U9749 (N_9749,N_5894,N_7198);
and U9750 (N_9750,N_7223,N_6164);
or U9751 (N_9751,N_5701,N_6334);
or U9752 (N_9752,N_6412,N_7004);
nand U9753 (N_9753,N_5254,N_6193);
or U9754 (N_9754,N_5366,N_7160);
or U9755 (N_9755,N_6012,N_5477);
nand U9756 (N_9756,N_6151,N_6144);
nor U9757 (N_9757,N_6727,N_7131);
and U9758 (N_9758,N_7358,N_6083);
nand U9759 (N_9759,N_6407,N_6768);
nand U9760 (N_9760,N_5556,N_6574);
nand U9761 (N_9761,N_5938,N_7360);
and U9762 (N_9762,N_5764,N_5371);
xnor U9763 (N_9763,N_6303,N_5598);
nor U9764 (N_9764,N_5707,N_6365);
nor U9765 (N_9765,N_6531,N_5270);
or U9766 (N_9766,N_5011,N_5704);
nand U9767 (N_9767,N_5560,N_6621);
nand U9768 (N_9768,N_6805,N_5258);
and U9769 (N_9769,N_6171,N_6504);
xor U9770 (N_9770,N_6560,N_5093);
xor U9771 (N_9771,N_6430,N_5782);
nor U9772 (N_9772,N_6866,N_7227);
or U9773 (N_9773,N_6617,N_6129);
nand U9774 (N_9774,N_5882,N_7080);
xor U9775 (N_9775,N_6829,N_5316);
xnor U9776 (N_9776,N_7110,N_5953);
nand U9777 (N_9777,N_6727,N_7281);
or U9778 (N_9778,N_5120,N_6923);
xnor U9779 (N_9779,N_7047,N_6700);
nor U9780 (N_9780,N_6888,N_7398);
or U9781 (N_9781,N_5259,N_6115);
and U9782 (N_9782,N_7348,N_5830);
nand U9783 (N_9783,N_6800,N_6092);
and U9784 (N_9784,N_5621,N_7330);
nor U9785 (N_9785,N_6695,N_6069);
nor U9786 (N_9786,N_6799,N_5766);
nor U9787 (N_9787,N_6537,N_6551);
or U9788 (N_9788,N_7381,N_7114);
nor U9789 (N_9789,N_6062,N_7253);
and U9790 (N_9790,N_5175,N_5503);
nand U9791 (N_9791,N_7229,N_7312);
nand U9792 (N_9792,N_7151,N_5390);
and U9793 (N_9793,N_6629,N_5479);
nor U9794 (N_9794,N_6084,N_5979);
nand U9795 (N_9795,N_7137,N_6102);
nand U9796 (N_9796,N_6008,N_6011);
xnor U9797 (N_9797,N_5663,N_6055);
xnor U9798 (N_9798,N_5933,N_5838);
xor U9799 (N_9799,N_5483,N_6155);
xnor U9800 (N_9800,N_7067,N_5933);
nor U9801 (N_9801,N_5470,N_7255);
or U9802 (N_9802,N_7167,N_5106);
nor U9803 (N_9803,N_5924,N_5139);
or U9804 (N_9804,N_6209,N_5361);
nor U9805 (N_9805,N_5886,N_5319);
nand U9806 (N_9806,N_6966,N_5917);
and U9807 (N_9807,N_6156,N_7108);
nand U9808 (N_9808,N_6904,N_6414);
nand U9809 (N_9809,N_6806,N_7167);
nand U9810 (N_9810,N_6899,N_5415);
or U9811 (N_9811,N_6161,N_5069);
or U9812 (N_9812,N_5342,N_7213);
nand U9813 (N_9813,N_5598,N_5775);
xor U9814 (N_9814,N_7018,N_5243);
nor U9815 (N_9815,N_6456,N_5142);
nand U9816 (N_9816,N_6741,N_7012);
and U9817 (N_9817,N_6384,N_7092);
nor U9818 (N_9818,N_7178,N_5184);
nand U9819 (N_9819,N_7231,N_5843);
or U9820 (N_9820,N_7297,N_7127);
and U9821 (N_9821,N_5241,N_5938);
and U9822 (N_9822,N_5097,N_5999);
xor U9823 (N_9823,N_7251,N_7394);
and U9824 (N_9824,N_6415,N_6286);
and U9825 (N_9825,N_7457,N_7177);
xnor U9826 (N_9826,N_5883,N_7248);
nand U9827 (N_9827,N_7315,N_5140);
nand U9828 (N_9828,N_5410,N_6683);
nand U9829 (N_9829,N_7377,N_6036);
xor U9830 (N_9830,N_6204,N_6228);
and U9831 (N_9831,N_7100,N_6811);
or U9832 (N_9832,N_7335,N_6065);
xor U9833 (N_9833,N_5895,N_5553);
or U9834 (N_9834,N_5048,N_6266);
nor U9835 (N_9835,N_7018,N_6320);
and U9836 (N_9836,N_6303,N_6404);
or U9837 (N_9837,N_5228,N_5394);
or U9838 (N_9838,N_7119,N_6013);
and U9839 (N_9839,N_7176,N_7391);
xnor U9840 (N_9840,N_6801,N_6114);
and U9841 (N_9841,N_6443,N_7480);
nand U9842 (N_9842,N_5463,N_6253);
nand U9843 (N_9843,N_5134,N_5646);
xor U9844 (N_9844,N_6405,N_5381);
xnor U9845 (N_9845,N_6495,N_6998);
xor U9846 (N_9846,N_6135,N_5203);
nand U9847 (N_9847,N_6281,N_6625);
nor U9848 (N_9848,N_5892,N_7296);
or U9849 (N_9849,N_7199,N_5833);
xnor U9850 (N_9850,N_5804,N_5872);
nor U9851 (N_9851,N_5782,N_6415);
or U9852 (N_9852,N_6733,N_5860);
xnor U9853 (N_9853,N_5889,N_6726);
or U9854 (N_9854,N_5067,N_6195);
and U9855 (N_9855,N_7174,N_6053);
xnor U9856 (N_9856,N_5125,N_6641);
xnor U9857 (N_9857,N_5806,N_5499);
or U9858 (N_9858,N_5723,N_7170);
xor U9859 (N_9859,N_6260,N_5569);
nand U9860 (N_9860,N_6277,N_5698);
or U9861 (N_9861,N_6494,N_6247);
and U9862 (N_9862,N_7121,N_6042);
nand U9863 (N_9863,N_5482,N_5484);
nor U9864 (N_9864,N_6571,N_6308);
or U9865 (N_9865,N_7304,N_5575);
nor U9866 (N_9866,N_5284,N_6421);
or U9867 (N_9867,N_5162,N_7042);
nor U9868 (N_9868,N_6662,N_6560);
and U9869 (N_9869,N_6628,N_7176);
xor U9870 (N_9870,N_5414,N_7325);
or U9871 (N_9871,N_5344,N_6792);
nor U9872 (N_9872,N_5924,N_5872);
xor U9873 (N_9873,N_7495,N_5356);
nand U9874 (N_9874,N_7196,N_7200);
and U9875 (N_9875,N_5601,N_5306);
nand U9876 (N_9876,N_6961,N_5814);
nor U9877 (N_9877,N_6936,N_6397);
nor U9878 (N_9878,N_6847,N_7067);
or U9879 (N_9879,N_7419,N_6009);
nand U9880 (N_9880,N_5637,N_5885);
nor U9881 (N_9881,N_6439,N_5626);
nand U9882 (N_9882,N_5573,N_6397);
nor U9883 (N_9883,N_5366,N_5073);
nor U9884 (N_9884,N_5040,N_7176);
xor U9885 (N_9885,N_6211,N_6797);
or U9886 (N_9886,N_6115,N_5996);
nand U9887 (N_9887,N_6136,N_5001);
nand U9888 (N_9888,N_5338,N_5260);
xnor U9889 (N_9889,N_7032,N_6871);
nor U9890 (N_9890,N_6124,N_7234);
or U9891 (N_9891,N_6025,N_6982);
xnor U9892 (N_9892,N_7320,N_5405);
xnor U9893 (N_9893,N_6069,N_6740);
nor U9894 (N_9894,N_5478,N_6058);
and U9895 (N_9895,N_5915,N_5003);
and U9896 (N_9896,N_7416,N_6872);
xnor U9897 (N_9897,N_6638,N_5396);
or U9898 (N_9898,N_6792,N_7481);
nand U9899 (N_9899,N_7483,N_6404);
nand U9900 (N_9900,N_6029,N_5002);
xnor U9901 (N_9901,N_6440,N_6348);
and U9902 (N_9902,N_7295,N_6159);
xnor U9903 (N_9903,N_7007,N_6295);
xor U9904 (N_9904,N_6845,N_7062);
xor U9905 (N_9905,N_5005,N_6226);
nor U9906 (N_9906,N_5881,N_5671);
or U9907 (N_9907,N_5655,N_7148);
or U9908 (N_9908,N_7147,N_6684);
nand U9909 (N_9909,N_5435,N_5035);
xnor U9910 (N_9910,N_5029,N_6894);
or U9911 (N_9911,N_7162,N_7010);
and U9912 (N_9912,N_6100,N_5936);
and U9913 (N_9913,N_5652,N_5846);
and U9914 (N_9914,N_7046,N_6939);
xnor U9915 (N_9915,N_5118,N_6922);
xor U9916 (N_9916,N_5005,N_6053);
xnor U9917 (N_9917,N_6451,N_5127);
and U9918 (N_9918,N_6513,N_6049);
nand U9919 (N_9919,N_6538,N_5190);
and U9920 (N_9920,N_5680,N_6564);
or U9921 (N_9921,N_7470,N_5993);
nor U9922 (N_9922,N_6315,N_6654);
nand U9923 (N_9923,N_6090,N_7104);
nand U9924 (N_9924,N_6011,N_6862);
nor U9925 (N_9925,N_7287,N_7142);
and U9926 (N_9926,N_6663,N_7008);
or U9927 (N_9927,N_5529,N_6568);
nor U9928 (N_9928,N_6125,N_5563);
nand U9929 (N_9929,N_5106,N_6539);
or U9930 (N_9930,N_6059,N_6953);
xor U9931 (N_9931,N_7415,N_6198);
nor U9932 (N_9932,N_5089,N_7366);
and U9933 (N_9933,N_7322,N_7489);
xnor U9934 (N_9934,N_5352,N_5044);
xnor U9935 (N_9935,N_6394,N_6410);
and U9936 (N_9936,N_6416,N_6644);
and U9937 (N_9937,N_5479,N_6016);
and U9938 (N_9938,N_5690,N_6914);
nand U9939 (N_9939,N_7105,N_5437);
or U9940 (N_9940,N_7001,N_7234);
and U9941 (N_9941,N_6029,N_6765);
and U9942 (N_9942,N_6693,N_5495);
nor U9943 (N_9943,N_7121,N_6775);
or U9944 (N_9944,N_6811,N_5505);
or U9945 (N_9945,N_5764,N_7103);
nor U9946 (N_9946,N_7278,N_5833);
or U9947 (N_9947,N_6257,N_7220);
or U9948 (N_9948,N_6374,N_5628);
xor U9949 (N_9949,N_5776,N_7414);
nor U9950 (N_9950,N_5271,N_7300);
nor U9951 (N_9951,N_6556,N_5110);
xnor U9952 (N_9952,N_6666,N_5071);
nor U9953 (N_9953,N_5510,N_7024);
and U9954 (N_9954,N_5801,N_6595);
nand U9955 (N_9955,N_6896,N_6564);
or U9956 (N_9956,N_6785,N_6597);
xnor U9957 (N_9957,N_7422,N_5038);
or U9958 (N_9958,N_6689,N_6254);
nor U9959 (N_9959,N_5949,N_6876);
nand U9960 (N_9960,N_6933,N_6400);
nand U9961 (N_9961,N_7273,N_6589);
nor U9962 (N_9962,N_5764,N_6737);
and U9963 (N_9963,N_7188,N_6827);
and U9964 (N_9964,N_5882,N_7259);
nor U9965 (N_9965,N_5529,N_6717);
or U9966 (N_9966,N_5535,N_5607);
or U9967 (N_9967,N_6316,N_6118);
and U9968 (N_9968,N_7008,N_6646);
and U9969 (N_9969,N_7075,N_5655);
or U9970 (N_9970,N_6756,N_7104);
xor U9971 (N_9971,N_6164,N_7021);
xor U9972 (N_9972,N_7272,N_6281);
and U9973 (N_9973,N_5028,N_5570);
and U9974 (N_9974,N_6714,N_6744);
nor U9975 (N_9975,N_5686,N_6670);
nand U9976 (N_9976,N_6190,N_7188);
and U9977 (N_9977,N_7019,N_5389);
and U9978 (N_9978,N_7109,N_6733);
nand U9979 (N_9979,N_6583,N_5227);
nor U9980 (N_9980,N_7412,N_5122);
nor U9981 (N_9981,N_6798,N_5811);
nor U9982 (N_9982,N_6245,N_5317);
nor U9983 (N_9983,N_5872,N_5697);
nor U9984 (N_9984,N_5053,N_7046);
nor U9985 (N_9985,N_5749,N_6833);
nor U9986 (N_9986,N_6210,N_6512);
or U9987 (N_9987,N_6695,N_7493);
xor U9988 (N_9988,N_6658,N_6635);
xnor U9989 (N_9989,N_5574,N_7319);
and U9990 (N_9990,N_6878,N_6996);
nor U9991 (N_9991,N_6722,N_5057);
nor U9992 (N_9992,N_5258,N_6561);
nor U9993 (N_9993,N_6799,N_6959);
or U9994 (N_9994,N_6958,N_5934);
xor U9995 (N_9995,N_5490,N_6985);
or U9996 (N_9996,N_7223,N_5492);
or U9997 (N_9997,N_5505,N_6963);
nand U9998 (N_9998,N_7159,N_6897);
and U9999 (N_9999,N_7406,N_5600);
or UO_0 (O_0,N_9681,N_9947);
xor UO_1 (O_1,N_9858,N_8955);
nor UO_2 (O_2,N_8155,N_8312);
nor UO_3 (O_3,N_9691,N_9563);
xnor UO_4 (O_4,N_7545,N_7750);
or UO_5 (O_5,N_8068,N_8833);
xor UO_6 (O_6,N_8033,N_9803);
nand UO_7 (O_7,N_9688,N_9569);
or UO_8 (O_8,N_7866,N_9540);
xnor UO_9 (O_9,N_8158,N_9825);
xor UO_10 (O_10,N_8794,N_8115);
nor UO_11 (O_11,N_9103,N_7851);
nand UO_12 (O_12,N_9822,N_8821);
xor UO_13 (O_13,N_8101,N_9793);
nor UO_14 (O_14,N_9228,N_8313);
xor UO_15 (O_15,N_8686,N_9602);
nor UO_16 (O_16,N_9152,N_8746);
xor UO_17 (O_17,N_9154,N_7671);
nor UO_18 (O_18,N_8924,N_9525);
nor UO_19 (O_19,N_9375,N_8301);
nor UO_20 (O_20,N_9489,N_8465);
nor UO_21 (O_21,N_9266,N_9246);
nand UO_22 (O_22,N_7767,N_7602);
xnor UO_23 (O_23,N_8580,N_7631);
nor UO_24 (O_24,N_7939,N_8407);
nor UO_25 (O_25,N_8729,N_8903);
and UO_26 (O_26,N_7892,N_9811);
nor UO_27 (O_27,N_8309,N_8829);
nor UO_28 (O_28,N_7787,N_9172);
nor UO_29 (O_29,N_9659,N_9021);
nor UO_30 (O_30,N_9801,N_8627);
and UO_31 (O_31,N_9049,N_8736);
xor UO_32 (O_32,N_9549,N_9961);
and UO_33 (O_33,N_9839,N_7789);
nor UO_34 (O_34,N_9787,N_9080);
xor UO_35 (O_35,N_9548,N_9881);
nor UO_36 (O_36,N_7670,N_8933);
nor UO_37 (O_37,N_7616,N_8269);
nand UO_38 (O_38,N_8731,N_8723);
and UO_39 (O_39,N_9215,N_8106);
nor UO_40 (O_40,N_9187,N_8725);
and UO_41 (O_41,N_7501,N_7676);
xnor UO_42 (O_42,N_8298,N_8786);
and UO_43 (O_43,N_8830,N_9868);
nor UO_44 (O_44,N_8140,N_8343);
nor UO_45 (O_45,N_7765,N_7887);
and UO_46 (O_46,N_9675,N_8180);
nor UO_47 (O_47,N_7998,N_8117);
nand UO_48 (O_48,N_7827,N_8275);
nor UO_49 (O_49,N_7831,N_9272);
nor UO_50 (O_50,N_8677,N_7589);
nor UO_51 (O_51,N_9227,N_9698);
nor UO_52 (O_52,N_8041,N_9427);
nor UO_53 (O_53,N_9934,N_8133);
and UO_54 (O_54,N_9762,N_7563);
nand UO_55 (O_55,N_8369,N_8753);
and UO_56 (O_56,N_7500,N_9888);
and UO_57 (O_57,N_7693,N_9977);
or UO_58 (O_58,N_8505,N_8459);
and UO_59 (O_59,N_9588,N_7697);
xnor UO_60 (O_60,N_7841,N_9848);
xnor UO_61 (O_61,N_8286,N_8433);
nor UO_62 (O_62,N_8705,N_9336);
or UO_63 (O_63,N_8449,N_8385);
nor UO_64 (O_64,N_7856,N_8314);
xor UO_65 (O_65,N_9339,N_8111);
nor UO_66 (O_66,N_9054,N_9164);
or UO_67 (O_67,N_8405,N_7511);
xnor UO_68 (O_68,N_7510,N_8108);
xor UO_69 (O_69,N_8240,N_8262);
or UO_70 (O_70,N_7538,N_9233);
xnor UO_71 (O_71,N_9895,N_8531);
and UO_72 (O_72,N_7885,N_9778);
nor UO_73 (O_73,N_7595,N_9689);
or UO_74 (O_74,N_8857,N_7592);
or UO_75 (O_75,N_7632,N_9897);
nor UO_76 (O_76,N_8763,N_7682);
and UO_77 (O_77,N_8475,N_8975);
or UO_78 (O_78,N_8048,N_7803);
nand UO_79 (O_79,N_8522,N_7521);
nor UO_80 (O_80,N_9704,N_8495);
nor UO_81 (O_81,N_7915,N_9160);
xor UO_82 (O_82,N_9867,N_8342);
or UO_83 (O_83,N_8053,N_8675);
nor UO_84 (O_84,N_8610,N_8875);
and UO_85 (O_85,N_8581,N_7959);
and UO_86 (O_86,N_8819,N_8141);
nand UO_87 (O_87,N_9917,N_9758);
and UO_88 (O_88,N_9327,N_8653);
xnor UO_89 (O_89,N_9679,N_8907);
xor UO_90 (O_90,N_9650,N_8318);
or UO_91 (O_91,N_9518,N_8595);
and UO_92 (O_92,N_8165,N_8303);
nor UO_93 (O_93,N_7869,N_9996);
nor UO_94 (O_94,N_9557,N_8509);
or UO_95 (O_95,N_9517,N_9311);
xor UO_96 (O_96,N_8174,N_9815);
or UO_97 (O_97,N_9425,N_7728);
xor UO_98 (O_98,N_7871,N_8254);
nand UO_99 (O_99,N_8925,N_7516);
nor UO_100 (O_100,N_9429,N_8018);
nor UO_101 (O_101,N_8144,N_7677);
xnor UO_102 (O_102,N_8056,N_9504);
nand UO_103 (O_103,N_9285,N_8386);
or UO_104 (O_104,N_8119,N_7834);
or UO_105 (O_105,N_8584,N_8344);
xor UO_106 (O_106,N_9404,N_9220);
xnor UO_107 (O_107,N_8513,N_9855);
nand UO_108 (O_108,N_7822,N_8596);
and UO_109 (O_109,N_9728,N_7786);
xor UO_110 (O_110,N_7839,N_9929);
xor UO_111 (O_111,N_8035,N_9723);
nand UO_112 (O_112,N_9715,N_9886);
or UO_113 (O_113,N_7580,N_7925);
and UO_114 (O_114,N_8276,N_9909);
nor UO_115 (O_115,N_9705,N_8058);
xor UO_116 (O_116,N_8952,N_7539);
or UO_117 (O_117,N_7977,N_7986);
nand UO_118 (O_118,N_9457,N_9510);
or UO_119 (O_119,N_8066,N_9774);
or UO_120 (O_120,N_7819,N_7854);
nand UO_121 (O_121,N_9256,N_8431);
nor UO_122 (O_122,N_8444,N_9890);
nand UO_123 (O_123,N_9841,N_9821);
and UO_124 (O_124,N_9648,N_8381);
nand UO_125 (O_125,N_8109,N_7738);
or UO_126 (O_126,N_9291,N_8561);
nand UO_127 (O_127,N_9133,N_7881);
nor UO_128 (O_128,N_7691,N_7953);
xnor UO_129 (O_129,N_9029,N_7864);
nand UO_130 (O_130,N_9824,N_8556);
and UO_131 (O_131,N_8355,N_8977);
or UO_132 (O_132,N_8926,N_8965);
xnor UO_133 (O_133,N_8899,N_8599);
nor UO_134 (O_134,N_7720,N_9150);
and UO_135 (O_135,N_9100,N_8420);
or UO_136 (O_136,N_9075,N_8236);
xnor UO_137 (O_137,N_9282,N_8929);
and UO_138 (O_138,N_8438,N_8796);
nor UO_139 (O_139,N_7911,N_9694);
nor UO_140 (O_140,N_9610,N_8204);
or UO_141 (O_141,N_8942,N_8370);
xnor UO_142 (O_142,N_9112,N_9614);
or UO_143 (O_143,N_9725,N_8797);
nand UO_144 (O_144,N_9853,N_9230);
or UO_145 (O_145,N_7759,N_9907);
nand UO_146 (O_146,N_9345,N_9837);
nor UO_147 (O_147,N_9885,N_9414);
and UO_148 (O_148,N_8644,N_7544);
nor UO_149 (O_149,N_8597,N_9322);
xor UO_150 (O_150,N_8608,N_9446);
nor UO_151 (O_151,N_8574,N_9896);
xnor UO_152 (O_152,N_8146,N_9204);
nor UO_153 (O_153,N_9562,N_8970);
nand UO_154 (O_154,N_7771,N_7583);
and UO_155 (O_155,N_8223,N_9248);
nand UO_156 (O_156,N_8060,N_8569);
nand UO_157 (O_157,N_9524,N_7665);
or UO_158 (O_158,N_8194,N_8422);
nor UO_159 (O_159,N_8974,N_8589);
and UO_160 (O_160,N_9786,N_9229);
or UO_161 (O_161,N_8493,N_8266);
and UO_162 (O_162,N_7681,N_9009);
nand UO_163 (O_163,N_8643,N_9799);
or UO_164 (O_164,N_9773,N_7833);
and UO_165 (O_165,N_7782,N_8095);
and UO_166 (O_166,N_7941,N_9948);
nor UO_167 (O_167,N_9503,N_8568);
nor UO_168 (O_168,N_9341,N_7740);
nor UO_169 (O_169,N_9206,N_7794);
xnor UO_170 (O_170,N_8326,N_8429);
and UO_171 (O_171,N_8798,N_8618);
nor UO_172 (O_172,N_8220,N_9102);
nand UO_173 (O_173,N_7991,N_9059);
nand UO_174 (O_174,N_7659,N_7503);
nand UO_175 (O_175,N_8480,N_8500);
nor UO_176 (O_176,N_8553,N_8594);
and UO_177 (O_177,N_9861,N_8019);
xnor UO_178 (O_178,N_7893,N_8305);
nand UO_179 (O_179,N_8417,N_8206);
nand UO_180 (O_180,N_8349,N_9436);
and UO_181 (O_181,N_8674,N_7725);
nand UO_182 (O_182,N_9241,N_8613);
and UO_183 (O_183,N_9697,N_8982);
nor UO_184 (O_184,N_8157,N_8319);
or UO_185 (O_185,N_8792,N_8916);
and UO_186 (O_186,N_9768,N_9739);
or UO_187 (O_187,N_8815,N_8352);
and UO_188 (O_188,N_7591,N_9915);
nor UO_189 (O_189,N_7652,N_7969);
or UO_190 (O_190,N_9651,N_8196);
and UO_191 (O_191,N_7684,N_8171);
or UO_192 (O_192,N_9987,N_7690);
or UO_193 (O_193,N_7791,N_7774);
xor UO_194 (O_194,N_8912,N_7612);
and UO_195 (O_195,N_9488,N_8441);
nand UO_196 (O_196,N_9533,N_8722);
or UO_197 (O_197,N_9329,N_8107);
nand UO_198 (O_198,N_9912,N_9388);
or UO_199 (O_199,N_8414,N_9349);
xor UO_200 (O_200,N_7624,N_8772);
xnor UO_201 (O_201,N_8691,N_8470);
and UO_202 (O_202,N_8813,N_8550);
or UO_203 (O_203,N_7811,N_8964);
xor UO_204 (O_204,N_8463,N_9876);
xor UO_205 (O_205,N_8538,N_9367);
nand UO_206 (O_206,N_7916,N_9817);
xnor UO_207 (O_207,N_7743,N_9485);
xor UO_208 (O_208,N_9321,N_7549);
nand UO_209 (O_209,N_9862,N_8192);
nand UO_210 (O_210,N_8235,N_9911);
and UO_211 (O_211,N_8800,N_9142);
nand UO_212 (O_212,N_8064,N_9840);
nand UO_213 (O_213,N_7711,N_8423);
nand UO_214 (O_214,N_8714,N_9596);
or UO_215 (O_215,N_9835,N_8898);
or UO_216 (O_216,N_9083,N_8951);
nand UO_217 (O_217,N_8418,N_7999);
or UO_218 (O_218,N_9555,N_8866);
xnor UO_219 (O_219,N_8743,N_7513);
or UO_220 (O_220,N_9324,N_9070);
and UO_221 (O_221,N_7872,N_8049);
and UO_222 (O_222,N_9406,N_8973);
and UO_223 (O_223,N_9137,N_9226);
nor UO_224 (O_224,N_8372,N_9472);
or UO_225 (O_225,N_7927,N_8577);
and UO_226 (O_226,N_9209,N_8211);
and UO_227 (O_227,N_9985,N_7603);
nand UO_228 (O_228,N_9041,N_7519);
and UO_229 (O_229,N_9258,N_7918);
nand UO_230 (O_230,N_7975,N_7657);
xor UO_231 (O_231,N_8208,N_8219);
or UO_232 (O_232,N_8408,N_8900);
nor UO_233 (O_233,N_8249,N_7989);
nand UO_234 (O_234,N_9318,N_8255);
nand UO_235 (O_235,N_9802,N_9666);
and UO_236 (O_236,N_9539,N_7783);
or UO_237 (O_237,N_7809,N_9465);
and UO_238 (O_238,N_9086,N_8928);
and UO_239 (O_239,N_9293,N_9298);
nor UO_240 (O_240,N_9808,N_9968);
or UO_241 (O_241,N_8440,N_9294);
xnor UO_242 (O_242,N_7674,N_8591);
xnor UO_243 (O_243,N_7560,N_9036);
nand UO_244 (O_244,N_9594,N_8914);
or UO_245 (O_245,N_7997,N_8619);
xor UO_246 (O_246,N_8320,N_9893);
and UO_247 (O_247,N_7920,N_9119);
nand UO_248 (O_248,N_8003,N_8265);
nor UO_249 (O_249,N_8991,N_8862);
nor UO_250 (O_250,N_8810,N_9529);
xor UO_251 (O_251,N_7609,N_9714);
xor UO_252 (O_252,N_8185,N_9898);
xor UO_253 (O_253,N_8410,N_9900);
and UO_254 (O_254,N_9267,N_7733);
xnor UO_255 (O_255,N_9496,N_8766);
or UO_256 (O_256,N_9450,N_8084);
or UO_257 (O_257,N_8832,N_9173);
and UO_258 (O_258,N_9222,N_8946);
nand UO_259 (O_259,N_9490,N_8274);
xnor UO_260 (O_260,N_8181,N_7847);
nand UO_261 (O_261,N_7857,N_9995);
nor UO_262 (O_262,N_8879,N_8524);
xor UO_263 (O_263,N_9129,N_8555);
nor UO_264 (O_264,N_7570,N_7830);
or UO_265 (O_265,N_9359,N_8374);
and UO_266 (O_266,N_9292,N_9672);
nor UO_267 (O_267,N_7944,N_7983);
and UO_268 (O_268,N_8085,N_7636);
xnor UO_269 (O_269,N_8008,N_8840);
and UO_270 (O_270,N_8452,N_7528);
or UO_271 (O_271,N_9491,N_9348);
or UO_272 (O_272,N_8878,N_9880);
xor UO_273 (O_273,N_9175,N_9783);
nor UO_274 (O_274,N_9988,N_8757);
and UO_275 (O_275,N_9850,N_8189);
xnor UO_276 (O_276,N_8915,N_9983);
or UO_277 (O_277,N_9597,N_9584);
nor UO_278 (O_278,N_8708,N_8486);
or UO_279 (O_279,N_9168,N_8567);
xnor UO_280 (O_280,N_8961,N_8506);
and UO_281 (O_281,N_8329,N_9068);
xor UO_282 (O_282,N_7930,N_7994);
nand UO_283 (O_283,N_8934,N_9012);
nor UO_284 (O_284,N_8570,N_8163);
nand UO_285 (O_285,N_8241,N_9665);
or UO_286 (O_286,N_7565,N_9386);
nor UO_287 (O_287,N_8790,N_8016);
and UO_288 (O_288,N_9473,N_9186);
nor UO_289 (O_289,N_8153,N_7810);
nor UO_290 (O_290,N_8215,N_9600);
nand UO_291 (O_291,N_9875,N_9605);
xor UO_292 (O_292,N_8649,N_8118);
and UO_293 (O_293,N_8761,N_9537);
nor UO_294 (O_294,N_9952,N_8838);
or UO_295 (O_295,N_9066,N_8175);
xnor UO_296 (O_296,N_9501,N_8113);
nor UO_297 (O_297,N_7561,N_9125);
xnor UO_298 (O_298,N_8436,N_7798);
xor UO_299 (O_299,N_8998,N_8017);
xor UO_300 (O_300,N_8997,N_8388);
nand UO_301 (O_301,N_7817,N_8213);
nor UO_302 (O_302,N_9956,N_8062);
nand UO_303 (O_303,N_8839,N_8404);
and UO_304 (O_304,N_8086,N_9883);
or UO_305 (O_305,N_8870,N_9521);
and UO_306 (O_306,N_8477,N_9140);
xnor UO_307 (O_307,N_9471,N_8874);
nand UO_308 (O_308,N_7796,N_8411);
and UO_309 (O_309,N_7522,N_7897);
or UO_310 (O_310,N_9249,N_8406);
xor UO_311 (O_311,N_7970,N_8563);
or UO_312 (O_312,N_8300,N_7568);
and UO_313 (O_313,N_9287,N_9239);
xnor UO_314 (O_314,N_7962,N_8657);
nor UO_315 (O_315,N_8642,N_9699);
nand UO_316 (O_316,N_8076,N_9097);
or UO_317 (O_317,N_7751,N_8047);
and UO_318 (O_318,N_8634,N_9586);
nand UO_319 (O_319,N_8353,N_8345);
nand UO_320 (O_320,N_8983,N_9735);
and UO_321 (O_321,N_8519,N_9146);
nor UO_322 (O_322,N_9500,N_8639);
nand UO_323 (O_323,N_8079,N_7715);
and UO_324 (O_324,N_9202,N_7553);
and UO_325 (O_325,N_9703,N_8995);
or UO_326 (O_326,N_9194,N_9957);
and UO_327 (O_327,N_8384,N_9244);
and UO_328 (O_328,N_7778,N_9312);
nor UO_329 (O_329,N_9523,N_8947);
nor UO_330 (O_330,N_9709,N_9116);
nand UO_331 (O_331,N_8132,N_9343);
nand UO_332 (O_332,N_7643,N_7950);
xor UO_333 (O_333,N_8605,N_7523);
and UO_334 (O_334,N_8718,N_9531);
nor UO_335 (O_335,N_8823,N_8549);
or UO_336 (O_336,N_7701,N_9409);
and UO_337 (O_337,N_7762,N_9663);
nor UO_338 (O_338,N_9148,N_8738);
nand UO_339 (O_339,N_9015,N_8304);
nand UO_340 (O_340,N_9891,N_9039);
nand UO_341 (O_341,N_8195,N_8492);
nor UO_342 (O_342,N_8566,N_7926);
nor UO_343 (O_343,N_7635,N_8861);
or UO_344 (O_344,N_9637,N_9147);
nand UO_345 (O_345,N_8336,N_9314);
xnor UO_346 (O_346,N_7517,N_7683);
and UO_347 (O_347,N_9829,N_9767);
nand UO_348 (O_348,N_8460,N_8337);
nor UO_349 (O_349,N_9437,N_9397);
or UO_350 (O_350,N_7928,N_8707);
nand UO_351 (O_351,N_9544,N_9509);
nor UO_352 (O_352,N_9719,N_8360);
or UO_353 (O_353,N_9538,N_7747);
and UO_354 (O_354,N_8854,N_9731);
xnor UO_355 (O_355,N_8376,N_7601);
nand UO_356 (O_356,N_9914,N_7859);
xnor UO_357 (O_357,N_8902,N_8789);
and UO_358 (O_358,N_8804,N_7895);
or UO_359 (O_359,N_8869,N_9374);
nor UO_360 (O_360,N_9284,N_8424);
nand UO_361 (O_361,N_7633,N_9000);
nor UO_362 (O_362,N_9331,N_7931);
and UO_363 (O_363,N_9989,N_8692);
nor UO_364 (O_364,N_9400,N_9274);
and UO_365 (O_365,N_8364,N_7900);
or UO_366 (O_366,N_8464,N_9692);
nand UO_367 (O_367,N_9683,N_9590);
or UO_368 (O_368,N_8072,N_7628);
nor UO_369 (O_369,N_9732,N_9480);
or UO_370 (O_370,N_8250,N_7863);
or UO_371 (O_371,N_9812,N_9117);
nand UO_372 (O_372,N_7692,N_9127);
nand UO_373 (O_373,N_8425,N_8122);
nor UO_374 (O_374,N_9408,N_8178);
nor UO_375 (O_375,N_8846,N_8092);
nand UO_376 (O_376,N_7706,N_7924);
nand UO_377 (O_377,N_9508,N_8745);
or UO_378 (O_378,N_9060,N_8373);
nand UO_379 (O_379,N_8400,N_8751);
nand UO_380 (O_380,N_7525,N_7566);
or UO_381 (O_381,N_8334,N_9846);
or UO_382 (O_382,N_7825,N_7978);
or UO_383 (O_383,N_7890,N_9892);
or UO_384 (O_384,N_8290,N_9960);
xor UO_385 (O_385,N_8537,N_8012);
or UO_386 (O_386,N_8901,N_7973);
and UO_387 (O_387,N_7907,N_9470);
and UO_388 (O_388,N_9208,N_7556);
and UO_389 (O_389,N_8979,N_8402);
and UO_390 (O_390,N_8698,N_8471);
nor UO_391 (O_391,N_7806,N_9564);
nand UO_392 (O_392,N_9165,N_9032);
or UO_393 (O_393,N_8490,N_9394);
and UO_394 (O_394,N_8831,N_8054);
and UO_395 (O_395,N_9664,N_7958);
nand UO_396 (O_396,N_7779,N_9753);
and UO_397 (O_397,N_8310,N_9608);
and UO_398 (O_398,N_9944,N_8264);
nand UO_399 (O_399,N_8484,N_8858);
xor UO_400 (O_400,N_9109,N_9695);
or UO_401 (O_401,N_8403,N_8014);
xnor UO_402 (O_402,N_9742,N_9347);
nand UO_403 (O_403,N_8325,N_7879);
nand UO_404 (O_404,N_9130,N_9099);
or UO_405 (O_405,N_9579,N_9644);
xor UO_406 (O_406,N_9746,N_9830);
or UO_407 (O_407,N_9082,N_8024);
xnor UO_408 (O_408,N_9928,N_9301);
or UO_409 (O_409,N_9118,N_9013);
nand UO_410 (O_410,N_9335,N_8881);
nand UO_411 (O_411,N_9669,N_7700);
xnor UO_412 (O_412,N_9071,N_9257);
xnor UO_413 (O_413,N_8281,N_7835);
nand UO_414 (O_414,N_9377,N_9877);
nor UO_415 (O_415,N_8702,N_8186);
xor UO_416 (O_416,N_7575,N_7564);
or UO_417 (O_417,N_8499,N_8046);
xnor UO_418 (O_418,N_9571,N_8988);
or UO_419 (O_419,N_9760,N_9833);
nand UO_420 (O_420,N_9219,N_9171);
and UO_421 (O_421,N_7672,N_8793);
and UO_422 (O_422,N_9747,N_9583);
nor UO_423 (O_423,N_9440,N_9556);
or UO_424 (O_424,N_9072,N_8527);
or UO_425 (O_425,N_7848,N_8151);
xnor UO_426 (O_426,N_8279,N_8367);
and UO_427 (O_427,N_8867,N_9804);
xor UO_428 (O_428,N_9483,N_8454);
and UO_429 (O_429,N_9474,N_9927);
or UO_430 (O_430,N_9031,N_7645);
or UO_431 (O_431,N_7878,N_7507);
nor UO_432 (O_432,N_9421,N_8205);
nand UO_433 (O_433,N_9048,N_9302);
nand UO_434 (O_434,N_9631,N_9999);
nor UO_435 (O_435,N_8532,N_9136);
nand UO_436 (O_436,N_7610,N_8612);
nand UO_437 (O_437,N_7760,N_9476);
nand UO_438 (O_438,N_9738,N_7651);
nand UO_439 (O_439,N_9477,N_8573);
xnor UO_440 (O_440,N_9213,N_8162);
xnor UO_441 (O_441,N_9764,N_8536);
nor UO_442 (O_442,N_9887,N_7813);
xnor UO_443 (O_443,N_8750,N_8713);
nand UO_444 (O_444,N_7955,N_8234);
nor UO_445 (O_445,N_9696,N_7764);
or UO_446 (O_446,N_7949,N_7730);
or UO_447 (O_447,N_8847,N_8347);
nor UO_448 (O_448,N_9613,N_8690);
and UO_449 (O_449,N_9591,N_8785);
nor UO_450 (O_450,N_9195,N_8603);
or UO_451 (O_451,N_8233,N_9744);
and UO_452 (O_452,N_7543,N_9676);
and UO_453 (O_453,N_8243,N_7736);
nor UO_454 (O_454,N_9445,N_9372);
and UO_455 (O_455,N_8629,N_8428);
nor UO_456 (O_456,N_9242,N_8292);
nand UO_457 (O_457,N_8699,N_7942);
and UO_458 (O_458,N_8138,N_8523);
nand UO_459 (O_459,N_8105,N_7917);
and UO_460 (O_460,N_9530,N_8020);
nor UO_461 (O_461,N_9678,N_9674);
xnor UO_462 (O_462,N_9297,N_8430);
and UO_463 (O_463,N_8371,N_9708);
or UO_464 (O_464,N_9874,N_8672);
and UO_465 (O_465,N_9288,N_9668);
or UO_466 (O_466,N_9149,N_9859);
nor UO_467 (O_467,N_9965,N_8863);
nand UO_468 (O_468,N_7638,N_9479);
and UO_469 (O_469,N_8882,N_8415);
nand UO_470 (O_470,N_8805,N_8010);
nor UO_471 (O_471,N_7552,N_8321);
or UO_472 (O_472,N_9765,N_9342);
and UO_473 (O_473,N_8356,N_9921);
nor UO_474 (O_474,N_9401,N_8395);
xnor UO_475 (O_475,N_8280,N_9502);
nor UO_476 (O_476,N_9693,N_8695);
nand UO_477 (O_477,N_8467,N_8980);
or UO_478 (O_478,N_8604,N_8198);
xnor UO_479 (O_479,N_9575,N_7712);
nor UO_480 (O_480,N_8892,N_8920);
and UO_481 (O_481,N_8501,N_8029);
and UO_482 (O_482,N_9972,N_9599);
xnor UO_483 (O_483,N_9951,N_9906);
xor UO_484 (O_484,N_8316,N_7727);
and UO_485 (O_485,N_7614,N_8957);
or UO_486 (O_486,N_7719,N_9499);
nand UO_487 (O_487,N_7888,N_8740);
xor UO_488 (O_488,N_9309,N_8450);
xnor UO_489 (O_489,N_9380,N_7828);
nand UO_490 (O_490,N_7948,N_8775);
xor UO_491 (O_491,N_8978,N_9869);
or UO_492 (O_492,N_9443,N_7874);
and UO_493 (O_493,N_8884,N_9441);
and UO_494 (O_494,N_7935,N_9300);
or UO_495 (O_495,N_9576,N_7667);
or UO_496 (O_496,N_8773,N_8607);
or UO_497 (O_497,N_8602,N_8038);
nor UO_498 (O_498,N_8311,N_9879);
and UO_499 (O_499,N_8363,N_7800);
nand UO_500 (O_500,N_9551,N_9356);
or UO_501 (O_501,N_8944,N_8658);
nand UO_502 (O_502,N_9459,N_9992);
xor UO_503 (O_503,N_8592,N_7607);
and UO_504 (O_504,N_9740,N_8525);
nor UO_505 (O_505,N_7627,N_9969);
nor UO_506 (O_506,N_7679,N_9317);
nand UO_507 (O_507,N_9831,N_7988);
nand UO_508 (O_508,N_7860,N_8401);
and UO_509 (O_509,N_7784,N_8593);
or UO_510 (O_510,N_9592,N_9950);
xnor UO_511 (O_511,N_8350,N_7703);
and UO_512 (O_512,N_7707,N_9203);
or UO_513 (O_513,N_7913,N_9135);
and UO_514 (O_514,N_9232,N_8724);
and UO_515 (O_515,N_9056,N_7721);
or UO_516 (O_516,N_8317,N_8073);
nand UO_517 (O_517,N_8479,N_9935);
nand UO_518 (O_518,N_7550,N_9937);
nand UO_519 (O_519,N_8295,N_8835);
nor UO_520 (O_520,N_9751,N_9998);
xnor UO_521 (O_521,N_8856,N_9816);
nand UO_522 (O_522,N_8950,N_9630);
or UO_523 (O_523,N_9276,N_8959);
and UO_524 (O_524,N_7896,N_8362);
xnor UO_525 (O_525,N_9749,N_9603);
xor UO_526 (O_526,N_8883,N_7613);
or UO_527 (O_527,N_8448,N_8859);
nand UO_528 (O_528,N_7723,N_9376);
or UO_529 (O_529,N_8943,N_8617);
nor UO_530 (O_530,N_8218,N_9494);
xor UO_531 (O_531,N_8891,N_7976);
nor UO_532 (O_532,N_8583,N_9076);
xor UO_533 (O_533,N_8742,N_9138);
and UO_534 (O_534,N_9657,N_9512);
xor UO_535 (O_535,N_7952,N_9990);
and UO_536 (O_536,N_8534,N_9254);
nor UO_537 (O_537,N_9418,N_9750);
xor UO_538 (O_538,N_7611,N_8447);
nor UO_539 (O_539,N_9090,N_7755);
and UO_540 (O_540,N_7634,N_7666);
and UO_541 (O_541,N_8528,N_8641);
nand UO_542 (O_542,N_8177,N_8392);
nand UO_543 (O_543,N_8055,N_8888);
nor UO_544 (O_544,N_9587,N_7982);
nand UO_545 (O_545,N_9338,N_9449);
or UO_546 (O_546,N_9104,N_8949);
nor UO_547 (O_547,N_7996,N_8307);
or UO_548 (O_548,N_9577,N_9007);
and UO_549 (O_549,N_9328,N_9702);
nor UO_550 (O_550,N_8202,N_9660);
nor UO_551 (O_551,N_9325,N_9279);
xor UO_552 (O_552,N_8268,N_9478);
xor UO_553 (O_553,N_8931,N_8783);
or UO_554 (O_554,N_9403,N_8004);
and UO_555 (O_555,N_8781,N_8445);
nand UO_556 (O_556,N_8094,N_8027);
nor UO_557 (O_557,N_9534,N_9210);
or UO_558 (O_558,N_9940,N_8278);
nor UO_559 (O_559,N_7938,N_8908);
nor UO_560 (O_560,N_9081,N_7618);
and UO_561 (O_561,N_8461,N_7731);
nand UO_562 (O_562,N_9889,N_7520);
xor UO_563 (O_563,N_8683,N_8396);
xnor UO_564 (O_564,N_8382,N_8131);
nor UO_565 (O_565,N_8922,N_8494);
xor UO_566 (O_566,N_8507,N_7702);
and UO_567 (O_567,N_9143,N_7630);
nor UO_568 (O_568,N_7621,N_8200);
or UO_569 (O_569,N_8668,N_8272);
xor UO_570 (O_570,N_9035,N_7669);
or UO_571 (O_571,N_7562,N_7752);
nand UO_572 (O_572,N_8709,N_8246);
nor UO_573 (O_573,N_8711,N_7619);
xor UO_574 (O_574,N_8535,N_9262);
nand UO_575 (O_575,N_8865,N_8379);
nand UO_576 (O_576,N_8811,N_8130);
and UO_577 (O_577,N_9273,N_9994);
or UO_578 (O_578,N_8985,N_9020);
or UO_579 (O_579,N_7815,N_7867);
and UO_580 (O_580,N_7967,N_7536);
nor UO_581 (O_581,N_9724,N_9981);
or UO_582 (O_582,N_8013,N_8663);
nor UO_583 (O_583,N_9286,N_9902);
nand UO_584 (O_584,N_8852,N_9532);
nor UO_585 (O_585,N_8727,N_7729);
xnor UO_586 (O_586,N_8207,N_9460);
and UO_587 (O_587,N_7546,N_9178);
and UO_588 (O_588,N_9759,N_9642);
and UO_589 (O_589,N_9792,N_9748);
xnor UO_590 (O_590,N_8121,N_8145);
and UO_591 (O_591,N_7773,N_7861);
nor UO_592 (O_592,N_9088,N_7537);
and UO_593 (O_593,N_9306,N_8728);
nor UO_594 (O_594,N_9685,N_9976);
and UO_595 (O_595,N_8466,N_9453);
and UO_596 (O_596,N_9016,N_7650);
nand UO_597 (O_597,N_7699,N_7776);
or UO_598 (O_598,N_9159,N_8080);
and UO_599 (O_599,N_7685,N_8496);
xnor UO_600 (O_600,N_9185,N_9238);
and UO_601 (O_601,N_7936,N_8816);
xor UO_602 (O_602,N_8588,N_8191);
nand UO_603 (O_603,N_9779,N_8161);
nand UO_604 (O_604,N_8147,N_9151);
nor UO_605 (O_605,N_9607,N_7987);
or UO_606 (O_606,N_9217,N_8614);
nor UO_607 (O_607,N_9495,N_9384);
and UO_608 (O_608,N_7576,N_7622);
xnor UO_609 (O_609,N_9701,N_8378);
or UO_610 (O_610,N_9098,N_9466);
xor UO_611 (O_611,N_7646,N_7688);
or UO_612 (O_612,N_9223,N_9924);
and UO_613 (O_613,N_9250,N_8576);
or UO_614 (O_614,N_9096,N_8911);
and UO_615 (O_615,N_9522,N_8253);
or UO_616 (O_616,N_7979,N_9733);
nand UO_617 (O_617,N_8606,N_8685);
nand UO_618 (O_618,N_9959,N_8427);
or UO_619 (O_619,N_7801,N_8628);
or UO_620 (O_620,N_9755,N_7649);
xor UO_621 (O_621,N_7937,N_8443);
or UO_622 (O_622,N_8067,N_9796);
or UO_623 (O_623,N_9212,N_8755);
nor UO_624 (O_624,N_9819,N_8232);
and UO_625 (O_625,N_8767,N_8023);
nand UO_626 (O_626,N_7640,N_9179);
or UO_627 (O_627,N_7947,N_9901);
or UO_628 (O_628,N_7742,N_8267);
and UO_629 (O_629,N_8328,N_9856);
or UO_630 (O_630,N_9568,N_7678);
xnor UO_631 (O_631,N_9237,N_9092);
nor UO_632 (O_632,N_8697,N_8229);
nand UO_633 (O_633,N_8116,N_8896);
nor UO_634 (O_634,N_8622,N_9923);
nand UO_635 (O_635,N_9355,N_8354);
and UO_636 (O_636,N_9444,N_9574);
and UO_637 (O_637,N_7637,N_9553);
or UO_638 (O_638,N_8633,N_9946);
xor UO_639 (O_639,N_7824,N_9006);
nor UO_640 (O_640,N_8764,N_8737);
nand UO_641 (O_641,N_9730,N_9645);
and UO_642 (O_642,N_9589,N_9757);
nand UO_643 (O_643,N_9176,N_8081);
nor UO_644 (O_644,N_8681,N_8179);
nor UO_645 (O_645,N_8917,N_7509);
and UO_646 (O_646,N_7814,N_8187);
nor UO_647 (O_647,N_7577,N_8601);
and UO_648 (O_648,N_8098,N_9844);
nor UO_649 (O_649,N_7724,N_9852);
and UO_650 (O_650,N_9871,N_9319);
and UO_651 (O_651,N_9926,N_9942);
xor UO_652 (O_652,N_7901,N_7797);
and UO_653 (O_653,N_8182,N_8779);
nor UO_654 (O_654,N_8769,N_8455);
nand UO_655 (O_655,N_8504,N_7506);
xor UO_656 (O_656,N_9908,N_8696);
xor UO_657 (O_657,N_8678,N_8842);
and UO_658 (O_658,N_8765,N_8817);
xor UO_659 (O_659,N_8542,N_9113);
and UO_660 (O_660,N_8011,N_7993);
nor UO_661 (O_661,N_9269,N_7541);
and UO_662 (O_662,N_8868,N_9834);
or UO_663 (O_663,N_7554,N_8530);
or UO_664 (O_664,N_8547,N_7573);
xnor UO_665 (O_665,N_8540,N_9188);
or UO_666 (O_666,N_7735,N_8197);
or UO_667 (O_667,N_9658,N_9818);
nand UO_668 (O_668,N_9617,N_8752);
or UO_669 (O_669,N_9463,N_8045);
and UO_670 (O_670,N_8700,N_9966);
or UO_671 (O_671,N_9128,N_8458);
nand UO_672 (O_672,N_8473,N_9554);
xor UO_673 (O_673,N_8887,N_9447);
and UO_674 (O_674,N_8483,N_8777);
xor UO_675 (O_675,N_8170,N_9430);
xnor UO_676 (O_676,N_9670,N_9017);
or UO_677 (O_677,N_9938,N_7608);
or UO_678 (O_678,N_7594,N_9925);
nor UO_679 (O_679,N_8733,N_9941);
and UO_680 (O_680,N_7593,N_7654);
nor UO_681 (O_681,N_9357,N_8061);
or UO_682 (O_682,N_8906,N_7853);
nor UO_683 (O_683,N_8097,N_9037);
and UO_684 (O_684,N_9438,N_9030);
nor UO_685 (O_685,N_9653,N_8102);
nand UO_686 (O_686,N_7992,N_7785);
nand UO_687 (O_687,N_9315,N_9431);
and UO_688 (O_688,N_9370,N_9550);
xnor UO_689 (O_689,N_8676,N_8956);
nor UO_690 (O_690,N_8638,N_8518);
nor UO_691 (O_691,N_8136,N_8771);
or UO_692 (O_692,N_9729,N_8758);
and UO_693 (O_693,N_8000,N_8843);
or UO_694 (O_694,N_7858,N_8167);
xor UO_695 (O_695,N_9560,N_9628);
nand UO_696 (O_696,N_8551,N_9727);
nand UO_697 (O_697,N_8341,N_9743);
or UO_698 (O_698,N_9800,N_9461);
xnor UO_699 (O_699,N_9105,N_8512);
and UO_700 (O_700,N_7909,N_7929);
nand UO_701 (O_701,N_9106,N_8621);
nor UO_702 (O_702,N_8877,N_7899);
xnor UO_703 (O_703,N_9079,N_9087);
and UO_704 (O_704,N_9667,N_8472);
nand UO_705 (O_705,N_8918,N_8383);
or UO_706 (O_706,N_8289,N_8989);
xnor UO_707 (O_707,N_8034,N_8930);
or UO_708 (O_708,N_9622,N_8335);
nor UO_709 (O_709,N_9484,N_9161);
or UO_710 (O_710,N_8245,N_8421);
nor UO_711 (O_711,N_9003,N_9391);
or UO_712 (O_712,N_8485,N_7821);
and UO_713 (O_713,N_8679,N_7551);
or UO_714 (O_714,N_7695,N_7623);
or UO_715 (O_715,N_9754,N_8582);
xnor UO_716 (O_716,N_7660,N_8508);
nand UO_717 (O_717,N_8966,N_8637);
xnor UO_718 (O_718,N_8071,N_9621);
or UO_719 (O_719,N_9620,N_9260);
xnor UO_720 (O_720,N_9611,N_9058);
and UO_721 (O_721,N_9177,N_8168);
or UO_722 (O_722,N_9638,N_9197);
nand UO_723 (O_723,N_9807,N_9791);
or UO_724 (O_724,N_8283,N_8780);
nand UO_725 (O_725,N_9413,N_9619);
or UO_726 (O_726,N_8225,N_9067);
nand UO_727 (O_727,N_9776,N_7673);
nor UO_728 (O_728,N_9798,N_7754);
nor UO_729 (O_729,N_8456,N_9094);
nor UO_730 (O_730,N_7661,N_7906);
and UO_731 (O_731,N_9402,N_8615);
or UO_732 (O_732,N_8426,N_8664);
nand UO_733 (O_733,N_8100,N_8776);
nor UO_734 (O_734,N_9606,N_7966);
and UO_735 (O_735,N_9687,N_9198);
or UO_736 (O_736,N_9050,N_9580);
xnor UO_737 (O_737,N_7772,N_7894);
xor UO_738 (O_738,N_9595,N_9713);
nor UO_739 (O_739,N_8324,N_7898);
nand UO_740 (O_740,N_8749,N_9332);
or UO_741 (O_741,N_8397,N_9493);
and UO_742 (O_742,N_8487,N_7656);
nand UO_743 (O_743,N_9955,N_9022);
nor UO_744 (O_744,N_8399,N_7763);
nand UO_745 (O_745,N_9381,N_9943);
nand UO_746 (O_746,N_9330,N_8539);
nor UO_747 (O_747,N_7956,N_8224);
and UO_748 (O_748,N_9930,N_8510);
nor UO_749 (O_749,N_8375,N_7555);
xnor UO_750 (O_750,N_9970,N_7795);
xor UO_751 (O_751,N_8822,N_7717);
or UO_752 (O_752,N_7504,N_8720);
and UO_753 (O_753,N_8688,N_8154);
nand UO_754 (O_754,N_9368,N_9221);
nand UO_755 (O_755,N_9395,N_8871);
xnor UO_756 (O_756,N_7696,N_8667);
xnor UO_757 (O_757,N_9827,N_8302);
or UO_758 (O_758,N_9905,N_8511);
nor UO_759 (O_759,N_9077,N_9064);
xnor UO_760 (O_760,N_8042,N_9310);
or UO_761 (O_761,N_7664,N_7689);
xor UO_762 (O_762,N_8394,N_7641);
nor UO_763 (O_763,N_7842,N_8416);
nor UO_764 (O_764,N_9647,N_8876);
or UO_765 (O_765,N_8704,N_9963);
xnor UO_766 (O_766,N_7642,N_7518);
xor UO_767 (O_767,N_8812,N_8666);
and UO_768 (O_768,N_7934,N_9305);
xor UO_769 (O_769,N_9468,N_7777);
nand UO_770 (O_770,N_8398,N_9024);
nand UO_771 (O_771,N_9639,N_9828);
nor UO_772 (O_772,N_7620,N_8609);
or UO_773 (O_773,N_8110,N_8600);
xnor UO_774 (O_774,N_8137,N_8488);
or UO_775 (O_775,N_8661,N_7832);
nor UO_776 (O_776,N_9385,N_9913);
or UO_777 (O_777,N_7886,N_9561);
or UO_778 (O_778,N_8271,N_9734);
nor UO_779 (O_779,N_8844,N_9643);
xor UO_780 (O_780,N_7816,N_8806);
nor UO_781 (O_781,N_7590,N_9492);
nor UO_782 (O_782,N_9462,N_8575);
nor UO_783 (O_783,N_8976,N_8129);
nand UO_784 (O_784,N_9775,N_9235);
and UO_785 (O_785,N_8824,N_8184);
nand UO_786 (O_786,N_7849,N_8560);
nor UO_787 (O_787,N_8760,N_8090);
and UO_788 (O_788,N_7877,N_8564);
and UO_789 (O_789,N_8331,N_9303);
and UO_790 (O_790,N_9573,N_8358);
nor UO_791 (O_791,N_9770,N_7968);
and UO_792 (O_792,N_9153,N_9253);
and UO_793 (O_793,N_9002,N_8074);
or UO_794 (O_794,N_9410,N_9190);
and UO_795 (O_795,N_8468,N_9565);
or UO_796 (O_796,N_7770,N_8193);
xor UO_797 (O_797,N_8377,N_8967);
nor UO_798 (O_798,N_8993,N_9974);
xnor UO_799 (O_799,N_8032,N_9464);
and UO_800 (O_800,N_9710,N_9252);
nor UO_801 (O_801,N_8717,N_8030);
xnor UO_802 (O_802,N_8669,N_8826);
nand UO_803 (O_803,N_7781,N_7574);
nand UO_804 (O_804,N_8124,N_7757);
xnor UO_805 (O_805,N_8216,N_7687);
nor UO_806 (O_806,N_9870,N_8557);
nand UO_807 (O_807,N_8057,N_9581);
nor UO_808 (O_808,N_8910,N_9014);
and UO_809 (O_809,N_7749,N_8127);
or UO_810 (O_810,N_9514,N_8203);
or UO_811 (O_811,N_9011,N_8489);
and UO_812 (O_812,N_8735,N_9601);
nand UO_813 (O_813,N_9847,N_7946);
nor UO_814 (O_814,N_9065,N_9527);
xor UO_815 (O_815,N_9726,N_9095);
nand UO_816 (O_816,N_9458,N_9326);
nand UO_817 (O_817,N_7995,N_7547);
nor UO_818 (O_818,N_9043,N_8732);
nand UO_819 (O_819,N_7605,N_9163);
or UO_820 (O_820,N_8655,N_8143);
xnor UO_821 (O_821,N_9123,N_7972);
nor UO_822 (O_822,N_9761,N_7596);
and UO_823 (O_823,N_9346,N_9369);
xor UO_824 (O_824,N_8149,N_8368);
or UO_825 (O_825,N_9982,N_7804);
or UO_826 (O_826,N_7903,N_7963);
nor UO_827 (O_827,N_8260,N_9189);
and UO_828 (O_828,N_9101,N_8624);
xnor UO_829 (O_829,N_7530,N_8172);
nand UO_830 (O_830,N_8288,N_8938);
and UO_831 (O_831,N_8026,N_7748);
or UO_832 (O_832,N_8784,N_8684);
and UO_833 (O_833,N_8257,N_9420);
and UO_834 (O_834,N_8972,N_9986);
or UO_835 (O_835,N_8359,N_9063);
and UO_836 (O_836,N_7737,N_7808);
nor UO_837 (O_837,N_7572,N_8277);
nor UO_838 (O_838,N_9842,N_7919);
nand UO_839 (O_839,N_7694,N_9307);
or UO_840 (O_840,N_9398,N_9181);
nand UO_841 (O_841,N_9199,N_9120);
nor UO_842 (O_842,N_7980,N_9763);
and UO_843 (O_843,N_9027,N_9091);
or UO_844 (O_844,N_8645,N_7606);
and UO_845 (O_845,N_9585,N_8091);
or UO_846 (O_846,N_7629,N_9813);
nand UO_847 (O_847,N_8693,N_9139);
nand UO_848 (O_848,N_8469,N_7584);
and UO_849 (O_849,N_9144,N_8820);
nand UO_850 (O_850,N_9967,N_7739);
or UO_851 (O_851,N_9456,N_8814);
nand UO_852 (O_852,N_9089,N_8715);
nand UO_853 (O_853,N_9157,N_9393);
and UO_854 (O_854,N_9487,N_9419);
xnor UO_855 (O_855,N_8927,N_8315);
or UO_856 (O_856,N_9004,N_7914);
or UO_857 (O_857,N_8936,N_9851);
or UO_858 (O_858,N_7984,N_8803);
xor UO_859 (O_859,N_9340,N_7883);
or UO_860 (O_860,N_8860,N_9993);
or UO_861 (O_861,N_8848,N_8293);
nor UO_862 (O_862,N_7582,N_7569);
nor UO_863 (O_863,N_9231,N_9781);
nand UO_864 (O_864,N_9823,N_9507);
and UO_865 (O_865,N_8893,N_8348);
nor UO_866 (O_866,N_8851,N_7514);
or UO_867 (O_867,N_7951,N_7905);
and UO_868 (O_868,N_9854,N_9107);
and UO_869 (O_869,N_8671,N_8873);
xor UO_870 (O_870,N_7807,N_8905);
nor UO_871 (O_871,N_9980,N_7882);
nand UO_872 (O_872,N_9467,N_8799);
or UO_873 (O_873,N_8571,N_9979);
nand UO_874 (O_874,N_9263,N_8515);
and UO_875 (O_875,N_9145,N_9649);
and UO_876 (O_876,N_8333,N_9434);
xor UO_877 (O_877,N_7617,N_8503);
or UO_878 (O_878,N_8330,N_8648);
and UO_879 (O_879,N_8770,N_8296);
or UO_880 (O_880,N_7921,N_9971);
xor UO_881 (O_881,N_8716,N_9038);
and UO_882 (O_882,N_8037,N_8183);
nand UO_883 (O_883,N_9114,N_8682);
xor UO_884 (O_884,N_8558,N_9224);
nor UO_885 (O_885,N_8754,N_8762);
or UO_886 (O_886,N_9741,N_9044);
and UO_887 (O_887,N_8994,N_9299);
nor UO_888 (O_888,N_9255,N_8992);
nand UO_889 (O_889,N_7578,N_9313);
nor UO_890 (O_890,N_9333,N_8015);
nor UO_891 (O_891,N_9899,N_7865);
and UO_892 (O_892,N_9865,N_9141);
nand UO_893 (O_893,N_8807,N_8339);
or UO_894 (O_894,N_9023,N_7585);
nor UO_895 (O_895,N_8545,N_9820);
nor UO_896 (O_896,N_7597,N_9766);
nand UO_897 (O_897,N_9520,N_8164);
nor UO_898 (O_898,N_9271,N_8482);
xnor UO_899 (O_899,N_8156,N_8730);
xnor UO_900 (O_900,N_9162,N_8457);
and UO_901 (O_901,N_8939,N_8897);
or UO_902 (O_902,N_8237,N_9001);
or UO_903 (O_903,N_8297,N_7838);
nor UO_904 (O_904,N_8650,N_9240);
nand UO_905 (O_905,N_9435,N_8050);
or UO_906 (O_906,N_9390,N_7756);
nand UO_907 (O_907,N_9546,N_8665);
and UO_908 (O_908,N_8969,N_7840);
and UO_909 (O_909,N_7524,N_8114);
xor UO_910 (O_910,N_8112,N_8239);
and UO_911 (O_911,N_8963,N_8841);
nor UO_912 (O_912,N_9782,N_8159);
xor UO_913 (O_913,N_9261,N_7829);
and UO_914 (O_914,N_9954,N_7775);
nor UO_915 (O_915,N_8712,N_7957);
and UO_916 (O_916,N_9234,N_8937);
nand UO_917 (O_917,N_8082,N_8028);
and UO_918 (O_918,N_8135,N_7532);
and UO_919 (O_919,N_8895,N_7653);
nand UO_920 (O_920,N_9364,N_8238);
xor UO_921 (O_921,N_8231,N_9910);
or UO_922 (O_922,N_7647,N_8825);
xor UO_923 (O_923,N_8476,N_8562);
nor UO_924 (O_924,N_8520,N_8446);
and UO_925 (O_925,N_8390,N_9797);
nand UO_926 (O_926,N_7709,N_9722);
or UO_927 (O_927,N_9170,N_9884);
and UO_928 (O_928,N_9396,N_9498);
nand UO_929 (O_929,N_9166,N_9428);
nand UO_930 (O_930,N_8894,N_7873);
xnor UO_931 (O_931,N_7716,N_8437);
nand UO_932 (O_932,N_7836,N_9218);
and UO_933 (O_933,N_9451,N_8652);
and UO_934 (O_934,N_9373,N_9057);
xnor UO_935 (O_935,N_9180,N_8774);
or UO_936 (O_936,N_8739,N_8726);
nand UO_937 (O_937,N_7964,N_9671);
or UO_938 (O_938,N_9184,N_9737);
nand UO_939 (O_939,N_9939,N_7548);
xor UO_940 (O_940,N_8904,N_9836);
xnor UO_941 (O_941,N_7726,N_8332);
nand UO_942 (O_942,N_9513,N_9916);
nand UO_943 (O_943,N_9872,N_8981);
nand UO_944 (O_944,N_9289,N_9352);
xnor UO_945 (O_945,N_7985,N_8282);
xnor UO_946 (O_946,N_8611,N_8270);
nor UO_947 (O_947,N_8498,N_9124);
and UO_948 (O_948,N_7734,N_9780);
nand UO_949 (O_949,N_9627,N_9864);
and UO_950 (O_950,N_9275,N_9806);
xnor UO_951 (O_951,N_8845,N_9365);
nor UO_952 (O_952,N_8598,N_8244);
xor UO_953 (O_953,N_8636,N_7846);
or UO_954 (O_954,N_8134,N_9200);
xnor UO_955 (O_955,N_7802,N_8230);
xnor UO_956 (O_956,N_7889,N_9363);
and UO_957 (O_957,N_8351,N_9062);
or UO_958 (O_958,N_7604,N_7588);
nand UO_959 (O_959,N_8941,N_7891);
xor UO_960 (O_960,N_9201,N_7710);
and UO_961 (O_961,N_9280,N_7529);
nand UO_962 (O_962,N_7615,N_9809);
and UO_963 (O_963,N_8005,N_9718);
nand UO_964 (O_964,N_9641,N_7704);
and UO_965 (O_965,N_8209,N_7820);
and UO_966 (O_966,N_8673,N_8478);
xor UO_967 (O_967,N_8357,N_9684);
xnor UO_968 (O_968,N_9010,N_8226);
or UO_969 (O_969,N_8710,N_8986);
xnor UO_970 (O_970,N_9482,N_9736);
and UO_971 (O_971,N_9958,N_9259);
and UO_972 (O_972,N_7558,N_8285);
nor UO_973 (O_973,N_8923,N_9281);
or UO_974 (O_974,N_8880,N_7686);
nand UO_975 (O_975,N_9618,N_8190);
xnor UO_976 (O_976,N_8340,N_8984);
nand UO_977 (O_977,N_8748,N_9268);
xnor UO_978 (O_978,N_9247,N_9903);
or UO_979 (O_979,N_8721,N_9110);
xor UO_980 (O_980,N_9706,N_8632);
or UO_981 (O_981,N_7527,N_8837);
nand UO_982 (O_982,N_7567,N_9720);
nand UO_983 (O_983,N_9379,N_9270);
nor UO_984 (O_984,N_9452,N_8391);
or UO_985 (O_985,N_9264,N_9158);
xor UO_986 (O_986,N_7843,N_8590);
nor UO_987 (O_987,N_8043,N_8631);
and UO_988 (O_988,N_8809,N_8474);
xor UO_989 (O_989,N_7868,N_9814);
or UO_990 (O_990,N_9785,N_8083);
nor UO_991 (O_991,N_9047,N_8909);
nor UO_992 (O_992,N_9680,N_7758);
or UO_993 (O_993,N_8258,N_9053);
xor UO_994 (O_994,N_8885,N_8380);
or UO_995 (O_995,N_8077,N_8259);
or UO_996 (O_996,N_7954,N_7766);
and UO_997 (O_997,N_8616,N_9034);
or UO_998 (O_998,N_9382,N_7876);
nor UO_999 (O_999,N_9405,N_9511);
nor UO_1000 (O_1000,N_9745,N_8913);
or UO_1001 (O_1001,N_8834,N_8166);
or UO_1002 (O_1002,N_7753,N_8960);
and UO_1003 (O_1003,N_8543,N_8210);
nand UO_1004 (O_1004,N_8123,N_9283);
xor UO_1005 (O_1005,N_8968,N_7508);
nand UO_1006 (O_1006,N_7744,N_8323);
nor UO_1007 (O_1007,N_7990,N_7981);
nand UO_1008 (O_1008,N_8572,N_7768);
xor UO_1009 (O_1009,N_7599,N_9122);
or UO_1010 (O_1010,N_7648,N_7932);
and UO_1011 (O_1011,N_8491,N_7850);
or UO_1012 (O_1012,N_9661,N_9919);
or UO_1013 (O_1013,N_9878,N_8808);
xor UO_1014 (O_1014,N_8529,N_8990);
nor UO_1015 (O_1015,N_7512,N_7761);
xnor UO_1016 (O_1016,N_9295,N_9353);
and UO_1017 (O_1017,N_9953,N_9997);
nand UO_1018 (O_1018,N_9169,N_7533);
nor UO_1019 (O_1019,N_8169,N_9354);
and UO_1020 (O_1020,N_9040,N_8818);
xor UO_1021 (O_1021,N_9922,N_8006);
nand UO_1022 (O_1022,N_8089,N_8855);
nor UO_1023 (O_1023,N_9975,N_9439);
and UO_1024 (O_1024,N_8251,N_8222);
xor UO_1025 (O_1025,N_9196,N_9634);
and UO_1026 (O_1026,N_7658,N_8248);
nand UO_1027 (O_1027,N_9567,N_9334);
nor UO_1028 (O_1028,N_9673,N_7745);
and UO_1029 (O_1029,N_8025,N_9304);
and UO_1030 (O_1030,N_9860,N_9132);
nor UO_1031 (O_1031,N_9784,N_8554);
and UO_1032 (O_1032,N_8836,N_8126);
xnor UO_1033 (O_1033,N_8199,N_9131);
and UO_1034 (O_1034,N_9028,N_9882);
or UO_1035 (O_1035,N_8227,N_8442);
nand UO_1036 (O_1036,N_7945,N_7908);
nor UO_1037 (O_1037,N_9415,N_7741);
xor UO_1038 (O_1038,N_8036,N_8212);
nand UO_1039 (O_1039,N_9826,N_9411);
nand UO_1040 (O_1040,N_8559,N_8214);
nand UO_1041 (O_1041,N_9857,N_9593);
xor UO_1042 (O_1042,N_9243,N_8120);
or UO_1043 (O_1043,N_8273,N_9843);
xor UO_1044 (O_1044,N_8327,N_9582);
nor UO_1045 (O_1045,N_7644,N_7526);
or UO_1046 (O_1046,N_8701,N_9362);
nor UO_1047 (O_1047,N_9399,N_9973);
or UO_1048 (O_1048,N_9051,N_9535);
or UO_1049 (O_1049,N_9069,N_9417);
and UO_1050 (O_1050,N_8694,N_8299);
nand UO_1051 (O_1051,N_9682,N_9541);
xnor UO_1052 (O_1052,N_8502,N_8768);
nand UO_1053 (O_1053,N_8338,N_9805);
xor UO_1054 (O_1054,N_9615,N_8096);
nor UO_1055 (O_1055,N_8791,N_9810);
xnor UO_1056 (O_1056,N_9290,N_7793);
and UO_1057 (O_1057,N_8007,N_9211);
xnor UO_1058 (O_1058,N_9045,N_8087);
xor UO_1059 (O_1059,N_7823,N_9486);
or UO_1060 (O_1060,N_9542,N_9863);
nor UO_1061 (O_1061,N_7655,N_8412);
xor UO_1062 (O_1062,N_8093,N_8889);
or UO_1063 (O_1063,N_8521,N_9931);
nand UO_1064 (O_1064,N_9646,N_9964);
nand UO_1065 (O_1065,N_8919,N_9716);
and UO_1066 (O_1066,N_8656,N_8160);
nor UO_1067 (O_1067,N_8291,N_8533);
or UO_1068 (O_1068,N_7626,N_9552);
nand UO_1069 (O_1069,N_8462,N_7531);
nor UO_1070 (O_1070,N_9026,N_8022);
or UO_1071 (O_1071,N_9635,N_8366);
nor UO_1072 (O_1072,N_8069,N_7845);
nand UO_1073 (O_1073,N_8052,N_7940);
xnor UO_1074 (O_1074,N_7884,N_9962);
xnor UO_1075 (O_1075,N_7625,N_8434);
nor UO_1076 (O_1076,N_9214,N_9025);
nor UO_1077 (O_1077,N_9018,N_8413);
nand UO_1078 (O_1078,N_9074,N_8587);
or UO_1079 (O_1079,N_9424,N_9629);
or UO_1080 (O_1080,N_8801,N_9371);
nor UO_1081 (O_1081,N_7675,N_7902);
xnor UO_1082 (O_1082,N_8263,N_8734);
xor UO_1083 (O_1083,N_7818,N_8747);
nor UO_1084 (O_1084,N_7587,N_8987);
and UO_1085 (O_1085,N_7974,N_7965);
xnor UO_1086 (O_1086,N_9771,N_9845);
and UO_1087 (O_1087,N_8439,N_9433);
or UO_1088 (O_1088,N_8128,N_9790);
nand UO_1089 (O_1089,N_9469,N_9700);
or UO_1090 (O_1090,N_8782,N_8962);
nand UO_1091 (O_1091,N_8544,N_8646);
nand UO_1092 (O_1092,N_9832,N_8065);
nor UO_1093 (O_1093,N_7870,N_8795);
nand UO_1094 (O_1094,N_9566,N_7790);
nand UO_1095 (O_1095,N_9624,N_8176);
nor UO_1096 (O_1096,N_9528,N_9155);
nand UO_1097 (O_1097,N_9655,N_9042);
nor UO_1098 (O_1098,N_7668,N_8039);
nor UO_1099 (O_1099,N_9920,N_8741);
nor UO_1100 (O_1100,N_8059,N_8640);
and UO_1101 (O_1101,N_9389,N_7505);
xnor UO_1102 (O_1102,N_9308,N_9111);
nor UO_1103 (O_1103,N_8481,N_8586);
or UO_1104 (O_1104,N_7598,N_9387);
nand UO_1105 (O_1105,N_7933,N_9788);
or UO_1106 (O_1106,N_7910,N_9121);
nand UO_1107 (O_1107,N_9078,N_8188);
xor UO_1108 (O_1108,N_7844,N_9265);
and UO_1109 (O_1109,N_8654,N_9416);
xnor UO_1110 (O_1110,N_7875,N_9033);
nand UO_1111 (O_1111,N_8009,N_9156);
nor UO_1112 (O_1112,N_8578,N_8031);
nor UO_1113 (O_1113,N_9205,N_9073);
xor UO_1114 (O_1114,N_7971,N_8308);
or UO_1115 (O_1115,N_7732,N_9216);
xnor UO_1116 (O_1116,N_9932,N_8565);
nor UO_1117 (O_1117,N_9126,N_8361);
or UO_1118 (O_1118,N_9904,N_9772);
and UO_1119 (O_1119,N_9115,N_8526);
nand UO_1120 (O_1120,N_8099,N_9085);
and UO_1121 (O_1121,N_8393,N_9008);
nand UO_1122 (O_1122,N_9712,N_9046);
and UO_1123 (O_1123,N_9351,N_8651);
or UO_1124 (O_1124,N_8886,N_8849);
nor UO_1125 (O_1125,N_7705,N_8802);
nor UO_1126 (O_1126,N_9350,N_9752);
or UO_1127 (O_1127,N_9505,N_8680);
nand UO_1128 (O_1128,N_9756,N_9654);
nand UO_1129 (O_1129,N_8635,N_7515);
nor UO_1130 (O_1130,N_8954,N_8228);
and UO_1131 (O_1131,N_9526,N_7639);
and UO_1132 (O_1132,N_8044,N_7960);
nand UO_1133 (O_1133,N_9360,N_9838);
and UO_1134 (O_1134,N_8284,N_8002);
nor UO_1135 (O_1135,N_9407,N_9769);
nand UO_1136 (O_1136,N_7852,N_7943);
xor UO_1137 (O_1137,N_7714,N_8497);
xnor UO_1138 (O_1138,N_9632,N_8148);
xor UO_1139 (O_1139,N_8935,N_9174);
xnor UO_1140 (O_1140,N_9949,N_7534);
or UO_1141 (O_1141,N_7792,N_9623);
nor UO_1142 (O_1142,N_9849,N_8419);
nand UO_1143 (O_1143,N_8217,N_8872);
nor UO_1144 (O_1144,N_8687,N_8853);
nor UO_1145 (O_1145,N_9193,N_8514);
nor UO_1146 (O_1146,N_7837,N_9598);
or UO_1147 (O_1147,N_8945,N_9225);
xnor UO_1148 (O_1148,N_8953,N_9423);
and UO_1149 (O_1149,N_8432,N_9545);
xor UO_1150 (O_1150,N_9358,N_9084);
and UO_1151 (O_1151,N_9093,N_9515);
nor UO_1152 (O_1152,N_9652,N_9690);
or UO_1153 (O_1153,N_9366,N_9636);
or UO_1154 (O_1154,N_8759,N_9677);
nor UO_1155 (O_1155,N_9656,N_9978);
and UO_1156 (O_1156,N_7542,N_9378);
and UO_1157 (O_1157,N_8620,N_9609);
or UO_1158 (O_1158,N_8201,N_8075);
and UO_1159 (O_1159,N_9519,N_8971);
nand UO_1160 (O_1160,N_9984,N_8630);
xnor UO_1161 (O_1161,N_9320,N_9426);
nand UO_1162 (O_1162,N_9625,N_9251);
nand UO_1163 (O_1163,N_9442,N_9455);
nand UO_1164 (O_1164,N_9167,N_9873);
nor UO_1165 (O_1165,N_9422,N_7581);
and UO_1166 (O_1166,N_8453,N_7571);
nand UO_1167 (O_1167,N_7722,N_7540);
or UO_1168 (O_1168,N_9717,N_7713);
nand UO_1169 (O_1169,N_8021,N_9711);
xor UO_1170 (O_1170,N_8546,N_7662);
nor UO_1171 (O_1171,N_9918,N_9794);
nand UO_1172 (O_1172,N_7769,N_9061);
nor UO_1173 (O_1173,N_9052,N_8051);
and UO_1174 (O_1174,N_9448,N_9707);
xor UO_1175 (O_1175,N_7904,N_8322);
nand UO_1176 (O_1176,N_9616,N_7698);
and UO_1177 (O_1177,N_8294,N_8828);
xnor UO_1178 (O_1178,N_8706,N_8864);
nand UO_1179 (O_1179,N_8365,N_8517);
or UO_1180 (O_1180,N_8139,N_9207);
nor UO_1181 (O_1181,N_9570,N_7663);
nor UO_1182 (O_1182,N_7502,N_7880);
xor UO_1183 (O_1183,N_9559,N_9936);
nand UO_1184 (O_1184,N_9191,N_8516);
nand UO_1185 (O_1185,N_8996,N_9134);
and UO_1186 (O_1186,N_7579,N_9894);
nor UO_1187 (O_1187,N_9055,N_7600);
and UO_1188 (O_1188,N_9432,N_8756);
and UO_1189 (O_1189,N_8152,N_8670);
xor UO_1190 (O_1190,N_8541,N_9795);
nand UO_1191 (O_1191,N_9640,N_9245);
xnor UO_1192 (O_1192,N_9578,N_9721);
and UO_1193 (O_1193,N_9412,N_9866);
or UO_1194 (O_1194,N_8247,N_9543);
or UO_1195 (O_1195,N_9236,N_8387);
nand UO_1196 (O_1196,N_7557,N_9633);
and UO_1197 (O_1197,N_9108,N_8078);
nor UO_1198 (O_1198,N_8850,N_9547);
and UO_1199 (O_1199,N_9945,N_7680);
xnor UO_1200 (O_1200,N_8626,N_9933);
nor UO_1201 (O_1201,N_8744,N_8150);
xnor UO_1202 (O_1202,N_9506,N_9777);
or UO_1203 (O_1203,N_9572,N_8719);
and UO_1204 (O_1204,N_8932,N_7746);
nand UO_1205 (O_1205,N_8623,N_8921);
nand UO_1206 (O_1206,N_9182,N_9019);
xor UO_1207 (O_1207,N_7922,N_9475);
xor UO_1208 (O_1208,N_9278,N_8662);
and UO_1209 (O_1209,N_8256,N_8070);
or UO_1210 (O_1210,N_9337,N_8660);
xor UO_1211 (O_1211,N_8346,N_7805);
or UO_1212 (O_1212,N_8088,N_8001);
xnor UO_1213 (O_1213,N_7718,N_7923);
or UO_1214 (O_1214,N_9296,N_8252);
xor UO_1215 (O_1215,N_8306,N_9481);
nand UO_1216 (O_1216,N_8552,N_9991);
or UO_1217 (O_1217,N_8242,N_8585);
xnor UO_1218 (O_1218,N_8040,N_9789);
xnor UO_1219 (O_1219,N_9662,N_8579);
and UO_1220 (O_1220,N_8103,N_8940);
or UO_1221 (O_1221,N_9516,N_8625);
and UO_1222 (O_1222,N_9686,N_7812);
xor UO_1223 (O_1223,N_9454,N_7799);
nand UO_1224 (O_1224,N_8788,N_9558);
xor UO_1225 (O_1225,N_8173,N_8125);
nand UO_1226 (O_1226,N_7780,N_9626);
nand UO_1227 (O_1227,N_8958,N_8948);
nand UO_1228 (O_1228,N_8787,N_9361);
and UO_1229 (O_1229,N_8142,N_8827);
or UO_1230 (O_1230,N_8451,N_9344);
nand UO_1231 (O_1231,N_9005,N_7559);
and UO_1232 (O_1232,N_8659,N_7862);
nor UO_1233 (O_1233,N_7855,N_9323);
or UO_1234 (O_1234,N_8890,N_7586);
and UO_1235 (O_1235,N_7826,N_9497);
or UO_1236 (O_1236,N_7708,N_9316);
or UO_1237 (O_1237,N_8409,N_8287);
and UO_1238 (O_1238,N_8221,N_8261);
and UO_1239 (O_1239,N_9383,N_9277);
and UO_1240 (O_1240,N_8389,N_7912);
or UO_1241 (O_1241,N_9536,N_8063);
xor UO_1242 (O_1242,N_8435,N_8689);
or UO_1243 (O_1243,N_9604,N_9183);
nor UO_1244 (O_1244,N_8104,N_8778);
nor UO_1245 (O_1245,N_7788,N_9392);
nand UO_1246 (O_1246,N_8647,N_7535);
or UO_1247 (O_1247,N_8548,N_9192);
nand UO_1248 (O_1248,N_9612,N_8703);
xnor UO_1249 (O_1249,N_7961,N_8999);
nor UO_1250 (O_1250,N_9749,N_9048);
or UO_1251 (O_1251,N_9240,N_7993);
or UO_1252 (O_1252,N_9100,N_8858);
nand UO_1253 (O_1253,N_9185,N_8899);
nand UO_1254 (O_1254,N_8019,N_8373);
or UO_1255 (O_1255,N_8597,N_7588);
nor UO_1256 (O_1256,N_9082,N_9218);
or UO_1257 (O_1257,N_9280,N_9265);
nand UO_1258 (O_1258,N_7929,N_9779);
and UO_1259 (O_1259,N_9169,N_9991);
and UO_1260 (O_1260,N_8191,N_8882);
or UO_1261 (O_1261,N_9741,N_8008);
nand UO_1262 (O_1262,N_8344,N_8601);
and UO_1263 (O_1263,N_7925,N_7951);
or UO_1264 (O_1264,N_8956,N_7695);
xor UO_1265 (O_1265,N_9374,N_9833);
or UO_1266 (O_1266,N_8258,N_9858);
xor UO_1267 (O_1267,N_9506,N_8565);
xor UO_1268 (O_1268,N_8523,N_7603);
nor UO_1269 (O_1269,N_8359,N_9042);
or UO_1270 (O_1270,N_9464,N_8575);
or UO_1271 (O_1271,N_7784,N_9706);
nor UO_1272 (O_1272,N_7740,N_9274);
nand UO_1273 (O_1273,N_9502,N_9734);
nand UO_1274 (O_1274,N_8412,N_7649);
nand UO_1275 (O_1275,N_8348,N_9776);
and UO_1276 (O_1276,N_8032,N_9418);
nor UO_1277 (O_1277,N_9952,N_8658);
and UO_1278 (O_1278,N_9062,N_9799);
and UO_1279 (O_1279,N_8307,N_7745);
xnor UO_1280 (O_1280,N_9970,N_9472);
nor UO_1281 (O_1281,N_8066,N_9753);
and UO_1282 (O_1282,N_9400,N_8361);
nand UO_1283 (O_1283,N_9858,N_9524);
and UO_1284 (O_1284,N_8337,N_7524);
nor UO_1285 (O_1285,N_8646,N_9745);
and UO_1286 (O_1286,N_7730,N_9704);
nor UO_1287 (O_1287,N_9668,N_9277);
and UO_1288 (O_1288,N_9778,N_7868);
xor UO_1289 (O_1289,N_8262,N_7504);
or UO_1290 (O_1290,N_7557,N_8048);
or UO_1291 (O_1291,N_9626,N_7782);
xor UO_1292 (O_1292,N_8775,N_7562);
and UO_1293 (O_1293,N_8775,N_9573);
nor UO_1294 (O_1294,N_9276,N_9719);
nand UO_1295 (O_1295,N_9574,N_9241);
nand UO_1296 (O_1296,N_9881,N_8139);
or UO_1297 (O_1297,N_9104,N_8148);
nand UO_1298 (O_1298,N_7936,N_8518);
or UO_1299 (O_1299,N_7942,N_9244);
xnor UO_1300 (O_1300,N_8666,N_7887);
or UO_1301 (O_1301,N_9455,N_9352);
nand UO_1302 (O_1302,N_9030,N_9168);
xnor UO_1303 (O_1303,N_7857,N_9572);
nand UO_1304 (O_1304,N_9380,N_8800);
xor UO_1305 (O_1305,N_8579,N_9374);
xnor UO_1306 (O_1306,N_8749,N_9510);
nor UO_1307 (O_1307,N_7926,N_8518);
nor UO_1308 (O_1308,N_7654,N_9144);
nand UO_1309 (O_1309,N_7790,N_9647);
nor UO_1310 (O_1310,N_8283,N_9841);
and UO_1311 (O_1311,N_9291,N_8583);
xor UO_1312 (O_1312,N_8856,N_8256);
nand UO_1313 (O_1313,N_9812,N_9420);
xor UO_1314 (O_1314,N_9063,N_8782);
and UO_1315 (O_1315,N_9827,N_9355);
nor UO_1316 (O_1316,N_7993,N_8468);
xor UO_1317 (O_1317,N_8266,N_9656);
nor UO_1318 (O_1318,N_8668,N_7569);
or UO_1319 (O_1319,N_7871,N_8654);
or UO_1320 (O_1320,N_9894,N_9130);
nor UO_1321 (O_1321,N_8248,N_8695);
nand UO_1322 (O_1322,N_9130,N_7750);
xnor UO_1323 (O_1323,N_8735,N_9571);
nand UO_1324 (O_1324,N_9883,N_8375);
or UO_1325 (O_1325,N_8416,N_9986);
and UO_1326 (O_1326,N_8044,N_8535);
nor UO_1327 (O_1327,N_9970,N_7986);
nand UO_1328 (O_1328,N_9393,N_7833);
nor UO_1329 (O_1329,N_7974,N_9401);
nor UO_1330 (O_1330,N_8477,N_9549);
xnor UO_1331 (O_1331,N_8992,N_9282);
or UO_1332 (O_1332,N_9559,N_9509);
xnor UO_1333 (O_1333,N_7716,N_7648);
or UO_1334 (O_1334,N_9651,N_8639);
or UO_1335 (O_1335,N_8485,N_9428);
nor UO_1336 (O_1336,N_9073,N_8551);
nor UO_1337 (O_1337,N_8140,N_8109);
and UO_1338 (O_1338,N_8805,N_8107);
xnor UO_1339 (O_1339,N_8247,N_9696);
and UO_1340 (O_1340,N_9247,N_7650);
nand UO_1341 (O_1341,N_7526,N_7577);
nand UO_1342 (O_1342,N_8938,N_7981);
xor UO_1343 (O_1343,N_7547,N_8016);
or UO_1344 (O_1344,N_8281,N_7577);
xnor UO_1345 (O_1345,N_9912,N_7573);
or UO_1346 (O_1346,N_9992,N_9268);
or UO_1347 (O_1347,N_9982,N_9139);
nor UO_1348 (O_1348,N_8319,N_8824);
or UO_1349 (O_1349,N_9321,N_9793);
xor UO_1350 (O_1350,N_7574,N_8579);
xnor UO_1351 (O_1351,N_8560,N_8268);
and UO_1352 (O_1352,N_8816,N_8407);
and UO_1353 (O_1353,N_8545,N_9189);
nor UO_1354 (O_1354,N_8333,N_8445);
nor UO_1355 (O_1355,N_8911,N_7505);
and UO_1356 (O_1356,N_9045,N_9633);
and UO_1357 (O_1357,N_9336,N_8174);
xnor UO_1358 (O_1358,N_8392,N_9204);
nand UO_1359 (O_1359,N_9642,N_7881);
and UO_1360 (O_1360,N_8713,N_9497);
and UO_1361 (O_1361,N_8055,N_9938);
or UO_1362 (O_1362,N_8947,N_7870);
nor UO_1363 (O_1363,N_9267,N_9484);
nor UO_1364 (O_1364,N_9937,N_7537);
nand UO_1365 (O_1365,N_7632,N_8943);
or UO_1366 (O_1366,N_9258,N_9492);
or UO_1367 (O_1367,N_8906,N_8059);
nand UO_1368 (O_1368,N_8550,N_8973);
xor UO_1369 (O_1369,N_9809,N_9557);
nor UO_1370 (O_1370,N_8008,N_9336);
or UO_1371 (O_1371,N_7979,N_8709);
and UO_1372 (O_1372,N_9698,N_8366);
and UO_1373 (O_1373,N_8346,N_9220);
nor UO_1374 (O_1374,N_8818,N_8590);
and UO_1375 (O_1375,N_9496,N_8416);
xnor UO_1376 (O_1376,N_9812,N_8295);
xnor UO_1377 (O_1377,N_7617,N_8768);
xor UO_1378 (O_1378,N_8993,N_9957);
and UO_1379 (O_1379,N_8751,N_7978);
and UO_1380 (O_1380,N_9373,N_8414);
nand UO_1381 (O_1381,N_7785,N_8042);
nand UO_1382 (O_1382,N_8191,N_8666);
and UO_1383 (O_1383,N_8507,N_8477);
xor UO_1384 (O_1384,N_7501,N_9150);
nor UO_1385 (O_1385,N_8475,N_8249);
xor UO_1386 (O_1386,N_8563,N_8258);
nand UO_1387 (O_1387,N_8204,N_9588);
and UO_1388 (O_1388,N_9743,N_8159);
nand UO_1389 (O_1389,N_7735,N_9012);
and UO_1390 (O_1390,N_8495,N_8806);
nor UO_1391 (O_1391,N_8180,N_9852);
xnor UO_1392 (O_1392,N_7582,N_9651);
nor UO_1393 (O_1393,N_9148,N_7893);
nor UO_1394 (O_1394,N_9144,N_9740);
nand UO_1395 (O_1395,N_9307,N_8047);
or UO_1396 (O_1396,N_9787,N_9421);
or UO_1397 (O_1397,N_7889,N_9366);
nand UO_1398 (O_1398,N_9756,N_9665);
nand UO_1399 (O_1399,N_9130,N_7570);
nand UO_1400 (O_1400,N_9412,N_9970);
xnor UO_1401 (O_1401,N_8706,N_9888);
nand UO_1402 (O_1402,N_9113,N_9587);
nor UO_1403 (O_1403,N_9562,N_9139);
or UO_1404 (O_1404,N_9511,N_8045);
nor UO_1405 (O_1405,N_8231,N_9449);
or UO_1406 (O_1406,N_7692,N_8098);
or UO_1407 (O_1407,N_9891,N_9593);
or UO_1408 (O_1408,N_9919,N_7590);
and UO_1409 (O_1409,N_9008,N_9391);
or UO_1410 (O_1410,N_7685,N_9984);
and UO_1411 (O_1411,N_8333,N_7700);
nand UO_1412 (O_1412,N_8452,N_9508);
and UO_1413 (O_1413,N_8754,N_8654);
nand UO_1414 (O_1414,N_8445,N_8223);
nor UO_1415 (O_1415,N_7878,N_9947);
xor UO_1416 (O_1416,N_7864,N_9652);
nand UO_1417 (O_1417,N_7767,N_9062);
or UO_1418 (O_1418,N_9090,N_9417);
and UO_1419 (O_1419,N_7704,N_9996);
nor UO_1420 (O_1420,N_8933,N_9245);
nand UO_1421 (O_1421,N_7776,N_7701);
or UO_1422 (O_1422,N_9596,N_8242);
nand UO_1423 (O_1423,N_7791,N_8976);
nand UO_1424 (O_1424,N_7980,N_8489);
nor UO_1425 (O_1425,N_8511,N_9394);
nor UO_1426 (O_1426,N_9653,N_8427);
or UO_1427 (O_1427,N_9529,N_8319);
nor UO_1428 (O_1428,N_8798,N_9710);
nor UO_1429 (O_1429,N_8562,N_8914);
nand UO_1430 (O_1430,N_8377,N_8794);
and UO_1431 (O_1431,N_9087,N_9197);
nand UO_1432 (O_1432,N_8005,N_9389);
xnor UO_1433 (O_1433,N_7557,N_7642);
and UO_1434 (O_1434,N_8497,N_9651);
and UO_1435 (O_1435,N_8712,N_8127);
xnor UO_1436 (O_1436,N_8895,N_8262);
and UO_1437 (O_1437,N_9670,N_7818);
xor UO_1438 (O_1438,N_9307,N_9323);
and UO_1439 (O_1439,N_8024,N_9932);
and UO_1440 (O_1440,N_7808,N_8340);
nor UO_1441 (O_1441,N_9301,N_8597);
or UO_1442 (O_1442,N_8894,N_9864);
xor UO_1443 (O_1443,N_9878,N_8386);
and UO_1444 (O_1444,N_8372,N_8808);
xor UO_1445 (O_1445,N_8529,N_9883);
or UO_1446 (O_1446,N_8092,N_9773);
nor UO_1447 (O_1447,N_8082,N_9331);
xnor UO_1448 (O_1448,N_9924,N_9935);
xor UO_1449 (O_1449,N_8161,N_7978);
nand UO_1450 (O_1450,N_9566,N_8329);
nor UO_1451 (O_1451,N_7672,N_9054);
and UO_1452 (O_1452,N_7919,N_7940);
nand UO_1453 (O_1453,N_8245,N_8850);
nand UO_1454 (O_1454,N_7733,N_9950);
and UO_1455 (O_1455,N_7928,N_7793);
xnor UO_1456 (O_1456,N_8020,N_8310);
and UO_1457 (O_1457,N_8874,N_8328);
or UO_1458 (O_1458,N_9602,N_9774);
or UO_1459 (O_1459,N_9361,N_9778);
or UO_1460 (O_1460,N_9275,N_8744);
or UO_1461 (O_1461,N_8644,N_9523);
xnor UO_1462 (O_1462,N_7668,N_9625);
nor UO_1463 (O_1463,N_9961,N_9758);
xnor UO_1464 (O_1464,N_7667,N_7517);
nor UO_1465 (O_1465,N_7568,N_8597);
nor UO_1466 (O_1466,N_8668,N_8720);
xnor UO_1467 (O_1467,N_9409,N_9718);
nor UO_1468 (O_1468,N_9548,N_8990);
or UO_1469 (O_1469,N_8950,N_8356);
or UO_1470 (O_1470,N_8310,N_9166);
xnor UO_1471 (O_1471,N_8567,N_9792);
and UO_1472 (O_1472,N_8671,N_8793);
nor UO_1473 (O_1473,N_7824,N_9081);
or UO_1474 (O_1474,N_9477,N_8453);
nand UO_1475 (O_1475,N_8777,N_8598);
nor UO_1476 (O_1476,N_7975,N_8834);
nor UO_1477 (O_1477,N_9606,N_8556);
nand UO_1478 (O_1478,N_8357,N_9057);
or UO_1479 (O_1479,N_9413,N_9066);
nand UO_1480 (O_1480,N_8133,N_8713);
nand UO_1481 (O_1481,N_9505,N_9010);
nor UO_1482 (O_1482,N_9056,N_8796);
nor UO_1483 (O_1483,N_8083,N_8907);
nand UO_1484 (O_1484,N_8136,N_9686);
and UO_1485 (O_1485,N_8364,N_8930);
and UO_1486 (O_1486,N_7820,N_8668);
or UO_1487 (O_1487,N_9578,N_8446);
nand UO_1488 (O_1488,N_9055,N_7960);
or UO_1489 (O_1489,N_9852,N_7626);
and UO_1490 (O_1490,N_8611,N_8003);
and UO_1491 (O_1491,N_9452,N_9271);
and UO_1492 (O_1492,N_8937,N_8307);
and UO_1493 (O_1493,N_7580,N_9867);
nor UO_1494 (O_1494,N_9622,N_8476);
xnor UO_1495 (O_1495,N_9129,N_8823);
nor UO_1496 (O_1496,N_9595,N_9061);
nor UO_1497 (O_1497,N_8503,N_7963);
and UO_1498 (O_1498,N_8910,N_9259);
and UO_1499 (O_1499,N_8879,N_9591);
endmodule