module basic_3000_30000_3500_6_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_1951,In_2649);
and U1 (N_1,In_99,In_2107);
or U2 (N_2,In_664,In_2716);
and U3 (N_3,In_2638,In_2346);
xor U4 (N_4,In_2465,In_1872);
nand U5 (N_5,In_2602,In_1858);
nand U6 (N_6,In_1026,In_2013);
xor U7 (N_7,In_2031,In_867);
nand U8 (N_8,In_1154,In_305);
and U9 (N_9,In_2614,In_417);
and U10 (N_10,In_791,In_27);
nand U11 (N_11,In_2805,In_1160);
or U12 (N_12,In_2367,In_866);
and U13 (N_13,In_2523,In_1931);
nand U14 (N_14,In_2934,In_19);
xnor U15 (N_15,In_2084,In_1933);
nor U16 (N_16,In_2237,In_2749);
and U17 (N_17,In_1962,In_1470);
nor U18 (N_18,In_2265,In_1192);
xor U19 (N_19,In_2697,In_336);
nor U20 (N_20,In_1000,In_2291);
nor U21 (N_21,In_792,In_2741);
nand U22 (N_22,In_359,In_2177);
nand U23 (N_23,In_236,In_961);
or U24 (N_24,In_2621,In_2894);
nand U25 (N_25,In_738,In_697);
nor U26 (N_26,In_2920,In_178);
nor U27 (N_27,In_1821,In_1723);
nor U28 (N_28,In_2005,In_2678);
nor U29 (N_29,In_2190,In_1417);
nand U30 (N_30,In_2924,In_2342);
nor U31 (N_31,In_2516,In_1393);
and U32 (N_32,In_592,In_2313);
and U33 (N_33,In_1698,In_2268);
and U34 (N_34,In_973,In_569);
nand U35 (N_35,In_2685,In_2592);
or U36 (N_36,In_1203,In_905);
nand U37 (N_37,In_79,In_2792);
or U38 (N_38,In_2832,In_606);
nor U39 (N_39,In_1819,In_123);
nand U40 (N_40,In_1349,In_2316);
nor U41 (N_41,In_1800,In_307);
and U42 (N_42,In_1104,In_223);
or U43 (N_43,In_2821,In_1469);
or U44 (N_44,In_140,In_1188);
xnor U45 (N_45,In_1381,In_921);
or U46 (N_46,In_580,In_1194);
nand U47 (N_47,In_2979,In_428);
nor U48 (N_48,In_2051,In_2955);
nand U49 (N_49,In_1182,In_1429);
nor U50 (N_50,In_2566,In_2677);
nor U51 (N_51,In_1528,In_1530);
and U52 (N_52,In_427,In_477);
nor U53 (N_53,In_795,In_1881);
and U54 (N_54,In_2002,In_1685);
and U55 (N_55,In_479,In_1444);
or U56 (N_56,In_1582,In_2085);
or U57 (N_57,In_2389,In_2088);
nor U58 (N_58,In_2132,In_2189);
and U59 (N_59,In_304,In_1700);
nor U60 (N_60,In_462,In_2992);
nor U61 (N_61,In_702,In_2562);
nor U62 (N_62,In_1015,In_370);
xor U63 (N_63,In_2783,In_2989);
nor U64 (N_64,In_1047,In_2670);
nand U65 (N_65,In_1190,In_2522);
nand U66 (N_66,In_2744,In_2674);
nor U67 (N_67,In_1979,In_1006);
xor U68 (N_68,In_1851,In_1930);
nand U69 (N_69,In_2248,In_1435);
nand U70 (N_70,In_208,In_2167);
xnor U71 (N_71,In_607,In_458);
nand U72 (N_72,In_2943,In_2405);
nand U73 (N_73,In_2683,In_2915);
and U74 (N_74,In_104,In_597);
and U75 (N_75,In_12,In_1892);
nand U76 (N_76,In_1361,In_555);
nor U77 (N_77,In_1603,In_967);
and U78 (N_78,In_1390,In_167);
or U79 (N_79,In_872,In_2066);
and U80 (N_80,In_1826,In_1277);
nor U81 (N_81,In_2143,In_1511);
nor U82 (N_82,In_2350,In_2220);
or U83 (N_83,In_719,In_1343);
nand U84 (N_84,In_2175,In_1988);
nand U85 (N_85,In_1012,In_2323);
or U86 (N_86,In_2283,In_810);
nand U87 (N_87,In_1082,In_2254);
or U88 (N_88,In_1269,In_1123);
nand U89 (N_89,In_940,In_2266);
nor U90 (N_90,In_2038,In_480);
or U91 (N_91,In_1344,In_2339);
nand U92 (N_92,In_249,In_2871);
or U93 (N_93,In_1611,In_471);
or U94 (N_94,In_168,In_988);
or U95 (N_95,In_668,In_920);
and U96 (N_96,In_1298,In_269);
xor U97 (N_97,In_882,In_2882);
nand U98 (N_98,In_913,In_1897);
and U99 (N_99,In_235,In_2988);
nor U100 (N_100,In_1706,In_2176);
or U101 (N_101,In_1455,In_784);
nand U102 (N_102,In_847,In_1790);
nand U103 (N_103,In_2462,In_239);
or U104 (N_104,In_112,In_2642);
nand U105 (N_105,In_2021,In_1338);
and U106 (N_106,In_2470,In_2327);
nand U107 (N_107,In_959,In_1620);
or U108 (N_108,In_1863,In_2489);
nand U109 (N_109,In_2635,In_133);
and U110 (N_110,In_2448,In_2954);
or U111 (N_111,In_274,In_1260);
nor U112 (N_112,In_2769,In_1337);
or U113 (N_113,In_1382,In_290);
nor U114 (N_114,In_1908,In_1735);
or U115 (N_115,In_2914,In_1447);
and U116 (N_116,In_2607,In_957);
nand U117 (N_117,In_2329,In_2536);
nor U118 (N_118,In_1781,In_553);
xnor U119 (N_119,In_338,In_2215);
nor U120 (N_120,In_86,In_677);
and U121 (N_121,In_2898,In_2588);
or U122 (N_122,In_296,In_1297);
and U123 (N_123,In_1063,In_2634);
nor U124 (N_124,In_1958,In_2491);
nor U125 (N_125,In_363,In_979);
and U126 (N_126,In_2969,In_2127);
nand U127 (N_127,In_789,In_895);
xor U128 (N_128,In_1596,In_1542);
and U129 (N_129,In_2715,In_92);
nand U130 (N_130,In_1887,In_651);
nand U131 (N_131,In_1374,In_2145);
nor U132 (N_132,In_2009,In_519);
and U133 (N_133,In_2856,In_453);
and U134 (N_134,In_466,In_2549);
nand U135 (N_135,In_2766,In_2723);
xnor U136 (N_136,In_575,In_2394);
or U137 (N_137,In_340,In_1757);
or U138 (N_138,In_1984,In_35);
and U139 (N_139,In_217,In_1276);
and U140 (N_140,In_284,In_253);
or U141 (N_141,In_134,In_1072);
xor U142 (N_142,In_1701,In_1245);
xnor U143 (N_143,In_467,In_1322);
nor U144 (N_144,In_2318,In_2192);
or U145 (N_145,In_1605,In_685);
and U146 (N_146,In_1546,In_2270);
nor U147 (N_147,In_1999,In_2324);
or U148 (N_148,In_1731,In_2016);
and U149 (N_149,In_2539,In_2358);
or U150 (N_150,In_1938,In_2960);
and U151 (N_151,In_1630,In_73);
and U152 (N_152,In_1064,In_2774);
or U153 (N_153,In_1873,In_507);
and U154 (N_154,In_489,In_2015);
nand U155 (N_155,In_1207,In_1778);
nand U156 (N_156,In_1849,In_2378);
xor U157 (N_157,In_1643,In_523);
and U158 (N_158,In_1783,In_2740);
nand U159 (N_159,In_2393,In_1848);
or U160 (N_160,In_2933,In_684);
nand U161 (N_161,In_1493,In_2935);
xor U162 (N_162,In_2633,In_2403);
nand U163 (N_163,In_308,In_2781);
or U164 (N_164,In_837,In_715);
and U165 (N_165,In_1810,In_2042);
nor U166 (N_166,In_82,In_2879);
or U167 (N_167,In_1717,In_823);
nand U168 (N_168,In_1220,In_2929);
and U169 (N_169,In_2250,In_1593);
nand U170 (N_170,In_2983,In_2593);
or U171 (N_171,In_1193,In_1299);
and U172 (N_172,In_77,In_2527);
and U173 (N_173,In_564,In_17);
nand U174 (N_174,In_209,In_444);
nand U175 (N_175,In_2867,In_566);
or U176 (N_176,In_412,In_889);
xor U177 (N_177,In_2807,In_2325);
nor U178 (N_178,In_549,In_909);
nand U179 (N_179,In_380,In_1023);
nor U180 (N_180,In_2278,In_716);
nor U181 (N_181,In_1882,In_2862);
and U182 (N_182,In_53,In_2753);
and U183 (N_183,In_232,In_741);
and U184 (N_184,In_2946,In_1041);
nor U185 (N_185,In_2353,In_590);
or U186 (N_186,In_1852,In_385);
and U187 (N_187,In_2654,In_583);
or U188 (N_188,In_171,In_2445);
nand U189 (N_189,In_1316,In_1574);
and U190 (N_190,In_1871,In_998);
nand U191 (N_191,In_2776,In_1215);
or U192 (N_192,In_2761,In_733);
or U193 (N_193,In_887,In_983);
nor U194 (N_194,In_2387,In_828);
nor U195 (N_195,In_54,In_577);
nor U196 (N_196,In_2736,In_1143);
nor U197 (N_197,In_2952,In_721);
xor U198 (N_198,In_2124,In_2440);
or U199 (N_199,In_2902,In_874);
xor U200 (N_200,In_917,In_1088);
or U201 (N_201,In_778,In_2599);
nor U202 (N_202,In_579,In_1742);
nand U203 (N_203,In_1949,In_2106);
nand U204 (N_204,In_306,In_1607);
or U205 (N_205,In_2974,In_1524);
and U206 (N_206,In_391,In_986);
and U207 (N_207,In_2354,In_1670);
and U208 (N_208,In_672,In_110);
nor U209 (N_209,In_2351,In_1782);
or U210 (N_210,In_1665,In_757);
or U211 (N_211,In_135,In_1902);
nor U212 (N_212,In_2560,In_1387);
nor U213 (N_213,In_1624,In_1895);
or U214 (N_214,In_1886,In_100);
or U215 (N_215,In_1773,In_2461);
and U216 (N_216,In_1971,In_500);
and U217 (N_217,In_1310,In_1446);
or U218 (N_218,In_1463,In_2721);
and U219 (N_219,In_491,In_2137);
nor U220 (N_220,In_2460,In_439);
xnor U221 (N_221,In_522,In_1237);
xnor U222 (N_222,In_1651,In_197);
and U223 (N_223,In_2398,In_871);
xor U224 (N_224,In_857,In_2108);
nand U225 (N_225,In_2950,In_1648);
xnor U226 (N_226,In_169,In_1081);
or U227 (N_227,In_2646,In_1549);
or U228 (N_228,In_2571,In_93);
or U229 (N_229,In_1021,In_2547);
nor U230 (N_230,In_2476,In_2280);
nor U231 (N_231,In_2391,In_573);
and U232 (N_232,In_87,In_1140);
nor U233 (N_233,In_1721,In_2857);
or U234 (N_234,In_2616,In_2964);
nand U235 (N_235,In_2511,In_1476);
and U236 (N_236,In_2851,In_1766);
and U237 (N_237,In_2415,In_855);
xor U238 (N_238,In_2503,In_506);
and U239 (N_239,In_517,In_226);
or U240 (N_240,In_145,In_1953);
and U241 (N_241,In_1924,In_455);
nor U242 (N_242,In_1947,In_885);
xor U243 (N_243,In_122,In_640);
nand U244 (N_244,In_854,In_215);
nand U245 (N_245,In_176,In_2409);
nor U246 (N_246,In_2453,In_2793);
or U247 (N_247,In_747,In_671);
and U248 (N_248,In_578,In_128);
and U249 (N_249,In_2225,In_1516);
xnor U250 (N_250,In_831,In_1442);
nor U251 (N_251,In_1765,In_2606);
or U252 (N_252,In_834,In_2153);
and U253 (N_253,In_1769,In_1481);
or U254 (N_254,In_755,In_746);
nor U255 (N_255,In_325,In_13);
nor U256 (N_256,In_1640,In_493);
nand U257 (N_257,In_2029,In_1535);
nor U258 (N_258,In_1108,In_273);
xnor U259 (N_259,In_2884,In_1919);
or U260 (N_260,In_2500,In_1366);
nor U261 (N_261,In_107,In_1234);
nand U262 (N_262,In_204,In_2800);
xnor U263 (N_263,In_930,In_2840);
and U264 (N_264,In_2348,In_423);
and U265 (N_265,In_1622,In_2008);
or U266 (N_266,In_2594,In_1289);
nand U267 (N_267,In_2033,In_334);
or U268 (N_268,In_1578,In_775);
or U269 (N_269,In_1279,In_1219);
xnor U270 (N_270,In_2151,In_2200);
and U271 (N_271,In_1649,In_2073);
xor U272 (N_272,In_648,In_1936);
or U273 (N_273,In_432,In_1208);
xor U274 (N_274,In_804,In_1818);
and U275 (N_275,In_413,In_2680);
and U276 (N_276,In_2385,In_229);
or U277 (N_277,In_2229,In_562);
nand U278 (N_278,In_1427,In_399);
nor U279 (N_279,In_2502,In_2247);
nor U280 (N_280,In_536,In_2994);
nor U281 (N_281,In_951,In_2519);
nor U282 (N_282,In_1018,In_1537);
and U283 (N_283,In_1167,In_928);
nor U284 (N_284,In_632,In_2427);
xnor U285 (N_285,In_908,In_1471);
or U286 (N_286,In_873,In_1084);
and U287 (N_287,In_1307,In_1967);
and U288 (N_288,In_749,In_2990);
xnor U289 (N_289,In_2058,In_939);
nand U290 (N_290,In_2298,In_1312);
nor U291 (N_291,In_1974,In_310);
nand U292 (N_292,In_976,In_311);
nor U293 (N_293,In_1691,In_29);
xor U294 (N_294,In_1392,In_618);
and U295 (N_295,In_2425,In_1532);
nor U296 (N_296,In_2657,In_1472);
or U297 (N_297,In_2624,In_1078);
and U298 (N_298,In_2217,In_2883);
nand U299 (N_299,In_2704,In_1166);
nand U300 (N_300,In_487,In_1761);
nor U301 (N_301,In_1106,In_510);
or U302 (N_302,In_2973,In_1907);
xor U303 (N_303,In_2839,In_954);
or U304 (N_304,In_1326,In_1645);
nand U305 (N_305,In_2640,In_159);
and U306 (N_306,In_2376,In_2352);
nand U307 (N_307,In_2302,In_1340);
nand U308 (N_308,In_2865,In_1294);
or U309 (N_309,In_730,In_2564);
nand U310 (N_310,In_2004,In_2942);
nand U311 (N_311,In_1384,In_1667);
nand U312 (N_312,In_674,In_2428);
and U313 (N_313,In_2396,In_266);
and U314 (N_314,In_720,In_1689);
and U315 (N_315,In_2173,In_1270);
nor U316 (N_316,In_431,In_2292);
or U317 (N_317,In_1341,In_881);
or U318 (N_318,In_2052,In_241);
nand U319 (N_319,In_2446,In_1466);
nand U320 (N_320,In_2402,In_2355);
nand U321 (N_321,In_964,In_1797);
or U322 (N_322,In_1929,In_1457);
nand U323 (N_323,In_2861,In_1856);
and U324 (N_324,In_2010,In_1705);
nor U325 (N_325,In_330,In_1816);
nor U326 (N_326,In_2538,In_2034);
and U327 (N_327,In_814,In_2320);
or U328 (N_328,In_1490,In_314);
or U329 (N_329,In_2876,In_260);
and U330 (N_330,In_2521,In_2639);
nand U331 (N_331,In_603,In_748);
nand U332 (N_332,In_2997,In_1432);
or U333 (N_333,In_904,In_761);
and U334 (N_334,In_1827,In_151);
and U335 (N_335,In_1504,In_1050);
nand U336 (N_336,In_395,In_1296);
nand U337 (N_337,In_2012,In_326);
nor U338 (N_338,In_2149,In_1776);
nor U339 (N_339,In_1865,In_1448);
nand U340 (N_340,In_827,In_1571);
and U341 (N_341,In_117,In_1687);
and U342 (N_342,In_806,In_2667);
xor U343 (N_343,In_699,In_138);
and U344 (N_344,In_824,In_1709);
nor U345 (N_345,In_916,In_1342);
nor U346 (N_346,In_1077,In_1495);
nand U347 (N_347,In_2507,In_1842);
nand U348 (N_348,In_1060,In_2494);
nor U349 (N_349,In_1673,In_1306);
nand U350 (N_350,In_2157,In_1346);
or U351 (N_351,In_240,In_196);
nor U352 (N_352,In_1257,In_418);
or U353 (N_353,In_335,In_2122);
xor U354 (N_354,In_1246,In_2183);
nand U355 (N_355,In_1889,In_1059);
xnor U356 (N_356,In_565,In_1066);
nand U357 (N_357,In_2650,In_96);
xnor U358 (N_358,In_1625,In_2510);
or U359 (N_359,In_2178,In_2758);
nand U360 (N_360,In_2155,In_1254);
or U361 (N_361,In_1132,In_2158);
nor U362 (N_362,In_2970,In_1421);
nand U363 (N_363,In_2032,In_525);
or U364 (N_364,In_2885,In_2238);
nand U365 (N_365,In_2362,In_2910);
nand U366 (N_366,In_2152,In_321);
or U367 (N_367,In_1811,In_2931);
nor U368 (N_368,In_1551,In_1362);
nor U369 (N_369,In_262,In_833);
nand U370 (N_370,In_275,In_820);
or U371 (N_371,In_1492,In_1225);
nand U372 (N_372,In_2431,In_1966);
xor U373 (N_373,In_2475,In_2813);
xor U374 (N_374,In_1868,In_392);
nand U375 (N_375,In_1556,In_1646);
or U376 (N_376,In_1692,In_2615);
nand U377 (N_377,In_2214,In_2858);
nand U378 (N_378,In_1049,In_2371);
nor U379 (N_379,In_2087,In_374);
and U380 (N_380,In_2919,In_840);
nand U381 (N_381,In_2868,In_68);
and U382 (N_382,In_102,In_1156);
and U383 (N_383,In_766,In_629);
and U384 (N_384,In_718,In_156);
nand U385 (N_385,In_2109,In_200);
nor U386 (N_386,In_1239,In_623);
nor U387 (N_387,In_201,In_55);
or U388 (N_388,In_2687,In_722);
nor U389 (N_389,In_2061,In_756);
and U390 (N_390,In_910,In_205);
nor U391 (N_391,In_1575,In_245);
or U392 (N_392,In_1029,In_1229);
nand U393 (N_393,In_1674,In_596);
and U394 (N_394,In_1621,In_1209);
and U395 (N_395,In_2819,In_644);
and U396 (N_396,In_2720,In_376);
nor U397 (N_397,In_1359,In_2976);
nand U398 (N_398,In_468,In_1459);
nand U399 (N_399,In_1976,In_2574);
or U400 (N_400,In_924,In_1354);
nand U401 (N_401,In_647,In_1584);
and U402 (N_402,In_2047,In_103);
nand U403 (N_403,In_160,In_767);
and U404 (N_404,In_2784,In_667);
nor U405 (N_405,In_341,In_2755);
or U406 (N_406,In_1367,In_2754);
xnor U407 (N_407,In_1468,In_2558);
nor U408 (N_408,In_852,In_1515);
and U409 (N_409,In_407,In_2811);
or U410 (N_410,In_978,In_187);
nand U411 (N_411,In_2568,In_680);
nor U412 (N_412,In_403,In_485);
and U413 (N_413,In_1750,In_2294);
and U414 (N_414,In_843,In_2307);
nor U415 (N_415,In_1775,In_2452);
or U416 (N_416,In_1870,In_1807);
or U417 (N_417,In_587,In_830);
nand U418 (N_418,In_595,In_1904);
nor U419 (N_419,In_688,In_2836);
and U420 (N_420,In_542,In_2386);
nand U421 (N_421,In_1096,In_353);
nor U422 (N_422,In_2748,In_2202);
or U423 (N_423,In_1615,In_605);
and U424 (N_424,In_2565,In_1200);
nand U425 (N_425,In_1682,In_776);
or U426 (N_426,In_2791,In_1631);
nor U427 (N_427,In_1512,In_2197);
nand U428 (N_428,In_11,In_2347);
nor U429 (N_429,In_676,In_2605);
and U430 (N_430,In_781,In_581);
or U431 (N_431,In_425,In_1869);
xnor U432 (N_432,In_348,In_221);
xnor U433 (N_433,In_2742,In_1116);
or U434 (N_434,In_281,In_2121);
or U435 (N_435,In_1487,In_1710);
nand U436 (N_436,In_2673,In_2543);
and U437 (N_437,In_1331,In_1025);
nand U438 (N_438,In_2552,In_842);
nand U439 (N_439,In_546,In_23);
and U440 (N_440,In_1564,In_1583);
nor U441 (N_441,In_1360,In_2222);
nor U442 (N_442,In_2728,In_787);
xor U443 (N_443,In_2421,In_2866);
or U444 (N_444,In_2810,In_768);
and U445 (N_445,In_1830,In_63);
or U446 (N_446,In_2414,In_1558);
nand U447 (N_447,In_2477,In_649);
or U448 (N_448,In_255,In_1035);
and U449 (N_449,In_433,In_2844);
nand U450 (N_450,In_1076,In_2799);
nor U451 (N_451,In_1725,In_2665);
nor U452 (N_452,In_1690,In_14);
nor U453 (N_453,In_965,In_2553);
xor U454 (N_454,In_2893,In_550);
nor U455 (N_455,In_2435,In_530);
and U456 (N_456,In_1879,In_292);
nor U457 (N_457,In_47,In_400);
nand U458 (N_458,In_533,In_1428);
nand U459 (N_459,In_2903,In_2583);
or U460 (N_460,In_276,In_2561);
nor U461 (N_461,In_84,In_2864);
or U462 (N_462,In_1880,In_2760);
xnor U463 (N_463,In_1676,In_626);
nor U464 (N_464,In_2656,In_1259);
nand U465 (N_465,In_1946,In_802);
nor U466 (N_466,In_2384,In_2762);
or U467 (N_467,In_101,In_270);
or U468 (N_468,In_858,In_1119);
nand U469 (N_469,In_1738,In_1204);
nand U470 (N_470,In_1244,In_1653);
and U471 (N_471,In_2366,In_2365);
nor U472 (N_472,In_1439,In_119);
nand U473 (N_473,In_1370,In_2636);
nor U474 (N_474,In_464,In_131);
or U475 (N_475,In_1832,In_696);
nand U476 (N_476,In_896,In_1732);
xor U477 (N_477,In_2257,In_687);
or U478 (N_478,In_1426,In_1008);
nor U479 (N_479,In_1960,In_278);
xor U480 (N_480,In_1695,In_2922);
nand U481 (N_481,In_848,In_2301);
or U482 (N_482,In_1825,In_2699);
xnor U483 (N_483,In_2095,In_454);
and U484 (N_484,In_2717,In_797);
and U485 (N_485,In_4,In_970);
nor U486 (N_486,In_2182,In_243);
nor U487 (N_487,In_202,In_61);
and U488 (N_488,In_1896,In_1386);
xnor U489 (N_489,In_1027,In_870);
and U490 (N_490,In_2060,In_2118);
nor U491 (N_491,In_2785,In_2514);
or U492 (N_492,In_2727,In_1718);
nand U493 (N_493,In_2056,In_2269);
nand U494 (N_494,In_157,In_1044);
and U495 (N_495,In_2901,In_1126);
and U496 (N_496,In_1975,In_1040);
or U497 (N_497,In_1996,In_1201);
nor U498 (N_498,In_233,In_1965);
and U499 (N_499,In_1068,In_2211);
or U500 (N_500,In_693,In_557);
and U501 (N_501,In_438,In_1350);
and U502 (N_502,In_815,In_2493);
nand U503 (N_503,In_1062,In_1763);
nand U504 (N_504,In_1402,In_1599);
nor U505 (N_505,In_925,In_461);
nand U506 (N_506,In_2408,In_146);
nand U507 (N_507,In_2530,In_1037);
nand U508 (N_508,In_2747,In_2105);
or U509 (N_509,In_446,In_195);
nor U510 (N_510,In_303,In_888);
nand U511 (N_511,In_1719,In_2773);
nor U512 (N_512,In_1683,In_1854);
and U513 (N_513,In_505,In_1022);
nor U514 (N_514,In_927,In_2300);
nand U515 (N_515,In_347,In_283);
nand U516 (N_516,In_2987,In_2891);
and U517 (N_517,In_2996,In_512);
and U518 (N_518,In_1510,In_1736);
or U519 (N_519,In_2570,In_191);
nand U520 (N_520,In_2967,In_2587);
or U521 (N_521,In_2698,In_2091);
nor U522 (N_522,In_2652,In_2125);
and U523 (N_523,In_173,In_2199);
or U524 (N_524,In_993,In_734);
and U525 (N_525,In_2490,In_2820);
and U526 (N_526,In_1061,In_2369);
and U527 (N_527,In_1952,In_944);
and U528 (N_528,In_657,In_2030);
nand U529 (N_529,In_938,In_421);
or U530 (N_530,In_864,In_1831);
nor U531 (N_531,In_673,In_437);
and U532 (N_532,In_349,In_1550);
nor U533 (N_533,In_182,In_953);
or U534 (N_534,In_1661,In_2046);
nand U535 (N_535,In_1642,In_631);
xor U536 (N_536,In_935,In_1085);
nand U537 (N_537,In_1232,In_378);
and U538 (N_538,In_1726,In_20);
nand U539 (N_539,In_992,In_2627);
nand U540 (N_540,In_456,In_2231);
or U541 (N_541,In_1594,In_2092);
and U542 (N_542,In_1369,In_2963);
or U543 (N_543,In_2732,In_822);
and U544 (N_544,In_2113,In_1998);
nand U545 (N_545,In_1989,In_495);
or U546 (N_546,In_1177,In_798);
or U547 (N_547,In_2923,In_2338);
and U548 (N_548,In_2442,In_198);
and U549 (N_549,In_877,In_2998);
and U550 (N_550,In_2383,In_1634);
nor U551 (N_551,In_469,In_120);
and U552 (N_552,In_1138,In_1454);
nand U553 (N_553,In_1679,In_2708);
nand U554 (N_554,In_2968,In_2416);
nor U555 (N_555,In_2028,In_2472);
and U556 (N_556,In_1993,In_876);
and U557 (N_557,In_1389,In_594);
nor U558 (N_558,In_2289,In_1655);
or U559 (N_559,In_520,In_361);
or U560 (N_560,In_2601,In_2567);
and U561 (N_561,In_1145,In_902);
or U562 (N_562,In_1329,In_1555);
nand U563 (N_563,In_1313,In_574);
nor U564 (N_564,In_2959,In_237);
nand U565 (N_565,In_2837,In_1236);
nand U566 (N_566,In_2406,In_801);
nor U567 (N_567,In_1489,In_934);
nand U568 (N_568,In_1149,In_58);
or U569 (N_569,In_1632,In_2644);
nand U570 (N_570,In_1748,In_1118);
nor U571 (N_571,In_2756,In_1514);
or U572 (N_572,In_1527,In_1371);
or U573 (N_573,In_1074,In_2925);
xor U574 (N_574,In_36,In_1434);
or U575 (N_575,In_2534,In_1823);
nand U576 (N_576,In_1416,In_132);
nand U577 (N_577,In_2326,In_1168);
or U578 (N_578,In_1176,In_496);
nor U579 (N_579,In_691,In_1635);
nand U580 (N_580,In_2279,In_1302);
xor U581 (N_581,In_2076,In_2201);
and U582 (N_582,In_1753,In_429);
and U583 (N_583,In_724,In_1292);
and U584 (N_584,In_2166,In_1983);
nand U585 (N_585,In_52,In_899);
and U586 (N_586,In_819,In_2123);
or U587 (N_587,In_231,In_1538);
nor U588 (N_588,In_799,In_1995);
and U589 (N_589,In_424,In_600);
nand U590 (N_590,In_113,In_1780);
or U591 (N_591,In_2713,In_1478);
or U592 (N_592,In_2572,In_1503);
nand U593 (N_593,In_1336,In_1668);
or U594 (N_594,In_1090,In_838);
or U595 (N_595,In_2563,In_2459);
nand U596 (N_596,In_2827,In_1315);
or U597 (N_597,In_2999,In_297);
nand U598 (N_598,In_2815,In_2055);
nor U599 (N_599,In_2763,In_2528);
nand U600 (N_600,In_2048,In_449);
or U601 (N_601,In_139,In_1660);
nor U602 (N_602,In_844,In_790);
nor U603 (N_603,In_2234,In_220);
or U604 (N_604,In_1205,In_524);
nand U605 (N_605,In_868,In_2418);
and U606 (N_606,In_1456,In_2335);
nand U607 (N_607,In_1186,In_2438);
nand U608 (N_608,In_1637,In_662);
nor U609 (N_609,In_545,In_2395);
xor U610 (N_610,In_1754,In_758);
or U611 (N_611,In_638,In_2277);
nand U612 (N_612,In_2613,In_1039);
nand U613 (N_613,In_946,In_154);
or U614 (N_614,In_484,In_1042);
and U615 (N_615,In_1227,In_1274);
nand U616 (N_616,In_1768,In_1170);
or U617 (N_617,In_862,In_2133);
nor U618 (N_618,In_1628,In_2172);
nor U619 (N_619,In_2743,In_1494);
or U620 (N_620,In_1058,In_912);
and U621 (N_621,In_937,In_1226);
nand U622 (N_622,In_703,In_2682);
nor U623 (N_623,In_279,In_440);
nand U624 (N_624,In_572,In_2496);
nor U625 (N_625,In_2411,In_1716);
xnor U626 (N_626,In_2545,In_2332);
xor U627 (N_627,In_322,In_2473);
nand U628 (N_628,In_2436,In_161);
and U629 (N_629,In_502,In_2317);
and U630 (N_630,In_177,In_2432);
nand U631 (N_631,In_650,In_2382);
or U632 (N_632,In_2870,In_1185);
and U633 (N_633,In_2018,In_179);
and U634 (N_634,In_288,In_2449);
or U635 (N_635,In_293,In_2114);
or U636 (N_636,In_898,In_1217);
nor U637 (N_637,In_955,In_2180);
or U638 (N_638,In_1334,In_2814);
or U639 (N_639,In_2185,In_1536);
and U640 (N_640,In_2647,In_2466);
xor U641 (N_641,In_2083,In_144);
and U642 (N_642,In_387,In_2207);
nor U643 (N_643,In_2424,In_65);
nor U644 (N_644,In_2,In_1534);
nand U645 (N_645,In_365,In_654);
or U646 (N_646,In_114,In_1100);
nand U647 (N_647,In_2093,In_1323);
and U648 (N_648,In_2945,In_2104);
and U649 (N_649,In_883,In_2196);
nand U650 (N_650,In_356,In_1715);
and U651 (N_651,In_254,In_116);
nor U652 (N_652,In_38,In_2757);
or U653 (N_653,In_2542,In_1057);
nor U654 (N_654,In_1752,In_2050);
nand U655 (N_655,In_2219,In_1496);
xor U656 (N_656,In_30,In_1388);
and U657 (N_657,In_949,In_2806);
and U658 (N_658,In_251,In_1400);
or U659 (N_659,In_1843,In_2399);
nand U660 (N_660,In_544,In_222);
and U661 (N_661,In_1650,In_2357);
nor U662 (N_662,In_1121,In_2099);
xnor U663 (N_663,In_1377,In_2306);
and U664 (N_664,In_1610,In_227);
nor U665 (N_665,In_2711,In_2159);
xnor U666 (N_666,In_762,In_148);
nand U667 (N_667,In_932,In_2900);
nand U668 (N_668,In_1948,In_1867);
nand U669 (N_669,In_1910,In_2778);
nor U670 (N_670,In_2360,In_1214);
xnor U671 (N_671,In_372,In_470);
nand U672 (N_672,In_2912,In_2916);
xnor U673 (N_673,In_2086,In_1609);
or U674 (N_674,In_2241,In_1301);
nor U675 (N_675,In_2193,In_2625);
xor U676 (N_676,In_2610,In_616);
nand U677 (N_677,In_1179,In_665);
nand U678 (N_678,In_1704,In_2433);
xor U679 (N_679,In_1189,In_731);
or U680 (N_680,In_420,In_2694);
or U681 (N_681,In_2223,In_450);
and U682 (N_682,In_2904,In_342);
or U683 (N_683,In_2710,In_947);
xnor U684 (N_684,In_2311,In_2730);
xor U685 (N_685,In_2469,In_865);
nor U686 (N_686,In_106,In_2256);
nand U687 (N_687,In_1702,In_1923);
nor U688 (N_688,In_1211,In_1834);
nand U689 (N_689,In_2260,In_2027);
nor U690 (N_690,In_742,In_1588);
nor U691 (N_691,In_1355,In_1547);
or U692 (N_692,In_1411,In_2794);
xor U693 (N_693,In_1320,In_2349);
or U694 (N_694,In_1985,In_2580);
and U695 (N_695,In_675,In_2729);
and U696 (N_696,In_1739,In_2859);
xor U697 (N_697,In_782,In_1922);
nor U698 (N_698,In_2823,In_206);
nor U699 (N_699,In_2689,In_2097);
nand U700 (N_700,In_918,In_371);
nand U701 (N_701,In_1488,In_825);
or U702 (N_702,In_1019,In_1791);
and U703 (N_703,In_974,In_901);
nor U704 (N_704,In_860,In_1169);
nand U705 (N_705,In_2596,In_1927);
nor U706 (N_706,In_436,In_2194);
or U707 (N_707,In_637,In_1364);
or U708 (N_708,In_2872,In_1069);
or U709 (N_709,In_1445,In_2848);
nor U710 (N_710,In_2874,In_1171);
nor U711 (N_711,In_692,In_2343);
xnor U712 (N_712,In_261,In_663);
and U713 (N_713,In_1333,In_1614);
xnor U714 (N_714,In_210,In_622);
or U715 (N_715,In_2102,In_511);
nand U716 (N_716,In_2262,In_999);
or U717 (N_717,In_2274,In_1174);
nand U718 (N_718,In_435,In_1513);
nand U719 (N_719,In_1707,In_2917);
and U720 (N_720,In_2972,In_1900);
nor U721 (N_721,In_1325,In_1912);
or U722 (N_722,In_1351,In_1142);
nor U723 (N_723,In_2853,In_2098);
and U724 (N_724,In_2171,In_194);
nand U725 (N_725,In_2331,In_2725);
nor U726 (N_726,In_763,In_926);
and U727 (N_727,In_2077,In_1916);
nand U728 (N_728,In_430,In_745);
and U729 (N_729,In_2750,In_1841);
xor U730 (N_730,In_1678,In_537);
xor U731 (N_731,In_2138,In_2255);
or U732 (N_732,In_2454,In_2873);
nand U733 (N_733,In_1557,In_1941);
xor U734 (N_734,In_1977,In_1124);
and U735 (N_735,In_175,In_891);
and U736 (N_736,In_2645,In_422);
nand U737 (N_737,In_2825,In_360);
or U738 (N_738,In_2535,In_1802);
nor U739 (N_739,In_2471,In_1267);
or U740 (N_740,In_1441,In_2938);
nor U741 (N_741,In_118,In_987);
nor U742 (N_742,In_2575,In_796);
and U743 (N_743,In_1275,In_2966);
nand U744 (N_744,In_2246,In_1569);
nand U745 (N_745,In_2112,In_2430);
xor U746 (N_746,In_2288,In_1114);
nor U747 (N_747,In_1449,In_1568);
xor U748 (N_748,In_1874,In_2796);
and U749 (N_749,In_1525,In_1278);
xnor U750 (N_750,In_1309,In_2410);
nor U751 (N_751,In_636,In_619);
and U752 (N_752,In_2263,In_599);
nand U753 (N_753,In_2632,In_2537);
or U754 (N_754,In_1083,In_1395);
nor U755 (N_755,In_2591,In_2019);
and U756 (N_756,In_401,In_460);
nor U757 (N_757,In_1945,In_1055);
nand U758 (N_758,In_2569,In_2737);
and U759 (N_759,In_31,In_1137);
and U760 (N_760,In_771,In_914);
and U761 (N_761,In_1828,In_2629);
nand U762 (N_762,In_2508,In_1353);
nor U763 (N_763,In_698,In_390);
and U764 (N_764,In_2457,In_783);
nor U765 (N_765,In_2532,In_2962);
nand U766 (N_766,In_551,In_465);
nor U767 (N_767,In_1010,In_1437);
nand U768 (N_768,In_1460,In_2531);
xor U769 (N_769,In_91,In_1348);
and U770 (N_770,In_2467,In_1767);
or U771 (N_771,In_80,In_1619);
nor U772 (N_772,In_547,In_1221);
and U773 (N_773,In_472,In_15);
and U774 (N_774,In_1885,In_966);
or U775 (N_775,In_2497,In_2714);
xor U776 (N_776,In_2426,In_1133);
nand U777 (N_777,In_1982,In_1862);
nand U778 (N_778,In_604,In_98);
and U779 (N_779,In_1864,In_1223);
or U780 (N_780,In_1795,In_2905);
nand U781 (N_781,In_354,In_318);
or U782 (N_782,In_2822,In_1693);
nor U783 (N_783,In_2096,In_661);
nor U784 (N_784,In_737,In_1198);
and U785 (N_785,In_2878,In_821);
and U786 (N_786,In_1708,In_2146);
or U787 (N_787,In_2209,In_1376);
nand U788 (N_788,In_1147,In_879);
xor U789 (N_789,In_1419,In_1838);
or U790 (N_790,In_1385,In_543);
nor U791 (N_791,In_2653,In_1373);
and U792 (N_792,In_2579,In_1002);
or U793 (N_793,In_1921,In_1243);
xor U794 (N_794,In_2608,In_2977);
nand U795 (N_795,In_1407,In_807);
or U796 (N_796,In_2770,In_441);
or U797 (N_797,In_2363,In_2513);
or U798 (N_798,In_1794,In_2341);
nand U799 (N_799,In_2011,In_1552);
nor U800 (N_800,In_1180,In_1680);
nand U801 (N_801,In_271,In_2078);
and U802 (N_802,In_1409,In_33);
xnor U803 (N_803,In_2506,In_1666);
and U804 (N_804,In_1639,In_710);
nand U805 (N_805,In_459,In_759);
and U806 (N_806,In_2210,In_2314);
and U807 (N_807,In_2499,In_1291);
nand U808 (N_808,In_2419,In_1418);
or U809 (N_809,In_1300,In_2829);
nor U810 (N_810,In_527,In_327);
or U811 (N_811,In_1383,In_2160);
nand U812 (N_812,In_1601,In_2828);
or U813 (N_813,In_713,In_2062);
and U814 (N_814,In_2734,In_2044);
nand U815 (N_815,In_2412,In_1303);
xor U816 (N_816,In_1266,In_2622);
xnor U817 (N_817,In_2928,In_331);
nand U818 (N_818,In_1153,In_863);
xor U819 (N_819,In_845,In_1436);
nor U820 (N_820,In_1860,In_1330);
or U821 (N_821,In_346,In_2686);
nor U822 (N_822,In_773,In_656);
nand U823 (N_823,In_1408,In_1175);
and U824 (N_824,In_2486,In_2559);
nor U825 (N_825,In_1671,In_7);
xor U826 (N_826,In_2128,In_1253);
and U827 (N_827,In_1627,In_1508);
or U828 (N_828,In_706,In_2668);
and U829 (N_829,In_1053,In_192);
and U830 (N_830,In_2162,In_903);
or U831 (N_831,In_1099,In_2150);
nand U832 (N_832,In_1617,In_1560);
or U833 (N_833,In_1152,In_2577);
nand U834 (N_834,In_1932,In_627);
nand U835 (N_835,In_2407,In_1847);
or U836 (N_836,In_739,In_977);
nand U837 (N_837,In_2782,In_2877);
and U838 (N_838,In_585,In_1561);
nand U839 (N_839,In_1755,In_832);
nand U840 (N_840,In_2941,In_1533);
nor U841 (N_841,In_1183,In_2374);
and U842 (N_842,In_1913,In_1506);
nand U843 (N_843,In_509,In_1075);
nor U844 (N_844,In_2035,In_1222);
or U845 (N_845,In_1523,In_2081);
nand U846 (N_846,In_1311,In_42);
and U847 (N_847,In_69,In_1937);
nand U848 (N_848,In_188,In_2980);
or U849 (N_849,In_1399,In_163);
nand U850 (N_850,In_2947,In_2359);
xor U851 (N_851,In_189,In_463);
nor U852 (N_852,In_1080,In_1939);
nor U853 (N_853,In_2589,In_526);
xnor U854 (N_854,In_2195,In_2595);
xor U855 (N_855,In_426,In_2478);
nor U856 (N_856,In_2380,In_1638);
nand U857 (N_857,In_2243,In_1282);
xor U858 (N_858,In_44,In_1034);
and U859 (N_859,In_190,In_124);
and U860 (N_860,In_714,In_1901);
nand U861 (N_861,In_2233,In_1453);
nand U862 (N_862,In_373,In_90);
nand U863 (N_863,In_655,In_108);
and U864 (N_864,In_1206,In_1120);
nor U865 (N_865,In_2681,In_1846);
nor U866 (N_866,In_2481,In_1317);
nor U867 (N_867,In_1694,In_2824);
and U868 (N_868,In_2637,In_990);
and U869 (N_869,In_39,In_2984);
or U870 (N_870,In_398,In_2337);
and U871 (N_871,In_991,In_2089);
nand U872 (N_872,In_1730,In_2482);
nand U873 (N_873,In_2336,In_504);
nand U874 (N_874,In_839,In_2285);
or U875 (N_875,In_121,In_1144);
or U876 (N_876,In_602,In_528);
nor U877 (N_877,In_2235,In_2244);
and U878 (N_878,In_2953,In_1191);
nand U879 (N_879,In_1728,In_1963);
or U880 (N_880,In_2304,In_434);
or U881 (N_881,In_2651,In_1151);
nand U882 (N_882,In_1013,In_764);
nand U883 (N_883,In_267,In_2140);
nand U884 (N_884,In_1817,In_2392);
nand U885 (N_885,In_1772,In_473);
nor U886 (N_886,In_315,In_2181);
or U887 (N_887,In_2726,In_382);
or U888 (N_888,In_2249,In_1554);
and U889 (N_889,In_1131,In_968);
nand U890 (N_890,In_2068,In_1917);
nor U891 (N_891,In_2709,In_141);
nand U892 (N_892,In_2264,In_1379);
or U893 (N_893,In_2100,In_2529);
or U894 (N_894,In_875,In_379);
nand U895 (N_895,In_170,In_1163);
or U896 (N_896,In_2434,In_2696);
or U897 (N_897,In_529,In_37);
or U898 (N_898,In_1,In_1696);
or U899 (N_899,In_2986,In_377);
and U900 (N_900,In_712,In_478);
or U901 (N_901,In_582,In_2258);
nor U902 (N_902,In_1230,In_2803);
and U903 (N_903,In_2939,In_850);
and U904 (N_904,In_2659,In_1711);
or U905 (N_905,In_1043,In_589);
nand U906 (N_906,In_150,In_1249);
or U907 (N_907,In_1497,In_1777);
and U908 (N_908,In_1484,In_2937);
xnor U909 (N_909,In_1212,In_185);
xor U910 (N_910,In_736,In_1727);
xor U911 (N_911,In_1380,In_620);
nor U912 (N_912,In_393,In_2921);
nor U913 (N_913,In_2648,In_2671);
and U914 (N_914,In_2609,In_300);
nor U915 (N_915,In_277,In_415);
nand U916 (N_916,In_2203,In_2790);
or U917 (N_917,In_1135,In_1256);
or U918 (N_918,In_408,In_1815);
nor U919 (N_919,In_2669,In_1591);
nand U920 (N_920,In_817,In_1906);
or U921 (N_921,In_339,In_2020);
or U922 (N_922,In_1779,In_1016);
xor U923 (N_923,In_351,In_958);
nand U924 (N_924,In_2186,In_298);
and U925 (N_925,In_1722,In_2437);
nor U926 (N_926,In_389,In_586);
nor U927 (N_927,In_2069,In_1806);
and U928 (N_928,In_474,In_1959);
nand U929 (N_929,In_76,In_1293);
or U930 (N_930,In_2487,In_1238);
nor U931 (N_931,In_669,In_2364);
and U932 (N_932,In_2312,In_1509);
xnor U933 (N_933,In_950,In_2333);
nor U934 (N_934,In_1375,In_1324);
xor U935 (N_935,In_1036,In_1652);
nor U936 (N_936,In_1866,In_2218);
xnor U937 (N_937,In_457,In_1878);
and U938 (N_938,In_1658,In_2041);
nor U939 (N_939,In_1699,In_2381);
nand U940 (N_940,In_2447,In_10);
xor U941 (N_941,In_317,In_2751);
or U942 (N_942,In_2206,In_1522);
xor U943 (N_943,In_2422,In_1567);
or U944 (N_944,In_1129,In_384);
nand U945 (N_945,In_1461,In_149);
nand U946 (N_946,In_64,In_2119);
and U947 (N_947,In_800,In_995);
or U948 (N_948,In_1287,In_1368);
or U949 (N_949,In_2847,In_1545);
xor U950 (N_950,In_1098,In_285);
or U951 (N_951,In_948,In_1224);
or U952 (N_952,In_1955,In_1352);
nor U953 (N_953,In_2957,In_1479);
and U954 (N_954,In_49,In_1032);
or U955 (N_955,In_1803,In_406);
nand U956 (N_956,In_2368,In_1475);
or U957 (N_957,In_166,In_559);
nor U958 (N_958,In_155,In_1592);
nor U959 (N_959,In_2739,In_2134);
and U960 (N_960,In_880,In_956);
and U961 (N_961,In_70,In_919);
or U962 (N_962,In_2930,In_1934);
nand U963 (N_963,In_2103,In_2345);
nand U964 (N_964,In_2174,In_2617);
and U965 (N_965,In_2413,In_2841);
or U966 (N_966,In_2544,In_563);
xnor U967 (N_967,In_1950,In_2148);
and U968 (N_968,In_1314,In_1796);
and U969 (N_969,In_1213,In_779);
nand U970 (N_970,In_1365,In_2000);
or U971 (N_971,In_1202,In_1729);
or U972 (N_972,In_1033,In_2443);
nor U973 (N_973,In_695,In_1681);
nor U974 (N_974,In_1271,In_770);
and U975 (N_975,In_1787,In_612);
nand U976 (N_976,In_264,In_214);
xor U977 (N_977,In_1519,In_2007);
xnor U978 (N_978,In_609,In_2474);
nand U979 (N_979,In_1961,In_2224);
xor U980 (N_980,In_816,In_1589);
nor U981 (N_981,In_2082,In_2808);
or U982 (N_982,In_238,In_2115);
and U983 (N_983,In_2718,In_659);
nor U984 (N_984,In_1130,In_2693);
and U985 (N_985,In_2932,In_299);
nand U986 (N_986,In_1647,In_1391);
nor U987 (N_987,In_294,In_2719);
nor U988 (N_988,In_1195,In_1134);
nor U989 (N_989,In_83,In_1986);
and U990 (N_990,In_711,In_1744);
xor U991 (N_991,In_2971,In_56);
or U992 (N_992,In_1559,In_2293);
or U993 (N_993,In_1837,In_1290);
nor U994 (N_994,In_88,In_443);
or U995 (N_995,In_2401,In_225);
xnor U996 (N_996,In_2147,In_1465);
and U997 (N_997,In_2631,In_552);
nand U998 (N_998,In_1957,In_181);
nor U999 (N_999,In_1150,In_1009);
or U1000 (N_1000,In_2764,In_1404);
or U1001 (N_1001,In_2745,In_642);
nor U1002 (N_1002,In_751,In_1406);
or U1003 (N_1003,In_1283,In_2948);
and U1004 (N_1004,In_811,In_147);
nor U1005 (N_1005,In_2040,In_2484);
and U1006 (N_1006,In_2251,In_1590);
nor U1007 (N_1007,In_2846,In_1051);
and U1008 (N_1008,In_1644,In_2842);
nor U1009 (N_1009,In_1462,In_2611);
nand U1010 (N_1010,In_345,In_890);
and U1011 (N_1011,In_1600,In_1295);
or U1012 (N_1012,In_367,In_394);
nand U1013 (N_1013,In_813,In_1491);
nand U1014 (N_1014,In_1629,In_2869);
or U1015 (N_1015,In_2361,In_332);
or U1016 (N_1016,In_960,In_2036);
xor U1017 (N_1017,In_2079,In_2356);
xor U1018 (N_1018,In_2191,In_535);
and U1019 (N_1019,In_2712,In_735);
nor U1020 (N_1020,In_1157,In_2282);
nor U1021 (N_1021,In_2658,In_1011);
nand U1022 (N_1022,In_2014,In_1940);
or U1023 (N_1023,In_1345,In_996);
xnor U1024 (N_1024,In_481,In_362);
or U1025 (N_1025,In_936,In_689);
nor U1026 (N_1026,In_1972,In_2586);
nand U1027 (N_1027,In_2309,In_617);
or U1028 (N_1028,In_788,In_774);
or U1029 (N_1029,In_2504,In_690);
or U1030 (N_1030,In_1501,In_2126);
nand U1031 (N_1031,In_2455,In_2144);
or U1032 (N_1032,In_2818,In_541);
nand U1033 (N_1033,In_452,In_2551);
nor U1034 (N_1034,In_969,In_1048);
and U1035 (N_1035,In_1285,In_1443);
nand U1036 (N_1036,In_1893,In_1094);
or U1037 (N_1037,In_803,In_386);
xnor U1038 (N_1038,In_447,In_2110);
and U1039 (N_1039,In_143,In_2090);
nand U1040 (N_1040,In_2170,In_2271);
and U1041 (N_1041,In_1944,In_2855);
and U1042 (N_1042,In_26,In_2692);
nand U1043 (N_1043,In_2468,In_2584);
nor U1044 (N_1044,In_634,In_2540);
and U1045 (N_1045,In_492,In_2666);
or U1046 (N_1046,In_2444,In_272);
nor U1047 (N_1047,In_835,In_717);
nor U1048 (N_1048,In_2129,In_639);
and U1049 (N_1049,In_212,In_109);
nand U1050 (N_1050,In_1273,In_1518);
xnor U1051 (N_1051,In_753,In_1233);
or U1052 (N_1052,In_1431,In_286);
or U1053 (N_1053,In_2252,In_2663);
nor U1054 (N_1054,In_1741,In_2897);
nand U1055 (N_1055,In_1543,In_531);
nand U1056 (N_1056,In_1987,In_2295);
nor U1057 (N_1057,In_1759,In_1857);
and U1058 (N_1058,In_2985,In_1544);
and U1059 (N_1059,In_1005,In_1883);
and U1060 (N_1060,In_2541,In_2187);
and U1061 (N_1061,In_1517,In_2679);
nand U1062 (N_1062,In_952,In_383);
and U1063 (N_1063,In_1764,In_1861);
or U1064 (N_1064,In_1541,In_1809);
nand U1065 (N_1065,In_1928,In_2515);
xor U1066 (N_1066,In_1641,In_2775);
or U1067 (N_1067,In_74,In_2768);
nor U1068 (N_1068,In_2833,In_1894);
or U1069 (N_1069,In_2330,In_2049);
nor U1070 (N_1070,In_1771,In_2944);
and U1071 (N_1071,In_614,In_381);
xnor U1072 (N_1072,In_2909,In_2281);
or U1073 (N_1073,In_532,In_1425);
nor U1074 (N_1074,In_2053,In_1606);
or U1075 (N_1075,In_911,In_2390);
or U1076 (N_1076,In_1920,In_1839);
nand U1077 (N_1077,In_2526,In_601);
nand U1078 (N_1078,In_1805,In_793);
and U1079 (N_1079,In_1565,In_1909);
nand U1080 (N_1080,In_1070,In_2045);
and U1081 (N_1081,In_893,In_2618);
nand U1082 (N_1082,In_316,In_2057);
and U1083 (N_1083,In_1164,In_1474);
nand U1084 (N_1084,In_41,In_333);
and U1085 (N_1085,In_252,In_2722);
nor U1086 (N_1086,In_1822,In_59);
xnor U1087 (N_1087,In_1968,In_242);
and U1088 (N_1088,In_851,In_1079);
or U1089 (N_1089,In_2501,In_2816);
or U1090 (N_1090,In_1196,In_51);
or U1091 (N_1091,In_234,In_2849);
or U1092 (N_1092,In_497,In_2597);
and U1093 (N_1093,In_1097,In_247);
nor U1094 (N_1094,In_67,In_291);
nor U1095 (N_1095,In_1562,In_1990);
or U1096 (N_1096,In_1507,In_518);
nor U1097 (N_1097,In_900,In_2080);
or U1098 (N_1098,In_1793,In_2272);
and U1099 (N_1099,In_1613,In_230);
and U1100 (N_1100,In_2787,In_1608);
or U1101 (N_1101,In_997,In_558);
and U1102 (N_1102,In_670,In_1720);
nand U1103 (N_1103,In_2117,In_2630);
or U1104 (N_1104,In_2101,In_448);
and U1105 (N_1105,In_1935,In_2156);
nor U1106 (N_1106,In_923,In_130);
and U1107 (N_1107,In_2212,In_2261);
nor U1108 (N_1108,In_350,In_1758);
or U1109 (N_1109,In_2978,In_1712);
or U1110 (N_1110,In_115,In_1268);
or U1111 (N_1111,In_1991,In_1813);
nand U1112 (N_1112,In_0,In_1844);
or U1113 (N_1113,In_2546,In_2850);
or U1114 (N_1114,In_388,In_513);
nand U1115 (N_1115,In_397,In_1394);
nor U1116 (N_1116,In_289,In_2037);
nor U1117 (N_1117,In_1786,In_2375);
or U1118 (N_1118,In_2094,In_1672);
and U1119 (N_1119,In_1785,In_158);
and U1120 (N_1120,In_1450,In_2834);
nor U1121 (N_1121,In_1911,In_1216);
and U1122 (N_1122,In_295,In_268);
nand U1123 (N_1123,In_301,In_193);
nor U1124 (N_1124,In_732,In_1413);
xor U1125 (N_1125,In_1056,In_943);
and U1126 (N_1126,In_136,In_1581);
and U1127 (N_1127,In_9,In_216);
or U1128 (N_1128,In_2626,In_2887);
or U1129 (N_1129,In_2888,In_2956);
nor U1130 (N_1130,In_414,In_1423);
nor U1131 (N_1131,In_2344,In_81);
nand U1132 (N_1132,In_2024,In_963);
xor U1133 (N_1133,In_856,In_2322);
or U1134 (N_1134,In_2205,In_929);
nor U1135 (N_1135,In_2063,In_246);
nand U1136 (N_1136,In_971,In_1473);
or U1137 (N_1137,In_1499,In_1548);
nand U1138 (N_1138,In_777,In_2731);
nand U1139 (N_1139,In_6,In_2845);
nand U1140 (N_1140,In_1762,In_2512);
and U1141 (N_1141,In_2141,In_2701);
nand U1142 (N_1142,In_1899,In_2221);
or U1143 (N_1143,In_1284,In_328);
nor U1144 (N_1144,In_750,In_416);
nand U1145 (N_1145,In_853,In_1859);
nor U1146 (N_1146,In_1467,In_1579);
nor U1147 (N_1147,In_2752,In_1158);
nand U1148 (N_1148,In_2026,In_2804);
or U1149 (N_1149,In_2483,In_71);
nand U1150 (N_1150,In_127,In_1978);
and U1151 (N_1151,In_2911,In_561);
and U1152 (N_1152,In_1789,In_302);
xor U1153 (N_1153,In_772,In_1770);
or U1154 (N_1154,In_2573,In_1181);
or U1155 (N_1155,In_343,In_490);
nor U1156 (N_1156,In_2798,In_508);
nor U1157 (N_1157,In_2981,In_1747);
nand U1158 (N_1158,In_613,In_2072);
or U1159 (N_1159,In_43,In_2065);
and U1160 (N_1160,In_498,In_2982);
and U1161 (N_1161,In_1812,In_915);
xnor U1162 (N_1162,In_2275,In_1272);
nand U1163 (N_1163,In_1992,In_1521);
nor U1164 (N_1164,In_2253,In_501);
or U1165 (N_1165,In_2951,In_2797);
and U1166 (N_1166,In_22,In_1636);
nor U1167 (N_1167,In_972,In_1089);
xor U1168 (N_1168,In_355,In_2664);
or U1169 (N_1169,In_1784,In_2927);
and U1170 (N_1170,In_2429,In_2735);
nand U1171 (N_1171,In_1563,In_1845);
and U1172 (N_1172,In_2860,In_686);
nand U1173 (N_1173,In_1876,In_2612);
nor U1174 (N_1174,In_2706,In_364);
or U1175 (N_1175,In_1675,In_1840);
nor U1176 (N_1176,In_2006,In_1107);
xor U1177 (N_1177,In_740,In_1240);
nor U1178 (N_1178,In_744,In_405);
and U1179 (N_1179,In_836,In_588);
or U1180 (N_1180,In_32,In_323);
nor U1181 (N_1181,In_1788,In_410);
or U1182 (N_1182,In_1888,In_931);
and U1183 (N_1183,In_554,In_402);
nand U1184 (N_1184,In_2464,In_259);
nand U1185 (N_1185,In_1657,In_2310);
nor U1186 (N_1186,In_2303,In_368);
and U1187 (N_1187,In_1148,In_2738);
nand U1188 (N_1188,In_945,In_1814);
nor U1189 (N_1189,In_1903,In_1440);
and U1190 (N_1190,In_994,In_666);
or U1191 (N_1191,In_1743,In_287);
nand U1192 (N_1192,In_576,In_1086);
and U1193 (N_1193,In_1677,In_2590);
or U1194 (N_1194,In_1502,In_2067);
nor U1195 (N_1195,In_818,In_2450);
or U1196 (N_1196,In_2071,In_2451);
nor U1197 (N_1197,In_1656,In_2703);
and U1198 (N_1198,In_24,In_1798);
nand U1199 (N_1199,In_1247,In_125);
nand U1200 (N_1200,In_869,In_878);
and U1201 (N_1201,In_2204,In_2603);
nor U1202 (N_1202,In_375,In_142);
nor U1203 (N_1203,In_570,In_2533);
nor U1204 (N_1204,In_1824,In_922);
nor U1205 (N_1205,In_1663,In_2881);
and U1206 (N_1206,In_2684,In_2377);
or U1207 (N_1207,In_1398,In_2498);
or U1208 (N_1208,In_358,In_2600);
or U1209 (N_1209,In_1031,In_2817);
nor U1210 (N_1210,In_593,In_89);
and U1211 (N_1211,In_539,In_2771);
nor U1212 (N_1212,In_1498,In_2672);
nor U1213 (N_1213,In_2688,In_2379);
nor U1214 (N_1214,In_2417,In_486);
nand U1215 (N_1215,In_2213,In_897);
nor U1216 (N_1216,In_514,In_46);
nor U1217 (N_1217,In_1482,In_258);
or U1218 (N_1218,In_1997,In_476);
nand U1219 (N_1219,In_1308,In_1242);
and U1220 (N_1220,In_729,In_1073);
nand U1221 (N_1221,In_475,In_105);
nor U1222 (N_1222,In_57,In_1251);
or U1223 (N_1223,In_2479,In_1363);
or U1224 (N_1224,In_1520,In_1804);
and U1225 (N_1225,In_211,In_1576);
nand U1226 (N_1226,In_812,In_2582);
or U1227 (N_1227,In_2154,In_2965);
and U1228 (N_1228,In_1401,In_2907);
and U1229 (N_1229,In_1703,In_1612);
and U1230 (N_1230,In_2707,In_2690);
and U1231 (N_1231,In_780,In_1464);
xor U1232 (N_1232,In_679,In_630);
nor U1233 (N_1233,In_2458,In_1280);
nand U1234 (N_1234,In_2135,In_975);
xor U1235 (N_1235,In_2854,In_34);
and U1236 (N_1236,In_1122,In_1597);
and U1237 (N_1237,In_366,In_1480);
and U1238 (N_1238,In_1101,In_1141);
or U1239 (N_1239,In_1540,In_2179);
or U1240 (N_1240,In_2801,In_2463);
xnor U1241 (N_1241,In_1697,In_320);
and U1242 (N_1242,In_2328,In_1969);
nor U1243 (N_1243,In_2242,In_2165);
or U1244 (N_1244,In_906,In_1103);
or U1245 (N_1245,In_2777,In_1914);
nor U1246 (N_1246,In_694,In_2628);
nand U1247 (N_1247,In_2441,In_1172);
or U1248 (N_1248,In_2691,In_2232);
nor U1249 (N_1249,In_1485,In_2456);
nand U1250 (N_1250,In_981,In_2554);
nor U1251 (N_1251,In_727,In_725);
and U1252 (N_1252,In_2555,In_2259);
nor U1253 (N_1253,In_2961,In_21);
xnor U1254 (N_1254,In_66,In_180);
nand U1255 (N_1255,In_700,In_2518);
and U1256 (N_1256,In_1925,In_2852);
nor U1257 (N_1257,In_1430,In_265);
xnor U1258 (N_1258,In_2188,In_1014);
and U1259 (N_1259,In_1105,In_282);
nand U1260 (N_1260,In_1420,In_660);
nand U1261 (N_1261,In_2139,In_2585);
nand U1262 (N_1262,In_2495,In_1112);
nand U1263 (N_1263,In_941,In_2142);
or U1264 (N_1264,In_645,In_1829);
nor U1265 (N_1265,In_2675,In_2895);
nand U1266 (N_1266,In_1003,In_1155);
and U1267 (N_1267,In_1109,In_2423);
and U1268 (N_1268,In_2896,In_1110);
nor U1269 (N_1269,In_111,In_1505);
or U1270 (N_1270,In_2245,In_1994);
xor U1271 (N_1271,In_1477,In_2643);
and U1272 (N_1272,In_2918,In_2505);
and U1273 (N_1273,In_2297,In_1028);
nor U1274 (N_1274,In_1305,In_1093);
nand U1275 (N_1275,In_1451,In_1335);
nand U1276 (N_1276,In_1618,In_2054);
nand U1277 (N_1277,In_892,In_499);
nand U1278 (N_1278,In_2908,In_164);
xor U1279 (N_1279,In_556,In_754);
nand U1280 (N_1280,In_2070,In_1410);
and U1281 (N_1281,In_219,In_2075);
or U1282 (N_1282,In_515,In_174);
nand U1283 (N_1283,In_2039,In_1146);
or U1284 (N_1284,In_1139,In_2524);
nor U1285 (N_1285,In_1127,In_1397);
and U1286 (N_1286,In_2604,In_2676);
and U1287 (N_1287,In_1372,In_2991);
nand U1288 (N_1288,In_1577,In_1095);
or U1289 (N_1289,In_2641,In_1286);
nor U1290 (N_1290,In_646,In_1570);
nor U1291 (N_1291,In_494,In_1801);
and U1292 (N_1292,In_256,In_186);
and U1293 (N_1293,In_1378,In_548);
and U1294 (N_1294,In_329,In_707);
nor U1295 (N_1295,In_2198,In_1714);
or U1296 (N_1296,In_2598,In_728);
nor U1297 (N_1297,In_2958,In_1414);
or U1298 (N_1298,In_1898,In_984);
or U1299 (N_1299,In_1572,In_538);
nor U1300 (N_1300,In_826,In_2880);
and U1301 (N_1301,In_1228,In_95);
nor U1302 (N_1302,In_786,In_2284);
and U1303 (N_1303,In_224,In_723);
nand U1304 (N_1304,In_50,In_1045);
and U1305 (N_1305,In_28,In_62);
nor U1306 (N_1306,In_1173,In_2759);
xor U1307 (N_1307,In_2520,In_1117);
or U1308 (N_1308,In_2276,In_2400);
nand U1309 (N_1309,In_2397,In_18);
and U1310 (N_1310,In_2767,In_1102);
nor U1311 (N_1311,In_94,In_643);
nor U1312 (N_1312,In_1347,In_726);
nor U1313 (N_1313,In_705,In_1598);
nand U1314 (N_1314,In_404,In_280);
or U1315 (N_1315,In_2556,In_1905);
or U1316 (N_1316,In_250,In_503);
nand U1317 (N_1317,In_2581,In_1531);
nor U1318 (N_1318,In_2003,In_2548);
or U1319 (N_1319,In_1745,In_1713);
nor U1320 (N_1320,In_571,In_199);
or U1321 (N_1321,In_704,In_1111);
xor U1322 (N_1322,In_794,In_907);
nand U1323 (N_1323,In_1321,In_2240);
or U1324 (N_1324,In_624,In_611);
xor U1325 (N_1325,In_841,In_1452);
nor U1326 (N_1326,In_1001,In_162);
or U1327 (N_1327,In_859,In_610);
and U1328 (N_1328,In_1184,In_1396);
nor U1329 (N_1329,In_1128,In_1054);
or U1330 (N_1330,In_1024,In_809);
and U1331 (N_1331,In_1926,In_1733);
nor U1332 (N_1332,In_708,In_608);
nand U1333 (N_1333,In_1422,In_1017);
and U1334 (N_1334,In_312,In_861);
nor U1335 (N_1335,In_1586,In_2226);
nor U1336 (N_1336,In_1595,In_1356);
and U1337 (N_1337,In_615,In_369);
or U1338 (N_1338,In_2169,In_2655);
nand U1339 (N_1339,In_534,In_1942);
or U1340 (N_1340,In_1734,In_760);
or U1341 (N_1341,In_701,In_1264);
or U1342 (N_1342,In_1973,In_396);
or U1343 (N_1343,In_2702,In_1438);
or U1344 (N_1344,In_2838,In_2863);
nor U1345 (N_1345,In_1724,In_2802);
nor U1346 (N_1346,In_483,In_244);
and U1347 (N_1347,In_1288,In_652);
or U1348 (N_1348,In_1030,In_1255);
nand U1349 (N_1349,In_962,In_584);
and U1350 (N_1350,In_1792,In_2940);
and U1351 (N_1351,In_2525,In_1756);
or U1352 (N_1352,In_2492,In_1890);
nor U1353 (N_1353,In_2550,In_1332);
nand U1354 (N_1354,In_1178,In_886);
and U1355 (N_1355,In_2949,In_805);
xnor U1356 (N_1356,In_1855,In_2830);
nand U1357 (N_1357,In_1052,In_172);
xor U1358 (N_1358,In_2130,In_1918);
and U1359 (N_1359,In_1405,In_1187);
xnor U1360 (N_1360,In_985,In_1970);
and U1361 (N_1361,In_337,In_1587);
nor U1362 (N_1362,In_2287,In_2788);
and U1363 (N_1363,In_1087,In_1424);
and U1364 (N_1364,In_591,In_45);
or U1365 (N_1365,In_5,In_2017);
nand U1366 (N_1366,In_2022,In_1357);
or U1367 (N_1367,In_1358,In_2305);
nand U1368 (N_1368,In_2290,In_2116);
or U1369 (N_1369,In_1737,In_2372);
nor U1370 (N_1370,In_2216,In_2236);
nor U1371 (N_1371,In_2120,In_2163);
or U1372 (N_1372,In_1964,In_152);
or U1373 (N_1373,In_635,In_2661);
or U1374 (N_1374,In_808,In_1573);
nand U1375 (N_1375,In_2321,In_1526);
nor U1376 (N_1376,In_2724,In_2886);
and U1377 (N_1377,In_2926,In_309);
and U1378 (N_1378,In_1820,In_2517);
or U1379 (N_1379,In_1218,In_2812);
and U1380 (N_1380,In_2208,In_1659);
or U1381 (N_1381,In_1046,In_48);
nand U1382 (N_1382,In_1664,In_442);
nor U1383 (N_1383,In_628,In_2993);
or U1384 (N_1384,In_1486,In_153);
xor U1385 (N_1385,In_678,In_2700);
and U1386 (N_1386,In_568,In_1004);
nor U1387 (N_1387,In_1115,In_2509);
xor U1388 (N_1388,In_1038,In_769);
xnor U1389 (N_1389,In_2043,In_2227);
nor U1390 (N_1390,In_129,In_1684);
nor U1391 (N_1391,In_1339,In_1836);
or U1392 (N_1392,In_1875,In_2835);
or U1393 (N_1393,In_1853,In_137);
nor U1394 (N_1394,In_409,In_184);
or U1395 (N_1395,In_846,In_2161);
nand U1396 (N_1396,In_357,In_1633);
or U1397 (N_1397,In_633,In_1210);
and U1398 (N_1398,In_451,In_2809);
and U1399 (N_1399,In_2315,In_2308);
and U1400 (N_1400,In_1850,In_344);
and U1401 (N_1401,In_1662,In_2025);
nor U1402 (N_1402,In_1529,In_2906);
nand U1403 (N_1403,In_1751,In_1235);
and U1404 (N_1404,In_16,In_521);
nand U1405 (N_1405,In_1162,In_213);
nand U1406 (N_1406,In_2831,In_1669);
and U1407 (N_1407,In_1616,In_2370);
or U1408 (N_1408,In_1458,In_621);
and U1409 (N_1409,In_1136,In_1248);
and U1410 (N_1410,In_1020,In_2228);
xor U1411 (N_1411,In_319,In_60);
xor U1412 (N_1412,In_97,In_1199);
nor U1413 (N_1413,In_75,In_1585);
nand U1414 (N_1414,In_1252,In_2889);
and U1415 (N_1415,In_445,In_752);
or U1416 (N_1416,In_2184,In_709);
or U1417 (N_1417,In_641,In_2480);
nand U1418 (N_1418,In_2733,In_1774);
nor U1419 (N_1419,In_419,In_681);
or U1420 (N_1420,In_743,In_207);
nor U1421 (N_1421,In_1604,In_516);
nor U1422 (N_1422,In_1433,In_2319);
xnor U1423 (N_1423,In_1318,In_1319);
nor U1424 (N_1424,In_1884,In_598);
and U1425 (N_1425,In_1602,In_1263);
and U1426 (N_1426,In_2439,In_1981);
nor U1427 (N_1427,In_1067,In_25);
nor U1428 (N_1428,In_2267,In_2899);
nand U1429 (N_1429,In_2557,In_2388);
nand U1430 (N_1430,In_1500,In_2786);
and U1431 (N_1431,In_2239,In_1980);
or U1432 (N_1432,In_2936,In_682);
or U1433 (N_1433,In_1623,In_1749);
nor U1434 (N_1434,In_1808,In_1161);
or U1435 (N_1435,In_1580,In_2001);
xor U1436 (N_1436,In_884,In_1943);
nand U1437 (N_1437,In_982,In_1553);
nand U1438 (N_1438,In_2485,In_2913);
or U1439 (N_1439,In_785,In_2780);
nor U1440 (N_1440,In_658,In_560);
nand U1441 (N_1441,In_2875,In_1403);
nand U1442 (N_1442,In_2340,In_1688);
or U1443 (N_1443,In_1415,In_2975);
nand U1444 (N_1444,In_1007,In_488);
or U1445 (N_1445,In_78,In_3);
and U1446 (N_1446,In_228,In_1954);
and U1447 (N_1447,In_1261,In_1626);
nand U1448 (N_1448,In_2576,In_2789);
nand U1449 (N_1449,In_1265,In_1833);
and U1450 (N_1450,In_2623,In_942);
or U1451 (N_1451,In_2074,In_625);
and U1452 (N_1452,In_1197,In_165);
nor U1453 (N_1453,In_2420,In_1891);
and U1454 (N_1454,In_683,In_126);
or U1455 (N_1455,In_1065,In_1835);
nor U1456 (N_1456,In_2892,In_849);
and U1457 (N_1457,In_2136,In_324);
and U1458 (N_1458,In_2111,In_2373);
or U1459 (N_1459,In_2064,In_72);
nand U1460 (N_1460,In_2795,In_1250);
and U1461 (N_1461,In_989,In_1539);
and U1462 (N_1462,In_85,In_1262);
nor U1463 (N_1463,In_653,In_1746);
or U1464 (N_1464,In_2995,In_829);
or U1465 (N_1465,In_2662,In_313);
or U1466 (N_1466,In_203,In_1159);
or U1467 (N_1467,In_1241,In_352);
and U1468 (N_1468,In_540,In_2843);
nor U1469 (N_1469,In_1281,In_2488);
xnor U1470 (N_1470,In_765,In_1165);
nand U1471 (N_1471,In_2131,In_1092);
or U1472 (N_1472,In_2695,In_2299);
or U1473 (N_1473,In_1091,In_2619);
or U1474 (N_1474,In_1231,In_8);
and U1475 (N_1475,In_1956,In_567);
nand U1476 (N_1476,In_2230,In_2705);
or U1477 (N_1477,In_2404,In_482);
or U1478 (N_1478,In_263,In_1877);
or U1479 (N_1479,In_248,In_2826);
or U1480 (N_1480,In_1483,In_2772);
nand U1481 (N_1481,In_2660,In_2578);
or U1482 (N_1482,In_2023,In_2890);
xor U1483 (N_1483,In_1125,In_1740);
or U1484 (N_1484,In_1799,In_2620);
nand U1485 (N_1485,In_933,In_2746);
and U1486 (N_1486,In_257,In_183);
and U1487 (N_1487,In_894,In_2273);
or U1488 (N_1488,In_1566,In_1654);
nand U1489 (N_1489,In_1760,In_2779);
and U1490 (N_1490,In_411,In_1328);
nand U1491 (N_1491,In_1686,In_2164);
nand U1492 (N_1492,In_1304,In_1327);
and U1493 (N_1493,In_2296,In_218);
and U1494 (N_1494,In_1258,In_1113);
nor U1495 (N_1495,In_2765,In_2334);
or U1496 (N_1496,In_1071,In_40);
nand U1497 (N_1497,In_2286,In_1915);
and U1498 (N_1498,In_2168,In_980);
xor U1499 (N_1499,In_1412,In_2059);
xnor U1500 (N_1500,In_179,In_2879);
nor U1501 (N_1501,In_861,In_2108);
or U1502 (N_1502,In_1692,In_359);
or U1503 (N_1503,In_234,In_1998);
or U1504 (N_1504,In_484,In_612);
xnor U1505 (N_1505,In_621,In_733);
nor U1506 (N_1506,In_2847,In_1844);
nor U1507 (N_1507,In_1252,In_826);
nand U1508 (N_1508,In_1063,In_564);
or U1509 (N_1509,In_1934,In_1673);
and U1510 (N_1510,In_2202,In_2696);
or U1511 (N_1511,In_1679,In_786);
nand U1512 (N_1512,In_1240,In_2313);
nor U1513 (N_1513,In_2451,In_2588);
nor U1514 (N_1514,In_106,In_1117);
nand U1515 (N_1515,In_1474,In_986);
xnor U1516 (N_1516,In_2900,In_1754);
or U1517 (N_1517,In_2738,In_1962);
or U1518 (N_1518,In_1566,In_1353);
xnor U1519 (N_1519,In_2903,In_434);
nor U1520 (N_1520,In_2046,In_2588);
nand U1521 (N_1521,In_2112,In_2517);
or U1522 (N_1522,In_1634,In_696);
and U1523 (N_1523,In_2331,In_360);
nand U1524 (N_1524,In_470,In_2655);
xnor U1525 (N_1525,In_2278,In_2518);
and U1526 (N_1526,In_944,In_2837);
nor U1527 (N_1527,In_40,In_2239);
nand U1528 (N_1528,In_747,In_1845);
nand U1529 (N_1529,In_1788,In_629);
nand U1530 (N_1530,In_352,In_1309);
nand U1531 (N_1531,In_196,In_1406);
xor U1532 (N_1532,In_327,In_1258);
and U1533 (N_1533,In_1889,In_2253);
xor U1534 (N_1534,In_1106,In_1411);
nor U1535 (N_1535,In_1732,In_2656);
and U1536 (N_1536,In_837,In_1892);
nand U1537 (N_1537,In_2921,In_101);
or U1538 (N_1538,In_873,In_2347);
and U1539 (N_1539,In_2840,In_1751);
and U1540 (N_1540,In_2532,In_717);
and U1541 (N_1541,In_2966,In_2448);
nand U1542 (N_1542,In_2264,In_1828);
xor U1543 (N_1543,In_901,In_2734);
or U1544 (N_1544,In_1448,In_1508);
or U1545 (N_1545,In_1896,In_2039);
and U1546 (N_1546,In_2483,In_951);
nand U1547 (N_1547,In_1710,In_1606);
nor U1548 (N_1548,In_56,In_318);
or U1549 (N_1549,In_2463,In_1509);
and U1550 (N_1550,In_515,In_845);
and U1551 (N_1551,In_167,In_2770);
and U1552 (N_1552,In_1747,In_2988);
nor U1553 (N_1553,In_1640,In_1960);
nor U1554 (N_1554,In_2175,In_1070);
nor U1555 (N_1555,In_2365,In_32);
nor U1556 (N_1556,In_1059,In_2685);
xor U1557 (N_1557,In_2153,In_1179);
or U1558 (N_1558,In_2578,In_34);
nand U1559 (N_1559,In_526,In_639);
or U1560 (N_1560,In_2903,In_2178);
and U1561 (N_1561,In_437,In_1891);
nand U1562 (N_1562,In_2950,In_1926);
nor U1563 (N_1563,In_2386,In_23);
nor U1564 (N_1564,In_1583,In_813);
nor U1565 (N_1565,In_984,In_1934);
nor U1566 (N_1566,In_1615,In_2292);
or U1567 (N_1567,In_253,In_2282);
nor U1568 (N_1568,In_146,In_2710);
nor U1569 (N_1569,In_1348,In_856);
nand U1570 (N_1570,In_54,In_2137);
nor U1571 (N_1571,In_848,In_2989);
or U1572 (N_1572,In_2618,In_680);
or U1573 (N_1573,In_1632,In_220);
nand U1574 (N_1574,In_1067,In_1246);
or U1575 (N_1575,In_955,In_1947);
nand U1576 (N_1576,In_2635,In_62);
nor U1577 (N_1577,In_482,In_2227);
nor U1578 (N_1578,In_1339,In_2705);
nand U1579 (N_1579,In_1736,In_2508);
or U1580 (N_1580,In_758,In_2487);
or U1581 (N_1581,In_2710,In_1321);
nor U1582 (N_1582,In_437,In_282);
and U1583 (N_1583,In_1442,In_1012);
and U1584 (N_1584,In_340,In_1740);
and U1585 (N_1585,In_45,In_1565);
nor U1586 (N_1586,In_1280,In_469);
nor U1587 (N_1587,In_1380,In_597);
nor U1588 (N_1588,In_2302,In_38);
and U1589 (N_1589,In_916,In_238);
and U1590 (N_1590,In_1655,In_2073);
and U1591 (N_1591,In_2033,In_2805);
and U1592 (N_1592,In_2049,In_2582);
and U1593 (N_1593,In_516,In_40);
or U1594 (N_1594,In_2504,In_420);
nor U1595 (N_1595,In_1155,In_172);
nand U1596 (N_1596,In_1601,In_498);
and U1597 (N_1597,In_2482,In_360);
nor U1598 (N_1598,In_706,In_273);
nand U1599 (N_1599,In_1449,In_2918);
or U1600 (N_1600,In_2998,In_2459);
or U1601 (N_1601,In_2814,In_681);
and U1602 (N_1602,In_216,In_187);
and U1603 (N_1603,In_1288,In_1810);
xor U1604 (N_1604,In_328,In_2623);
and U1605 (N_1605,In_930,In_354);
nand U1606 (N_1606,In_2997,In_2750);
nand U1607 (N_1607,In_942,In_1688);
nand U1608 (N_1608,In_2798,In_1374);
or U1609 (N_1609,In_1966,In_2406);
xor U1610 (N_1610,In_1752,In_2260);
and U1611 (N_1611,In_1915,In_2974);
xnor U1612 (N_1612,In_2932,In_2028);
nor U1613 (N_1613,In_2773,In_2202);
xnor U1614 (N_1614,In_1159,In_1272);
or U1615 (N_1615,In_704,In_2017);
and U1616 (N_1616,In_2941,In_1565);
or U1617 (N_1617,In_2595,In_2148);
nor U1618 (N_1618,In_67,In_2519);
nor U1619 (N_1619,In_174,In_632);
nor U1620 (N_1620,In_862,In_1905);
or U1621 (N_1621,In_1724,In_1691);
or U1622 (N_1622,In_1163,In_547);
nor U1623 (N_1623,In_2160,In_2431);
and U1624 (N_1624,In_2309,In_2567);
nor U1625 (N_1625,In_2797,In_507);
and U1626 (N_1626,In_818,In_2130);
nor U1627 (N_1627,In_2681,In_781);
and U1628 (N_1628,In_2799,In_1240);
nor U1629 (N_1629,In_599,In_1337);
and U1630 (N_1630,In_7,In_47);
or U1631 (N_1631,In_1691,In_941);
nand U1632 (N_1632,In_1430,In_1549);
nand U1633 (N_1633,In_2759,In_781);
and U1634 (N_1634,In_1545,In_2793);
or U1635 (N_1635,In_1317,In_2529);
or U1636 (N_1636,In_2610,In_2547);
and U1637 (N_1637,In_2503,In_1596);
nor U1638 (N_1638,In_732,In_585);
or U1639 (N_1639,In_2858,In_563);
xor U1640 (N_1640,In_1438,In_1871);
and U1641 (N_1641,In_34,In_842);
and U1642 (N_1642,In_442,In_1206);
or U1643 (N_1643,In_379,In_2183);
xnor U1644 (N_1644,In_1700,In_2158);
nor U1645 (N_1645,In_1450,In_724);
and U1646 (N_1646,In_479,In_2924);
nor U1647 (N_1647,In_1386,In_2462);
nor U1648 (N_1648,In_755,In_2457);
or U1649 (N_1649,In_530,In_1768);
nand U1650 (N_1650,In_1985,In_1789);
nand U1651 (N_1651,In_1124,In_2521);
or U1652 (N_1652,In_2656,In_1941);
and U1653 (N_1653,In_2424,In_1174);
nor U1654 (N_1654,In_1005,In_1252);
or U1655 (N_1655,In_801,In_2951);
and U1656 (N_1656,In_63,In_2901);
nor U1657 (N_1657,In_1096,In_2282);
nand U1658 (N_1658,In_2220,In_2771);
or U1659 (N_1659,In_263,In_1466);
and U1660 (N_1660,In_1509,In_2593);
or U1661 (N_1661,In_1946,In_1980);
xnor U1662 (N_1662,In_531,In_383);
xnor U1663 (N_1663,In_1780,In_2654);
and U1664 (N_1664,In_690,In_226);
or U1665 (N_1665,In_674,In_2811);
nor U1666 (N_1666,In_1841,In_707);
or U1667 (N_1667,In_2934,In_1022);
and U1668 (N_1668,In_766,In_1129);
nand U1669 (N_1669,In_1273,In_1543);
nor U1670 (N_1670,In_1016,In_617);
and U1671 (N_1671,In_1085,In_693);
nand U1672 (N_1672,In_881,In_518);
and U1673 (N_1673,In_657,In_171);
or U1674 (N_1674,In_406,In_2804);
or U1675 (N_1675,In_2645,In_142);
and U1676 (N_1676,In_1758,In_99);
nand U1677 (N_1677,In_2906,In_775);
nor U1678 (N_1678,In_1441,In_901);
or U1679 (N_1679,In_1277,In_1593);
or U1680 (N_1680,In_1123,In_353);
or U1681 (N_1681,In_1297,In_2002);
and U1682 (N_1682,In_618,In_1158);
xor U1683 (N_1683,In_2466,In_464);
or U1684 (N_1684,In_2038,In_2290);
nor U1685 (N_1685,In_1755,In_1925);
nand U1686 (N_1686,In_34,In_2556);
and U1687 (N_1687,In_2897,In_1653);
and U1688 (N_1688,In_954,In_2171);
and U1689 (N_1689,In_778,In_1196);
and U1690 (N_1690,In_1999,In_2932);
or U1691 (N_1691,In_592,In_2954);
nor U1692 (N_1692,In_1528,In_1733);
or U1693 (N_1693,In_1060,In_665);
or U1694 (N_1694,In_2358,In_2072);
xor U1695 (N_1695,In_350,In_1085);
and U1696 (N_1696,In_2463,In_1420);
or U1697 (N_1697,In_1892,In_67);
or U1698 (N_1698,In_67,In_1595);
and U1699 (N_1699,In_1701,In_1377);
nor U1700 (N_1700,In_1317,In_2646);
and U1701 (N_1701,In_1926,In_2463);
and U1702 (N_1702,In_50,In_1940);
nor U1703 (N_1703,In_2998,In_58);
xor U1704 (N_1704,In_889,In_1001);
nand U1705 (N_1705,In_2670,In_201);
nand U1706 (N_1706,In_663,In_2758);
or U1707 (N_1707,In_2918,In_602);
and U1708 (N_1708,In_1799,In_2200);
or U1709 (N_1709,In_2388,In_2304);
nor U1710 (N_1710,In_2213,In_1491);
and U1711 (N_1711,In_663,In_1328);
or U1712 (N_1712,In_858,In_2774);
xnor U1713 (N_1713,In_2068,In_823);
and U1714 (N_1714,In_188,In_1719);
or U1715 (N_1715,In_1651,In_1728);
nor U1716 (N_1716,In_1945,In_534);
or U1717 (N_1717,In_2412,In_48);
and U1718 (N_1718,In_2158,In_292);
nand U1719 (N_1719,In_1355,In_1060);
nand U1720 (N_1720,In_2090,In_1668);
nor U1721 (N_1721,In_2862,In_96);
and U1722 (N_1722,In_268,In_743);
xor U1723 (N_1723,In_709,In_157);
nor U1724 (N_1724,In_91,In_2497);
and U1725 (N_1725,In_76,In_46);
or U1726 (N_1726,In_1901,In_1905);
nor U1727 (N_1727,In_2475,In_1894);
and U1728 (N_1728,In_1420,In_748);
and U1729 (N_1729,In_1241,In_208);
or U1730 (N_1730,In_541,In_2788);
and U1731 (N_1731,In_2297,In_1647);
or U1732 (N_1732,In_185,In_1714);
or U1733 (N_1733,In_1670,In_2832);
xor U1734 (N_1734,In_996,In_2793);
or U1735 (N_1735,In_2000,In_662);
and U1736 (N_1736,In_617,In_2287);
or U1737 (N_1737,In_1585,In_2479);
xnor U1738 (N_1738,In_1951,In_2424);
xnor U1739 (N_1739,In_755,In_2315);
or U1740 (N_1740,In_2210,In_293);
xor U1741 (N_1741,In_1359,In_604);
or U1742 (N_1742,In_1430,In_1589);
nand U1743 (N_1743,In_506,In_2261);
or U1744 (N_1744,In_2063,In_2072);
nor U1745 (N_1745,In_2483,In_2980);
and U1746 (N_1746,In_2051,In_2756);
or U1747 (N_1747,In_2970,In_824);
xor U1748 (N_1748,In_857,In_2822);
nand U1749 (N_1749,In_1162,In_365);
nor U1750 (N_1750,In_2342,In_1512);
nand U1751 (N_1751,In_572,In_2078);
nand U1752 (N_1752,In_1826,In_1288);
and U1753 (N_1753,In_2660,In_821);
or U1754 (N_1754,In_1226,In_883);
nor U1755 (N_1755,In_459,In_1720);
and U1756 (N_1756,In_1137,In_1166);
nand U1757 (N_1757,In_1903,In_763);
nor U1758 (N_1758,In_2095,In_209);
or U1759 (N_1759,In_151,In_804);
or U1760 (N_1760,In_1201,In_1311);
nand U1761 (N_1761,In_1049,In_1197);
and U1762 (N_1762,In_2270,In_1755);
nand U1763 (N_1763,In_1500,In_2963);
nand U1764 (N_1764,In_2228,In_2148);
or U1765 (N_1765,In_1708,In_276);
xnor U1766 (N_1766,In_1866,In_680);
and U1767 (N_1767,In_818,In_1614);
or U1768 (N_1768,In_2350,In_103);
nand U1769 (N_1769,In_1620,In_946);
and U1770 (N_1770,In_1839,In_2615);
and U1771 (N_1771,In_712,In_964);
nand U1772 (N_1772,In_2089,In_8);
xor U1773 (N_1773,In_2868,In_978);
and U1774 (N_1774,In_2690,In_2033);
and U1775 (N_1775,In_2974,In_2002);
nand U1776 (N_1776,In_1065,In_1274);
and U1777 (N_1777,In_543,In_838);
or U1778 (N_1778,In_2624,In_2560);
and U1779 (N_1779,In_64,In_1805);
or U1780 (N_1780,In_387,In_2254);
nand U1781 (N_1781,In_2646,In_1666);
nand U1782 (N_1782,In_683,In_1886);
nand U1783 (N_1783,In_2568,In_973);
and U1784 (N_1784,In_2886,In_2191);
and U1785 (N_1785,In_417,In_666);
nor U1786 (N_1786,In_1599,In_1407);
nor U1787 (N_1787,In_1396,In_1179);
and U1788 (N_1788,In_2427,In_2333);
nand U1789 (N_1789,In_2707,In_2620);
nor U1790 (N_1790,In_2866,In_2355);
or U1791 (N_1791,In_906,In_2450);
nand U1792 (N_1792,In_1653,In_460);
or U1793 (N_1793,In_2378,In_2121);
nor U1794 (N_1794,In_909,In_1353);
and U1795 (N_1795,In_474,In_1727);
xor U1796 (N_1796,In_1951,In_2248);
nor U1797 (N_1797,In_893,In_803);
nand U1798 (N_1798,In_1434,In_46);
nand U1799 (N_1799,In_2861,In_2054);
nor U1800 (N_1800,In_2593,In_1985);
and U1801 (N_1801,In_2943,In_2933);
or U1802 (N_1802,In_1090,In_1996);
or U1803 (N_1803,In_2342,In_226);
nand U1804 (N_1804,In_2913,In_1682);
nand U1805 (N_1805,In_2495,In_2025);
xnor U1806 (N_1806,In_2391,In_2195);
nand U1807 (N_1807,In_1782,In_1027);
and U1808 (N_1808,In_1784,In_999);
nand U1809 (N_1809,In_2953,In_1893);
nor U1810 (N_1810,In_827,In_1792);
xor U1811 (N_1811,In_1191,In_1074);
or U1812 (N_1812,In_2739,In_468);
nand U1813 (N_1813,In_173,In_2846);
and U1814 (N_1814,In_1382,In_293);
or U1815 (N_1815,In_2661,In_682);
nand U1816 (N_1816,In_2996,In_1923);
nor U1817 (N_1817,In_1071,In_1228);
nor U1818 (N_1818,In_467,In_1635);
nand U1819 (N_1819,In_1516,In_2077);
xnor U1820 (N_1820,In_922,In_2095);
nand U1821 (N_1821,In_1208,In_411);
nand U1822 (N_1822,In_2221,In_334);
nand U1823 (N_1823,In_1534,In_1214);
nor U1824 (N_1824,In_2486,In_2369);
nand U1825 (N_1825,In_303,In_1787);
and U1826 (N_1826,In_2628,In_2684);
nor U1827 (N_1827,In_2091,In_2259);
and U1828 (N_1828,In_1671,In_1155);
nor U1829 (N_1829,In_2159,In_1630);
or U1830 (N_1830,In_428,In_326);
nand U1831 (N_1831,In_889,In_1987);
nor U1832 (N_1832,In_2203,In_2690);
nand U1833 (N_1833,In_2431,In_1760);
and U1834 (N_1834,In_541,In_1380);
and U1835 (N_1835,In_25,In_706);
xor U1836 (N_1836,In_456,In_933);
or U1837 (N_1837,In_2067,In_369);
or U1838 (N_1838,In_838,In_421);
and U1839 (N_1839,In_2381,In_2227);
nor U1840 (N_1840,In_2077,In_473);
and U1841 (N_1841,In_345,In_2868);
nor U1842 (N_1842,In_157,In_1436);
and U1843 (N_1843,In_170,In_1746);
nand U1844 (N_1844,In_700,In_1787);
and U1845 (N_1845,In_1213,In_2091);
nor U1846 (N_1846,In_1273,In_2080);
nand U1847 (N_1847,In_1213,In_66);
and U1848 (N_1848,In_198,In_2067);
nand U1849 (N_1849,In_590,In_1781);
nand U1850 (N_1850,In_1740,In_2485);
and U1851 (N_1851,In_1756,In_2757);
or U1852 (N_1852,In_605,In_1713);
nor U1853 (N_1853,In_2604,In_1373);
nor U1854 (N_1854,In_461,In_1206);
nor U1855 (N_1855,In_720,In_1341);
nand U1856 (N_1856,In_493,In_484);
xnor U1857 (N_1857,In_2589,In_2432);
or U1858 (N_1858,In_1488,In_1545);
or U1859 (N_1859,In_1393,In_2552);
or U1860 (N_1860,In_502,In_2876);
xor U1861 (N_1861,In_672,In_2563);
nor U1862 (N_1862,In_1201,In_1450);
xnor U1863 (N_1863,In_956,In_1475);
and U1864 (N_1864,In_537,In_1356);
nor U1865 (N_1865,In_1717,In_652);
or U1866 (N_1866,In_1534,In_815);
and U1867 (N_1867,In_774,In_1441);
and U1868 (N_1868,In_1996,In_728);
and U1869 (N_1869,In_1755,In_1993);
nor U1870 (N_1870,In_1163,In_840);
or U1871 (N_1871,In_2427,In_1059);
nand U1872 (N_1872,In_713,In_2477);
or U1873 (N_1873,In_2389,In_324);
and U1874 (N_1874,In_2119,In_1198);
and U1875 (N_1875,In_2427,In_175);
nor U1876 (N_1876,In_1529,In_935);
or U1877 (N_1877,In_960,In_529);
xor U1878 (N_1878,In_813,In_490);
and U1879 (N_1879,In_1469,In_2183);
nor U1880 (N_1880,In_2745,In_197);
nor U1881 (N_1881,In_263,In_1068);
and U1882 (N_1882,In_1638,In_683);
and U1883 (N_1883,In_2658,In_2078);
nand U1884 (N_1884,In_1225,In_712);
and U1885 (N_1885,In_660,In_2389);
nor U1886 (N_1886,In_1925,In_2230);
nand U1887 (N_1887,In_1308,In_31);
nand U1888 (N_1888,In_824,In_1469);
xor U1889 (N_1889,In_810,In_435);
or U1890 (N_1890,In_776,In_2510);
xor U1891 (N_1891,In_545,In_2541);
xnor U1892 (N_1892,In_2980,In_2338);
nor U1893 (N_1893,In_1388,In_1015);
nor U1894 (N_1894,In_206,In_631);
nor U1895 (N_1895,In_2629,In_1495);
nor U1896 (N_1896,In_953,In_1099);
nor U1897 (N_1897,In_1736,In_2172);
nand U1898 (N_1898,In_2625,In_793);
and U1899 (N_1899,In_2784,In_2062);
nor U1900 (N_1900,In_2162,In_396);
xor U1901 (N_1901,In_2496,In_2545);
nand U1902 (N_1902,In_628,In_2779);
or U1903 (N_1903,In_1275,In_2999);
and U1904 (N_1904,In_2767,In_784);
or U1905 (N_1905,In_1042,In_1998);
or U1906 (N_1906,In_2639,In_1475);
and U1907 (N_1907,In_1267,In_1810);
xor U1908 (N_1908,In_383,In_1616);
and U1909 (N_1909,In_1420,In_418);
and U1910 (N_1910,In_2935,In_268);
nor U1911 (N_1911,In_2145,In_2685);
and U1912 (N_1912,In_286,In_2248);
nor U1913 (N_1913,In_2725,In_2643);
nor U1914 (N_1914,In_2610,In_813);
and U1915 (N_1915,In_1357,In_2448);
nor U1916 (N_1916,In_2179,In_1787);
or U1917 (N_1917,In_2187,In_1421);
nand U1918 (N_1918,In_644,In_1267);
nor U1919 (N_1919,In_1743,In_2901);
and U1920 (N_1920,In_1555,In_1540);
or U1921 (N_1921,In_896,In_2722);
nor U1922 (N_1922,In_2416,In_2687);
nand U1923 (N_1923,In_621,In_2823);
nand U1924 (N_1924,In_1385,In_2721);
nor U1925 (N_1925,In_981,In_1970);
and U1926 (N_1926,In_1404,In_1014);
and U1927 (N_1927,In_20,In_262);
nand U1928 (N_1928,In_1804,In_379);
or U1929 (N_1929,In_981,In_1067);
and U1930 (N_1930,In_121,In_940);
or U1931 (N_1931,In_2330,In_478);
or U1932 (N_1932,In_1140,In_2192);
nand U1933 (N_1933,In_2507,In_1479);
or U1934 (N_1934,In_2897,In_1230);
nand U1935 (N_1935,In_2338,In_2190);
nor U1936 (N_1936,In_2144,In_555);
or U1937 (N_1937,In_1256,In_411);
nand U1938 (N_1938,In_1826,In_852);
or U1939 (N_1939,In_2873,In_1734);
nor U1940 (N_1940,In_101,In_794);
and U1941 (N_1941,In_2389,In_1634);
nor U1942 (N_1942,In_795,In_504);
nor U1943 (N_1943,In_2062,In_2915);
and U1944 (N_1944,In_2887,In_853);
nor U1945 (N_1945,In_2141,In_1105);
nor U1946 (N_1946,In_509,In_1649);
nand U1947 (N_1947,In_1892,In_2327);
nor U1948 (N_1948,In_691,In_754);
or U1949 (N_1949,In_1035,In_353);
or U1950 (N_1950,In_2159,In_477);
nand U1951 (N_1951,In_1430,In_453);
nand U1952 (N_1952,In_1668,In_2214);
nand U1953 (N_1953,In_803,In_2075);
nor U1954 (N_1954,In_550,In_2265);
and U1955 (N_1955,In_2984,In_1151);
nor U1956 (N_1956,In_2660,In_1848);
nand U1957 (N_1957,In_1898,In_877);
nand U1958 (N_1958,In_2870,In_1456);
and U1959 (N_1959,In_754,In_2913);
and U1960 (N_1960,In_2996,In_495);
nor U1961 (N_1961,In_2750,In_2388);
nand U1962 (N_1962,In_1537,In_2008);
nand U1963 (N_1963,In_1977,In_2123);
nand U1964 (N_1964,In_736,In_891);
nor U1965 (N_1965,In_2148,In_2792);
nand U1966 (N_1966,In_1340,In_358);
or U1967 (N_1967,In_2603,In_2649);
nor U1968 (N_1968,In_451,In_2126);
or U1969 (N_1969,In_1886,In_2086);
xor U1970 (N_1970,In_680,In_1792);
nor U1971 (N_1971,In_66,In_2648);
nor U1972 (N_1972,In_1903,In_2509);
or U1973 (N_1973,In_1758,In_2114);
nand U1974 (N_1974,In_2339,In_2896);
or U1975 (N_1975,In_2749,In_2899);
nor U1976 (N_1976,In_510,In_1967);
nor U1977 (N_1977,In_2241,In_803);
or U1978 (N_1978,In_736,In_1311);
nor U1979 (N_1979,In_191,In_1940);
or U1980 (N_1980,In_2639,In_335);
and U1981 (N_1981,In_2109,In_1553);
xnor U1982 (N_1982,In_2896,In_890);
nand U1983 (N_1983,In_2939,In_1900);
and U1984 (N_1984,In_1870,In_2698);
or U1985 (N_1985,In_314,In_1172);
nand U1986 (N_1986,In_1219,In_772);
nand U1987 (N_1987,In_171,In_1095);
nand U1988 (N_1988,In_2698,In_34);
and U1989 (N_1989,In_1348,In_226);
nor U1990 (N_1990,In_279,In_1028);
and U1991 (N_1991,In_2665,In_2575);
nor U1992 (N_1992,In_1125,In_2969);
and U1993 (N_1993,In_763,In_1226);
nor U1994 (N_1994,In_1845,In_794);
and U1995 (N_1995,In_2975,In_1124);
xnor U1996 (N_1996,In_958,In_2799);
nand U1997 (N_1997,In_2940,In_2690);
and U1998 (N_1998,In_1209,In_364);
nand U1999 (N_1999,In_2900,In_632);
nor U2000 (N_2000,In_2026,In_914);
nor U2001 (N_2001,In_2597,In_1527);
and U2002 (N_2002,In_1268,In_68);
or U2003 (N_2003,In_332,In_1660);
nor U2004 (N_2004,In_1369,In_2884);
or U2005 (N_2005,In_1969,In_1089);
nand U2006 (N_2006,In_1816,In_2661);
and U2007 (N_2007,In_2901,In_1303);
nor U2008 (N_2008,In_1645,In_1850);
nand U2009 (N_2009,In_2615,In_510);
and U2010 (N_2010,In_723,In_1028);
nand U2011 (N_2011,In_1009,In_1285);
xnor U2012 (N_2012,In_1225,In_2015);
and U2013 (N_2013,In_2766,In_2148);
xnor U2014 (N_2014,In_1934,In_418);
nor U2015 (N_2015,In_2892,In_1854);
nand U2016 (N_2016,In_1146,In_344);
and U2017 (N_2017,In_654,In_1056);
nor U2018 (N_2018,In_2575,In_538);
nor U2019 (N_2019,In_2351,In_1794);
nor U2020 (N_2020,In_2752,In_2749);
nor U2021 (N_2021,In_1548,In_2094);
and U2022 (N_2022,In_1519,In_2396);
nand U2023 (N_2023,In_2645,In_1356);
xnor U2024 (N_2024,In_2556,In_405);
and U2025 (N_2025,In_1701,In_2419);
and U2026 (N_2026,In_2460,In_1680);
nor U2027 (N_2027,In_2477,In_846);
nand U2028 (N_2028,In_500,In_649);
nor U2029 (N_2029,In_848,In_695);
or U2030 (N_2030,In_1816,In_1164);
nand U2031 (N_2031,In_1195,In_1465);
or U2032 (N_2032,In_2302,In_2014);
and U2033 (N_2033,In_266,In_1968);
xnor U2034 (N_2034,In_876,In_1759);
nand U2035 (N_2035,In_1300,In_2990);
and U2036 (N_2036,In_1067,In_2122);
xnor U2037 (N_2037,In_2062,In_654);
nor U2038 (N_2038,In_589,In_2139);
or U2039 (N_2039,In_524,In_2198);
and U2040 (N_2040,In_828,In_2984);
nor U2041 (N_2041,In_501,In_2409);
and U2042 (N_2042,In_2529,In_1612);
nand U2043 (N_2043,In_2295,In_1387);
nand U2044 (N_2044,In_2152,In_658);
xor U2045 (N_2045,In_2095,In_2333);
and U2046 (N_2046,In_1707,In_1352);
nand U2047 (N_2047,In_2084,In_2039);
xnor U2048 (N_2048,In_2446,In_629);
nor U2049 (N_2049,In_2534,In_666);
nor U2050 (N_2050,In_678,In_2929);
or U2051 (N_2051,In_1288,In_1184);
nor U2052 (N_2052,In_2741,In_2263);
nand U2053 (N_2053,In_2844,In_2289);
nand U2054 (N_2054,In_427,In_778);
nand U2055 (N_2055,In_2341,In_1993);
or U2056 (N_2056,In_2415,In_114);
xnor U2057 (N_2057,In_2408,In_2918);
or U2058 (N_2058,In_910,In_999);
nor U2059 (N_2059,In_869,In_1458);
nor U2060 (N_2060,In_660,In_1605);
nor U2061 (N_2061,In_118,In_1810);
nor U2062 (N_2062,In_1041,In_2347);
and U2063 (N_2063,In_675,In_371);
xor U2064 (N_2064,In_1451,In_2549);
xnor U2065 (N_2065,In_2186,In_2209);
xor U2066 (N_2066,In_1389,In_2684);
xnor U2067 (N_2067,In_2735,In_2476);
nand U2068 (N_2068,In_381,In_1135);
nor U2069 (N_2069,In_2322,In_162);
nor U2070 (N_2070,In_147,In_2931);
or U2071 (N_2071,In_702,In_235);
or U2072 (N_2072,In_2069,In_30);
and U2073 (N_2073,In_588,In_2579);
nand U2074 (N_2074,In_2953,In_941);
or U2075 (N_2075,In_2177,In_1556);
xnor U2076 (N_2076,In_718,In_2232);
nand U2077 (N_2077,In_446,In_2093);
and U2078 (N_2078,In_1467,In_529);
or U2079 (N_2079,In_2007,In_1736);
nand U2080 (N_2080,In_1654,In_182);
xor U2081 (N_2081,In_652,In_2557);
or U2082 (N_2082,In_590,In_2212);
or U2083 (N_2083,In_2169,In_1478);
nor U2084 (N_2084,In_1368,In_811);
xnor U2085 (N_2085,In_2995,In_1605);
xnor U2086 (N_2086,In_626,In_2536);
nor U2087 (N_2087,In_2708,In_1910);
xnor U2088 (N_2088,In_739,In_2176);
and U2089 (N_2089,In_652,In_781);
or U2090 (N_2090,In_517,In_808);
or U2091 (N_2091,In_822,In_332);
xor U2092 (N_2092,In_290,In_510);
nand U2093 (N_2093,In_2607,In_1903);
and U2094 (N_2094,In_1132,In_478);
or U2095 (N_2095,In_1463,In_624);
or U2096 (N_2096,In_568,In_1366);
nand U2097 (N_2097,In_1781,In_1772);
xor U2098 (N_2098,In_1982,In_1764);
nand U2099 (N_2099,In_1285,In_3);
and U2100 (N_2100,In_1978,In_41);
and U2101 (N_2101,In_1998,In_952);
or U2102 (N_2102,In_2173,In_1716);
or U2103 (N_2103,In_2964,In_990);
nand U2104 (N_2104,In_1302,In_2612);
or U2105 (N_2105,In_1461,In_1053);
nor U2106 (N_2106,In_2210,In_728);
and U2107 (N_2107,In_171,In_2897);
nand U2108 (N_2108,In_2015,In_2970);
or U2109 (N_2109,In_1770,In_860);
and U2110 (N_2110,In_2343,In_2866);
or U2111 (N_2111,In_2921,In_2014);
nor U2112 (N_2112,In_2172,In_2730);
or U2113 (N_2113,In_2510,In_2745);
or U2114 (N_2114,In_2867,In_1643);
or U2115 (N_2115,In_1810,In_2344);
or U2116 (N_2116,In_1820,In_838);
or U2117 (N_2117,In_886,In_1778);
nand U2118 (N_2118,In_2183,In_761);
nor U2119 (N_2119,In_2394,In_930);
or U2120 (N_2120,In_1781,In_1997);
nor U2121 (N_2121,In_1251,In_659);
and U2122 (N_2122,In_221,In_647);
xor U2123 (N_2123,In_413,In_2382);
or U2124 (N_2124,In_1433,In_2639);
and U2125 (N_2125,In_919,In_2384);
nand U2126 (N_2126,In_2982,In_2360);
nor U2127 (N_2127,In_572,In_642);
nor U2128 (N_2128,In_2992,In_2019);
and U2129 (N_2129,In_2643,In_1331);
and U2130 (N_2130,In_1394,In_2917);
or U2131 (N_2131,In_2157,In_775);
xnor U2132 (N_2132,In_749,In_1480);
nor U2133 (N_2133,In_2290,In_1168);
and U2134 (N_2134,In_1342,In_2064);
nand U2135 (N_2135,In_199,In_1967);
nor U2136 (N_2136,In_1300,In_2822);
xnor U2137 (N_2137,In_121,In_2596);
or U2138 (N_2138,In_265,In_2752);
or U2139 (N_2139,In_1953,In_1453);
and U2140 (N_2140,In_443,In_2572);
and U2141 (N_2141,In_395,In_2399);
nand U2142 (N_2142,In_2546,In_1420);
nand U2143 (N_2143,In_2403,In_1735);
or U2144 (N_2144,In_1003,In_822);
or U2145 (N_2145,In_585,In_444);
nor U2146 (N_2146,In_1237,In_1356);
and U2147 (N_2147,In_1960,In_1863);
nand U2148 (N_2148,In_1579,In_1383);
and U2149 (N_2149,In_2962,In_2717);
or U2150 (N_2150,In_694,In_937);
nand U2151 (N_2151,In_2477,In_165);
nand U2152 (N_2152,In_1543,In_1748);
xnor U2153 (N_2153,In_2525,In_728);
nor U2154 (N_2154,In_2382,In_2595);
and U2155 (N_2155,In_1682,In_406);
and U2156 (N_2156,In_872,In_2684);
or U2157 (N_2157,In_1129,In_1814);
nand U2158 (N_2158,In_2886,In_352);
nand U2159 (N_2159,In_1390,In_389);
and U2160 (N_2160,In_417,In_1571);
nand U2161 (N_2161,In_1371,In_1917);
nor U2162 (N_2162,In_809,In_821);
nor U2163 (N_2163,In_685,In_1868);
or U2164 (N_2164,In_2392,In_2739);
and U2165 (N_2165,In_2990,In_1996);
xnor U2166 (N_2166,In_312,In_533);
xor U2167 (N_2167,In_1510,In_615);
nand U2168 (N_2168,In_2471,In_2558);
nor U2169 (N_2169,In_794,In_77);
nor U2170 (N_2170,In_434,In_1527);
and U2171 (N_2171,In_1390,In_1580);
or U2172 (N_2172,In_1103,In_94);
and U2173 (N_2173,In_1712,In_1391);
or U2174 (N_2174,In_2439,In_2498);
or U2175 (N_2175,In_1688,In_2857);
nor U2176 (N_2176,In_1934,In_234);
and U2177 (N_2177,In_1337,In_1592);
or U2178 (N_2178,In_1991,In_331);
and U2179 (N_2179,In_2014,In_2853);
nand U2180 (N_2180,In_2661,In_1006);
nor U2181 (N_2181,In_1249,In_2876);
nor U2182 (N_2182,In_2696,In_993);
or U2183 (N_2183,In_2752,In_420);
nor U2184 (N_2184,In_826,In_48);
nor U2185 (N_2185,In_2115,In_1656);
or U2186 (N_2186,In_81,In_1601);
nor U2187 (N_2187,In_676,In_1332);
nor U2188 (N_2188,In_1418,In_336);
nand U2189 (N_2189,In_705,In_2764);
or U2190 (N_2190,In_839,In_1666);
and U2191 (N_2191,In_1991,In_22);
or U2192 (N_2192,In_850,In_1742);
nor U2193 (N_2193,In_2190,In_2012);
or U2194 (N_2194,In_1661,In_449);
nand U2195 (N_2195,In_294,In_1366);
or U2196 (N_2196,In_2893,In_1679);
or U2197 (N_2197,In_2434,In_1581);
or U2198 (N_2198,In_2327,In_12);
nand U2199 (N_2199,In_2510,In_959);
nor U2200 (N_2200,In_2584,In_1608);
xor U2201 (N_2201,In_2555,In_1508);
or U2202 (N_2202,In_2794,In_1803);
nor U2203 (N_2203,In_2497,In_553);
or U2204 (N_2204,In_624,In_2955);
or U2205 (N_2205,In_840,In_1285);
xnor U2206 (N_2206,In_1539,In_697);
nand U2207 (N_2207,In_1760,In_11);
or U2208 (N_2208,In_582,In_2382);
or U2209 (N_2209,In_1992,In_1909);
nand U2210 (N_2210,In_1945,In_202);
and U2211 (N_2211,In_921,In_434);
nor U2212 (N_2212,In_2309,In_602);
and U2213 (N_2213,In_655,In_2331);
or U2214 (N_2214,In_1334,In_328);
or U2215 (N_2215,In_1143,In_2085);
nand U2216 (N_2216,In_843,In_618);
or U2217 (N_2217,In_2140,In_2085);
nor U2218 (N_2218,In_2766,In_2150);
xor U2219 (N_2219,In_88,In_471);
or U2220 (N_2220,In_1488,In_130);
or U2221 (N_2221,In_1137,In_259);
nor U2222 (N_2222,In_2115,In_1651);
nor U2223 (N_2223,In_679,In_2933);
nand U2224 (N_2224,In_2561,In_2487);
nor U2225 (N_2225,In_1745,In_2781);
and U2226 (N_2226,In_572,In_1000);
and U2227 (N_2227,In_2168,In_2149);
or U2228 (N_2228,In_1685,In_2783);
and U2229 (N_2229,In_2156,In_192);
or U2230 (N_2230,In_2299,In_2392);
nor U2231 (N_2231,In_2604,In_525);
or U2232 (N_2232,In_1595,In_764);
and U2233 (N_2233,In_921,In_1752);
and U2234 (N_2234,In_514,In_2501);
and U2235 (N_2235,In_117,In_47);
nor U2236 (N_2236,In_1357,In_2189);
nor U2237 (N_2237,In_1146,In_1620);
nand U2238 (N_2238,In_2057,In_1737);
and U2239 (N_2239,In_307,In_14);
or U2240 (N_2240,In_2902,In_2847);
or U2241 (N_2241,In_1362,In_1008);
and U2242 (N_2242,In_536,In_1317);
nor U2243 (N_2243,In_1258,In_1070);
nand U2244 (N_2244,In_870,In_2624);
and U2245 (N_2245,In_428,In_1474);
nand U2246 (N_2246,In_2823,In_645);
or U2247 (N_2247,In_1733,In_2623);
xnor U2248 (N_2248,In_610,In_920);
or U2249 (N_2249,In_2348,In_1350);
nor U2250 (N_2250,In_1311,In_551);
nand U2251 (N_2251,In_2625,In_2577);
and U2252 (N_2252,In_2197,In_1245);
nor U2253 (N_2253,In_703,In_2055);
or U2254 (N_2254,In_268,In_1146);
or U2255 (N_2255,In_1650,In_679);
and U2256 (N_2256,In_1650,In_1600);
and U2257 (N_2257,In_743,In_2982);
nor U2258 (N_2258,In_2166,In_77);
or U2259 (N_2259,In_2650,In_1952);
and U2260 (N_2260,In_2651,In_2398);
nand U2261 (N_2261,In_1705,In_1680);
and U2262 (N_2262,In_1541,In_2253);
and U2263 (N_2263,In_136,In_1409);
xnor U2264 (N_2264,In_2655,In_176);
xor U2265 (N_2265,In_2645,In_2787);
xnor U2266 (N_2266,In_846,In_612);
xnor U2267 (N_2267,In_64,In_2071);
nand U2268 (N_2268,In_1291,In_371);
nor U2269 (N_2269,In_826,In_273);
nor U2270 (N_2270,In_2939,In_2200);
nand U2271 (N_2271,In_2281,In_2136);
and U2272 (N_2272,In_2895,In_356);
xnor U2273 (N_2273,In_2738,In_1613);
nor U2274 (N_2274,In_510,In_2889);
or U2275 (N_2275,In_1357,In_925);
nand U2276 (N_2276,In_919,In_915);
nand U2277 (N_2277,In_2805,In_962);
and U2278 (N_2278,In_1121,In_2573);
nor U2279 (N_2279,In_870,In_1913);
and U2280 (N_2280,In_2323,In_2607);
nor U2281 (N_2281,In_1689,In_313);
nor U2282 (N_2282,In_2106,In_661);
nor U2283 (N_2283,In_2376,In_950);
and U2284 (N_2284,In_2551,In_2389);
nand U2285 (N_2285,In_2736,In_1992);
nor U2286 (N_2286,In_1535,In_2755);
xnor U2287 (N_2287,In_1697,In_722);
nand U2288 (N_2288,In_381,In_794);
and U2289 (N_2289,In_2655,In_41);
nand U2290 (N_2290,In_1937,In_873);
or U2291 (N_2291,In_1473,In_413);
nand U2292 (N_2292,In_2136,In_321);
nand U2293 (N_2293,In_406,In_2066);
or U2294 (N_2294,In_1391,In_2105);
or U2295 (N_2295,In_2981,In_1567);
nor U2296 (N_2296,In_2008,In_1935);
nor U2297 (N_2297,In_1452,In_411);
or U2298 (N_2298,In_2605,In_704);
nand U2299 (N_2299,In_1921,In_1911);
nand U2300 (N_2300,In_1912,In_498);
and U2301 (N_2301,In_2218,In_2923);
nand U2302 (N_2302,In_233,In_2941);
and U2303 (N_2303,In_1468,In_412);
and U2304 (N_2304,In_795,In_714);
nand U2305 (N_2305,In_969,In_51);
and U2306 (N_2306,In_1678,In_1603);
nand U2307 (N_2307,In_1212,In_49);
and U2308 (N_2308,In_281,In_728);
nor U2309 (N_2309,In_1796,In_2126);
nor U2310 (N_2310,In_1620,In_2976);
nor U2311 (N_2311,In_1391,In_714);
and U2312 (N_2312,In_2613,In_1979);
nor U2313 (N_2313,In_1261,In_89);
nor U2314 (N_2314,In_2722,In_2523);
nor U2315 (N_2315,In_1009,In_2383);
or U2316 (N_2316,In_2500,In_953);
nand U2317 (N_2317,In_806,In_1632);
nand U2318 (N_2318,In_781,In_2890);
and U2319 (N_2319,In_2185,In_563);
and U2320 (N_2320,In_1413,In_1709);
nand U2321 (N_2321,In_13,In_1908);
and U2322 (N_2322,In_2586,In_975);
nand U2323 (N_2323,In_2112,In_1575);
nor U2324 (N_2324,In_1184,In_797);
nor U2325 (N_2325,In_639,In_112);
or U2326 (N_2326,In_1913,In_420);
nand U2327 (N_2327,In_2467,In_907);
nand U2328 (N_2328,In_58,In_2246);
and U2329 (N_2329,In_2621,In_654);
xnor U2330 (N_2330,In_2951,In_2288);
and U2331 (N_2331,In_2855,In_1424);
and U2332 (N_2332,In_2549,In_574);
or U2333 (N_2333,In_497,In_529);
or U2334 (N_2334,In_1728,In_2001);
or U2335 (N_2335,In_1578,In_2145);
xnor U2336 (N_2336,In_297,In_603);
or U2337 (N_2337,In_1851,In_1832);
nor U2338 (N_2338,In_1809,In_2740);
nand U2339 (N_2339,In_1768,In_1668);
or U2340 (N_2340,In_871,In_2454);
nand U2341 (N_2341,In_2830,In_401);
or U2342 (N_2342,In_870,In_2035);
nor U2343 (N_2343,In_1151,In_353);
nand U2344 (N_2344,In_2996,In_2369);
nor U2345 (N_2345,In_972,In_73);
nand U2346 (N_2346,In_2651,In_187);
and U2347 (N_2347,In_1222,In_1812);
nor U2348 (N_2348,In_2187,In_1044);
nor U2349 (N_2349,In_946,In_702);
or U2350 (N_2350,In_2876,In_2346);
and U2351 (N_2351,In_2015,In_2157);
and U2352 (N_2352,In_496,In_2320);
nand U2353 (N_2353,In_682,In_209);
nand U2354 (N_2354,In_1336,In_107);
nor U2355 (N_2355,In_1040,In_2958);
nor U2356 (N_2356,In_2619,In_1842);
nor U2357 (N_2357,In_2753,In_541);
nor U2358 (N_2358,In_1968,In_2017);
nor U2359 (N_2359,In_2322,In_1379);
and U2360 (N_2360,In_2260,In_1612);
or U2361 (N_2361,In_341,In_2865);
nand U2362 (N_2362,In_2671,In_464);
nor U2363 (N_2363,In_1607,In_72);
xor U2364 (N_2364,In_545,In_2148);
or U2365 (N_2365,In_1061,In_1959);
nor U2366 (N_2366,In_2396,In_2166);
nand U2367 (N_2367,In_1332,In_1826);
nand U2368 (N_2368,In_1821,In_2392);
nand U2369 (N_2369,In_921,In_1263);
and U2370 (N_2370,In_824,In_1399);
or U2371 (N_2371,In_1354,In_281);
or U2372 (N_2372,In_1172,In_262);
or U2373 (N_2373,In_2392,In_388);
nor U2374 (N_2374,In_361,In_2892);
nor U2375 (N_2375,In_2731,In_1218);
or U2376 (N_2376,In_2246,In_1093);
and U2377 (N_2377,In_1242,In_627);
and U2378 (N_2378,In_2460,In_2152);
or U2379 (N_2379,In_1570,In_1308);
xnor U2380 (N_2380,In_541,In_271);
and U2381 (N_2381,In_2949,In_621);
xnor U2382 (N_2382,In_750,In_1884);
xor U2383 (N_2383,In_2792,In_294);
nand U2384 (N_2384,In_660,In_1825);
and U2385 (N_2385,In_276,In_2022);
or U2386 (N_2386,In_1806,In_2852);
and U2387 (N_2387,In_175,In_438);
nor U2388 (N_2388,In_2807,In_2481);
or U2389 (N_2389,In_1972,In_1811);
nor U2390 (N_2390,In_1692,In_2579);
nor U2391 (N_2391,In_787,In_2420);
nand U2392 (N_2392,In_30,In_2433);
nand U2393 (N_2393,In_706,In_651);
and U2394 (N_2394,In_1629,In_2401);
nor U2395 (N_2395,In_2811,In_683);
and U2396 (N_2396,In_1951,In_1096);
and U2397 (N_2397,In_2006,In_1047);
nor U2398 (N_2398,In_2928,In_2249);
and U2399 (N_2399,In_698,In_2690);
and U2400 (N_2400,In_252,In_1044);
nand U2401 (N_2401,In_2036,In_207);
nor U2402 (N_2402,In_1413,In_215);
nor U2403 (N_2403,In_614,In_671);
nand U2404 (N_2404,In_2314,In_2043);
or U2405 (N_2405,In_2628,In_1695);
nor U2406 (N_2406,In_2549,In_596);
nor U2407 (N_2407,In_620,In_410);
nand U2408 (N_2408,In_1999,In_998);
and U2409 (N_2409,In_1044,In_1570);
or U2410 (N_2410,In_2171,In_1465);
nor U2411 (N_2411,In_412,In_354);
or U2412 (N_2412,In_1998,In_2136);
and U2413 (N_2413,In_403,In_1795);
or U2414 (N_2414,In_1599,In_1);
xnor U2415 (N_2415,In_2117,In_2444);
nand U2416 (N_2416,In_918,In_1308);
and U2417 (N_2417,In_1126,In_1858);
nor U2418 (N_2418,In_1953,In_1108);
and U2419 (N_2419,In_2310,In_113);
nand U2420 (N_2420,In_2826,In_2509);
or U2421 (N_2421,In_2386,In_1301);
nor U2422 (N_2422,In_818,In_1299);
and U2423 (N_2423,In_1403,In_1648);
nor U2424 (N_2424,In_239,In_1732);
xor U2425 (N_2425,In_205,In_1629);
and U2426 (N_2426,In_2037,In_1205);
xor U2427 (N_2427,In_736,In_860);
xor U2428 (N_2428,In_1621,In_608);
and U2429 (N_2429,In_1618,In_1186);
and U2430 (N_2430,In_1549,In_766);
xor U2431 (N_2431,In_1441,In_1932);
nand U2432 (N_2432,In_2136,In_1375);
xnor U2433 (N_2433,In_2976,In_109);
or U2434 (N_2434,In_2312,In_1492);
nand U2435 (N_2435,In_450,In_1461);
nor U2436 (N_2436,In_148,In_4);
nor U2437 (N_2437,In_137,In_1070);
nand U2438 (N_2438,In_1255,In_57);
nand U2439 (N_2439,In_108,In_1592);
nor U2440 (N_2440,In_2559,In_1761);
nor U2441 (N_2441,In_2886,In_451);
nand U2442 (N_2442,In_1327,In_1565);
nand U2443 (N_2443,In_11,In_2627);
and U2444 (N_2444,In_944,In_1964);
and U2445 (N_2445,In_2383,In_793);
and U2446 (N_2446,In_2735,In_1351);
or U2447 (N_2447,In_508,In_187);
and U2448 (N_2448,In_2502,In_2248);
nand U2449 (N_2449,In_915,In_2175);
nand U2450 (N_2450,In_2662,In_810);
or U2451 (N_2451,In_1346,In_1187);
nand U2452 (N_2452,In_1148,In_84);
nand U2453 (N_2453,In_2594,In_1003);
nor U2454 (N_2454,In_1450,In_2272);
nor U2455 (N_2455,In_1410,In_1726);
nor U2456 (N_2456,In_1547,In_63);
nor U2457 (N_2457,In_1186,In_719);
or U2458 (N_2458,In_2182,In_591);
nor U2459 (N_2459,In_2277,In_1134);
and U2460 (N_2460,In_165,In_357);
and U2461 (N_2461,In_2789,In_2518);
nand U2462 (N_2462,In_1217,In_974);
nor U2463 (N_2463,In_2183,In_84);
nand U2464 (N_2464,In_1989,In_2895);
and U2465 (N_2465,In_1265,In_119);
nor U2466 (N_2466,In_2674,In_2821);
nor U2467 (N_2467,In_1848,In_1744);
or U2468 (N_2468,In_702,In_494);
nand U2469 (N_2469,In_292,In_853);
nand U2470 (N_2470,In_2996,In_555);
nor U2471 (N_2471,In_2975,In_1561);
nor U2472 (N_2472,In_671,In_553);
and U2473 (N_2473,In_433,In_987);
nand U2474 (N_2474,In_1687,In_101);
and U2475 (N_2475,In_1305,In_251);
nor U2476 (N_2476,In_59,In_655);
and U2477 (N_2477,In_2897,In_925);
and U2478 (N_2478,In_363,In_1868);
and U2479 (N_2479,In_2755,In_1292);
nor U2480 (N_2480,In_2724,In_465);
xnor U2481 (N_2481,In_2844,In_1455);
xnor U2482 (N_2482,In_1663,In_364);
nand U2483 (N_2483,In_634,In_2338);
nor U2484 (N_2484,In_2661,In_545);
or U2485 (N_2485,In_2976,In_472);
and U2486 (N_2486,In_1181,In_793);
nor U2487 (N_2487,In_2944,In_2685);
xnor U2488 (N_2488,In_890,In_928);
nor U2489 (N_2489,In_47,In_1362);
nor U2490 (N_2490,In_1935,In_1576);
nand U2491 (N_2491,In_2258,In_2661);
xor U2492 (N_2492,In_887,In_605);
or U2493 (N_2493,In_1715,In_2337);
nor U2494 (N_2494,In_62,In_1827);
nand U2495 (N_2495,In_296,In_1653);
or U2496 (N_2496,In_2345,In_1626);
nor U2497 (N_2497,In_1814,In_591);
nor U2498 (N_2498,In_2295,In_2496);
and U2499 (N_2499,In_1417,In_2511);
nand U2500 (N_2500,In_753,In_1725);
xor U2501 (N_2501,In_1477,In_1842);
nand U2502 (N_2502,In_44,In_1880);
and U2503 (N_2503,In_76,In_2896);
nor U2504 (N_2504,In_1685,In_453);
nor U2505 (N_2505,In_979,In_897);
nand U2506 (N_2506,In_391,In_515);
nor U2507 (N_2507,In_2579,In_1118);
and U2508 (N_2508,In_2536,In_243);
nor U2509 (N_2509,In_2574,In_1073);
and U2510 (N_2510,In_918,In_11);
xor U2511 (N_2511,In_1407,In_534);
or U2512 (N_2512,In_2408,In_378);
and U2513 (N_2513,In_2996,In_1548);
and U2514 (N_2514,In_2391,In_430);
or U2515 (N_2515,In_2704,In_2491);
or U2516 (N_2516,In_1633,In_2499);
nand U2517 (N_2517,In_1158,In_1046);
nor U2518 (N_2518,In_2756,In_404);
nor U2519 (N_2519,In_1789,In_263);
nand U2520 (N_2520,In_1370,In_941);
and U2521 (N_2521,In_126,In_640);
and U2522 (N_2522,In_1435,In_1362);
nand U2523 (N_2523,In_1634,In_807);
nor U2524 (N_2524,In_2242,In_358);
nand U2525 (N_2525,In_360,In_1828);
nor U2526 (N_2526,In_1773,In_30);
or U2527 (N_2527,In_1251,In_2783);
or U2528 (N_2528,In_462,In_687);
nand U2529 (N_2529,In_2502,In_31);
nor U2530 (N_2530,In_583,In_1072);
or U2531 (N_2531,In_2698,In_1150);
and U2532 (N_2532,In_2832,In_1471);
or U2533 (N_2533,In_2333,In_243);
nand U2534 (N_2534,In_2188,In_1506);
nand U2535 (N_2535,In_14,In_577);
nand U2536 (N_2536,In_1654,In_2211);
nor U2537 (N_2537,In_1124,In_1546);
and U2538 (N_2538,In_1196,In_1673);
nand U2539 (N_2539,In_869,In_629);
nand U2540 (N_2540,In_294,In_552);
and U2541 (N_2541,In_1741,In_1393);
nor U2542 (N_2542,In_788,In_2448);
and U2543 (N_2543,In_989,In_2216);
nand U2544 (N_2544,In_22,In_1645);
and U2545 (N_2545,In_1568,In_1037);
and U2546 (N_2546,In_2400,In_2481);
and U2547 (N_2547,In_46,In_1121);
or U2548 (N_2548,In_1704,In_2961);
xnor U2549 (N_2549,In_1262,In_576);
or U2550 (N_2550,In_874,In_54);
and U2551 (N_2551,In_670,In_900);
nand U2552 (N_2552,In_210,In_1284);
nor U2553 (N_2553,In_2058,In_1234);
or U2554 (N_2554,In_428,In_271);
xnor U2555 (N_2555,In_710,In_2509);
nor U2556 (N_2556,In_84,In_1035);
nor U2557 (N_2557,In_2158,In_841);
nor U2558 (N_2558,In_2398,In_2694);
and U2559 (N_2559,In_1680,In_207);
or U2560 (N_2560,In_602,In_2105);
nor U2561 (N_2561,In_355,In_663);
nand U2562 (N_2562,In_783,In_471);
and U2563 (N_2563,In_361,In_493);
and U2564 (N_2564,In_1744,In_793);
or U2565 (N_2565,In_714,In_18);
and U2566 (N_2566,In_551,In_1728);
and U2567 (N_2567,In_1816,In_2061);
xnor U2568 (N_2568,In_775,In_218);
and U2569 (N_2569,In_2325,In_2256);
and U2570 (N_2570,In_1105,In_166);
nor U2571 (N_2571,In_2799,In_2703);
xnor U2572 (N_2572,In_1326,In_1728);
nand U2573 (N_2573,In_1252,In_3);
and U2574 (N_2574,In_2367,In_1984);
nand U2575 (N_2575,In_1342,In_2371);
and U2576 (N_2576,In_1561,In_1879);
nand U2577 (N_2577,In_2082,In_1790);
and U2578 (N_2578,In_1474,In_1524);
xnor U2579 (N_2579,In_629,In_2868);
or U2580 (N_2580,In_1628,In_1213);
or U2581 (N_2581,In_2992,In_1714);
nand U2582 (N_2582,In_768,In_1037);
xnor U2583 (N_2583,In_737,In_182);
nor U2584 (N_2584,In_0,In_59);
or U2585 (N_2585,In_1941,In_263);
or U2586 (N_2586,In_906,In_1545);
nand U2587 (N_2587,In_2160,In_1433);
nor U2588 (N_2588,In_1861,In_381);
nor U2589 (N_2589,In_1091,In_2806);
nand U2590 (N_2590,In_197,In_1708);
nand U2591 (N_2591,In_607,In_1961);
nand U2592 (N_2592,In_668,In_535);
nor U2593 (N_2593,In_1016,In_2503);
nor U2594 (N_2594,In_2012,In_1144);
or U2595 (N_2595,In_482,In_1745);
or U2596 (N_2596,In_371,In_2257);
and U2597 (N_2597,In_2427,In_1583);
or U2598 (N_2598,In_35,In_372);
or U2599 (N_2599,In_923,In_2789);
nand U2600 (N_2600,In_55,In_2604);
xor U2601 (N_2601,In_1852,In_2927);
nor U2602 (N_2602,In_1538,In_80);
or U2603 (N_2603,In_1065,In_407);
nor U2604 (N_2604,In_1803,In_801);
and U2605 (N_2605,In_2508,In_752);
xor U2606 (N_2606,In_1489,In_2033);
nor U2607 (N_2607,In_746,In_522);
nand U2608 (N_2608,In_1851,In_96);
nor U2609 (N_2609,In_2343,In_130);
or U2610 (N_2610,In_243,In_1137);
or U2611 (N_2611,In_2643,In_663);
nand U2612 (N_2612,In_2298,In_216);
nand U2613 (N_2613,In_279,In_2278);
and U2614 (N_2614,In_29,In_2754);
nor U2615 (N_2615,In_1406,In_1879);
nor U2616 (N_2616,In_1516,In_2137);
and U2617 (N_2617,In_397,In_45);
or U2618 (N_2618,In_2517,In_1138);
nand U2619 (N_2619,In_143,In_2907);
nor U2620 (N_2620,In_1680,In_2354);
or U2621 (N_2621,In_2997,In_901);
xor U2622 (N_2622,In_697,In_547);
or U2623 (N_2623,In_147,In_1341);
or U2624 (N_2624,In_2073,In_119);
and U2625 (N_2625,In_1634,In_2281);
and U2626 (N_2626,In_1577,In_462);
nor U2627 (N_2627,In_77,In_1100);
or U2628 (N_2628,In_752,In_832);
or U2629 (N_2629,In_2928,In_753);
nor U2630 (N_2630,In_2751,In_1206);
and U2631 (N_2631,In_699,In_144);
nand U2632 (N_2632,In_2434,In_2547);
and U2633 (N_2633,In_24,In_289);
and U2634 (N_2634,In_1489,In_1987);
and U2635 (N_2635,In_2721,In_2387);
nand U2636 (N_2636,In_2949,In_2213);
nor U2637 (N_2637,In_202,In_1906);
or U2638 (N_2638,In_2778,In_10);
nor U2639 (N_2639,In_601,In_854);
and U2640 (N_2640,In_1385,In_79);
nand U2641 (N_2641,In_2247,In_1990);
nand U2642 (N_2642,In_2207,In_2773);
or U2643 (N_2643,In_198,In_1836);
or U2644 (N_2644,In_1916,In_1742);
or U2645 (N_2645,In_1498,In_456);
xor U2646 (N_2646,In_1795,In_2306);
or U2647 (N_2647,In_2100,In_664);
and U2648 (N_2648,In_2976,In_11);
xor U2649 (N_2649,In_1393,In_1480);
nand U2650 (N_2650,In_1377,In_838);
or U2651 (N_2651,In_449,In_177);
and U2652 (N_2652,In_1795,In_95);
or U2653 (N_2653,In_1672,In_636);
nand U2654 (N_2654,In_1833,In_864);
and U2655 (N_2655,In_2715,In_1898);
nand U2656 (N_2656,In_1215,In_2153);
or U2657 (N_2657,In_1735,In_1759);
and U2658 (N_2658,In_1198,In_772);
nor U2659 (N_2659,In_1718,In_262);
and U2660 (N_2660,In_2793,In_2590);
or U2661 (N_2661,In_1879,In_632);
xnor U2662 (N_2662,In_1869,In_2016);
xor U2663 (N_2663,In_1242,In_2376);
xor U2664 (N_2664,In_2700,In_1356);
and U2665 (N_2665,In_2352,In_163);
nor U2666 (N_2666,In_1174,In_1571);
or U2667 (N_2667,In_2528,In_2284);
nor U2668 (N_2668,In_2453,In_2753);
or U2669 (N_2669,In_595,In_1032);
or U2670 (N_2670,In_214,In_1671);
and U2671 (N_2671,In_1210,In_1827);
and U2672 (N_2672,In_2974,In_854);
and U2673 (N_2673,In_1750,In_2398);
or U2674 (N_2674,In_527,In_603);
xor U2675 (N_2675,In_774,In_2454);
nor U2676 (N_2676,In_2240,In_281);
and U2677 (N_2677,In_1738,In_16);
nor U2678 (N_2678,In_2770,In_2071);
nor U2679 (N_2679,In_1235,In_1594);
nand U2680 (N_2680,In_1701,In_1022);
nand U2681 (N_2681,In_1987,In_2130);
or U2682 (N_2682,In_2884,In_1224);
and U2683 (N_2683,In_570,In_611);
and U2684 (N_2684,In_936,In_2485);
nor U2685 (N_2685,In_518,In_2264);
and U2686 (N_2686,In_990,In_352);
nor U2687 (N_2687,In_82,In_181);
or U2688 (N_2688,In_154,In_2108);
and U2689 (N_2689,In_785,In_1352);
and U2690 (N_2690,In_2038,In_301);
nor U2691 (N_2691,In_1200,In_2239);
and U2692 (N_2692,In_1920,In_908);
or U2693 (N_2693,In_1354,In_1176);
and U2694 (N_2694,In_764,In_1841);
and U2695 (N_2695,In_1247,In_1287);
nand U2696 (N_2696,In_1490,In_2401);
nand U2697 (N_2697,In_612,In_2461);
nand U2698 (N_2698,In_2111,In_208);
nor U2699 (N_2699,In_2773,In_2654);
nor U2700 (N_2700,In_831,In_169);
or U2701 (N_2701,In_74,In_846);
nor U2702 (N_2702,In_834,In_2248);
or U2703 (N_2703,In_1764,In_2551);
xnor U2704 (N_2704,In_1415,In_437);
and U2705 (N_2705,In_1140,In_1589);
nor U2706 (N_2706,In_2444,In_768);
and U2707 (N_2707,In_1784,In_1229);
and U2708 (N_2708,In_910,In_1728);
nor U2709 (N_2709,In_1243,In_1701);
nand U2710 (N_2710,In_2730,In_239);
xor U2711 (N_2711,In_1559,In_2199);
nand U2712 (N_2712,In_2097,In_2062);
or U2713 (N_2713,In_2446,In_42);
or U2714 (N_2714,In_2841,In_2972);
and U2715 (N_2715,In_2420,In_2276);
and U2716 (N_2716,In_209,In_75);
and U2717 (N_2717,In_1722,In_934);
nor U2718 (N_2718,In_614,In_2813);
and U2719 (N_2719,In_2959,In_2635);
and U2720 (N_2720,In_313,In_1115);
nor U2721 (N_2721,In_918,In_1185);
and U2722 (N_2722,In_936,In_1598);
nand U2723 (N_2723,In_2924,In_1679);
xor U2724 (N_2724,In_1189,In_2928);
and U2725 (N_2725,In_2878,In_925);
nor U2726 (N_2726,In_2522,In_2906);
nand U2727 (N_2727,In_1400,In_2443);
and U2728 (N_2728,In_701,In_866);
or U2729 (N_2729,In_2865,In_1689);
or U2730 (N_2730,In_1898,In_1017);
nor U2731 (N_2731,In_1435,In_2039);
nor U2732 (N_2732,In_1505,In_2223);
nand U2733 (N_2733,In_1321,In_2241);
and U2734 (N_2734,In_2289,In_86);
nand U2735 (N_2735,In_889,In_1217);
nor U2736 (N_2736,In_648,In_477);
and U2737 (N_2737,In_763,In_1169);
and U2738 (N_2738,In_1479,In_657);
or U2739 (N_2739,In_404,In_599);
nand U2740 (N_2740,In_465,In_2746);
nand U2741 (N_2741,In_77,In_2886);
nand U2742 (N_2742,In_1056,In_820);
or U2743 (N_2743,In_1112,In_1505);
nor U2744 (N_2744,In_2358,In_462);
and U2745 (N_2745,In_2361,In_2304);
nor U2746 (N_2746,In_2199,In_827);
nand U2747 (N_2747,In_2008,In_1071);
nor U2748 (N_2748,In_59,In_2273);
and U2749 (N_2749,In_307,In_894);
nor U2750 (N_2750,In_90,In_605);
and U2751 (N_2751,In_1348,In_1625);
xnor U2752 (N_2752,In_1113,In_942);
and U2753 (N_2753,In_1725,In_1527);
and U2754 (N_2754,In_1316,In_210);
or U2755 (N_2755,In_1446,In_1721);
and U2756 (N_2756,In_1526,In_2464);
and U2757 (N_2757,In_1925,In_2866);
or U2758 (N_2758,In_2298,In_1525);
nand U2759 (N_2759,In_2443,In_815);
and U2760 (N_2760,In_896,In_781);
or U2761 (N_2761,In_2781,In_321);
nand U2762 (N_2762,In_1717,In_2403);
or U2763 (N_2763,In_2299,In_1538);
nand U2764 (N_2764,In_1141,In_593);
or U2765 (N_2765,In_331,In_1728);
and U2766 (N_2766,In_2853,In_518);
nor U2767 (N_2767,In_691,In_1279);
or U2768 (N_2768,In_2262,In_573);
nand U2769 (N_2769,In_542,In_2832);
and U2770 (N_2770,In_41,In_1502);
or U2771 (N_2771,In_1502,In_1290);
or U2772 (N_2772,In_2599,In_1195);
or U2773 (N_2773,In_2211,In_1896);
nor U2774 (N_2774,In_63,In_2842);
and U2775 (N_2775,In_1336,In_1412);
nor U2776 (N_2776,In_1706,In_680);
or U2777 (N_2777,In_2296,In_658);
and U2778 (N_2778,In_303,In_2262);
nand U2779 (N_2779,In_1730,In_2536);
and U2780 (N_2780,In_124,In_2076);
or U2781 (N_2781,In_2052,In_260);
or U2782 (N_2782,In_754,In_302);
or U2783 (N_2783,In_1173,In_567);
or U2784 (N_2784,In_1266,In_1031);
xnor U2785 (N_2785,In_2712,In_2032);
nand U2786 (N_2786,In_315,In_850);
nand U2787 (N_2787,In_2390,In_1472);
and U2788 (N_2788,In_1147,In_2254);
or U2789 (N_2789,In_271,In_1268);
nor U2790 (N_2790,In_405,In_580);
and U2791 (N_2791,In_934,In_904);
xor U2792 (N_2792,In_154,In_1768);
nand U2793 (N_2793,In_753,In_1362);
and U2794 (N_2794,In_764,In_1717);
nand U2795 (N_2795,In_2074,In_2778);
or U2796 (N_2796,In_166,In_1719);
or U2797 (N_2797,In_2705,In_538);
or U2798 (N_2798,In_1472,In_268);
xnor U2799 (N_2799,In_1160,In_1928);
xor U2800 (N_2800,In_2359,In_1799);
and U2801 (N_2801,In_1419,In_2112);
nand U2802 (N_2802,In_2890,In_2221);
or U2803 (N_2803,In_1943,In_1158);
or U2804 (N_2804,In_2175,In_1110);
nor U2805 (N_2805,In_1196,In_1638);
xnor U2806 (N_2806,In_770,In_513);
nor U2807 (N_2807,In_973,In_143);
and U2808 (N_2808,In_1526,In_1054);
and U2809 (N_2809,In_237,In_1875);
nor U2810 (N_2810,In_2350,In_1755);
nor U2811 (N_2811,In_1473,In_2194);
nor U2812 (N_2812,In_1015,In_584);
or U2813 (N_2813,In_1380,In_1098);
and U2814 (N_2814,In_2239,In_905);
and U2815 (N_2815,In_1242,In_2048);
and U2816 (N_2816,In_759,In_2334);
and U2817 (N_2817,In_1254,In_2191);
or U2818 (N_2818,In_1770,In_2803);
or U2819 (N_2819,In_103,In_2715);
nand U2820 (N_2820,In_2993,In_615);
and U2821 (N_2821,In_1142,In_2677);
nor U2822 (N_2822,In_2284,In_2470);
nand U2823 (N_2823,In_2375,In_2449);
nor U2824 (N_2824,In_1895,In_1811);
and U2825 (N_2825,In_1173,In_1444);
and U2826 (N_2826,In_2574,In_2163);
and U2827 (N_2827,In_1375,In_933);
nor U2828 (N_2828,In_2874,In_1222);
nand U2829 (N_2829,In_1381,In_45);
or U2830 (N_2830,In_1223,In_2516);
or U2831 (N_2831,In_2355,In_505);
and U2832 (N_2832,In_966,In_1487);
or U2833 (N_2833,In_2023,In_112);
and U2834 (N_2834,In_2047,In_706);
xor U2835 (N_2835,In_2379,In_1221);
or U2836 (N_2836,In_1413,In_78);
and U2837 (N_2837,In_603,In_582);
and U2838 (N_2838,In_157,In_486);
or U2839 (N_2839,In_2672,In_1598);
and U2840 (N_2840,In_1517,In_1001);
nor U2841 (N_2841,In_411,In_826);
nor U2842 (N_2842,In_2590,In_773);
and U2843 (N_2843,In_126,In_1122);
nor U2844 (N_2844,In_1576,In_1060);
nand U2845 (N_2845,In_446,In_129);
xnor U2846 (N_2846,In_2565,In_2005);
or U2847 (N_2847,In_1736,In_124);
nor U2848 (N_2848,In_2148,In_177);
or U2849 (N_2849,In_2156,In_383);
nor U2850 (N_2850,In_2465,In_382);
nand U2851 (N_2851,In_2834,In_180);
nor U2852 (N_2852,In_1671,In_181);
nor U2853 (N_2853,In_2738,In_2499);
nor U2854 (N_2854,In_1936,In_1454);
nor U2855 (N_2855,In_1404,In_1491);
xor U2856 (N_2856,In_1569,In_1671);
nor U2857 (N_2857,In_2484,In_74);
nand U2858 (N_2858,In_1841,In_1456);
nand U2859 (N_2859,In_2530,In_0);
nor U2860 (N_2860,In_567,In_1648);
nor U2861 (N_2861,In_2555,In_2537);
xor U2862 (N_2862,In_777,In_1190);
and U2863 (N_2863,In_2197,In_2808);
nand U2864 (N_2864,In_1162,In_2022);
nand U2865 (N_2865,In_2007,In_1320);
nor U2866 (N_2866,In_1472,In_219);
and U2867 (N_2867,In_994,In_1140);
nor U2868 (N_2868,In_1591,In_1991);
nand U2869 (N_2869,In_7,In_1499);
nor U2870 (N_2870,In_712,In_176);
nor U2871 (N_2871,In_527,In_1754);
and U2872 (N_2872,In_1218,In_1981);
nor U2873 (N_2873,In_1253,In_165);
or U2874 (N_2874,In_2172,In_1765);
or U2875 (N_2875,In_2934,In_1845);
nor U2876 (N_2876,In_2252,In_1256);
or U2877 (N_2877,In_1502,In_531);
nor U2878 (N_2878,In_245,In_930);
xnor U2879 (N_2879,In_1517,In_2331);
xnor U2880 (N_2880,In_345,In_1894);
nand U2881 (N_2881,In_962,In_1824);
or U2882 (N_2882,In_361,In_2443);
xor U2883 (N_2883,In_2387,In_2810);
xor U2884 (N_2884,In_536,In_2841);
and U2885 (N_2885,In_42,In_748);
nand U2886 (N_2886,In_228,In_1821);
nor U2887 (N_2887,In_24,In_1085);
nand U2888 (N_2888,In_556,In_1911);
or U2889 (N_2889,In_801,In_2944);
and U2890 (N_2890,In_2596,In_0);
xnor U2891 (N_2891,In_831,In_1387);
and U2892 (N_2892,In_1120,In_2914);
nor U2893 (N_2893,In_2601,In_2945);
and U2894 (N_2894,In_2146,In_2917);
or U2895 (N_2895,In_397,In_1837);
xnor U2896 (N_2896,In_196,In_353);
nor U2897 (N_2897,In_2669,In_1179);
nor U2898 (N_2898,In_1703,In_1327);
nor U2899 (N_2899,In_1975,In_2671);
nand U2900 (N_2900,In_2676,In_1245);
and U2901 (N_2901,In_1243,In_2875);
nand U2902 (N_2902,In_2558,In_861);
nand U2903 (N_2903,In_2434,In_2219);
or U2904 (N_2904,In_1609,In_1685);
nor U2905 (N_2905,In_1074,In_1105);
xor U2906 (N_2906,In_527,In_959);
nor U2907 (N_2907,In_1591,In_1231);
xnor U2908 (N_2908,In_830,In_2406);
or U2909 (N_2909,In_852,In_202);
or U2910 (N_2910,In_592,In_1716);
nand U2911 (N_2911,In_377,In_2799);
or U2912 (N_2912,In_822,In_2834);
and U2913 (N_2913,In_168,In_546);
nand U2914 (N_2914,In_17,In_2051);
nor U2915 (N_2915,In_1671,In_2324);
or U2916 (N_2916,In_804,In_1279);
nor U2917 (N_2917,In_2577,In_154);
and U2918 (N_2918,In_836,In_962);
xnor U2919 (N_2919,In_157,In_2136);
xnor U2920 (N_2920,In_1399,In_114);
nand U2921 (N_2921,In_2603,In_826);
or U2922 (N_2922,In_514,In_1052);
and U2923 (N_2923,In_2265,In_1108);
nor U2924 (N_2924,In_2750,In_1801);
nor U2925 (N_2925,In_1533,In_1615);
and U2926 (N_2926,In_459,In_1141);
nand U2927 (N_2927,In_1357,In_2789);
nor U2928 (N_2928,In_2053,In_286);
nor U2929 (N_2929,In_261,In_2506);
nand U2930 (N_2930,In_2815,In_2443);
nor U2931 (N_2931,In_628,In_1621);
nor U2932 (N_2932,In_2921,In_2642);
nand U2933 (N_2933,In_2935,In_1506);
or U2934 (N_2934,In_2889,In_1882);
and U2935 (N_2935,In_1984,In_1461);
or U2936 (N_2936,In_96,In_425);
xor U2937 (N_2937,In_1989,In_1985);
nand U2938 (N_2938,In_2611,In_1404);
nor U2939 (N_2939,In_2115,In_180);
or U2940 (N_2940,In_2791,In_2623);
and U2941 (N_2941,In_215,In_498);
and U2942 (N_2942,In_1325,In_269);
or U2943 (N_2943,In_2984,In_517);
or U2944 (N_2944,In_1546,In_2407);
or U2945 (N_2945,In_2691,In_2384);
and U2946 (N_2946,In_2522,In_2042);
nand U2947 (N_2947,In_2896,In_2974);
nand U2948 (N_2948,In_2626,In_1633);
nor U2949 (N_2949,In_100,In_75);
nor U2950 (N_2950,In_2873,In_1804);
nand U2951 (N_2951,In_1946,In_1778);
nand U2952 (N_2952,In_2224,In_591);
and U2953 (N_2953,In_1866,In_136);
nand U2954 (N_2954,In_806,In_2471);
nor U2955 (N_2955,In_2965,In_1854);
nor U2956 (N_2956,In_216,In_1682);
and U2957 (N_2957,In_1719,In_1230);
nor U2958 (N_2958,In_216,In_740);
xnor U2959 (N_2959,In_649,In_487);
nand U2960 (N_2960,In_1980,In_1418);
xor U2961 (N_2961,In_636,In_1434);
or U2962 (N_2962,In_1669,In_2579);
nand U2963 (N_2963,In_2046,In_1122);
or U2964 (N_2964,In_2654,In_129);
or U2965 (N_2965,In_2236,In_65);
nor U2966 (N_2966,In_1057,In_893);
nor U2967 (N_2967,In_2284,In_2956);
nand U2968 (N_2968,In_427,In_558);
nor U2969 (N_2969,In_2089,In_1491);
nor U2970 (N_2970,In_1555,In_2642);
and U2971 (N_2971,In_2972,In_1290);
or U2972 (N_2972,In_758,In_739);
nand U2973 (N_2973,In_2797,In_2654);
nand U2974 (N_2974,In_2097,In_2748);
xor U2975 (N_2975,In_261,In_2025);
nor U2976 (N_2976,In_1608,In_779);
nor U2977 (N_2977,In_1320,In_2177);
nand U2978 (N_2978,In_1048,In_596);
nand U2979 (N_2979,In_813,In_1805);
nand U2980 (N_2980,In_480,In_2550);
and U2981 (N_2981,In_1646,In_2353);
or U2982 (N_2982,In_485,In_1065);
or U2983 (N_2983,In_2872,In_475);
and U2984 (N_2984,In_713,In_172);
or U2985 (N_2985,In_2313,In_1336);
or U2986 (N_2986,In_1599,In_439);
or U2987 (N_2987,In_2304,In_1920);
nor U2988 (N_2988,In_1104,In_262);
nand U2989 (N_2989,In_1231,In_488);
nor U2990 (N_2990,In_519,In_1230);
or U2991 (N_2991,In_1040,In_2095);
nand U2992 (N_2992,In_101,In_1412);
nand U2993 (N_2993,In_2438,In_1831);
or U2994 (N_2994,In_913,In_1201);
nand U2995 (N_2995,In_682,In_1294);
nor U2996 (N_2996,In_886,In_751);
nand U2997 (N_2997,In_809,In_111);
and U2998 (N_2998,In_2984,In_1660);
nor U2999 (N_2999,In_1724,In_2818);
and U3000 (N_3000,In_652,In_1219);
nand U3001 (N_3001,In_406,In_1611);
and U3002 (N_3002,In_1097,In_1915);
xnor U3003 (N_3003,In_403,In_2030);
nand U3004 (N_3004,In_2727,In_2145);
nor U3005 (N_3005,In_2236,In_2898);
and U3006 (N_3006,In_1049,In_707);
nand U3007 (N_3007,In_1242,In_97);
nor U3008 (N_3008,In_2483,In_2169);
nand U3009 (N_3009,In_150,In_2262);
nand U3010 (N_3010,In_156,In_1044);
and U3011 (N_3011,In_473,In_1141);
and U3012 (N_3012,In_1598,In_2151);
and U3013 (N_3013,In_2032,In_1136);
nor U3014 (N_3014,In_160,In_87);
xnor U3015 (N_3015,In_2508,In_472);
nand U3016 (N_3016,In_2005,In_2290);
nand U3017 (N_3017,In_525,In_1502);
or U3018 (N_3018,In_2465,In_1011);
or U3019 (N_3019,In_2132,In_2927);
xor U3020 (N_3020,In_2098,In_1923);
nor U3021 (N_3021,In_336,In_1492);
or U3022 (N_3022,In_1901,In_2688);
xnor U3023 (N_3023,In_2199,In_2597);
xor U3024 (N_3024,In_496,In_1496);
nor U3025 (N_3025,In_1316,In_385);
and U3026 (N_3026,In_71,In_1168);
xnor U3027 (N_3027,In_249,In_756);
and U3028 (N_3028,In_816,In_328);
nand U3029 (N_3029,In_1211,In_2917);
and U3030 (N_3030,In_910,In_1387);
and U3031 (N_3031,In_2111,In_404);
nor U3032 (N_3032,In_2012,In_247);
nor U3033 (N_3033,In_9,In_1290);
and U3034 (N_3034,In_2206,In_819);
nor U3035 (N_3035,In_1607,In_939);
nor U3036 (N_3036,In_2481,In_1849);
nand U3037 (N_3037,In_1086,In_1872);
and U3038 (N_3038,In_2517,In_378);
nor U3039 (N_3039,In_1488,In_649);
nor U3040 (N_3040,In_1699,In_2486);
xnor U3041 (N_3041,In_2825,In_1931);
or U3042 (N_3042,In_813,In_1352);
nor U3043 (N_3043,In_2621,In_1415);
nor U3044 (N_3044,In_2763,In_1304);
and U3045 (N_3045,In_610,In_1546);
nor U3046 (N_3046,In_2699,In_2559);
nand U3047 (N_3047,In_2643,In_820);
and U3048 (N_3048,In_2695,In_56);
nand U3049 (N_3049,In_901,In_2404);
or U3050 (N_3050,In_723,In_339);
or U3051 (N_3051,In_2118,In_1534);
and U3052 (N_3052,In_2216,In_646);
nor U3053 (N_3053,In_2294,In_1932);
and U3054 (N_3054,In_1109,In_988);
or U3055 (N_3055,In_2379,In_2145);
nand U3056 (N_3056,In_2419,In_2335);
nand U3057 (N_3057,In_817,In_2009);
or U3058 (N_3058,In_1131,In_267);
and U3059 (N_3059,In_669,In_2590);
and U3060 (N_3060,In_1987,In_501);
nor U3061 (N_3061,In_787,In_76);
or U3062 (N_3062,In_2650,In_2991);
xor U3063 (N_3063,In_2044,In_2701);
or U3064 (N_3064,In_2050,In_1704);
nor U3065 (N_3065,In_592,In_2051);
or U3066 (N_3066,In_1772,In_511);
nand U3067 (N_3067,In_1305,In_1471);
xor U3068 (N_3068,In_987,In_2399);
and U3069 (N_3069,In_112,In_105);
nand U3070 (N_3070,In_900,In_2786);
nand U3071 (N_3071,In_1551,In_826);
nor U3072 (N_3072,In_607,In_445);
or U3073 (N_3073,In_41,In_348);
or U3074 (N_3074,In_1326,In_1503);
and U3075 (N_3075,In_1728,In_7);
or U3076 (N_3076,In_2176,In_2436);
xnor U3077 (N_3077,In_845,In_1886);
and U3078 (N_3078,In_1372,In_328);
or U3079 (N_3079,In_1616,In_2349);
and U3080 (N_3080,In_1066,In_674);
and U3081 (N_3081,In_2832,In_1982);
or U3082 (N_3082,In_2321,In_174);
nor U3083 (N_3083,In_2978,In_462);
nor U3084 (N_3084,In_343,In_2574);
nor U3085 (N_3085,In_72,In_2754);
or U3086 (N_3086,In_760,In_1380);
xor U3087 (N_3087,In_1041,In_1539);
xnor U3088 (N_3088,In_2810,In_387);
nor U3089 (N_3089,In_1084,In_2243);
nand U3090 (N_3090,In_2727,In_1845);
nand U3091 (N_3091,In_1051,In_2737);
and U3092 (N_3092,In_1209,In_518);
xor U3093 (N_3093,In_1577,In_524);
nor U3094 (N_3094,In_1552,In_1963);
nand U3095 (N_3095,In_2899,In_1923);
nor U3096 (N_3096,In_2873,In_942);
nor U3097 (N_3097,In_1438,In_1627);
nor U3098 (N_3098,In_99,In_1474);
and U3099 (N_3099,In_865,In_366);
nor U3100 (N_3100,In_2043,In_16);
nand U3101 (N_3101,In_2242,In_695);
and U3102 (N_3102,In_2414,In_2224);
nand U3103 (N_3103,In_1188,In_2099);
xnor U3104 (N_3104,In_2517,In_2330);
nand U3105 (N_3105,In_2488,In_1640);
nor U3106 (N_3106,In_99,In_1640);
or U3107 (N_3107,In_233,In_351);
nor U3108 (N_3108,In_1927,In_192);
nor U3109 (N_3109,In_1383,In_709);
nor U3110 (N_3110,In_2392,In_600);
nand U3111 (N_3111,In_428,In_497);
nor U3112 (N_3112,In_1162,In_2209);
and U3113 (N_3113,In_2132,In_2896);
or U3114 (N_3114,In_1428,In_163);
or U3115 (N_3115,In_2802,In_2256);
and U3116 (N_3116,In_56,In_2604);
nand U3117 (N_3117,In_207,In_1204);
or U3118 (N_3118,In_2273,In_2336);
nor U3119 (N_3119,In_2058,In_1272);
nor U3120 (N_3120,In_809,In_422);
or U3121 (N_3121,In_1684,In_2393);
and U3122 (N_3122,In_1223,In_1496);
nand U3123 (N_3123,In_2632,In_1397);
nand U3124 (N_3124,In_388,In_2537);
or U3125 (N_3125,In_2575,In_1380);
and U3126 (N_3126,In_2985,In_2167);
or U3127 (N_3127,In_1692,In_2601);
nand U3128 (N_3128,In_1048,In_2730);
nand U3129 (N_3129,In_1835,In_2022);
nor U3130 (N_3130,In_44,In_1307);
and U3131 (N_3131,In_446,In_1162);
or U3132 (N_3132,In_2029,In_2143);
and U3133 (N_3133,In_633,In_1837);
xnor U3134 (N_3134,In_1069,In_736);
and U3135 (N_3135,In_2002,In_221);
nor U3136 (N_3136,In_846,In_2824);
nand U3137 (N_3137,In_735,In_1939);
nor U3138 (N_3138,In_1631,In_2288);
or U3139 (N_3139,In_933,In_1722);
or U3140 (N_3140,In_1929,In_579);
nand U3141 (N_3141,In_19,In_1606);
and U3142 (N_3142,In_719,In_2757);
nor U3143 (N_3143,In_54,In_272);
or U3144 (N_3144,In_2815,In_2784);
and U3145 (N_3145,In_45,In_1816);
nor U3146 (N_3146,In_1620,In_353);
nand U3147 (N_3147,In_800,In_1003);
or U3148 (N_3148,In_996,In_2726);
nand U3149 (N_3149,In_2023,In_1028);
nand U3150 (N_3150,In_852,In_812);
nor U3151 (N_3151,In_492,In_1457);
or U3152 (N_3152,In_2940,In_2863);
and U3153 (N_3153,In_2477,In_354);
and U3154 (N_3154,In_2659,In_2700);
and U3155 (N_3155,In_1821,In_1437);
nand U3156 (N_3156,In_2611,In_1175);
or U3157 (N_3157,In_1037,In_806);
or U3158 (N_3158,In_23,In_1739);
nor U3159 (N_3159,In_1853,In_2738);
nor U3160 (N_3160,In_755,In_835);
nand U3161 (N_3161,In_1464,In_949);
nor U3162 (N_3162,In_1982,In_2894);
and U3163 (N_3163,In_1509,In_2309);
or U3164 (N_3164,In_1289,In_682);
xor U3165 (N_3165,In_2402,In_126);
or U3166 (N_3166,In_1024,In_2661);
xnor U3167 (N_3167,In_83,In_1744);
nand U3168 (N_3168,In_1632,In_2757);
nor U3169 (N_3169,In_2568,In_455);
nand U3170 (N_3170,In_1942,In_819);
nand U3171 (N_3171,In_24,In_111);
nand U3172 (N_3172,In_1392,In_2939);
and U3173 (N_3173,In_1449,In_845);
nand U3174 (N_3174,In_2928,In_2873);
nand U3175 (N_3175,In_2931,In_1816);
or U3176 (N_3176,In_2860,In_2203);
nand U3177 (N_3177,In_1223,In_40);
nand U3178 (N_3178,In_293,In_1699);
xor U3179 (N_3179,In_476,In_2574);
xor U3180 (N_3180,In_2128,In_46);
or U3181 (N_3181,In_770,In_91);
nand U3182 (N_3182,In_2385,In_291);
nand U3183 (N_3183,In_2340,In_2315);
nor U3184 (N_3184,In_2166,In_1164);
xnor U3185 (N_3185,In_2358,In_2144);
or U3186 (N_3186,In_2405,In_2885);
nand U3187 (N_3187,In_1649,In_555);
nor U3188 (N_3188,In_502,In_1491);
or U3189 (N_3189,In_1112,In_1188);
nand U3190 (N_3190,In_2015,In_2581);
nor U3191 (N_3191,In_1639,In_785);
or U3192 (N_3192,In_1597,In_2571);
nor U3193 (N_3193,In_2389,In_2538);
nor U3194 (N_3194,In_1173,In_2723);
nor U3195 (N_3195,In_969,In_1414);
nand U3196 (N_3196,In_1818,In_959);
nand U3197 (N_3197,In_655,In_2705);
nor U3198 (N_3198,In_1701,In_962);
and U3199 (N_3199,In_141,In_598);
nor U3200 (N_3200,In_2190,In_1721);
nor U3201 (N_3201,In_1457,In_1661);
or U3202 (N_3202,In_667,In_1643);
nor U3203 (N_3203,In_1297,In_2073);
or U3204 (N_3204,In_2255,In_2372);
and U3205 (N_3205,In_399,In_1980);
nor U3206 (N_3206,In_2524,In_1394);
or U3207 (N_3207,In_2436,In_1322);
or U3208 (N_3208,In_212,In_156);
or U3209 (N_3209,In_2431,In_796);
xnor U3210 (N_3210,In_67,In_2046);
nand U3211 (N_3211,In_2422,In_1424);
or U3212 (N_3212,In_136,In_1208);
and U3213 (N_3213,In_527,In_652);
nand U3214 (N_3214,In_2552,In_2063);
xor U3215 (N_3215,In_26,In_2217);
and U3216 (N_3216,In_2328,In_2325);
and U3217 (N_3217,In_1914,In_1027);
xor U3218 (N_3218,In_2222,In_1571);
nor U3219 (N_3219,In_658,In_437);
nand U3220 (N_3220,In_1987,In_325);
nand U3221 (N_3221,In_2702,In_32);
nor U3222 (N_3222,In_2037,In_1137);
or U3223 (N_3223,In_2888,In_492);
and U3224 (N_3224,In_715,In_678);
xor U3225 (N_3225,In_2087,In_553);
or U3226 (N_3226,In_701,In_2936);
and U3227 (N_3227,In_2832,In_2493);
and U3228 (N_3228,In_1565,In_2047);
nor U3229 (N_3229,In_824,In_284);
xnor U3230 (N_3230,In_2602,In_2305);
xor U3231 (N_3231,In_870,In_426);
and U3232 (N_3232,In_511,In_2412);
or U3233 (N_3233,In_2807,In_2038);
nor U3234 (N_3234,In_101,In_2355);
nor U3235 (N_3235,In_1178,In_519);
nor U3236 (N_3236,In_1737,In_357);
and U3237 (N_3237,In_1734,In_2853);
or U3238 (N_3238,In_2014,In_810);
nor U3239 (N_3239,In_2371,In_1041);
or U3240 (N_3240,In_189,In_2426);
nor U3241 (N_3241,In_1618,In_2485);
or U3242 (N_3242,In_1508,In_1193);
nand U3243 (N_3243,In_1933,In_2341);
and U3244 (N_3244,In_2730,In_606);
nor U3245 (N_3245,In_741,In_877);
or U3246 (N_3246,In_702,In_387);
nor U3247 (N_3247,In_1035,In_1795);
or U3248 (N_3248,In_2360,In_553);
or U3249 (N_3249,In_2263,In_2692);
or U3250 (N_3250,In_774,In_278);
xor U3251 (N_3251,In_2474,In_2128);
nor U3252 (N_3252,In_2881,In_1042);
and U3253 (N_3253,In_2380,In_2807);
and U3254 (N_3254,In_2079,In_1674);
nand U3255 (N_3255,In_2,In_1708);
nand U3256 (N_3256,In_1749,In_519);
or U3257 (N_3257,In_2160,In_1486);
nand U3258 (N_3258,In_2167,In_229);
nand U3259 (N_3259,In_2750,In_816);
nand U3260 (N_3260,In_1808,In_2455);
or U3261 (N_3261,In_1016,In_130);
nor U3262 (N_3262,In_2502,In_728);
nor U3263 (N_3263,In_1339,In_1723);
nor U3264 (N_3264,In_1099,In_371);
and U3265 (N_3265,In_1835,In_2162);
nor U3266 (N_3266,In_1757,In_1761);
nor U3267 (N_3267,In_2919,In_2844);
or U3268 (N_3268,In_1933,In_729);
and U3269 (N_3269,In_479,In_1163);
or U3270 (N_3270,In_1677,In_2749);
or U3271 (N_3271,In_1807,In_2074);
nand U3272 (N_3272,In_1738,In_1722);
nor U3273 (N_3273,In_2439,In_448);
and U3274 (N_3274,In_395,In_2186);
and U3275 (N_3275,In_1672,In_650);
xor U3276 (N_3276,In_10,In_2893);
and U3277 (N_3277,In_1884,In_234);
and U3278 (N_3278,In_2830,In_1074);
nand U3279 (N_3279,In_2177,In_88);
and U3280 (N_3280,In_2888,In_2178);
nand U3281 (N_3281,In_1891,In_1869);
nand U3282 (N_3282,In_1442,In_1996);
xor U3283 (N_3283,In_1779,In_1641);
nor U3284 (N_3284,In_181,In_2023);
nand U3285 (N_3285,In_695,In_321);
or U3286 (N_3286,In_292,In_630);
and U3287 (N_3287,In_2530,In_412);
xor U3288 (N_3288,In_172,In_613);
nor U3289 (N_3289,In_1296,In_1850);
or U3290 (N_3290,In_1143,In_955);
nor U3291 (N_3291,In_2141,In_726);
nor U3292 (N_3292,In_803,In_619);
or U3293 (N_3293,In_29,In_2595);
nand U3294 (N_3294,In_629,In_264);
or U3295 (N_3295,In_2635,In_1327);
and U3296 (N_3296,In_2822,In_2720);
and U3297 (N_3297,In_2141,In_1020);
nor U3298 (N_3298,In_2423,In_2594);
and U3299 (N_3299,In_221,In_625);
or U3300 (N_3300,In_372,In_1609);
nand U3301 (N_3301,In_1448,In_1517);
and U3302 (N_3302,In_1766,In_700);
nand U3303 (N_3303,In_2780,In_1100);
nor U3304 (N_3304,In_28,In_2646);
and U3305 (N_3305,In_1192,In_1437);
nor U3306 (N_3306,In_628,In_810);
and U3307 (N_3307,In_2838,In_734);
or U3308 (N_3308,In_1689,In_2989);
xnor U3309 (N_3309,In_378,In_1646);
nor U3310 (N_3310,In_2682,In_791);
nand U3311 (N_3311,In_2025,In_2200);
and U3312 (N_3312,In_2741,In_1840);
nand U3313 (N_3313,In_969,In_2095);
nor U3314 (N_3314,In_289,In_2);
and U3315 (N_3315,In_632,In_1276);
xor U3316 (N_3316,In_2517,In_1256);
nor U3317 (N_3317,In_2970,In_2025);
and U3318 (N_3318,In_2496,In_2063);
or U3319 (N_3319,In_2716,In_1143);
nand U3320 (N_3320,In_202,In_520);
and U3321 (N_3321,In_367,In_2644);
or U3322 (N_3322,In_340,In_2906);
and U3323 (N_3323,In_85,In_1241);
xor U3324 (N_3324,In_2263,In_1733);
and U3325 (N_3325,In_2152,In_2383);
xor U3326 (N_3326,In_782,In_2415);
and U3327 (N_3327,In_2740,In_592);
nand U3328 (N_3328,In_1171,In_985);
nor U3329 (N_3329,In_702,In_1916);
nand U3330 (N_3330,In_0,In_754);
and U3331 (N_3331,In_582,In_167);
nor U3332 (N_3332,In_1227,In_2455);
xor U3333 (N_3333,In_658,In_330);
or U3334 (N_3334,In_2702,In_1036);
nor U3335 (N_3335,In_733,In_2207);
nand U3336 (N_3336,In_2807,In_1373);
xnor U3337 (N_3337,In_112,In_711);
nand U3338 (N_3338,In_933,In_1261);
nor U3339 (N_3339,In_2579,In_1516);
nor U3340 (N_3340,In_1428,In_996);
or U3341 (N_3341,In_2233,In_1718);
xor U3342 (N_3342,In_2374,In_455);
or U3343 (N_3343,In_2335,In_445);
nand U3344 (N_3344,In_40,In_1896);
and U3345 (N_3345,In_1034,In_741);
and U3346 (N_3346,In_2374,In_744);
and U3347 (N_3347,In_225,In_1018);
nand U3348 (N_3348,In_1019,In_484);
or U3349 (N_3349,In_2233,In_2248);
or U3350 (N_3350,In_734,In_609);
or U3351 (N_3351,In_2453,In_1426);
and U3352 (N_3352,In_301,In_1097);
xor U3353 (N_3353,In_2661,In_2342);
and U3354 (N_3354,In_1835,In_1464);
and U3355 (N_3355,In_481,In_1186);
and U3356 (N_3356,In_1164,In_1889);
nor U3357 (N_3357,In_143,In_1586);
xor U3358 (N_3358,In_183,In_1361);
nor U3359 (N_3359,In_347,In_2381);
and U3360 (N_3360,In_2595,In_535);
or U3361 (N_3361,In_1470,In_454);
nand U3362 (N_3362,In_1404,In_163);
nand U3363 (N_3363,In_2679,In_2384);
or U3364 (N_3364,In_2349,In_2894);
nand U3365 (N_3365,In_234,In_2241);
and U3366 (N_3366,In_2979,In_403);
and U3367 (N_3367,In_113,In_1417);
and U3368 (N_3368,In_341,In_264);
nand U3369 (N_3369,In_2002,In_1078);
nand U3370 (N_3370,In_2430,In_546);
nand U3371 (N_3371,In_2610,In_2549);
nor U3372 (N_3372,In_810,In_1555);
and U3373 (N_3373,In_1464,In_72);
nand U3374 (N_3374,In_2840,In_1335);
or U3375 (N_3375,In_2166,In_453);
and U3376 (N_3376,In_657,In_437);
or U3377 (N_3377,In_1443,In_1367);
and U3378 (N_3378,In_1994,In_2782);
and U3379 (N_3379,In_2680,In_2072);
nor U3380 (N_3380,In_1713,In_1324);
xor U3381 (N_3381,In_2185,In_2168);
and U3382 (N_3382,In_1707,In_1243);
nand U3383 (N_3383,In_1212,In_2130);
and U3384 (N_3384,In_2567,In_2126);
nand U3385 (N_3385,In_1313,In_544);
or U3386 (N_3386,In_667,In_989);
nor U3387 (N_3387,In_1821,In_2914);
nand U3388 (N_3388,In_1271,In_440);
nor U3389 (N_3389,In_975,In_1540);
nor U3390 (N_3390,In_770,In_1109);
nor U3391 (N_3391,In_1863,In_1369);
and U3392 (N_3392,In_2882,In_2875);
nor U3393 (N_3393,In_2346,In_450);
nand U3394 (N_3394,In_1542,In_1113);
nand U3395 (N_3395,In_1417,In_2647);
nor U3396 (N_3396,In_2241,In_2501);
and U3397 (N_3397,In_1115,In_2128);
nor U3398 (N_3398,In_2115,In_1379);
nor U3399 (N_3399,In_236,In_2641);
xnor U3400 (N_3400,In_2491,In_499);
xor U3401 (N_3401,In_236,In_1796);
nor U3402 (N_3402,In_2115,In_1410);
nor U3403 (N_3403,In_2235,In_589);
or U3404 (N_3404,In_2940,In_848);
nand U3405 (N_3405,In_1485,In_1662);
and U3406 (N_3406,In_1240,In_1233);
nand U3407 (N_3407,In_753,In_2973);
nor U3408 (N_3408,In_872,In_23);
and U3409 (N_3409,In_2192,In_2975);
nor U3410 (N_3410,In_2721,In_1894);
and U3411 (N_3411,In_159,In_1308);
nand U3412 (N_3412,In_1155,In_2806);
nor U3413 (N_3413,In_88,In_1689);
nand U3414 (N_3414,In_1303,In_1668);
or U3415 (N_3415,In_716,In_1748);
nor U3416 (N_3416,In_2024,In_862);
nand U3417 (N_3417,In_565,In_2949);
nand U3418 (N_3418,In_2422,In_2200);
or U3419 (N_3419,In_2462,In_1718);
or U3420 (N_3420,In_2476,In_1535);
or U3421 (N_3421,In_403,In_902);
or U3422 (N_3422,In_1639,In_188);
and U3423 (N_3423,In_2539,In_75);
and U3424 (N_3424,In_1323,In_2816);
nor U3425 (N_3425,In_2776,In_966);
nand U3426 (N_3426,In_1445,In_2001);
and U3427 (N_3427,In_1824,In_2346);
nand U3428 (N_3428,In_2411,In_1972);
or U3429 (N_3429,In_1439,In_1604);
nor U3430 (N_3430,In_538,In_830);
or U3431 (N_3431,In_582,In_1806);
nand U3432 (N_3432,In_1193,In_1855);
nand U3433 (N_3433,In_2605,In_20);
and U3434 (N_3434,In_97,In_1978);
xnor U3435 (N_3435,In_1165,In_445);
nor U3436 (N_3436,In_549,In_1458);
nand U3437 (N_3437,In_1952,In_1206);
or U3438 (N_3438,In_1152,In_710);
nand U3439 (N_3439,In_1526,In_2630);
and U3440 (N_3440,In_2196,In_951);
or U3441 (N_3441,In_2549,In_1459);
nor U3442 (N_3442,In_562,In_2025);
xor U3443 (N_3443,In_269,In_497);
xnor U3444 (N_3444,In_925,In_586);
nor U3445 (N_3445,In_928,In_2346);
nor U3446 (N_3446,In_1607,In_2705);
or U3447 (N_3447,In_753,In_2453);
nand U3448 (N_3448,In_2770,In_697);
nor U3449 (N_3449,In_2881,In_2655);
nand U3450 (N_3450,In_1160,In_1297);
nor U3451 (N_3451,In_1742,In_1489);
and U3452 (N_3452,In_611,In_2416);
nand U3453 (N_3453,In_860,In_151);
or U3454 (N_3454,In_158,In_91);
nor U3455 (N_3455,In_1626,In_449);
xnor U3456 (N_3456,In_1527,In_14);
or U3457 (N_3457,In_2772,In_2575);
nand U3458 (N_3458,In_644,In_2510);
and U3459 (N_3459,In_1270,In_2819);
nand U3460 (N_3460,In_914,In_248);
nor U3461 (N_3461,In_1087,In_2686);
nor U3462 (N_3462,In_2605,In_997);
nor U3463 (N_3463,In_780,In_658);
and U3464 (N_3464,In_231,In_448);
nor U3465 (N_3465,In_895,In_2975);
nor U3466 (N_3466,In_50,In_2057);
nand U3467 (N_3467,In_687,In_2075);
or U3468 (N_3468,In_1482,In_2789);
and U3469 (N_3469,In_906,In_1236);
and U3470 (N_3470,In_1278,In_514);
and U3471 (N_3471,In_2523,In_1509);
and U3472 (N_3472,In_2795,In_452);
and U3473 (N_3473,In_260,In_2018);
and U3474 (N_3474,In_2395,In_1728);
nand U3475 (N_3475,In_632,In_757);
nor U3476 (N_3476,In_643,In_718);
or U3477 (N_3477,In_2842,In_1897);
nand U3478 (N_3478,In_1593,In_783);
nand U3479 (N_3479,In_428,In_275);
or U3480 (N_3480,In_2278,In_1189);
and U3481 (N_3481,In_2336,In_1569);
nor U3482 (N_3482,In_2241,In_2459);
nand U3483 (N_3483,In_2785,In_1566);
and U3484 (N_3484,In_391,In_53);
or U3485 (N_3485,In_2410,In_1107);
and U3486 (N_3486,In_1449,In_1403);
nor U3487 (N_3487,In_2244,In_2125);
xnor U3488 (N_3488,In_1451,In_526);
nor U3489 (N_3489,In_2166,In_2569);
and U3490 (N_3490,In_1389,In_1879);
nor U3491 (N_3491,In_1340,In_2770);
and U3492 (N_3492,In_2707,In_2456);
or U3493 (N_3493,In_1812,In_1172);
nor U3494 (N_3494,In_2316,In_1953);
nand U3495 (N_3495,In_1059,In_1280);
xor U3496 (N_3496,In_1600,In_1669);
nand U3497 (N_3497,In_2196,In_2067);
and U3498 (N_3498,In_2276,In_829);
nor U3499 (N_3499,In_1679,In_2802);
nor U3500 (N_3500,In_165,In_2268);
nand U3501 (N_3501,In_1828,In_581);
or U3502 (N_3502,In_2092,In_1583);
nand U3503 (N_3503,In_2502,In_1649);
nor U3504 (N_3504,In_978,In_103);
xor U3505 (N_3505,In_1898,In_2630);
nand U3506 (N_3506,In_1265,In_777);
or U3507 (N_3507,In_1264,In_1021);
and U3508 (N_3508,In_2222,In_811);
nor U3509 (N_3509,In_1497,In_1572);
nor U3510 (N_3510,In_2918,In_853);
or U3511 (N_3511,In_1943,In_2072);
or U3512 (N_3512,In_2473,In_333);
nor U3513 (N_3513,In_2921,In_2418);
or U3514 (N_3514,In_2045,In_2730);
and U3515 (N_3515,In_35,In_67);
nand U3516 (N_3516,In_7,In_2283);
nor U3517 (N_3517,In_299,In_2209);
nand U3518 (N_3518,In_1861,In_1646);
nor U3519 (N_3519,In_1912,In_2230);
nor U3520 (N_3520,In_2729,In_1454);
xnor U3521 (N_3521,In_2158,In_2886);
nand U3522 (N_3522,In_3,In_2318);
xnor U3523 (N_3523,In_1257,In_50);
nand U3524 (N_3524,In_104,In_595);
and U3525 (N_3525,In_471,In_450);
nand U3526 (N_3526,In_2969,In_839);
and U3527 (N_3527,In_1456,In_1637);
or U3528 (N_3528,In_668,In_554);
or U3529 (N_3529,In_530,In_776);
and U3530 (N_3530,In_2298,In_2032);
xnor U3531 (N_3531,In_1450,In_2716);
or U3532 (N_3532,In_2996,In_2251);
and U3533 (N_3533,In_2265,In_2500);
or U3534 (N_3534,In_973,In_762);
and U3535 (N_3535,In_1277,In_1994);
and U3536 (N_3536,In_1429,In_2309);
nand U3537 (N_3537,In_953,In_2916);
nor U3538 (N_3538,In_304,In_2981);
or U3539 (N_3539,In_2723,In_2099);
and U3540 (N_3540,In_136,In_1151);
nand U3541 (N_3541,In_920,In_712);
or U3542 (N_3542,In_1382,In_28);
or U3543 (N_3543,In_1126,In_386);
nor U3544 (N_3544,In_2633,In_2594);
xor U3545 (N_3545,In_477,In_850);
nor U3546 (N_3546,In_225,In_1984);
nand U3547 (N_3547,In_520,In_1074);
or U3548 (N_3548,In_849,In_1860);
nand U3549 (N_3549,In_2008,In_2583);
and U3550 (N_3550,In_126,In_450);
and U3551 (N_3551,In_2132,In_1008);
and U3552 (N_3552,In_881,In_2494);
or U3553 (N_3553,In_1383,In_152);
or U3554 (N_3554,In_1935,In_2821);
nand U3555 (N_3555,In_920,In_201);
and U3556 (N_3556,In_1990,In_1835);
nand U3557 (N_3557,In_277,In_907);
nand U3558 (N_3558,In_1576,In_1029);
nand U3559 (N_3559,In_2015,In_1367);
nor U3560 (N_3560,In_1963,In_2540);
and U3561 (N_3561,In_2133,In_1341);
or U3562 (N_3562,In_1316,In_2106);
and U3563 (N_3563,In_100,In_2852);
and U3564 (N_3564,In_932,In_728);
nor U3565 (N_3565,In_1282,In_2844);
and U3566 (N_3566,In_958,In_1573);
or U3567 (N_3567,In_63,In_2476);
or U3568 (N_3568,In_2273,In_649);
nand U3569 (N_3569,In_1256,In_1227);
nand U3570 (N_3570,In_257,In_642);
nor U3571 (N_3571,In_2885,In_438);
and U3572 (N_3572,In_2244,In_2520);
or U3573 (N_3573,In_2558,In_1395);
nor U3574 (N_3574,In_2420,In_905);
or U3575 (N_3575,In_2326,In_1675);
nand U3576 (N_3576,In_1367,In_2993);
xor U3577 (N_3577,In_1725,In_77);
nor U3578 (N_3578,In_2635,In_2400);
nor U3579 (N_3579,In_2440,In_892);
xor U3580 (N_3580,In_445,In_2995);
and U3581 (N_3581,In_1612,In_299);
xnor U3582 (N_3582,In_1767,In_496);
nor U3583 (N_3583,In_267,In_1931);
and U3584 (N_3584,In_151,In_167);
and U3585 (N_3585,In_153,In_1311);
or U3586 (N_3586,In_2913,In_2140);
nand U3587 (N_3587,In_1034,In_2273);
or U3588 (N_3588,In_1947,In_654);
nor U3589 (N_3589,In_1822,In_1716);
or U3590 (N_3590,In_2791,In_1792);
nor U3591 (N_3591,In_2267,In_78);
nor U3592 (N_3592,In_2087,In_1912);
nand U3593 (N_3593,In_2068,In_702);
or U3594 (N_3594,In_2476,In_1696);
nand U3595 (N_3595,In_538,In_2643);
or U3596 (N_3596,In_474,In_91);
or U3597 (N_3597,In_1669,In_2066);
nor U3598 (N_3598,In_2678,In_1420);
or U3599 (N_3599,In_2389,In_2076);
nand U3600 (N_3600,In_1686,In_783);
nand U3601 (N_3601,In_2931,In_2726);
nand U3602 (N_3602,In_1791,In_570);
xor U3603 (N_3603,In_1769,In_2572);
xor U3604 (N_3604,In_2959,In_1777);
nor U3605 (N_3605,In_1089,In_767);
nand U3606 (N_3606,In_1677,In_2820);
and U3607 (N_3607,In_480,In_25);
nor U3608 (N_3608,In_2209,In_759);
nor U3609 (N_3609,In_1277,In_1860);
and U3610 (N_3610,In_2539,In_2309);
xor U3611 (N_3611,In_2712,In_1193);
nor U3612 (N_3612,In_1729,In_187);
nand U3613 (N_3613,In_496,In_2474);
nor U3614 (N_3614,In_2635,In_2973);
or U3615 (N_3615,In_845,In_1891);
xor U3616 (N_3616,In_2881,In_2299);
and U3617 (N_3617,In_1203,In_2521);
nor U3618 (N_3618,In_2621,In_315);
nor U3619 (N_3619,In_1988,In_1668);
or U3620 (N_3620,In_535,In_1980);
or U3621 (N_3621,In_2069,In_1633);
nor U3622 (N_3622,In_2912,In_566);
and U3623 (N_3623,In_1467,In_1985);
nor U3624 (N_3624,In_405,In_655);
and U3625 (N_3625,In_2339,In_1144);
and U3626 (N_3626,In_1060,In_94);
nand U3627 (N_3627,In_14,In_2985);
and U3628 (N_3628,In_1636,In_2269);
nor U3629 (N_3629,In_2063,In_2557);
xor U3630 (N_3630,In_2634,In_2705);
and U3631 (N_3631,In_1067,In_593);
and U3632 (N_3632,In_2615,In_1861);
or U3633 (N_3633,In_2166,In_2973);
nor U3634 (N_3634,In_2814,In_2884);
and U3635 (N_3635,In_1625,In_2170);
or U3636 (N_3636,In_831,In_2695);
and U3637 (N_3637,In_496,In_666);
and U3638 (N_3638,In_2765,In_891);
nor U3639 (N_3639,In_1359,In_443);
or U3640 (N_3640,In_2913,In_2318);
nand U3641 (N_3641,In_2555,In_2986);
nand U3642 (N_3642,In_1380,In_1701);
and U3643 (N_3643,In_2185,In_1174);
or U3644 (N_3644,In_797,In_2449);
nor U3645 (N_3645,In_2827,In_1106);
and U3646 (N_3646,In_290,In_1848);
nand U3647 (N_3647,In_315,In_1548);
nand U3648 (N_3648,In_1848,In_1089);
nand U3649 (N_3649,In_1254,In_1663);
or U3650 (N_3650,In_2495,In_2424);
nor U3651 (N_3651,In_2382,In_2097);
and U3652 (N_3652,In_2398,In_128);
xor U3653 (N_3653,In_1976,In_1353);
and U3654 (N_3654,In_310,In_1090);
nor U3655 (N_3655,In_1813,In_2923);
or U3656 (N_3656,In_1432,In_563);
nor U3657 (N_3657,In_1438,In_1713);
nand U3658 (N_3658,In_2590,In_2170);
nand U3659 (N_3659,In_1883,In_2939);
or U3660 (N_3660,In_177,In_1250);
nor U3661 (N_3661,In_1900,In_613);
nand U3662 (N_3662,In_2791,In_151);
or U3663 (N_3663,In_2381,In_731);
nand U3664 (N_3664,In_2104,In_2316);
and U3665 (N_3665,In_2360,In_1884);
nor U3666 (N_3666,In_2988,In_369);
nor U3667 (N_3667,In_1832,In_2662);
and U3668 (N_3668,In_389,In_30);
nand U3669 (N_3669,In_2091,In_1483);
nor U3670 (N_3670,In_2233,In_1640);
nor U3671 (N_3671,In_2972,In_1866);
and U3672 (N_3672,In_2274,In_2178);
and U3673 (N_3673,In_718,In_178);
or U3674 (N_3674,In_573,In_2077);
nor U3675 (N_3675,In_83,In_888);
or U3676 (N_3676,In_2203,In_2427);
nand U3677 (N_3677,In_1373,In_50);
nor U3678 (N_3678,In_2121,In_740);
nor U3679 (N_3679,In_1631,In_2112);
and U3680 (N_3680,In_2461,In_2680);
or U3681 (N_3681,In_1499,In_2177);
nand U3682 (N_3682,In_2172,In_1871);
nor U3683 (N_3683,In_741,In_759);
or U3684 (N_3684,In_1849,In_1156);
nor U3685 (N_3685,In_1537,In_2330);
nand U3686 (N_3686,In_2814,In_1542);
or U3687 (N_3687,In_1927,In_1338);
nand U3688 (N_3688,In_1907,In_846);
xnor U3689 (N_3689,In_1376,In_577);
or U3690 (N_3690,In_2210,In_2317);
xnor U3691 (N_3691,In_1350,In_1573);
xor U3692 (N_3692,In_1460,In_1911);
and U3693 (N_3693,In_693,In_1532);
xnor U3694 (N_3694,In_1178,In_1857);
nand U3695 (N_3695,In_2519,In_258);
or U3696 (N_3696,In_2017,In_1034);
nor U3697 (N_3697,In_2670,In_1485);
nor U3698 (N_3698,In_256,In_613);
nand U3699 (N_3699,In_2861,In_977);
or U3700 (N_3700,In_1521,In_787);
nor U3701 (N_3701,In_1328,In_284);
and U3702 (N_3702,In_438,In_2447);
and U3703 (N_3703,In_1988,In_335);
or U3704 (N_3704,In_2853,In_1713);
xnor U3705 (N_3705,In_1808,In_2237);
nand U3706 (N_3706,In_1307,In_2553);
nor U3707 (N_3707,In_746,In_1313);
nand U3708 (N_3708,In_2917,In_2979);
and U3709 (N_3709,In_87,In_107);
or U3710 (N_3710,In_1442,In_203);
nand U3711 (N_3711,In_2297,In_1670);
and U3712 (N_3712,In_170,In_1130);
nor U3713 (N_3713,In_4,In_837);
nor U3714 (N_3714,In_2492,In_1076);
or U3715 (N_3715,In_1532,In_1355);
nand U3716 (N_3716,In_517,In_2001);
or U3717 (N_3717,In_2578,In_2555);
and U3718 (N_3718,In_2323,In_1673);
nor U3719 (N_3719,In_1516,In_1351);
and U3720 (N_3720,In_518,In_311);
nor U3721 (N_3721,In_1541,In_140);
xor U3722 (N_3722,In_1661,In_1025);
nor U3723 (N_3723,In_1988,In_2361);
xor U3724 (N_3724,In_1473,In_2957);
nor U3725 (N_3725,In_691,In_166);
nand U3726 (N_3726,In_1813,In_1711);
nor U3727 (N_3727,In_1166,In_2603);
or U3728 (N_3728,In_1077,In_2039);
and U3729 (N_3729,In_586,In_1144);
nor U3730 (N_3730,In_2547,In_2722);
nand U3731 (N_3731,In_135,In_991);
nand U3732 (N_3732,In_830,In_924);
nand U3733 (N_3733,In_2211,In_71);
nand U3734 (N_3734,In_1431,In_653);
and U3735 (N_3735,In_1993,In_457);
or U3736 (N_3736,In_1576,In_2749);
and U3737 (N_3737,In_359,In_2295);
or U3738 (N_3738,In_1036,In_1018);
nand U3739 (N_3739,In_574,In_2688);
or U3740 (N_3740,In_639,In_236);
nand U3741 (N_3741,In_2702,In_786);
or U3742 (N_3742,In_740,In_805);
nor U3743 (N_3743,In_35,In_869);
nand U3744 (N_3744,In_2269,In_1222);
nor U3745 (N_3745,In_840,In_982);
and U3746 (N_3746,In_1920,In_1121);
or U3747 (N_3747,In_1342,In_2160);
nand U3748 (N_3748,In_293,In_2328);
and U3749 (N_3749,In_783,In_508);
nand U3750 (N_3750,In_2817,In_2025);
or U3751 (N_3751,In_2111,In_281);
nand U3752 (N_3752,In_1702,In_1034);
and U3753 (N_3753,In_2217,In_16);
nand U3754 (N_3754,In_97,In_855);
xor U3755 (N_3755,In_690,In_810);
nor U3756 (N_3756,In_2114,In_1325);
or U3757 (N_3757,In_1505,In_602);
xor U3758 (N_3758,In_1943,In_448);
xor U3759 (N_3759,In_1413,In_2510);
xor U3760 (N_3760,In_1653,In_1991);
nor U3761 (N_3761,In_853,In_336);
or U3762 (N_3762,In_531,In_2410);
or U3763 (N_3763,In_757,In_421);
nand U3764 (N_3764,In_2938,In_2124);
and U3765 (N_3765,In_1000,In_1577);
or U3766 (N_3766,In_1182,In_538);
xnor U3767 (N_3767,In_470,In_1271);
nor U3768 (N_3768,In_420,In_1351);
nand U3769 (N_3769,In_381,In_597);
nand U3770 (N_3770,In_1735,In_2477);
xnor U3771 (N_3771,In_1203,In_2950);
and U3772 (N_3772,In_1796,In_1588);
xnor U3773 (N_3773,In_2138,In_599);
and U3774 (N_3774,In_736,In_2606);
and U3775 (N_3775,In_26,In_1061);
and U3776 (N_3776,In_1217,In_2089);
nand U3777 (N_3777,In_1297,In_2416);
xor U3778 (N_3778,In_2697,In_2779);
or U3779 (N_3779,In_562,In_146);
nor U3780 (N_3780,In_2986,In_1556);
or U3781 (N_3781,In_2163,In_2376);
or U3782 (N_3782,In_1650,In_1088);
xor U3783 (N_3783,In_593,In_1929);
nor U3784 (N_3784,In_2638,In_1375);
and U3785 (N_3785,In_230,In_1386);
xor U3786 (N_3786,In_2032,In_210);
xnor U3787 (N_3787,In_1373,In_1143);
and U3788 (N_3788,In_2733,In_2925);
or U3789 (N_3789,In_367,In_2743);
nor U3790 (N_3790,In_2356,In_2898);
nor U3791 (N_3791,In_2117,In_1119);
and U3792 (N_3792,In_2273,In_1997);
nor U3793 (N_3793,In_2080,In_132);
or U3794 (N_3794,In_664,In_2612);
nor U3795 (N_3795,In_1810,In_94);
nor U3796 (N_3796,In_928,In_372);
nand U3797 (N_3797,In_889,In_1186);
nand U3798 (N_3798,In_2255,In_627);
nor U3799 (N_3799,In_48,In_1890);
or U3800 (N_3800,In_200,In_2772);
and U3801 (N_3801,In_2966,In_1948);
nand U3802 (N_3802,In_2332,In_2359);
and U3803 (N_3803,In_1555,In_122);
nand U3804 (N_3804,In_2514,In_1092);
or U3805 (N_3805,In_1550,In_1789);
nor U3806 (N_3806,In_1221,In_1902);
and U3807 (N_3807,In_2034,In_1869);
or U3808 (N_3808,In_781,In_1413);
nand U3809 (N_3809,In_705,In_5);
and U3810 (N_3810,In_250,In_2416);
xor U3811 (N_3811,In_2461,In_1635);
xnor U3812 (N_3812,In_2375,In_1132);
and U3813 (N_3813,In_2981,In_1113);
nand U3814 (N_3814,In_2565,In_512);
nand U3815 (N_3815,In_2637,In_2592);
nand U3816 (N_3816,In_912,In_455);
and U3817 (N_3817,In_2886,In_1379);
or U3818 (N_3818,In_628,In_115);
or U3819 (N_3819,In_2090,In_2429);
nand U3820 (N_3820,In_782,In_2321);
nand U3821 (N_3821,In_1730,In_2033);
or U3822 (N_3822,In_22,In_2197);
nand U3823 (N_3823,In_1411,In_418);
xnor U3824 (N_3824,In_1108,In_2407);
and U3825 (N_3825,In_1973,In_2910);
or U3826 (N_3826,In_716,In_1890);
or U3827 (N_3827,In_485,In_815);
and U3828 (N_3828,In_1112,In_599);
and U3829 (N_3829,In_942,In_2013);
nor U3830 (N_3830,In_2215,In_2064);
and U3831 (N_3831,In_1345,In_1987);
xnor U3832 (N_3832,In_2670,In_1694);
or U3833 (N_3833,In_227,In_2397);
and U3834 (N_3834,In_774,In_1715);
and U3835 (N_3835,In_1549,In_1072);
or U3836 (N_3836,In_2986,In_2010);
and U3837 (N_3837,In_2576,In_1919);
and U3838 (N_3838,In_740,In_406);
nand U3839 (N_3839,In_979,In_2182);
nand U3840 (N_3840,In_1340,In_2733);
or U3841 (N_3841,In_830,In_1072);
nor U3842 (N_3842,In_958,In_1493);
or U3843 (N_3843,In_1146,In_481);
nand U3844 (N_3844,In_2946,In_2370);
or U3845 (N_3845,In_1095,In_305);
nor U3846 (N_3846,In_1660,In_85);
nor U3847 (N_3847,In_2668,In_1172);
and U3848 (N_3848,In_2373,In_705);
xnor U3849 (N_3849,In_1543,In_2118);
nand U3850 (N_3850,In_2356,In_1347);
xnor U3851 (N_3851,In_1243,In_189);
nand U3852 (N_3852,In_376,In_1435);
nand U3853 (N_3853,In_2446,In_152);
xor U3854 (N_3854,In_1964,In_666);
and U3855 (N_3855,In_1153,In_756);
or U3856 (N_3856,In_1344,In_1942);
and U3857 (N_3857,In_1192,In_277);
nor U3858 (N_3858,In_873,In_1565);
and U3859 (N_3859,In_1658,In_460);
xor U3860 (N_3860,In_2050,In_2524);
and U3861 (N_3861,In_1659,In_2395);
nor U3862 (N_3862,In_392,In_197);
nor U3863 (N_3863,In_2340,In_912);
and U3864 (N_3864,In_349,In_404);
nand U3865 (N_3865,In_1069,In_804);
or U3866 (N_3866,In_2103,In_1464);
nand U3867 (N_3867,In_1047,In_2594);
and U3868 (N_3868,In_2678,In_1746);
nor U3869 (N_3869,In_503,In_1605);
nor U3870 (N_3870,In_732,In_2182);
and U3871 (N_3871,In_1560,In_1338);
nand U3872 (N_3872,In_745,In_125);
xor U3873 (N_3873,In_2174,In_2447);
nand U3874 (N_3874,In_831,In_2506);
or U3875 (N_3875,In_1066,In_1094);
xor U3876 (N_3876,In_400,In_1910);
xnor U3877 (N_3877,In_1175,In_1626);
or U3878 (N_3878,In_301,In_2321);
xor U3879 (N_3879,In_914,In_2173);
nand U3880 (N_3880,In_1902,In_50);
or U3881 (N_3881,In_2548,In_2487);
or U3882 (N_3882,In_359,In_1027);
or U3883 (N_3883,In_2654,In_818);
xor U3884 (N_3884,In_522,In_397);
nor U3885 (N_3885,In_726,In_2918);
or U3886 (N_3886,In_607,In_2993);
nand U3887 (N_3887,In_1553,In_1743);
or U3888 (N_3888,In_1825,In_2426);
nor U3889 (N_3889,In_1493,In_1340);
nand U3890 (N_3890,In_831,In_1956);
or U3891 (N_3891,In_406,In_1743);
nor U3892 (N_3892,In_227,In_2027);
or U3893 (N_3893,In_894,In_763);
and U3894 (N_3894,In_2781,In_2855);
nand U3895 (N_3895,In_2638,In_2459);
nand U3896 (N_3896,In_2402,In_1562);
nor U3897 (N_3897,In_2720,In_1172);
xnor U3898 (N_3898,In_2958,In_2452);
and U3899 (N_3899,In_176,In_328);
xor U3900 (N_3900,In_625,In_251);
or U3901 (N_3901,In_2869,In_2951);
nor U3902 (N_3902,In_2980,In_176);
or U3903 (N_3903,In_2109,In_2542);
nor U3904 (N_3904,In_2709,In_497);
and U3905 (N_3905,In_1023,In_1759);
nand U3906 (N_3906,In_826,In_2376);
nor U3907 (N_3907,In_2449,In_423);
or U3908 (N_3908,In_2973,In_1024);
nor U3909 (N_3909,In_687,In_315);
nand U3910 (N_3910,In_2069,In_100);
nand U3911 (N_3911,In_2947,In_2024);
or U3912 (N_3912,In_2186,In_53);
and U3913 (N_3913,In_736,In_872);
nand U3914 (N_3914,In_708,In_1047);
nor U3915 (N_3915,In_2638,In_1419);
and U3916 (N_3916,In_2975,In_2633);
or U3917 (N_3917,In_1669,In_966);
nand U3918 (N_3918,In_2749,In_142);
or U3919 (N_3919,In_959,In_1812);
and U3920 (N_3920,In_1033,In_1298);
nor U3921 (N_3921,In_2085,In_52);
nor U3922 (N_3922,In_235,In_2207);
and U3923 (N_3923,In_1003,In_159);
and U3924 (N_3924,In_2136,In_1766);
or U3925 (N_3925,In_2705,In_2287);
and U3926 (N_3926,In_2322,In_2420);
nand U3927 (N_3927,In_27,In_2202);
nor U3928 (N_3928,In_1456,In_878);
and U3929 (N_3929,In_2759,In_2558);
and U3930 (N_3930,In_2508,In_2510);
or U3931 (N_3931,In_795,In_1679);
xor U3932 (N_3932,In_1432,In_1246);
and U3933 (N_3933,In_385,In_219);
or U3934 (N_3934,In_502,In_1142);
and U3935 (N_3935,In_532,In_1152);
nor U3936 (N_3936,In_1808,In_2597);
nand U3937 (N_3937,In_288,In_2276);
or U3938 (N_3938,In_1934,In_2441);
or U3939 (N_3939,In_1752,In_1341);
nand U3940 (N_3940,In_2444,In_1546);
and U3941 (N_3941,In_1866,In_2209);
nor U3942 (N_3942,In_2205,In_2751);
nand U3943 (N_3943,In_672,In_1805);
nor U3944 (N_3944,In_2464,In_2024);
or U3945 (N_3945,In_2392,In_1171);
nand U3946 (N_3946,In_1537,In_79);
nand U3947 (N_3947,In_436,In_428);
xnor U3948 (N_3948,In_1987,In_2408);
or U3949 (N_3949,In_751,In_2876);
xnor U3950 (N_3950,In_2140,In_594);
nor U3951 (N_3951,In_2017,In_2550);
nand U3952 (N_3952,In_2633,In_206);
xnor U3953 (N_3953,In_1665,In_2651);
and U3954 (N_3954,In_2875,In_1272);
and U3955 (N_3955,In_201,In_607);
and U3956 (N_3956,In_1749,In_1207);
and U3957 (N_3957,In_293,In_2973);
nor U3958 (N_3958,In_2422,In_2917);
nand U3959 (N_3959,In_2917,In_1328);
nor U3960 (N_3960,In_1262,In_1391);
or U3961 (N_3961,In_586,In_2737);
and U3962 (N_3962,In_47,In_601);
and U3963 (N_3963,In_1463,In_1956);
nor U3964 (N_3964,In_1988,In_133);
and U3965 (N_3965,In_691,In_116);
nor U3966 (N_3966,In_162,In_2151);
nor U3967 (N_3967,In_1371,In_1350);
xor U3968 (N_3968,In_2791,In_880);
and U3969 (N_3969,In_1714,In_1327);
nor U3970 (N_3970,In_532,In_2913);
and U3971 (N_3971,In_107,In_1069);
nor U3972 (N_3972,In_2290,In_1410);
nor U3973 (N_3973,In_90,In_2595);
xor U3974 (N_3974,In_573,In_438);
nand U3975 (N_3975,In_463,In_2391);
or U3976 (N_3976,In_422,In_1897);
and U3977 (N_3977,In_1456,In_345);
and U3978 (N_3978,In_2979,In_1951);
or U3979 (N_3979,In_2636,In_2766);
and U3980 (N_3980,In_1536,In_1260);
xor U3981 (N_3981,In_202,In_559);
or U3982 (N_3982,In_593,In_2078);
nand U3983 (N_3983,In_2894,In_2506);
xnor U3984 (N_3984,In_2369,In_675);
nor U3985 (N_3985,In_1476,In_912);
nor U3986 (N_3986,In_2679,In_45);
nand U3987 (N_3987,In_1427,In_110);
xnor U3988 (N_3988,In_201,In_721);
nand U3989 (N_3989,In_2021,In_2663);
or U3990 (N_3990,In_742,In_459);
or U3991 (N_3991,In_28,In_1655);
or U3992 (N_3992,In_952,In_166);
xnor U3993 (N_3993,In_1360,In_2867);
and U3994 (N_3994,In_2780,In_609);
nand U3995 (N_3995,In_2929,In_1979);
nand U3996 (N_3996,In_399,In_2643);
or U3997 (N_3997,In_495,In_2648);
or U3998 (N_3998,In_1988,In_9);
nor U3999 (N_3999,In_2348,In_2282);
nand U4000 (N_4000,In_750,In_2837);
nor U4001 (N_4001,In_1546,In_1680);
nor U4002 (N_4002,In_2896,In_2010);
or U4003 (N_4003,In_1026,In_2958);
xor U4004 (N_4004,In_30,In_829);
nand U4005 (N_4005,In_985,In_349);
nor U4006 (N_4006,In_1649,In_1560);
or U4007 (N_4007,In_388,In_809);
nand U4008 (N_4008,In_2452,In_1364);
nor U4009 (N_4009,In_1575,In_961);
nor U4010 (N_4010,In_827,In_1910);
xor U4011 (N_4011,In_1933,In_494);
nand U4012 (N_4012,In_2294,In_1011);
xor U4013 (N_4013,In_1881,In_2594);
nand U4014 (N_4014,In_2731,In_2596);
and U4015 (N_4015,In_1093,In_18);
or U4016 (N_4016,In_2525,In_259);
or U4017 (N_4017,In_347,In_890);
and U4018 (N_4018,In_1122,In_1458);
and U4019 (N_4019,In_969,In_3);
nor U4020 (N_4020,In_634,In_2571);
and U4021 (N_4021,In_1460,In_732);
or U4022 (N_4022,In_437,In_471);
nand U4023 (N_4023,In_406,In_2644);
nand U4024 (N_4024,In_421,In_1869);
nor U4025 (N_4025,In_2736,In_1901);
and U4026 (N_4026,In_2579,In_713);
and U4027 (N_4027,In_807,In_2700);
or U4028 (N_4028,In_702,In_2593);
xor U4029 (N_4029,In_2726,In_2552);
and U4030 (N_4030,In_1001,In_2310);
xnor U4031 (N_4031,In_2608,In_637);
nand U4032 (N_4032,In_2697,In_2463);
nand U4033 (N_4033,In_1798,In_280);
and U4034 (N_4034,In_2221,In_2883);
or U4035 (N_4035,In_2055,In_2083);
or U4036 (N_4036,In_2576,In_1181);
or U4037 (N_4037,In_624,In_2880);
nand U4038 (N_4038,In_759,In_26);
nand U4039 (N_4039,In_1581,In_756);
or U4040 (N_4040,In_1027,In_919);
nand U4041 (N_4041,In_1193,In_2931);
xor U4042 (N_4042,In_258,In_2341);
nand U4043 (N_4043,In_1910,In_2911);
nor U4044 (N_4044,In_2565,In_2198);
and U4045 (N_4045,In_1082,In_632);
nand U4046 (N_4046,In_1884,In_2290);
and U4047 (N_4047,In_1298,In_2220);
nand U4048 (N_4048,In_532,In_2929);
or U4049 (N_4049,In_60,In_677);
nor U4050 (N_4050,In_2161,In_828);
or U4051 (N_4051,In_622,In_2196);
xor U4052 (N_4052,In_2847,In_980);
nand U4053 (N_4053,In_2488,In_1069);
xor U4054 (N_4054,In_587,In_1082);
nand U4055 (N_4055,In_2353,In_206);
or U4056 (N_4056,In_2272,In_260);
nor U4057 (N_4057,In_2927,In_2079);
and U4058 (N_4058,In_2515,In_2902);
nor U4059 (N_4059,In_2277,In_2478);
nor U4060 (N_4060,In_888,In_1476);
or U4061 (N_4061,In_1228,In_883);
or U4062 (N_4062,In_1650,In_1968);
or U4063 (N_4063,In_2323,In_2043);
and U4064 (N_4064,In_1639,In_1886);
and U4065 (N_4065,In_187,In_730);
xnor U4066 (N_4066,In_1745,In_2621);
and U4067 (N_4067,In_2583,In_9);
or U4068 (N_4068,In_2091,In_2815);
xnor U4069 (N_4069,In_2387,In_2933);
xnor U4070 (N_4070,In_798,In_1143);
or U4071 (N_4071,In_809,In_1076);
nand U4072 (N_4072,In_1902,In_1411);
nand U4073 (N_4073,In_1031,In_2459);
nand U4074 (N_4074,In_2853,In_1546);
and U4075 (N_4075,In_2321,In_2882);
or U4076 (N_4076,In_498,In_916);
or U4077 (N_4077,In_1712,In_556);
and U4078 (N_4078,In_1692,In_1957);
or U4079 (N_4079,In_1271,In_1760);
and U4080 (N_4080,In_2470,In_767);
nand U4081 (N_4081,In_244,In_1492);
nor U4082 (N_4082,In_476,In_495);
nor U4083 (N_4083,In_1075,In_2158);
or U4084 (N_4084,In_2381,In_18);
nor U4085 (N_4085,In_1750,In_730);
nor U4086 (N_4086,In_1080,In_235);
nand U4087 (N_4087,In_677,In_621);
or U4088 (N_4088,In_75,In_2749);
nand U4089 (N_4089,In_1020,In_145);
nor U4090 (N_4090,In_1235,In_2498);
xor U4091 (N_4091,In_2088,In_2465);
nand U4092 (N_4092,In_2324,In_1955);
nand U4093 (N_4093,In_1537,In_2326);
nor U4094 (N_4094,In_2648,In_2150);
nand U4095 (N_4095,In_997,In_1941);
or U4096 (N_4096,In_529,In_342);
xnor U4097 (N_4097,In_1418,In_266);
nand U4098 (N_4098,In_387,In_526);
nand U4099 (N_4099,In_333,In_2272);
or U4100 (N_4100,In_2183,In_2017);
xnor U4101 (N_4101,In_2659,In_171);
and U4102 (N_4102,In_309,In_1592);
xnor U4103 (N_4103,In_188,In_1016);
and U4104 (N_4104,In_2312,In_2884);
and U4105 (N_4105,In_2976,In_2024);
and U4106 (N_4106,In_138,In_2224);
nor U4107 (N_4107,In_2007,In_2735);
and U4108 (N_4108,In_866,In_2705);
or U4109 (N_4109,In_617,In_770);
or U4110 (N_4110,In_41,In_2620);
and U4111 (N_4111,In_699,In_2983);
and U4112 (N_4112,In_1710,In_2899);
nor U4113 (N_4113,In_1142,In_984);
nand U4114 (N_4114,In_1345,In_2706);
nor U4115 (N_4115,In_664,In_775);
xor U4116 (N_4116,In_2946,In_1553);
or U4117 (N_4117,In_1216,In_603);
and U4118 (N_4118,In_1033,In_1415);
nand U4119 (N_4119,In_1378,In_289);
and U4120 (N_4120,In_142,In_214);
nand U4121 (N_4121,In_551,In_1144);
xor U4122 (N_4122,In_524,In_927);
and U4123 (N_4123,In_1049,In_2304);
nand U4124 (N_4124,In_2956,In_2317);
or U4125 (N_4125,In_2384,In_2044);
or U4126 (N_4126,In_2670,In_1354);
nor U4127 (N_4127,In_771,In_1931);
or U4128 (N_4128,In_1300,In_2455);
nor U4129 (N_4129,In_2474,In_151);
and U4130 (N_4130,In_2636,In_678);
and U4131 (N_4131,In_2439,In_2862);
and U4132 (N_4132,In_1922,In_1401);
nor U4133 (N_4133,In_462,In_1461);
or U4134 (N_4134,In_1396,In_2573);
nand U4135 (N_4135,In_2152,In_2218);
xnor U4136 (N_4136,In_63,In_1996);
nor U4137 (N_4137,In_28,In_227);
and U4138 (N_4138,In_34,In_909);
xnor U4139 (N_4139,In_587,In_2404);
or U4140 (N_4140,In_424,In_2513);
nand U4141 (N_4141,In_844,In_748);
or U4142 (N_4142,In_1301,In_2676);
or U4143 (N_4143,In_2402,In_506);
or U4144 (N_4144,In_1582,In_967);
or U4145 (N_4145,In_1427,In_1426);
or U4146 (N_4146,In_2576,In_188);
or U4147 (N_4147,In_2125,In_2595);
or U4148 (N_4148,In_1014,In_2928);
nand U4149 (N_4149,In_767,In_998);
nand U4150 (N_4150,In_58,In_116);
or U4151 (N_4151,In_470,In_2349);
xnor U4152 (N_4152,In_2255,In_1936);
and U4153 (N_4153,In_2079,In_1809);
nor U4154 (N_4154,In_2141,In_2593);
nor U4155 (N_4155,In_2352,In_1104);
nor U4156 (N_4156,In_2637,In_1903);
or U4157 (N_4157,In_2343,In_2898);
nor U4158 (N_4158,In_2588,In_2286);
and U4159 (N_4159,In_105,In_1805);
and U4160 (N_4160,In_1153,In_803);
and U4161 (N_4161,In_839,In_934);
nand U4162 (N_4162,In_2315,In_679);
and U4163 (N_4163,In_1061,In_2204);
nor U4164 (N_4164,In_1569,In_2615);
nor U4165 (N_4165,In_905,In_1284);
xor U4166 (N_4166,In_2262,In_1523);
and U4167 (N_4167,In_2124,In_481);
nand U4168 (N_4168,In_989,In_445);
and U4169 (N_4169,In_837,In_951);
xnor U4170 (N_4170,In_1926,In_464);
xnor U4171 (N_4171,In_835,In_2074);
and U4172 (N_4172,In_988,In_2998);
nor U4173 (N_4173,In_2559,In_2524);
nor U4174 (N_4174,In_2928,In_911);
xnor U4175 (N_4175,In_997,In_2178);
nand U4176 (N_4176,In_2344,In_171);
nand U4177 (N_4177,In_501,In_1304);
or U4178 (N_4178,In_2689,In_894);
or U4179 (N_4179,In_212,In_1163);
and U4180 (N_4180,In_390,In_821);
and U4181 (N_4181,In_1510,In_2926);
xnor U4182 (N_4182,In_1271,In_980);
or U4183 (N_4183,In_1010,In_378);
nor U4184 (N_4184,In_453,In_260);
nor U4185 (N_4185,In_2761,In_15);
and U4186 (N_4186,In_2017,In_1049);
nand U4187 (N_4187,In_1727,In_1057);
nor U4188 (N_4188,In_202,In_910);
or U4189 (N_4189,In_389,In_1410);
or U4190 (N_4190,In_227,In_2124);
nand U4191 (N_4191,In_255,In_1759);
nor U4192 (N_4192,In_2363,In_1144);
or U4193 (N_4193,In_1366,In_2568);
nand U4194 (N_4194,In_2,In_1986);
or U4195 (N_4195,In_2570,In_1687);
nand U4196 (N_4196,In_2930,In_1483);
nor U4197 (N_4197,In_92,In_2836);
nand U4198 (N_4198,In_2200,In_284);
nor U4199 (N_4199,In_1530,In_1029);
or U4200 (N_4200,In_855,In_489);
and U4201 (N_4201,In_2966,In_272);
or U4202 (N_4202,In_884,In_1246);
nand U4203 (N_4203,In_2444,In_1818);
nand U4204 (N_4204,In_2226,In_1655);
nor U4205 (N_4205,In_2687,In_2817);
nor U4206 (N_4206,In_309,In_2537);
or U4207 (N_4207,In_327,In_654);
nand U4208 (N_4208,In_2939,In_2070);
or U4209 (N_4209,In_169,In_351);
nor U4210 (N_4210,In_1619,In_248);
or U4211 (N_4211,In_349,In_2686);
xor U4212 (N_4212,In_845,In_1410);
nand U4213 (N_4213,In_2358,In_1604);
nor U4214 (N_4214,In_1866,In_1652);
nand U4215 (N_4215,In_2594,In_454);
or U4216 (N_4216,In_1098,In_2409);
and U4217 (N_4217,In_1066,In_1268);
and U4218 (N_4218,In_1825,In_2446);
nor U4219 (N_4219,In_125,In_825);
and U4220 (N_4220,In_2420,In_504);
nor U4221 (N_4221,In_533,In_419);
and U4222 (N_4222,In_761,In_2458);
xor U4223 (N_4223,In_2721,In_1611);
or U4224 (N_4224,In_936,In_119);
xnor U4225 (N_4225,In_165,In_2090);
nor U4226 (N_4226,In_2760,In_1140);
nand U4227 (N_4227,In_570,In_1951);
xor U4228 (N_4228,In_2869,In_1359);
nor U4229 (N_4229,In_1083,In_1495);
or U4230 (N_4230,In_1022,In_2428);
and U4231 (N_4231,In_4,In_1969);
or U4232 (N_4232,In_2687,In_1195);
xor U4233 (N_4233,In_1036,In_662);
or U4234 (N_4234,In_1882,In_1865);
or U4235 (N_4235,In_1778,In_1476);
and U4236 (N_4236,In_2878,In_1054);
xor U4237 (N_4237,In_862,In_2294);
xor U4238 (N_4238,In_892,In_574);
nor U4239 (N_4239,In_2444,In_2950);
and U4240 (N_4240,In_1732,In_2012);
nand U4241 (N_4241,In_2469,In_1172);
nand U4242 (N_4242,In_234,In_760);
and U4243 (N_4243,In_2004,In_2897);
and U4244 (N_4244,In_1565,In_1432);
or U4245 (N_4245,In_416,In_2922);
or U4246 (N_4246,In_2080,In_1989);
nand U4247 (N_4247,In_276,In_1127);
nand U4248 (N_4248,In_290,In_74);
nor U4249 (N_4249,In_2774,In_930);
and U4250 (N_4250,In_2723,In_2527);
nor U4251 (N_4251,In_2139,In_1904);
xnor U4252 (N_4252,In_2372,In_2669);
xnor U4253 (N_4253,In_2127,In_241);
or U4254 (N_4254,In_315,In_126);
nor U4255 (N_4255,In_2119,In_477);
nand U4256 (N_4256,In_2686,In_2165);
nor U4257 (N_4257,In_186,In_110);
nand U4258 (N_4258,In_1084,In_18);
or U4259 (N_4259,In_407,In_1679);
nor U4260 (N_4260,In_2420,In_1987);
or U4261 (N_4261,In_1035,In_1271);
nor U4262 (N_4262,In_535,In_826);
or U4263 (N_4263,In_1218,In_407);
nand U4264 (N_4264,In_1077,In_1364);
or U4265 (N_4265,In_193,In_729);
or U4266 (N_4266,In_881,In_993);
nand U4267 (N_4267,In_1406,In_662);
nand U4268 (N_4268,In_2998,In_259);
and U4269 (N_4269,In_1816,In_1395);
nor U4270 (N_4270,In_792,In_1708);
and U4271 (N_4271,In_910,In_2857);
nand U4272 (N_4272,In_1233,In_1714);
and U4273 (N_4273,In_1082,In_152);
or U4274 (N_4274,In_529,In_2699);
nor U4275 (N_4275,In_2825,In_2192);
or U4276 (N_4276,In_448,In_2519);
nand U4277 (N_4277,In_1537,In_895);
or U4278 (N_4278,In_1478,In_661);
or U4279 (N_4279,In_635,In_2935);
nand U4280 (N_4280,In_2407,In_862);
or U4281 (N_4281,In_733,In_1111);
nor U4282 (N_4282,In_626,In_533);
nand U4283 (N_4283,In_810,In_844);
xnor U4284 (N_4284,In_2790,In_415);
nand U4285 (N_4285,In_2425,In_2898);
and U4286 (N_4286,In_2888,In_420);
nor U4287 (N_4287,In_860,In_1130);
and U4288 (N_4288,In_449,In_1433);
and U4289 (N_4289,In_2096,In_2027);
nor U4290 (N_4290,In_958,In_2087);
nor U4291 (N_4291,In_362,In_2597);
nor U4292 (N_4292,In_1356,In_176);
nand U4293 (N_4293,In_2370,In_2563);
nand U4294 (N_4294,In_426,In_12);
nor U4295 (N_4295,In_849,In_1782);
nor U4296 (N_4296,In_350,In_1821);
and U4297 (N_4297,In_1472,In_442);
nor U4298 (N_4298,In_1517,In_284);
or U4299 (N_4299,In_1492,In_992);
nor U4300 (N_4300,In_487,In_2978);
nor U4301 (N_4301,In_2864,In_523);
or U4302 (N_4302,In_847,In_390);
xnor U4303 (N_4303,In_2734,In_1649);
nor U4304 (N_4304,In_2844,In_2725);
nor U4305 (N_4305,In_2831,In_1685);
or U4306 (N_4306,In_1760,In_2437);
or U4307 (N_4307,In_111,In_2792);
or U4308 (N_4308,In_2065,In_1151);
and U4309 (N_4309,In_2652,In_2962);
nand U4310 (N_4310,In_1486,In_2042);
nor U4311 (N_4311,In_2706,In_190);
nor U4312 (N_4312,In_164,In_2496);
nand U4313 (N_4313,In_1070,In_822);
or U4314 (N_4314,In_2387,In_1735);
nor U4315 (N_4315,In_2897,In_2928);
and U4316 (N_4316,In_1464,In_1184);
or U4317 (N_4317,In_318,In_2033);
nand U4318 (N_4318,In_1477,In_2082);
and U4319 (N_4319,In_1616,In_2163);
nor U4320 (N_4320,In_2530,In_1245);
nand U4321 (N_4321,In_2855,In_1049);
and U4322 (N_4322,In_366,In_2693);
nand U4323 (N_4323,In_1612,In_1086);
nand U4324 (N_4324,In_1870,In_1488);
or U4325 (N_4325,In_2862,In_2460);
nand U4326 (N_4326,In_579,In_356);
and U4327 (N_4327,In_2142,In_8);
nor U4328 (N_4328,In_2269,In_2113);
nor U4329 (N_4329,In_1846,In_2080);
or U4330 (N_4330,In_698,In_745);
nor U4331 (N_4331,In_1722,In_752);
nor U4332 (N_4332,In_841,In_1800);
nor U4333 (N_4333,In_2719,In_1928);
xnor U4334 (N_4334,In_1747,In_1260);
xnor U4335 (N_4335,In_600,In_2565);
nand U4336 (N_4336,In_1817,In_2032);
or U4337 (N_4337,In_232,In_2938);
and U4338 (N_4338,In_1977,In_586);
and U4339 (N_4339,In_278,In_1181);
nor U4340 (N_4340,In_2061,In_306);
xnor U4341 (N_4341,In_657,In_1442);
and U4342 (N_4342,In_1459,In_2056);
and U4343 (N_4343,In_2914,In_1438);
or U4344 (N_4344,In_2398,In_69);
nor U4345 (N_4345,In_763,In_1518);
nand U4346 (N_4346,In_2150,In_2015);
nand U4347 (N_4347,In_518,In_534);
or U4348 (N_4348,In_31,In_1921);
nor U4349 (N_4349,In_1090,In_2995);
xor U4350 (N_4350,In_1008,In_1245);
xor U4351 (N_4351,In_372,In_1244);
nand U4352 (N_4352,In_686,In_1432);
xor U4353 (N_4353,In_1405,In_1781);
or U4354 (N_4354,In_2602,In_1375);
or U4355 (N_4355,In_403,In_975);
nand U4356 (N_4356,In_1326,In_643);
nand U4357 (N_4357,In_276,In_1006);
nor U4358 (N_4358,In_2399,In_1081);
xnor U4359 (N_4359,In_274,In_249);
nand U4360 (N_4360,In_295,In_1593);
nand U4361 (N_4361,In_954,In_1104);
nand U4362 (N_4362,In_1953,In_1254);
xor U4363 (N_4363,In_818,In_1782);
nor U4364 (N_4364,In_2726,In_1741);
nor U4365 (N_4365,In_522,In_1513);
nor U4366 (N_4366,In_2735,In_909);
nor U4367 (N_4367,In_2236,In_2758);
xor U4368 (N_4368,In_1779,In_782);
xor U4369 (N_4369,In_2108,In_2042);
or U4370 (N_4370,In_2735,In_1718);
and U4371 (N_4371,In_1371,In_235);
and U4372 (N_4372,In_172,In_2058);
and U4373 (N_4373,In_100,In_1670);
nor U4374 (N_4374,In_2542,In_1943);
nand U4375 (N_4375,In_1419,In_2136);
nand U4376 (N_4376,In_2558,In_495);
nand U4377 (N_4377,In_1529,In_2246);
nor U4378 (N_4378,In_369,In_2153);
or U4379 (N_4379,In_494,In_1409);
nor U4380 (N_4380,In_426,In_2319);
nand U4381 (N_4381,In_781,In_1949);
or U4382 (N_4382,In_2813,In_954);
xor U4383 (N_4383,In_2968,In_256);
xnor U4384 (N_4384,In_1667,In_1363);
nor U4385 (N_4385,In_2834,In_296);
and U4386 (N_4386,In_1470,In_474);
and U4387 (N_4387,In_1860,In_1736);
nor U4388 (N_4388,In_1409,In_2010);
or U4389 (N_4389,In_2166,In_2028);
or U4390 (N_4390,In_2143,In_2655);
nor U4391 (N_4391,In_1264,In_2651);
nand U4392 (N_4392,In_702,In_629);
nor U4393 (N_4393,In_2036,In_982);
nand U4394 (N_4394,In_2948,In_2814);
nand U4395 (N_4395,In_1108,In_2145);
nand U4396 (N_4396,In_755,In_2411);
or U4397 (N_4397,In_1239,In_1669);
or U4398 (N_4398,In_1868,In_1558);
and U4399 (N_4399,In_1138,In_1133);
or U4400 (N_4400,In_168,In_1346);
and U4401 (N_4401,In_185,In_2019);
xnor U4402 (N_4402,In_430,In_1933);
nand U4403 (N_4403,In_2801,In_19);
nor U4404 (N_4404,In_497,In_908);
nand U4405 (N_4405,In_618,In_592);
or U4406 (N_4406,In_1214,In_1418);
or U4407 (N_4407,In_740,In_1060);
or U4408 (N_4408,In_2525,In_2582);
nor U4409 (N_4409,In_547,In_557);
or U4410 (N_4410,In_409,In_1476);
or U4411 (N_4411,In_2440,In_2714);
nor U4412 (N_4412,In_1624,In_1366);
xnor U4413 (N_4413,In_984,In_1913);
and U4414 (N_4414,In_543,In_540);
or U4415 (N_4415,In_796,In_2930);
nor U4416 (N_4416,In_2381,In_1288);
nand U4417 (N_4417,In_1480,In_2959);
xor U4418 (N_4418,In_232,In_520);
and U4419 (N_4419,In_2587,In_477);
nor U4420 (N_4420,In_501,In_2671);
nand U4421 (N_4421,In_401,In_1143);
or U4422 (N_4422,In_2943,In_2603);
or U4423 (N_4423,In_1814,In_1311);
nand U4424 (N_4424,In_903,In_2827);
and U4425 (N_4425,In_265,In_364);
and U4426 (N_4426,In_103,In_2292);
nor U4427 (N_4427,In_1393,In_2900);
and U4428 (N_4428,In_2604,In_324);
nand U4429 (N_4429,In_2816,In_986);
xnor U4430 (N_4430,In_1234,In_2782);
nand U4431 (N_4431,In_9,In_1596);
nor U4432 (N_4432,In_107,In_782);
nor U4433 (N_4433,In_755,In_2696);
nand U4434 (N_4434,In_2875,In_692);
nor U4435 (N_4435,In_2004,In_2716);
xnor U4436 (N_4436,In_2836,In_750);
or U4437 (N_4437,In_1228,In_1837);
and U4438 (N_4438,In_273,In_415);
nor U4439 (N_4439,In_146,In_367);
and U4440 (N_4440,In_1772,In_1188);
nand U4441 (N_4441,In_2797,In_2316);
nand U4442 (N_4442,In_310,In_10);
xnor U4443 (N_4443,In_580,In_1894);
nor U4444 (N_4444,In_593,In_1287);
xor U4445 (N_4445,In_262,In_2834);
and U4446 (N_4446,In_1241,In_1233);
xnor U4447 (N_4447,In_1860,In_754);
nor U4448 (N_4448,In_2221,In_723);
nand U4449 (N_4449,In_212,In_699);
and U4450 (N_4450,In_1564,In_533);
and U4451 (N_4451,In_865,In_503);
or U4452 (N_4452,In_931,In_285);
nand U4453 (N_4453,In_2477,In_2879);
and U4454 (N_4454,In_1431,In_1143);
and U4455 (N_4455,In_563,In_2952);
nor U4456 (N_4456,In_1188,In_864);
or U4457 (N_4457,In_2640,In_813);
or U4458 (N_4458,In_148,In_2298);
or U4459 (N_4459,In_1017,In_606);
or U4460 (N_4460,In_1756,In_1475);
and U4461 (N_4461,In_1275,In_245);
or U4462 (N_4462,In_2069,In_1198);
and U4463 (N_4463,In_1567,In_1335);
nor U4464 (N_4464,In_2420,In_1381);
and U4465 (N_4465,In_1552,In_2964);
or U4466 (N_4466,In_2747,In_2304);
nor U4467 (N_4467,In_2524,In_450);
nor U4468 (N_4468,In_2405,In_1545);
nor U4469 (N_4469,In_2118,In_2420);
nor U4470 (N_4470,In_613,In_95);
nand U4471 (N_4471,In_2100,In_2308);
nand U4472 (N_4472,In_1658,In_2279);
nor U4473 (N_4473,In_1389,In_2196);
and U4474 (N_4474,In_2682,In_2872);
and U4475 (N_4475,In_2438,In_2226);
and U4476 (N_4476,In_2036,In_2145);
nand U4477 (N_4477,In_669,In_2707);
nand U4478 (N_4478,In_2340,In_2422);
nor U4479 (N_4479,In_1307,In_2779);
and U4480 (N_4480,In_255,In_1259);
and U4481 (N_4481,In_2205,In_1092);
xnor U4482 (N_4482,In_2605,In_2441);
nand U4483 (N_4483,In_1156,In_2800);
and U4484 (N_4484,In_2376,In_2229);
or U4485 (N_4485,In_864,In_1657);
nor U4486 (N_4486,In_54,In_1732);
xor U4487 (N_4487,In_135,In_1283);
xnor U4488 (N_4488,In_1989,In_2880);
and U4489 (N_4489,In_345,In_480);
nand U4490 (N_4490,In_1856,In_1105);
nand U4491 (N_4491,In_547,In_1687);
nor U4492 (N_4492,In_2920,In_1417);
nor U4493 (N_4493,In_2386,In_1751);
xnor U4494 (N_4494,In_2868,In_682);
nor U4495 (N_4495,In_2285,In_736);
and U4496 (N_4496,In_2410,In_1884);
and U4497 (N_4497,In_2861,In_1420);
nand U4498 (N_4498,In_2576,In_930);
nor U4499 (N_4499,In_455,In_488);
xnor U4500 (N_4500,In_2214,In_2160);
xor U4501 (N_4501,In_2960,In_1662);
nor U4502 (N_4502,In_220,In_1267);
nor U4503 (N_4503,In_400,In_1022);
and U4504 (N_4504,In_2630,In_2223);
nor U4505 (N_4505,In_293,In_679);
and U4506 (N_4506,In_51,In_1283);
nand U4507 (N_4507,In_732,In_1028);
nor U4508 (N_4508,In_471,In_1721);
and U4509 (N_4509,In_355,In_463);
or U4510 (N_4510,In_504,In_36);
xor U4511 (N_4511,In_2594,In_2847);
or U4512 (N_4512,In_1621,In_30);
or U4513 (N_4513,In_799,In_667);
nand U4514 (N_4514,In_1967,In_7);
nand U4515 (N_4515,In_167,In_2789);
or U4516 (N_4516,In_639,In_937);
nor U4517 (N_4517,In_405,In_1343);
nand U4518 (N_4518,In_2469,In_1157);
or U4519 (N_4519,In_2981,In_1462);
and U4520 (N_4520,In_1211,In_2606);
or U4521 (N_4521,In_1564,In_242);
nor U4522 (N_4522,In_1560,In_1096);
nand U4523 (N_4523,In_678,In_1884);
or U4524 (N_4524,In_1360,In_2635);
nand U4525 (N_4525,In_2797,In_404);
nand U4526 (N_4526,In_193,In_292);
nand U4527 (N_4527,In_591,In_1443);
or U4528 (N_4528,In_963,In_2427);
nand U4529 (N_4529,In_2078,In_2228);
and U4530 (N_4530,In_1309,In_482);
nor U4531 (N_4531,In_2396,In_1658);
nor U4532 (N_4532,In_2656,In_2801);
nand U4533 (N_4533,In_147,In_779);
nand U4534 (N_4534,In_1284,In_1636);
nand U4535 (N_4535,In_2336,In_2934);
nand U4536 (N_4536,In_2118,In_2275);
nor U4537 (N_4537,In_1325,In_1177);
or U4538 (N_4538,In_2399,In_82);
nand U4539 (N_4539,In_2436,In_991);
and U4540 (N_4540,In_1535,In_2595);
and U4541 (N_4541,In_463,In_1001);
xnor U4542 (N_4542,In_189,In_2696);
nand U4543 (N_4543,In_1546,In_2622);
or U4544 (N_4544,In_227,In_1725);
or U4545 (N_4545,In_2368,In_502);
nor U4546 (N_4546,In_857,In_449);
or U4547 (N_4547,In_1064,In_46);
nand U4548 (N_4548,In_1530,In_1389);
nor U4549 (N_4549,In_2808,In_2440);
nor U4550 (N_4550,In_2886,In_533);
or U4551 (N_4551,In_1812,In_624);
nand U4552 (N_4552,In_296,In_68);
nand U4553 (N_4553,In_2470,In_2);
or U4554 (N_4554,In_2819,In_749);
or U4555 (N_4555,In_1765,In_1141);
and U4556 (N_4556,In_1756,In_2684);
nor U4557 (N_4557,In_2652,In_1908);
or U4558 (N_4558,In_2126,In_1005);
and U4559 (N_4559,In_890,In_2658);
xor U4560 (N_4560,In_2956,In_570);
nor U4561 (N_4561,In_2415,In_1890);
or U4562 (N_4562,In_1206,In_1086);
or U4563 (N_4563,In_276,In_1267);
or U4564 (N_4564,In_1765,In_2424);
or U4565 (N_4565,In_2719,In_2948);
and U4566 (N_4566,In_1516,In_1533);
xnor U4567 (N_4567,In_347,In_895);
nor U4568 (N_4568,In_346,In_2032);
xnor U4569 (N_4569,In_477,In_2105);
nand U4570 (N_4570,In_2948,In_1238);
or U4571 (N_4571,In_651,In_1565);
or U4572 (N_4572,In_1850,In_540);
or U4573 (N_4573,In_477,In_1034);
and U4574 (N_4574,In_1334,In_1989);
nand U4575 (N_4575,In_2094,In_2311);
or U4576 (N_4576,In_2819,In_2351);
nand U4577 (N_4577,In_617,In_2392);
xor U4578 (N_4578,In_2250,In_1111);
or U4579 (N_4579,In_1643,In_2080);
or U4580 (N_4580,In_2299,In_2037);
and U4581 (N_4581,In_1396,In_902);
or U4582 (N_4582,In_1553,In_1943);
or U4583 (N_4583,In_2251,In_2939);
nor U4584 (N_4584,In_941,In_1186);
or U4585 (N_4585,In_1982,In_1814);
xor U4586 (N_4586,In_2856,In_2428);
xnor U4587 (N_4587,In_2522,In_2404);
nand U4588 (N_4588,In_2423,In_1805);
or U4589 (N_4589,In_2769,In_2176);
nor U4590 (N_4590,In_593,In_950);
nand U4591 (N_4591,In_1237,In_2367);
and U4592 (N_4592,In_1444,In_665);
or U4593 (N_4593,In_2961,In_993);
xnor U4594 (N_4594,In_1066,In_2722);
nor U4595 (N_4595,In_1507,In_2661);
or U4596 (N_4596,In_934,In_1985);
and U4597 (N_4597,In_604,In_2248);
and U4598 (N_4598,In_1161,In_2931);
xor U4599 (N_4599,In_2774,In_2752);
nor U4600 (N_4600,In_81,In_1784);
nand U4601 (N_4601,In_556,In_2029);
and U4602 (N_4602,In_1835,In_1852);
or U4603 (N_4603,In_958,In_1680);
nor U4604 (N_4604,In_177,In_1309);
nand U4605 (N_4605,In_1891,In_2688);
xnor U4606 (N_4606,In_2635,In_2457);
and U4607 (N_4607,In_2708,In_755);
and U4608 (N_4608,In_130,In_1539);
nand U4609 (N_4609,In_45,In_1064);
xnor U4610 (N_4610,In_321,In_2312);
or U4611 (N_4611,In_2865,In_2646);
nor U4612 (N_4612,In_2565,In_2023);
or U4613 (N_4613,In_1986,In_2611);
nor U4614 (N_4614,In_1636,In_894);
or U4615 (N_4615,In_2842,In_438);
and U4616 (N_4616,In_1942,In_803);
xnor U4617 (N_4617,In_1482,In_551);
and U4618 (N_4618,In_683,In_2416);
or U4619 (N_4619,In_2641,In_943);
nand U4620 (N_4620,In_1711,In_298);
nand U4621 (N_4621,In_343,In_1081);
nor U4622 (N_4622,In_1771,In_2373);
and U4623 (N_4623,In_1791,In_1157);
nor U4624 (N_4624,In_953,In_738);
nand U4625 (N_4625,In_2889,In_300);
nand U4626 (N_4626,In_2297,In_910);
or U4627 (N_4627,In_1829,In_410);
nor U4628 (N_4628,In_2396,In_2067);
nand U4629 (N_4629,In_2227,In_1513);
nand U4630 (N_4630,In_238,In_578);
nor U4631 (N_4631,In_2693,In_2658);
nand U4632 (N_4632,In_738,In_1273);
nand U4633 (N_4633,In_598,In_104);
nand U4634 (N_4634,In_2917,In_1056);
nand U4635 (N_4635,In_2010,In_2027);
and U4636 (N_4636,In_2639,In_2188);
and U4637 (N_4637,In_1191,In_2803);
xnor U4638 (N_4638,In_1441,In_1119);
nor U4639 (N_4639,In_704,In_1839);
or U4640 (N_4640,In_2636,In_2048);
or U4641 (N_4641,In_2524,In_2509);
nand U4642 (N_4642,In_2182,In_712);
nor U4643 (N_4643,In_1374,In_30);
or U4644 (N_4644,In_1315,In_1464);
nor U4645 (N_4645,In_259,In_890);
nor U4646 (N_4646,In_931,In_1896);
or U4647 (N_4647,In_2876,In_2776);
and U4648 (N_4648,In_1152,In_620);
or U4649 (N_4649,In_2629,In_603);
nand U4650 (N_4650,In_1534,In_1527);
xnor U4651 (N_4651,In_1749,In_1529);
and U4652 (N_4652,In_1448,In_2920);
and U4653 (N_4653,In_1493,In_165);
or U4654 (N_4654,In_2190,In_2905);
nor U4655 (N_4655,In_2259,In_1583);
and U4656 (N_4656,In_1499,In_2851);
nand U4657 (N_4657,In_2730,In_1273);
nand U4658 (N_4658,In_592,In_2061);
nor U4659 (N_4659,In_1344,In_2908);
or U4660 (N_4660,In_115,In_1943);
nor U4661 (N_4661,In_2999,In_988);
nor U4662 (N_4662,In_2587,In_1534);
xor U4663 (N_4663,In_1027,In_1493);
or U4664 (N_4664,In_312,In_243);
nand U4665 (N_4665,In_2376,In_1973);
nor U4666 (N_4666,In_2960,In_1929);
nor U4667 (N_4667,In_1139,In_2487);
or U4668 (N_4668,In_605,In_1050);
nand U4669 (N_4669,In_1259,In_2299);
xnor U4670 (N_4670,In_752,In_345);
or U4671 (N_4671,In_2564,In_1033);
nand U4672 (N_4672,In_6,In_2169);
nand U4673 (N_4673,In_658,In_2541);
nor U4674 (N_4674,In_476,In_1634);
nand U4675 (N_4675,In_785,In_2753);
and U4676 (N_4676,In_86,In_363);
nand U4677 (N_4677,In_2720,In_1733);
and U4678 (N_4678,In_2503,In_2667);
or U4679 (N_4679,In_579,In_804);
or U4680 (N_4680,In_1821,In_675);
nand U4681 (N_4681,In_797,In_2312);
xor U4682 (N_4682,In_330,In_1586);
nor U4683 (N_4683,In_992,In_1777);
or U4684 (N_4684,In_1430,In_1086);
nand U4685 (N_4685,In_151,In_2741);
and U4686 (N_4686,In_2580,In_12);
nand U4687 (N_4687,In_2341,In_568);
or U4688 (N_4688,In_1563,In_2941);
or U4689 (N_4689,In_1634,In_1460);
or U4690 (N_4690,In_1942,In_1463);
nand U4691 (N_4691,In_2687,In_66);
or U4692 (N_4692,In_534,In_1117);
or U4693 (N_4693,In_2012,In_1792);
and U4694 (N_4694,In_1444,In_763);
nand U4695 (N_4695,In_239,In_1880);
nor U4696 (N_4696,In_2294,In_1822);
or U4697 (N_4697,In_256,In_1762);
nor U4698 (N_4698,In_2573,In_1205);
or U4699 (N_4699,In_2634,In_2659);
nor U4700 (N_4700,In_2086,In_1244);
nand U4701 (N_4701,In_714,In_2101);
and U4702 (N_4702,In_103,In_1049);
nor U4703 (N_4703,In_1289,In_1431);
and U4704 (N_4704,In_1740,In_2834);
nor U4705 (N_4705,In_1405,In_101);
or U4706 (N_4706,In_2953,In_2570);
nand U4707 (N_4707,In_501,In_2712);
and U4708 (N_4708,In_1779,In_2556);
and U4709 (N_4709,In_1017,In_2207);
or U4710 (N_4710,In_205,In_2269);
nor U4711 (N_4711,In_2463,In_1252);
or U4712 (N_4712,In_1990,In_1744);
xor U4713 (N_4713,In_2233,In_1978);
nand U4714 (N_4714,In_2345,In_1242);
nand U4715 (N_4715,In_2027,In_2547);
and U4716 (N_4716,In_492,In_831);
or U4717 (N_4717,In_321,In_574);
nor U4718 (N_4718,In_2167,In_1860);
and U4719 (N_4719,In_2895,In_1189);
xnor U4720 (N_4720,In_1206,In_2700);
nand U4721 (N_4721,In_592,In_322);
and U4722 (N_4722,In_1958,In_164);
nor U4723 (N_4723,In_1946,In_1502);
or U4724 (N_4724,In_1945,In_1104);
and U4725 (N_4725,In_171,In_412);
nor U4726 (N_4726,In_2787,In_1639);
nand U4727 (N_4727,In_2427,In_831);
nand U4728 (N_4728,In_1552,In_2218);
and U4729 (N_4729,In_2756,In_417);
and U4730 (N_4730,In_927,In_2942);
nand U4731 (N_4731,In_1101,In_1646);
and U4732 (N_4732,In_857,In_744);
nor U4733 (N_4733,In_159,In_485);
or U4734 (N_4734,In_1066,In_1801);
nor U4735 (N_4735,In_2435,In_2342);
xor U4736 (N_4736,In_574,In_1739);
nor U4737 (N_4737,In_1489,In_750);
nand U4738 (N_4738,In_1023,In_2101);
and U4739 (N_4739,In_1994,In_1887);
and U4740 (N_4740,In_2710,In_231);
or U4741 (N_4741,In_184,In_23);
nand U4742 (N_4742,In_1772,In_190);
or U4743 (N_4743,In_1087,In_2066);
and U4744 (N_4744,In_1655,In_1379);
and U4745 (N_4745,In_512,In_503);
and U4746 (N_4746,In_2075,In_2878);
xnor U4747 (N_4747,In_1303,In_349);
and U4748 (N_4748,In_1724,In_491);
nand U4749 (N_4749,In_1263,In_264);
and U4750 (N_4750,In_2766,In_1121);
nor U4751 (N_4751,In_1089,In_1352);
nand U4752 (N_4752,In_505,In_2120);
and U4753 (N_4753,In_866,In_2739);
nor U4754 (N_4754,In_353,In_2463);
or U4755 (N_4755,In_1158,In_2976);
nand U4756 (N_4756,In_893,In_1513);
and U4757 (N_4757,In_406,In_2918);
nand U4758 (N_4758,In_670,In_1999);
nor U4759 (N_4759,In_2413,In_934);
nand U4760 (N_4760,In_2628,In_632);
nor U4761 (N_4761,In_152,In_329);
nand U4762 (N_4762,In_2429,In_768);
nor U4763 (N_4763,In_76,In_1497);
nor U4764 (N_4764,In_873,In_2059);
or U4765 (N_4765,In_2950,In_886);
xor U4766 (N_4766,In_2101,In_1220);
nor U4767 (N_4767,In_1771,In_73);
nor U4768 (N_4768,In_1115,In_700);
and U4769 (N_4769,In_517,In_1175);
nand U4770 (N_4770,In_189,In_1492);
and U4771 (N_4771,In_2116,In_657);
nand U4772 (N_4772,In_792,In_386);
and U4773 (N_4773,In_588,In_2830);
nand U4774 (N_4774,In_2483,In_91);
or U4775 (N_4775,In_373,In_2644);
nor U4776 (N_4776,In_2936,In_98);
or U4777 (N_4777,In_1011,In_2642);
nand U4778 (N_4778,In_2900,In_1282);
and U4779 (N_4779,In_1833,In_1897);
nor U4780 (N_4780,In_2987,In_35);
nor U4781 (N_4781,In_127,In_332);
and U4782 (N_4782,In_1297,In_1168);
or U4783 (N_4783,In_1268,In_232);
xor U4784 (N_4784,In_1480,In_13);
nor U4785 (N_4785,In_2089,In_1335);
or U4786 (N_4786,In_877,In_1645);
nor U4787 (N_4787,In_1032,In_1179);
and U4788 (N_4788,In_1632,In_803);
or U4789 (N_4789,In_492,In_1862);
nand U4790 (N_4790,In_2256,In_517);
xnor U4791 (N_4791,In_1901,In_1462);
or U4792 (N_4792,In_625,In_715);
xnor U4793 (N_4793,In_1786,In_1037);
or U4794 (N_4794,In_2746,In_1842);
nand U4795 (N_4795,In_972,In_2034);
nor U4796 (N_4796,In_814,In_2678);
or U4797 (N_4797,In_2875,In_2727);
and U4798 (N_4798,In_249,In_117);
nand U4799 (N_4799,In_1901,In_524);
and U4800 (N_4800,In_1086,In_586);
nor U4801 (N_4801,In_655,In_74);
nand U4802 (N_4802,In_2302,In_2225);
nand U4803 (N_4803,In_521,In_1126);
or U4804 (N_4804,In_2149,In_568);
or U4805 (N_4805,In_2875,In_1856);
or U4806 (N_4806,In_2878,In_2625);
and U4807 (N_4807,In_2043,In_96);
or U4808 (N_4808,In_750,In_320);
nand U4809 (N_4809,In_2628,In_945);
and U4810 (N_4810,In_1355,In_1046);
nand U4811 (N_4811,In_1197,In_2169);
nor U4812 (N_4812,In_835,In_410);
and U4813 (N_4813,In_77,In_706);
or U4814 (N_4814,In_741,In_2376);
nor U4815 (N_4815,In_1896,In_702);
nand U4816 (N_4816,In_1399,In_582);
xnor U4817 (N_4817,In_1771,In_2611);
nor U4818 (N_4818,In_2790,In_1834);
nand U4819 (N_4819,In_658,In_518);
nor U4820 (N_4820,In_1239,In_833);
and U4821 (N_4821,In_1274,In_2858);
xnor U4822 (N_4822,In_908,In_1321);
or U4823 (N_4823,In_918,In_2084);
or U4824 (N_4824,In_907,In_615);
nand U4825 (N_4825,In_2019,In_1662);
or U4826 (N_4826,In_1257,In_422);
or U4827 (N_4827,In_117,In_536);
or U4828 (N_4828,In_2449,In_2611);
or U4829 (N_4829,In_291,In_1302);
nor U4830 (N_4830,In_1417,In_2605);
nand U4831 (N_4831,In_814,In_2536);
nor U4832 (N_4832,In_176,In_1086);
nand U4833 (N_4833,In_162,In_1185);
nor U4834 (N_4834,In_2340,In_1535);
xor U4835 (N_4835,In_1160,In_1706);
nand U4836 (N_4836,In_752,In_434);
nand U4837 (N_4837,In_1717,In_2170);
and U4838 (N_4838,In_411,In_1703);
or U4839 (N_4839,In_177,In_2645);
and U4840 (N_4840,In_2615,In_917);
and U4841 (N_4841,In_2618,In_419);
nor U4842 (N_4842,In_1839,In_1090);
and U4843 (N_4843,In_816,In_2546);
and U4844 (N_4844,In_818,In_2001);
nand U4845 (N_4845,In_1477,In_865);
nor U4846 (N_4846,In_646,In_2527);
or U4847 (N_4847,In_164,In_242);
xnor U4848 (N_4848,In_2338,In_2896);
nor U4849 (N_4849,In_2960,In_156);
nor U4850 (N_4850,In_910,In_2793);
or U4851 (N_4851,In_860,In_743);
or U4852 (N_4852,In_288,In_1903);
or U4853 (N_4853,In_1683,In_2379);
and U4854 (N_4854,In_2772,In_1463);
nand U4855 (N_4855,In_2318,In_2103);
nor U4856 (N_4856,In_609,In_1069);
nor U4857 (N_4857,In_1981,In_655);
nand U4858 (N_4858,In_804,In_1497);
or U4859 (N_4859,In_1607,In_272);
nand U4860 (N_4860,In_2558,In_997);
or U4861 (N_4861,In_452,In_1611);
or U4862 (N_4862,In_2317,In_718);
or U4863 (N_4863,In_2042,In_1470);
nand U4864 (N_4864,In_2977,In_1507);
nand U4865 (N_4865,In_435,In_319);
or U4866 (N_4866,In_839,In_2);
and U4867 (N_4867,In_2900,In_2548);
and U4868 (N_4868,In_415,In_2144);
nor U4869 (N_4869,In_1774,In_1982);
nand U4870 (N_4870,In_206,In_2014);
and U4871 (N_4871,In_707,In_2834);
nand U4872 (N_4872,In_2801,In_567);
nor U4873 (N_4873,In_1790,In_1051);
nor U4874 (N_4874,In_1700,In_777);
or U4875 (N_4875,In_347,In_253);
or U4876 (N_4876,In_1339,In_781);
nand U4877 (N_4877,In_1392,In_389);
or U4878 (N_4878,In_1979,In_2052);
and U4879 (N_4879,In_394,In_2094);
and U4880 (N_4880,In_2130,In_124);
nand U4881 (N_4881,In_2734,In_894);
and U4882 (N_4882,In_465,In_1469);
and U4883 (N_4883,In_1773,In_212);
nor U4884 (N_4884,In_2395,In_293);
nor U4885 (N_4885,In_66,In_879);
and U4886 (N_4886,In_727,In_790);
nand U4887 (N_4887,In_2168,In_2238);
or U4888 (N_4888,In_2881,In_1148);
nand U4889 (N_4889,In_2499,In_2816);
or U4890 (N_4890,In_810,In_288);
nand U4891 (N_4891,In_2686,In_777);
and U4892 (N_4892,In_1113,In_2982);
nor U4893 (N_4893,In_26,In_1400);
and U4894 (N_4894,In_2787,In_373);
nand U4895 (N_4895,In_1416,In_2385);
nand U4896 (N_4896,In_785,In_2841);
and U4897 (N_4897,In_1707,In_97);
and U4898 (N_4898,In_2376,In_1205);
nand U4899 (N_4899,In_1269,In_756);
nand U4900 (N_4900,In_2885,In_1714);
or U4901 (N_4901,In_262,In_669);
nor U4902 (N_4902,In_1578,In_345);
nand U4903 (N_4903,In_1367,In_2474);
xnor U4904 (N_4904,In_2142,In_176);
nand U4905 (N_4905,In_161,In_349);
and U4906 (N_4906,In_1374,In_134);
nor U4907 (N_4907,In_2151,In_342);
xor U4908 (N_4908,In_439,In_2082);
and U4909 (N_4909,In_736,In_1278);
nand U4910 (N_4910,In_2766,In_720);
or U4911 (N_4911,In_1880,In_1600);
nor U4912 (N_4912,In_2126,In_316);
nand U4913 (N_4913,In_1935,In_1943);
nand U4914 (N_4914,In_2062,In_1103);
or U4915 (N_4915,In_1158,In_1405);
nand U4916 (N_4916,In_1342,In_1608);
nand U4917 (N_4917,In_2948,In_1629);
or U4918 (N_4918,In_2774,In_383);
and U4919 (N_4919,In_122,In_2427);
nor U4920 (N_4920,In_2641,In_2684);
nand U4921 (N_4921,In_1681,In_1771);
and U4922 (N_4922,In_2150,In_1602);
nor U4923 (N_4923,In_1850,In_1048);
xnor U4924 (N_4924,In_1514,In_1395);
or U4925 (N_4925,In_2628,In_567);
and U4926 (N_4926,In_57,In_1397);
or U4927 (N_4927,In_642,In_2385);
nor U4928 (N_4928,In_1184,In_1868);
nor U4929 (N_4929,In_2526,In_2271);
or U4930 (N_4930,In_2381,In_1356);
nor U4931 (N_4931,In_1908,In_2550);
xor U4932 (N_4932,In_1677,In_1226);
and U4933 (N_4933,In_2751,In_1373);
nand U4934 (N_4934,In_396,In_2683);
nand U4935 (N_4935,In_1680,In_696);
or U4936 (N_4936,In_1061,In_2291);
nor U4937 (N_4937,In_2195,In_2812);
nand U4938 (N_4938,In_2579,In_1465);
or U4939 (N_4939,In_236,In_929);
nand U4940 (N_4940,In_2552,In_2273);
nor U4941 (N_4941,In_1164,In_1801);
nor U4942 (N_4942,In_2932,In_916);
nand U4943 (N_4943,In_1030,In_1694);
and U4944 (N_4944,In_1329,In_2814);
or U4945 (N_4945,In_2059,In_628);
or U4946 (N_4946,In_787,In_2106);
nand U4947 (N_4947,In_1274,In_945);
nand U4948 (N_4948,In_1099,In_1258);
and U4949 (N_4949,In_2131,In_2870);
nor U4950 (N_4950,In_1052,In_80);
or U4951 (N_4951,In_861,In_234);
or U4952 (N_4952,In_742,In_1513);
nand U4953 (N_4953,In_1016,In_2317);
or U4954 (N_4954,In_1323,In_213);
nor U4955 (N_4955,In_1690,In_2880);
nand U4956 (N_4956,In_568,In_2581);
xor U4957 (N_4957,In_2538,In_936);
nand U4958 (N_4958,In_2470,In_1465);
or U4959 (N_4959,In_1100,In_2203);
or U4960 (N_4960,In_1130,In_2619);
and U4961 (N_4961,In_943,In_1950);
nor U4962 (N_4962,In_2196,In_316);
or U4963 (N_4963,In_1511,In_2897);
and U4964 (N_4964,In_2301,In_1499);
nand U4965 (N_4965,In_1911,In_1132);
nor U4966 (N_4966,In_807,In_2490);
nor U4967 (N_4967,In_1371,In_1952);
or U4968 (N_4968,In_691,In_2864);
xor U4969 (N_4969,In_635,In_2533);
and U4970 (N_4970,In_2402,In_298);
or U4971 (N_4971,In_1517,In_1093);
xor U4972 (N_4972,In_2619,In_596);
or U4973 (N_4973,In_1025,In_1243);
or U4974 (N_4974,In_2048,In_432);
nand U4975 (N_4975,In_1164,In_659);
nor U4976 (N_4976,In_1770,In_978);
nand U4977 (N_4977,In_285,In_817);
or U4978 (N_4978,In_2382,In_2144);
nand U4979 (N_4979,In_273,In_1334);
and U4980 (N_4980,In_2764,In_974);
nand U4981 (N_4981,In_595,In_885);
or U4982 (N_4982,In_2261,In_1576);
and U4983 (N_4983,In_759,In_2737);
nor U4984 (N_4984,In_932,In_2999);
xor U4985 (N_4985,In_1802,In_2342);
xor U4986 (N_4986,In_110,In_140);
and U4987 (N_4987,In_1047,In_137);
or U4988 (N_4988,In_1485,In_941);
nor U4989 (N_4989,In_737,In_891);
xor U4990 (N_4990,In_2177,In_1035);
nor U4991 (N_4991,In_2683,In_546);
and U4992 (N_4992,In_1496,In_632);
nand U4993 (N_4993,In_2725,In_2330);
or U4994 (N_4994,In_2352,In_1388);
or U4995 (N_4995,In_1124,In_172);
nor U4996 (N_4996,In_2102,In_1228);
or U4997 (N_4997,In_2249,In_1523);
or U4998 (N_4998,In_882,In_987);
nand U4999 (N_4999,In_2475,In_835);
nand U5000 (N_5000,N_2864,N_1219);
nor U5001 (N_5001,N_4987,N_1862);
or U5002 (N_5002,N_806,N_967);
and U5003 (N_5003,N_3908,N_1919);
and U5004 (N_5004,N_1851,N_2236);
and U5005 (N_5005,N_4029,N_4452);
or U5006 (N_5006,N_1645,N_2138);
nand U5007 (N_5007,N_1194,N_2609);
nor U5008 (N_5008,N_2939,N_1001);
nor U5009 (N_5009,N_879,N_3560);
nand U5010 (N_5010,N_1594,N_1244);
or U5011 (N_5011,N_1382,N_4084);
or U5012 (N_5012,N_3638,N_2847);
or U5013 (N_5013,N_3054,N_4828);
and U5014 (N_5014,N_4106,N_4576);
or U5015 (N_5015,N_2608,N_2200);
and U5016 (N_5016,N_4259,N_2308);
nor U5017 (N_5017,N_485,N_1271);
or U5018 (N_5018,N_647,N_1928);
nand U5019 (N_5019,N_4254,N_977);
xor U5020 (N_5020,N_238,N_2181);
nor U5021 (N_5021,N_3048,N_2105);
nand U5022 (N_5022,N_341,N_3804);
nor U5023 (N_5023,N_1886,N_2361);
nor U5024 (N_5024,N_4581,N_540);
nor U5025 (N_5025,N_1225,N_972);
nand U5026 (N_5026,N_1958,N_3898);
and U5027 (N_5027,N_764,N_4024);
or U5028 (N_5028,N_1245,N_1107);
and U5029 (N_5029,N_2971,N_2371);
or U5030 (N_5030,N_4966,N_563);
or U5031 (N_5031,N_940,N_4922);
nor U5032 (N_5032,N_2733,N_3374);
or U5033 (N_5033,N_82,N_2123);
nand U5034 (N_5034,N_338,N_1946);
nand U5035 (N_5035,N_1033,N_3372);
nand U5036 (N_5036,N_4070,N_462);
or U5037 (N_5037,N_2402,N_4339);
xnor U5038 (N_5038,N_3650,N_1854);
nand U5039 (N_5039,N_2849,N_263);
nor U5040 (N_5040,N_4709,N_992);
and U5041 (N_5041,N_4234,N_2285);
or U5042 (N_5042,N_1050,N_4596);
nor U5043 (N_5043,N_1307,N_245);
or U5044 (N_5044,N_3931,N_2839);
nor U5045 (N_5045,N_4474,N_2401);
and U5046 (N_5046,N_4522,N_609);
nand U5047 (N_5047,N_3718,N_67);
nand U5048 (N_5048,N_4951,N_3841);
nor U5049 (N_5049,N_646,N_3617);
nand U5050 (N_5050,N_631,N_291);
nor U5051 (N_5051,N_2202,N_4607);
and U5052 (N_5052,N_968,N_1653);
nor U5053 (N_5053,N_4209,N_3499);
or U5054 (N_5054,N_4134,N_2955);
nand U5055 (N_5055,N_4739,N_2342);
xnor U5056 (N_5056,N_4066,N_3000);
nand U5057 (N_5057,N_4756,N_347);
and U5058 (N_5058,N_3849,N_1455);
nand U5059 (N_5059,N_1343,N_2912);
nand U5060 (N_5060,N_4257,N_991);
and U5061 (N_5061,N_2390,N_785);
nor U5062 (N_5062,N_4701,N_4569);
or U5063 (N_5063,N_449,N_2273);
nand U5064 (N_5064,N_1908,N_2859);
and U5065 (N_5065,N_3683,N_1168);
nor U5066 (N_5066,N_1735,N_1896);
nor U5067 (N_5067,N_699,N_1598);
nor U5068 (N_5068,N_3798,N_3042);
or U5069 (N_5069,N_1777,N_2662);
and U5070 (N_5070,N_3118,N_3583);
or U5071 (N_5071,N_1736,N_1709);
nor U5072 (N_5072,N_3209,N_2570);
nand U5073 (N_5073,N_2850,N_2149);
or U5074 (N_5074,N_2998,N_225);
or U5075 (N_5075,N_2504,N_3641);
or U5076 (N_5076,N_3434,N_2016);
nand U5077 (N_5077,N_3356,N_745);
and U5078 (N_5078,N_3396,N_3445);
nand U5079 (N_5079,N_2799,N_613);
xor U5080 (N_5080,N_4003,N_639);
and U5081 (N_5081,N_3390,N_2428);
nand U5082 (N_5082,N_859,N_1938);
nor U5083 (N_5083,N_1404,N_507);
nand U5084 (N_5084,N_1446,N_4861);
nand U5085 (N_5085,N_3015,N_4348);
or U5086 (N_5086,N_4353,N_1296);
or U5087 (N_5087,N_796,N_3814);
nor U5088 (N_5088,N_3240,N_2623);
nand U5089 (N_5089,N_1883,N_1581);
and U5090 (N_5090,N_3738,N_1092);
or U5091 (N_5091,N_4717,N_4967);
nand U5092 (N_5092,N_3123,N_1534);
or U5093 (N_5093,N_800,N_2145);
and U5094 (N_5094,N_4042,N_3388);
nor U5095 (N_5095,N_545,N_4456);
nand U5096 (N_5096,N_1066,N_1876);
nand U5097 (N_5097,N_3187,N_2446);
or U5098 (N_5098,N_4376,N_3690);
or U5099 (N_5099,N_2812,N_1286);
nor U5100 (N_5100,N_111,N_1700);
nand U5101 (N_5101,N_2685,N_4732);
or U5102 (N_5102,N_2600,N_2590);
nor U5103 (N_5103,N_3518,N_1985);
or U5104 (N_5104,N_4696,N_1131);
and U5105 (N_5105,N_1879,N_576);
nand U5106 (N_5106,N_936,N_3364);
nor U5107 (N_5107,N_4008,N_508);
nand U5108 (N_5108,N_3485,N_265);
and U5109 (N_5109,N_4885,N_2040);
nand U5110 (N_5110,N_675,N_2742);
and U5111 (N_5111,N_1114,N_2238);
xnor U5112 (N_5112,N_1759,N_1556);
xor U5113 (N_5113,N_122,N_3360);
nor U5114 (N_5114,N_4934,N_2916);
and U5115 (N_5115,N_4074,N_4163);
or U5116 (N_5116,N_4505,N_3647);
or U5117 (N_5117,N_4453,N_4538);
xor U5118 (N_5118,N_155,N_3822);
or U5119 (N_5119,N_2922,N_2459);
nand U5120 (N_5120,N_3021,N_4905);
nor U5121 (N_5121,N_1885,N_4245);
nor U5122 (N_5122,N_3018,N_2044);
and U5123 (N_5123,N_1062,N_3864);
and U5124 (N_5124,N_131,N_1921);
or U5125 (N_5125,N_2545,N_2887);
or U5126 (N_5126,N_2081,N_4892);
nor U5127 (N_5127,N_2862,N_3632);
or U5128 (N_5128,N_3805,N_3443);
and U5129 (N_5129,N_4034,N_2874);
and U5130 (N_5130,N_1022,N_4817);
and U5131 (N_5131,N_1280,N_2247);
nand U5132 (N_5132,N_2317,N_270);
and U5133 (N_5133,N_4304,N_565);
and U5134 (N_5134,N_4473,N_4557);
nor U5135 (N_5135,N_4691,N_3155);
nor U5136 (N_5136,N_2786,N_531);
nor U5137 (N_5137,N_234,N_4285);
or U5138 (N_5138,N_414,N_4663);
nor U5139 (N_5139,N_1877,N_853);
or U5140 (N_5140,N_3252,N_2487);
nand U5141 (N_5141,N_2429,N_3208);
nand U5142 (N_5142,N_3929,N_2036);
or U5143 (N_5143,N_603,N_4387);
nand U5144 (N_5144,N_4032,N_2163);
and U5145 (N_5145,N_3793,N_103);
or U5146 (N_5146,N_1787,N_496);
nand U5147 (N_5147,N_2813,N_3838);
or U5148 (N_5148,N_3921,N_1095);
or U5149 (N_5149,N_1159,N_2048);
nor U5150 (N_5150,N_3397,N_3667);
and U5151 (N_5151,N_2303,N_3633);
or U5152 (N_5152,N_682,N_714);
or U5153 (N_5153,N_1354,N_4333);
nand U5154 (N_5154,N_599,N_62);
xnor U5155 (N_5155,N_1243,N_2577);
nand U5156 (N_5156,N_1375,N_1496);
nor U5157 (N_5157,N_1997,N_4238);
and U5158 (N_5158,N_815,N_1111);
nand U5159 (N_5159,N_2985,N_3528);
and U5160 (N_5160,N_2548,N_1264);
nand U5161 (N_5161,N_1656,N_3287);
and U5162 (N_5162,N_84,N_2251);
and U5163 (N_5163,N_333,N_1403);
nand U5164 (N_5164,N_4909,N_3450);
nand U5165 (N_5165,N_19,N_3681);
nor U5166 (N_5166,N_3669,N_3501);
nand U5167 (N_5167,N_1955,N_1843);
and U5168 (N_5168,N_2152,N_2219);
or U5169 (N_5169,N_4840,N_4266);
nor U5170 (N_5170,N_2496,N_4476);
nor U5171 (N_5171,N_2403,N_4422);
nor U5172 (N_5172,N_2766,N_712);
or U5173 (N_5173,N_4526,N_871);
nand U5174 (N_5174,N_917,N_3712);
nor U5175 (N_5175,N_23,N_4423);
nor U5176 (N_5176,N_4762,N_3810);
and U5177 (N_5177,N_2783,N_4095);
nor U5178 (N_5178,N_137,N_1423);
nand U5179 (N_5179,N_3612,N_3757);
or U5180 (N_5180,N_1930,N_4484);
nor U5181 (N_5181,N_380,N_2982);
nand U5182 (N_5182,N_4960,N_4436);
and U5183 (N_5183,N_4420,N_2738);
nor U5184 (N_5184,N_4736,N_2903);
nor U5185 (N_5185,N_592,N_4716);
nand U5186 (N_5186,N_2283,N_962);
or U5187 (N_5187,N_1449,N_3089);
nand U5188 (N_5188,N_4994,N_1756);
nor U5189 (N_5189,N_2926,N_1628);
or U5190 (N_5190,N_627,N_4779);
nand U5191 (N_5191,N_4938,N_6);
and U5192 (N_5192,N_4202,N_3271);
or U5193 (N_5193,N_4170,N_1075);
or U5194 (N_5194,N_2382,N_3164);
nor U5195 (N_5195,N_1504,N_1918);
and U5196 (N_5196,N_3590,N_2690);
xnor U5197 (N_5197,N_113,N_3473);
nor U5198 (N_5198,N_2215,N_2104);
or U5199 (N_5199,N_4690,N_1234);
xor U5200 (N_5200,N_2727,N_756);
nor U5201 (N_5201,N_2058,N_392);
nand U5202 (N_5202,N_2527,N_3367);
nand U5203 (N_5203,N_2954,N_2789);
and U5204 (N_5204,N_4150,N_163);
or U5205 (N_5205,N_348,N_1348);
and U5206 (N_5206,N_3602,N_3621);
nand U5207 (N_5207,N_66,N_1542);
nand U5208 (N_5208,N_3185,N_4454);
or U5209 (N_5209,N_3500,N_3503);
or U5210 (N_5210,N_3437,N_896);
and U5211 (N_5211,N_4835,N_1603);
or U5212 (N_5212,N_2996,N_551);
nand U5213 (N_5213,N_1697,N_3512);
nand U5214 (N_5214,N_1817,N_2097);
and U5215 (N_5215,N_4511,N_2881);
nand U5216 (N_5216,N_621,N_334);
and U5217 (N_5217,N_1256,N_1277);
xnor U5218 (N_5218,N_424,N_1056);
or U5219 (N_5219,N_537,N_2935);
nor U5220 (N_5220,N_520,N_2415);
nand U5221 (N_5221,N_2945,N_1755);
nor U5222 (N_5222,N_4860,N_897);
nand U5223 (N_5223,N_568,N_1472);
nor U5224 (N_5224,N_2516,N_886);
or U5225 (N_5225,N_4377,N_126);
nor U5226 (N_5226,N_3327,N_3279);
nand U5227 (N_5227,N_4881,N_1391);
nand U5228 (N_5228,N_3221,N_2355);
nor U5229 (N_5229,N_4046,N_1304);
nor U5230 (N_5230,N_472,N_3657);
xor U5231 (N_5231,N_1861,N_1574);
nand U5232 (N_5232,N_1940,N_4337);
and U5233 (N_5233,N_4528,N_1721);
nand U5234 (N_5234,N_4880,N_2556);
xnor U5235 (N_5235,N_3458,N_3300);
nand U5236 (N_5236,N_560,N_2424);
nand U5237 (N_5237,N_276,N_884);
nand U5238 (N_5238,N_2573,N_4652);
nor U5239 (N_5239,N_116,N_835);
xnor U5240 (N_5240,N_4954,N_4407);
and U5241 (N_5241,N_3978,N_1566);
nand U5242 (N_5242,N_1913,N_1714);
or U5243 (N_5243,N_4187,N_497);
nand U5244 (N_5244,N_2858,N_458);
and U5245 (N_5245,N_3312,N_642);
or U5246 (N_5246,N_3698,N_3919);
nor U5247 (N_5247,N_2805,N_2808);
and U5248 (N_5248,N_1763,N_4253);
or U5249 (N_5249,N_4524,N_2065);
xor U5250 (N_5250,N_4913,N_198);
and U5251 (N_5251,N_4281,N_662);
or U5252 (N_5252,N_4800,N_2185);
and U5253 (N_5253,N_279,N_1462);
nor U5254 (N_5254,N_1715,N_1482);
and U5255 (N_5255,N_3609,N_1591);
nor U5256 (N_5256,N_3147,N_309);
nand U5257 (N_5257,N_3333,N_426);
nor U5258 (N_5258,N_2763,N_41);
and U5259 (N_5259,N_194,N_422);
nor U5260 (N_5260,N_3469,N_4115);
nand U5261 (N_5261,N_700,N_60);
nor U5262 (N_5262,N_2790,N_3525);
or U5263 (N_5263,N_499,N_2677);
nand U5264 (N_5264,N_3523,N_4211);
xor U5265 (N_5265,N_1298,N_1327);
and U5266 (N_5266,N_2328,N_3383);
and U5267 (N_5267,N_1698,N_241);
nand U5268 (N_5268,N_809,N_3951);
or U5269 (N_5269,N_3012,N_4737);
and U5270 (N_5270,N_4059,N_3070);
and U5271 (N_5271,N_2218,N_2363);
nand U5272 (N_5272,N_4445,N_2077);
xor U5273 (N_5273,N_595,N_2171);
xnor U5274 (N_5274,N_425,N_1903);
nor U5275 (N_5275,N_2452,N_1021);
and U5276 (N_5276,N_4513,N_3161);
nor U5277 (N_5277,N_4232,N_1559);
or U5278 (N_5278,N_3131,N_1352);
and U5279 (N_5279,N_1150,N_1179);
nand U5280 (N_5280,N_4590,N_2442);
and U5281 (N_5281,N_1098,N_4598);
nand U5282 (N_5282,N_3836,N_4834);
or U5283 (N_5283,N_4137,N_2759);
xnor U5284 (N_5284,N_3758,N_1405);
or U5285 (N_5285,N_1029,N_908);
and U5286 (N_5286,N_2351,N_3283);
nand U5287 (N_5287,N_2172,N_858);
and U5288 (N_5288,N_2417,N_661);
or U5289 (N_5289,N_1740,N_1690);
or U5290 (N_5290,N_1431,N_1729);
and U5291 (N_5291,N_1905,N_1646);
nor U5292 (N_5292,N_3477,N_1670);
nor U5293 (N_5293,N_794,N_4208);
nand U5294 (N_5294,N_4441,N_3069);
nand U5295 (N_5295,N_2932,N_4323);
nor U5296 (N_5296,N_1276,N_3225);
nor U5297 (N_5297,N_754,N_168);
nand U5298 (N_5298,N_3791,N_2760);
and U5299 (N_5299,N_640,N_2453);
nand U5300 (N_5300,N_4133,N_1710);
or U5301 (N_5301,N_4306,N_1595);
nand U5302 (N_5302,N_856,N_4749);
or U5303 (N_5303,N_3153,N_1223);
nand U5304 (N_5304,N_1228,N_4470);
or U5305 (N_5305,N_1959,N_4279);
nor U5306 (N_5306,N_1198,N_1082);
nor U5307 (N_5307,N_2892,N_4969);
or U5308 (N_5308,N_4096,N_92);
or U5309 (N_5309,N_4290,N_2716);
and U5310 (N_5310,N_4342,N_2663);
and U5311 (N_5311,N_4444,N_813);
and U5312 (N_5312,N_2230,N_1520);
xnor U5313 (N_5313,N_3552,N_4174);
xor U5314 (N_5314,N_1667,N_1568);
and U5315 (N_5315,N_1464,N_2474);
nor U5316 (N_5316,N_3113,N_4111);
nor U5317 (N_5317,N_1068,N_984);
and U5318 (N_5318,N_1932,N_3395);
or U5319 (N_5319,N_2116,N_7);
and U5320 (N_5320,N_1943,N_3946);
and U5321 (N_5321,N_4993,N_3341);
xnor U5322 (N_5322,N_74,N_2937);
or U5323 (N_5323,N_211,N_2774);
or U5324 (N_5324,N_1782,N_1119);
nand U5325 (N_5325,N_4023,N_834);
or U5326 (N_5326,N_1535,N_2306);
nor U5327 (N_5327,N_4125,N_2997);
nand U5328 (N_5328,N_3906,N_183);
xnor U5329 (N_5329,N_1575,N_1407);
or U5330 (N_5330,N_3739,N_3977);
or U5331 (N_5331,N_1696,N_881);
or U5332 (N_5332,N_2602,N_3441);
xor U5333 (N_5333,N_372,N_2906);
nor U5334 (N_5334,N_47,N_159);
nor U5335 (N_5335,N_2193,N_3128);
nor U5336 (N_5336,N_726,N_1703);
xnor U5337 (N_5337,N_1406,N_4918);
and U5338 (N_5338,N_522,N_1996);
xor U5339 (N_5339,N_955,N_352);
or U5340 (N_5340,N_4862,N_4225);
xor U5341 (N_5341,N_4519,N_3868);
or U5342 (N_5342,N_38,N_1726);
and U5343 (N_5343,N_3858,N_1840);
xnor U5344 (N_5344,N_3890,N_3080);
and U5345 (N_5345,N_1383,N_482);
nand U5346 (N_5346,N_1920,N_1013);
and U5347 (N_5347,N_3142,N_2778);
nand U5348 (N_5348,N_518,N_795);
nand U5349 (N_5349,N_1080,N_4108);
and U5350 (N_5350,N_4078,N_3444);
and U5351 (N_5351,N_4038,N_1683);
and U5352 (N_5352,N_1576,N_1505);
or U5353 (N_5353,N_4713,N_4532);
nor U5354 (N_5354,N_2529,N_1866);
and U5355 (N_5355,N_1483,N_3453);
nand U5356 (N_5356,N_4357,N_3220);
and U5357 (N_5357,N_822,N_423);
nand U5358 (N_5358,N_3675,N_2753);
or U5359 (N_5359,N_4567,N_4375);
nor U5360 (N_5360,N_573,N_1160);
and U5361 (N_5361,N_3817,N_2636);
xnor U5362 (N_5362,N_3997,N_68);
nor U5363 (N_5363,N_4801,N_1229);
nand U5364 (N_5364,N_1065,N_4571);
xor U5365 (N_5365,N_4260,N_1799);
nor U5366 (N_5366,N_624,N_611);
or U5367 (N_5367,N_1084,N_618);
and U5368 (N_5368,N_468,N_648);
xnor U5369 (N_5369,N_1000,N_4492);
and U5370 (N_5370,N_3756,N_4400);
nor U5371 (N_5371,N_513,N_1724);
and U5372 (N_5372,N_4248,N_4523);
and U5373 (N_5373,N_1516,N_2398);
and U5374 (N_5374,N_901,N_824);
nor U5375 (N_5375,N_546,N_2338);
or U5376 (N_5376,N_2824,N_3861);
nor U5377 (N_5377,N_2539,N_3957);
nand U5378 (N_5378,N_4916,N_3309);
or U5379 (N_5379,N_3926,N_3373);
and U5380 (N_5380,N_2167,N_2457);
xor U5381 (N_5381,N_3830,N_3952);
nand U5382 (N_5382,N_2223,N_4130);
and U5383 (N_5383,N_3570,N_4241);
and U5384 (N_5384,N_4823,N_21);
or U5385 (N_5385,N_747,N_3120);
or U5386 (N_5386,N_1402,N_3677);
nand U5387 (N_5387,N_4933,N_1509);
nand U5388 (N_5388,N_3983,N_50);
and U5389 (N_5389,N_838,N_1273);
and U5390 (N_5390,N_1239,N_4907);
and U5391 (N_5391,N_805,N_3410);
or U5392 (N_5392,N_4151,N_3857);
nor U5393 (N_5393,N_2706,N_777);
nor U5394 (N_5394,N_2080,N_4575);
and U5395 (N_5395,N_4228,N_3066);
nand U5396 (N_5396,N_4276,N_914);
nand U5397 (N_5397,N_3622,N_3363);
nor U5398 (N_5398,N_3806,N_4043);
nor U5399 (N_5399,N_857,N_3121);
nand U5400 (N_5400,N_1947,N_550);
nor U5401 (N_5401,N_3203,N_4446);
nand U5402 (N_5402,N_3246,N_4251);
nand U5403 (N_5403,N_3627,N_369);
and U5404 (N_5404,N_2035,N_3947);
or U5405 (N_5405,N_2369,N_1832);
nand U5406 (N_5406,N_4540,N_4612);
or U5407 (N_5407,N_4838,N_749);
and U5408 (N_5408,N_464,N_2125);
nor U5409 (N_5409,N_4846,N_1731);
nand U5410 (N_5410,N_2465,N_2427);
and U5411 (N_5411,N_4551,N_2173);
or U5412 (N_5412,N_4010,N_1328);
nand U5413 (N_5413,N_134,N_1676);
nand U5414 (N_5414,N_1481,N_3186);
nor U5415 (N_5415,N_4827,N_3331);
nor U5416 (N_5416,N_79,N_3234);
and U5417 (N_5417,N_2603,N_4468);
nor U5418 (N_5418,N_1798,N_827);
nor U5419 (N_5419,N_3495,N_4961);
or U5420 (N_5420,N_4483,N_1643);
nor U5421 (N_5421,N_1567,N_2066);
xor U5422 (N_5422,N_2454,N_2099);
nand U5423 (N_5423,N_1816,N_680);
or U5424 (N_5424,N_1378,N_4247);
nand U5425 (N_5425,N_1424,N_1887);
nor U5426 (N_5426,N_3050,N_511);
nor U5427 (N_5427,N_1781,N_3435);
and U5428 (N_5428,N_4056,N_3330);
and U5429 (N_5429,N_2003,N_3476);
nor U5430 (N_5430,N_4644,N_3965);
or U5431 (N_5431,N_3299,N_1802);
and U5432 (N_5432,N_2549,N_633);
or U5433 (N_5433,N_1240,N_1162);
and U5434 (N_5434,N_2846,N_4466);
and U5435 (N_5435,N_252,N_4327);
nand U5436 (N_5436,N_1976,N_2803);
nand U5437 (N_5437,N_2784,N_3726);
nor U5438 (N_5438,N_3124,N_538);
nand U5439 (N_5439,N_620,N_2661);
nand U5440 (N_5440,N_4844,N_2501);
nand U5441 (N_5441,N_3903,N_4272);
nand U5442 (N_5442,N_4591,N_4660);
or U5443 (N_5443,N_626,N_2626);
nand U5444 (N_5444,N_4689,N_4877);
xnor U5445 (N_5445,N_2005,N_539);
or U5446 (N_5446,N_678,N_2143);
or U5447 (N_5447,N_1599,N_1102);
nor U5448 (N_5448,N_1360,N_1425);
and U5449 (N_5449,N_1143,N_3201);
nor U5450 (N_5450,N_2168,N_1129);
xor U5451 (N_5451,N_2814,N_898);
nor U5452 (N_5452,N_3544,N_156);
and U5453 (N_5453,N_2358,N_401);
and U5454 (N_5454,N_1904,N_2221);
nand U5455 (N_5455,N_3532,N_514);
nor U5456 (N_5456,N_810,N_1990);
nor U5457 (N_5457,N_4711,N_2385);
nand U5458 (N_5458,N_2232,N_3884);
or U5459 (N_5459,N_1372,N_1408);
nand U5460 (N_5460,N_575,N_3945);
nand U5461 (N_5461,N_3183,N_3350);
or U5462 (N_5462,N_1701,N_952);
or U5463 (N_5463,N_3216,N_1644);
nand U5464 (N_5464,N_1476,N_2581);
or U5465 (N_5465,N_3338,N_3016);
nand U5466 (N_5466,N_4434,N_4282);
nor U5467 (N_5467,N_2000,N_922);
and U5468 (N_5468,N_1350,N_4890);
nor U5469 (N_5469,N_933,N_1569);
nor U5470 (N_5470,N_3024,N_3087);
xor U5471 (N_5471,N_1565,N_2828);
xor U5472 (N_5472,N_3274,N_3212);
or U5473 (N_5473,N_4600,N_4138);
nor U5474 (N_5474,N_2708,N_2816);
nand U5475 (N_5475,N_3031,N_1176);
or U5476 (N_5476,N_3723,N_1422);
nor U5477 (N_5477,N_3852,N_148);
nand U5478 (N_5478,N_1834,N_304);
nor U5479 (N_5479,N_344,N_2121);
or U5480 (N_5480,N_2550,N_1260);
or U5481 (N_5481,N_205,N_1563);
or U5482 (N_5482,N_3956,N_4288);
and U5483 (N_5483,N_250,N_85);
nor U5484 (N_5484,N_3497,N_990);
and U5485 (N_5485,N_2695,N_1460);
nand U5486 (N_5486,N_3874,N_3684);
nand U5487 (N_5487,N_3750,N_1553);
and U5488 (N_5488,N_4797,N_2141);
nand U5489 (N_5489,N_4325,N_128);
xnor U5490 (N_5490,N_2615,N_2295);
or U5491 (N_5491,N_3569,N_4169);
xnor U5492 (N_5492,N_3178,N_4667);
nor U5493 (N_5493,N_873,N_3056);
or U5494 (N_5494,N_287,N_3081);
nor U5495 (N_5495,N_2340,N_214);
nor U5496 (N_5496,N_2830,N_4794);
or U5497 (N_5497,N_3809,N_3301);
xnor U5498 (N_5498,N_3752,N_891);
nand U5499 (N_5499,N_1823,N_2473);
and U5500 (N_5500,N_3154,N_4005);
nor U5501 (N_5501,N_4390,N_4770);
xnor U5502 (N_5502,N_3953,N_1078);
or U5503 (N_5503,N_4087,N_4536);
nor U5504 (N_5504,N_3238,N_3691);
xor U5505 (N_5505,N_2378,N_3037);
nand U5506 (N_5506,N_2068,N_889);
and U5507 (N_5507,N_3589,N_654);
nor U5508 (N_5508,N_1537,N_559);
nor U5509 (N_5509,N_2072,N_619);
nor U5510 (N_5510,N_269,N_2157);
nand U5511 (N_5511,N_1253,N_336);
and U5512 (N_5512,N_3916,N_3559);
nor U5513 (N_5513,N_3470,N_4776);
nor U5514 (N_5514,N_2462,N_2884);
nor U5515 (N_5515,N_2055,N_3454);
xor U5516 (N_5516,N_2112,N_799);
and U5517 (N_5517,N_2201,N_2481);
and U5518 (N_5518,N_2210,N_707);
and U5519 (N_5519,N_1786,N_2523);
and U5520 (N_5520,N_4784,N_4635);
xnor U5521 (N_5521,N_1430,N_4315);
or U5522 (N_5522,N_324,N_4714);
and U5523 (N_5523,N_4610,N_2394);
nor U5524 (N_5524,N_2995,N_3888);
nor U5525 (N_5525,N_2848,N_3992);
nor U5526 (N_5526,N_3659,N_3315);
nand U5527 (N_5527,N_1133,N_3175);
and U5528 (N_5528,N_2655,N_3053);
xor U5529 (N_5529,N_4177,N_281);
or U5530 (N_5530,N_4,N_870);
xnor U5531 (N_5531,N_3839,N_4839);
xor U5532 (N_5532,N_4808,N_4803);
nor U5533 (N_5533,N_1337,N_3872);
nor U5534 (N_5534,N_2861,N_365);
nand U5535 (N_5535,N_4022,N_1181);
or U5536 (N_5536,N_1587,N_1517);
nor U5537 (N_5537,N_2377,N_2633);
xor U5538 (N_5538,N_2019,N_4027);
or U5539 (N_5539,N_4584,N_30);
and U5540 (N_5540,N_25,N_3424);
and U5541 (N_5541,N_114,N_4299);
nand U5542 (N_5542,N_4123,N_4221);
or U5543 (N_5543,N_2469,N_311);
xor U5544 (N_5544,N_2804,N_3352);
or U5545 (N_5545,N_4975,N_1858);
or U5546 (N_5546,N_143,N_4408);
nand U5547 (N_5547,N_461,N_1805);
and U5548 (N_5548,N_3111,N_1043);
xor U5549 (N_5549,N_4608,N_3880);
nand U5550 (N_5550,N_3244,N_2126);
or U5551 (N_5551,N_2261,N_2853);
nor U5552 (N_5552,N_2082,N_2946);
nand U5553 (N_5553,N_902,N_681);
or U5554 (N_5554,N_3819,N_2237);
or U5555 (N_5555,N_3672,N_4307);
nand U5556 (N_5556,N_2924,N_4751);
nand U5557 (N_5557,N_4167,N_1027);
nor U5558 (N_5558,N_803,N_3755);
or U5559 (N_5559,N_3136,N_3150);
nor U5560 (N_5560,N_1088,N_4508);
and U5561 (N_5561,N_1158,N_2129);
nor U5562 (N_5562,N_4274,N_2522);
and U5563 (N_5563,N_581,N_3975);
or U5564 (N_5564,N_4903,N_190);
and U5565 (N_5565,N_1801,N_4521);
nand U5566 (N_5566,N_2255,N_811);
and U5567 (N_5567,N_258,N_3766);
xnor U5568 (N_5568,N_299,N_2497);
nor U5569 (N_5569,N_665,N_1140);
and U5570 (N_5570,N_1982,N_22);
or U5571 (N_5571,N_2046,N_3597);
nand U5572 (N_5572,N_2572,N_552);
nand U5573 (N_5573,N_2645,N_1640);
nor U5574 (N_5574,N_4802,N_1077);
nand U5575 (N_5575,N_2779,N_701);
and U5576 (N_5576,N_2037,N_3002);
nand U5577 (N_5577,N_110,N_2400);
and U5578 (N_5578,N_1901,N_1708);
and U5579 (N_5579,N_3505,N_2967);
nand U5580 (N_5580,N_2478,N_4659);
and U5581 (N_5581,N_437,N_3236);
nor U5582 (N_5582,N_288,N_517);
and U5583 (N_5583,N_1197,N_597);
or U5584 (N_5584,N_2724,N_2153);
nor U5585 (N_5585,N_2692,N_188);
nor U5586 (N_5586,N_2854,N_3889);
or U5587 (N_5587,N_4184,N_3480);
nor U5588 (N_5588,N_2930,N_4688);
nand U5589 (N_5589,N_1992,N_2011);
and U5590 (N_5590,N_487,N_4585);
xnor U5591 (N_5591,N_179,N_3114);
nand U5592 (N_5592,N_2687,N_1771);
and U5593 (N_5593,N_363,N_3353);
or U5594 (N_5594,N_4772,N_1468);
nor U5595 (N_5595,N_3662,N_2697);
or U5596 (N_5596,N_4546,N_3546);
and U5597 (N_5597,N_602,N_1008);
nor U5598 (N_5598,N_169,N_453);
nand U5599 (N_5599,N_4780,N_1467);
or U5600 (N_5600,N_1130,N_2710);
or U5601 (N_5601,N_2386,N_4147);
nor U5602 (N_5602,N_2533,N_2564);
nor U5603 (N_5603,N_443,N_2898);
nor U5604 (N_5604,N_1776,N_2961);
nor U5605 (N_5605,N_1837,N_4421);
or U5606 (N_5606,N_4563,N_3658);
xnor U5607 (N_5607,N_247,N_2594);
and U5608 (N_5608,N_4369,N_4592);
xnor U5609 (N_5609,N_4017,N_4603);
or U5610 (N_5610,N_2815,N_4425);
nor U5611 (N_5611,N_4866,N_1325);
nand U5612 (N_5612,N_3467,N_1463);
and U5613 (N_5613,N_3379,N_2674);
xnor U5614 (N_5614,N_4236,N_2617);
nor U5615 (N_5615,N_3522,N_4578);
and U5616 (N_5616,N_1981,N_1262);
xnor U5617 (N_5617,N_2512,N_2648);
and U5618 (N_5618,N_3253,N_4116);
or U5619 (N_5619,N_2640,N_1550);
nor U5620 (N_5620,N_2693,N_236);
or U5621 (N_5621,N_3526,N_1580);
xnor U5622 (N_5622,N_1110,N_1942);
nand U5623 (N_5623,N_4380,N_1549);
or U5624 (N_5624,N_1370,N_3571);
nand U5625 (N_5625,N_1766,N_2370);
or U5626 (N_5626,N_524,N_1730);
and U5627 (N_5627,N_3170,N_651);
or U5628 (N_5628,N_894,N_361);
xor U5629 (N_5629,N_4235,N_2353);
xnor U5630 (N_5630,N_1259,N_4925);
nand U5631 (N_5631,N_4856,N_3040);
and U5632 (N_5632,N_1597,N_3862);
or U5633 (N_5633,N_1518,N_752);
and U5634 (N_5634,N_863,N_3896);
and U5635 (N_5635,N_1410,N_96);
nor U5636 (N_5636,N_448,N_3222);
and U5637 (N_5637,N_1583,N_3905);
and U5638 (N_5638,N_1164,N_379);
nor U5639 (N_5639,N_2135,N_3387);
nor U5640 (N_5640,N_1344,N_1917);
nor U5641 (N_5641,N_880,N_4873);
nand U5642 (N_5642,N_4386,N_3654);
or U5643 (N_5643,N_833,N_3696);
and U5644 (N_5644,N_4388,N_2580);
and U5645 (N_5645,N_727,N_142);
nand U5646 (N_5646,N_2975,N_899);
or U5647 (N_5647,N_2493,N_1437);
xor U5648 (N_5648,N_2807,N_319);
and U5649 (N_5649,N_2162,N_650);
nand U5650 (N_5650,N_3129,N_3574);
xor U5651 (N_5651,N_2204,N_2981);
or U5652 (N_5652,N_1466,N_4082);
nor U5653 (N_5653,N_4593,N_1532);
or U5654 (N_5654,N_1732,N_4601);
or U5655 (N_5655,N_2764,N_1945);
or U5656 (N_5656,N_4609,N_1833);
or U5657 (N_5657,N_135,N_200);
xor U5658 (N_5658,N_4648,N_956);
and U5659 (N_5659,N_1261,N_3109);
or U5660 (N_5660,N_4155,N_2448);
and U5661 (N_5661,N_1389,N_1039);
or U5662 (N_5662,N_3047,N_2240);
and U5663 (N_5663,N_4746,N_1141);
nor U5664 (N_5664,N_4291,N_1285);
nor U5665 (N_5665,N_2021,N_3734);
and U5666 (N_5666,N_2387,N_1931);
and U5667 (N_5667,N_1663,N_643);
nand U5668 (N_5668,N_1282,N_3648);
nor U5669 (N_5669,N_757,N_3823);
nand U5670 (N_5670,N_2851,N_720);
and U5671 (N_5671,N_191,N_3744);
and U5672 (N_5672,N_948,N_1070);
nor U5673 (N_5673,N_2823,N_4850);
nand U5674 (N_5674,N_2653,N_2091);
nor U5675 (N_5675,N_596,N_3101);
and U5676 (N_5676,N_1807,N_544);
nand U5677 (N_5677,N_2307,N_1845);
and U5678 (N_5678,N_3585,N_2284);
nor U5679 (N_5679,N_4703,N_3117);
nand U5680 (N_5680,N_2672,N_848);
nor U5681 (N_5681,N_4308,N_2542);
or U5682 (N_5682,N_1956,N_1508);
nand U5683 (N_5683,N_1381,N_455);
nor U5684 (N_5684,N_4171,N_1555);
nand U5685 (N_5685,N_2977,N_2656);
or U5686 (N_5686,N_2301,N_4331);
or U5687 (N_5687,N_950,N_320);
and U5688 (N_5688,N_4588,N_4851);
nor U5689 (N_5689,N_571,N_3097);
nor U5690 (N_5690,N_3918,N_2405);
or U5691 (N_5691,N_4863,N_3886);
or U5692 (N_5692,N_3761,N_4162);
and U5693 (N_5693,N_3732,N_1138);
and U5694 (N_5694,N_4643,N_2668);
nand U5695 (N_5695,N_16,N_4200);
or U5696 (N_5696,N_4296,N_2913);
or U5697 (N_5697,N_2318,N_816);
or U5698 (N_5698,N_4481,N_193);
nand U5699 (N_5699,N_242,N_3032);
nand U5700 (N_5700,N_877,N_2467);
and U5701 (N_5701,N_1157,N_2878);
or U5702 (N_5702,N_206,N_1806);
and U5703 (N_5703,N_3515,N_3656);
and U5704 (N_5704,N_3915,N_3248);
nor U5705 (N_5705,N_3984,N_2793);
or U5706 (N_5706,N_478,N_768);
nand U5707 (N_5707,N_3165,N_852);
nand U5708 (N_5708,N_11,N_3082);
nor U5709 (N_5709,N_906,N_2726);
and U5710 (N_5710,N_3751,N_3263);
or U5711 (N_5711,N_4439,N_153);
nor U5712 (N_5712,N_3892,N_2611);
or U5713 (N_5713,N_4902,N_1452);
or U5714 (N_5714,N_2025,N_4520);
and U5715 (N_5715,N_4970,N_3239);
xnor U5716 (N_5716,N_2357,N_186);
nand U5717 (N_5717,N_2897,N_4706);
nor U5718 (N_5718,N_4054,N_2443);
xnor U5719 (N_5719,N_4356,N_4389);
nor U5720 (N_5720,N_3711,N_3736);
nand U5721 (N_5721,N_574,N_1752);
nor U5722 (N_5722,N_1944,N_585);
and U5723 (N_5723,N_88,N_2746);
or U5724 (N_5724,N_4275,N_2147);
nor U5725 (N_5725,N_2253,N_4352);
and U5726 (N_5726,N_2928,N_1744);
and U5727 (N_5727,N_4677,N_4071);
nand U5728 (N_5728,N_1911,N_2298);
and U5729 (N_5729,N_3088,N_4819);
nor U5730 (N_5730,N_2392,N_616);
nor U5731 (N_5731,N_2744,N_4152);
and U5732 (N_5732,N_915,N_2736);
or U5733 (N_5733,N_1478,N_2563);
nor U5734 (N_5734,N_3769,N_3140);
nand U5735 (N_5735,N_1011,N_4870);
or U5736 (N_5736,N_1651,N_1613);
and U5737 (N_5737,N_3763,N_1682);
and U5738 (N_5738,N_735,N_1333);
nand U5739 (N_5739,N_3573,N_1356);
nor U5740 (N_5740,N_3634,N_711);
nand U5741 (N_5741,N_3673,N_4730);
nor U5742 (N_5742,N_532,N_705);
and U5743 (N_5743,N_172,N_3829);
nor U5744 (N_5744,N_1175,N_2811);
and U5745 (N_5745,N_1134,N_431);
nand U5746 (N_5746,N_4795,N_1647);
nor U5747 (N_5747,N_2735,N_3620);
nor U5748 (N_5748,N_175,N_3368);
nor U5749 (N_5749,N_4496,N_1395);
and U5750 (N_5750,N_1543,N_1605);
or U5751 (N_5751,N_4658,N_608);
and U5752 (N_5752,N_2324,N_937);
and U5753 (N_5753,N_1617,N_1018);
nand U5754 (N_5754,N_2666,N_350);
and U5755 (N_5755,N_3972,N_3533);
or U5756 (N_5756,N_1186,N_849);
and U5757 (N_5757,N_529,N_4514);
or U5758 (N_5758,N_4579,N_1725);
nor U5759 (N_5759,N_4028,N_1925);
xnor U5760 (N_5760,N_4666,N_2343);
and U5761 (N_5761,N_4629,N_1737);
and U5762 (N_5762,N_3130,N_3455);
and U5763 (N_5763,N_2341,N_4940);
and U5764 (N_5764,N_2364,N_3325);
nand U5765 (N_5765,N_2749,N_1723);
and U5766 (N_5766,N_3489,N_2734);
or U5767 (N_5767,N_1436,N_2389);
and U5768 (N_5768,N_1954,N_3014);
nor U5769 (N_5769,N_2148,N_1185);
and U5770 (N_5770,N_1991,N_2503);
nand U5771 (N_5771,N_2407,N_4813);
nand U5772 (N_5772,N_1053,N_895);
nand U5773 (N_5773,N_2725,N_4981);
xor U5774 (N_5774,N_4239,N_1914);
nand U5775 (N_5775,N_3232,N_3025);
and U5776 (N_5776,N_3653,N_2605);
or U5777 (N_5777,N_4638,N_4294);
nor U5778 (N_5778,N_2027,N_2175);
or U5779 (N_5779,N_3466,N_3297);
xnor U5780 (N_5780,N_2923,N_2543);
and U5781 (N_5781,N_3762,N_4415);
and U5782 (N_5782,N_932,N_1503);
nor U5783 (N_5783,N_4215,N_1118);
xnor U5784 (N_5784,N_4252,N_2472);
xnor U5785 (N_5785,N_4855,N_2616);
and U5786 (N_5786,N_109,N_150);
nand U5787 (N_5787,N_2120,N_4820);
nand U5788 (N_5788,N_4678,N_634);
and U5789 (N_5789,N_36,N_2090);
nor U5790 (N_5790,N_370,N_2638);
or U5791 (N_5791,N_2559,N_4486);
xor U5792 (N_5792,N_33,N_1124);
nand U5793 (N_5793,N_1457,N_1864);
nor U5794 (N_5794,N_1216,N_490);
and U5795 (N_5795,N_2393,N_2032);
nand U5796 (N_5796,N_2321,N_1623);
nor U5797 (N_5797,N_3019,N_492);
and U5798 (N_5798,N_541,N_1355);
xor U5799 (N_5799,N_2291,N_1025);
and U5800 (N_5800,N_1187,N_1222);
and U5801 (N_5801,N_3507,N_3358);
or U5802 (N_5802,N_2918,N_2630);
or U5803 (N_5803,N_1902,N_1633);
nor U5804 (N_5804,N_1177,N_1828);
and U5805 (N_5805,N_584,N_1872);
nand U5806 (N_5806,N_1188,N_3558);
nand U5807 (N_5807,N_629,N_164);
or U5808 (N_5808,N_2160,N_2972);
or U5809 (N_5809,N_4755,N_430);
or U5810 (N_5810,N_3035,N_1213);
and U5811 (N_5811,N_4504,N_4894);
nand U5812 (N_5812,N_1975,N_2411);
and U5813 (N_5813,N_2676,N_1804);
nand U5814 (N_5814,N_2511,N_4695);
and U5815 (N_5815,N_4748,N_4222);
or U5816 (N_5816,N_3959,N_2568);
nand U5817 (N_5817,N_3378,N_543);
nand U5818 (N_5818,N_3071,N_4611);
nand U5819 (N_5819,N_463,N_15);
nand U5820 (N_5820,N_502,N_3588);
xor U5821 (N_5821,N_1525,N_2319);
nand U5822 (N_5822,N_526,N_178);
xnor U5823 (N_5823,N_3548,N_4103);
nand U5824 (N_5824,N_3943,N_4061);
and U5825 (N_5825,N_641,N_1836);
or U5826 (N_5826,N_3451,N_2541);
or U5827 (N_5827,N_4384,N_2604);
nand U5828 (N_5828,N_1960,N_3530);
or U5829 (N_5829,N_4060,N_1632);
and U5830 (N_5830,N_1868,N_4429);
xor U5831 (N_5831,N_261,N_2372);
xnor U5832 (N_5832,N_4766,N_3679);
xor U5833 (N_5833,N_4487,N_104);
and U5834 (N_5834,N_2907,N_152);
xnor U5835 (N_5835,N_2436,N_3777);
or U5836 (N_5836,N_670,N_1322);
nor U5837 (N_5837,N_4119,N_1358);
nand U5838 (N_5838,N_120,N_4782);
nor U5839 (N_5839,N_2199,N_4080);
nor U5840 (N_5840,N_326,N_2277);
or U5841 (N_5841,N_3639,N_1637);
nand U5842 (N_5842,N_2991,N_2711);
and U5843 (N_5843,N_1512,N_436);
xnor U5844 (N_5844,N_2499,N_2988);
nor U5845 (N_5845,N_3020,N_3365);
and U5846 (N_5846,N_4604,N_3556);
nand U5847 (N_5847,N_4343,N_325);
nor U5848 (N_5848,N_1631,N_1671);
xor U5849 (N_5849,N_450,N_2339);
nand U5850 (N_5850,N_530,N_4411);
nor U5851 (N_5851,N_3345,N_4895);
nand U5852 (N_5852,N_3270,N_4530);
and U5853 (N_5853,N_4745,N_1953);
nand U5854 (N_5854,N_3979,N_495);
nand U5855 (N_5855,N_1047,N_1346);
nand U5856 (N_5856,N_912,N_2519);
nand U5857 (N_5857,N_980,N_949);
nor U5858 (N_5858,N_81,N_2546);
and U5859 (N_5859,N_3816,N_147);
nand U5860 (N_5860,N_2592,N_2484);
nor U5861 (N_5861,N_0,N_2004);
or U5862 (N_5862,N_2280,N_4460);
nand U5863 (N_5863,N_4107,N_1783);
and U5864 (N_5864,N_2151,N_841);
and U5865 (N_5865,N_4219,N_535);
or U5866 (N_5866,N_4668,N_3870);
nand U5867 (N_5867,N_1906,N_2045);
or U5868 (N_5868,N_3423,N_2263);
nand U5869 (N_5869,N_2624,N_2041);
and U5870 (N_5870,N_623,N_4930);
and U5871 (N_5871,N_1681,N_3614);
nand U5872 (N_5872,N_1849,N_2226);
nor U5873 (N_5873,N_2883,N_3431);
nor U5874 (N_5874,N_666,N_407);
nor U5875 (N_5875,N_758,N_4495);
and U5876 (N_5876,N_1939,N_3651);
and U5877 (N_5877,N_695,N_3776);
nand U5878 (N_5878,N_2409,N_2601);
nor U5879 (N_5879,N_3033,N_1009);
nand U5880 (N_5880,N_1558,N_2567);
or U5881 (N_5881,N_4565,N_1146);
xnor U5882 (N_5882,N_237,N_3964);
or U5883 (N_5883,N_3256,N_579);
and U5884 (N_5884,N_3875,N_2801);
nand U5885 (N_5885,N_3433,N_393);
or U5886 (N_5886,N_3421,N_2258);
nor U5887 (N_5887,N_3250,N_3567);
xnor U5888 (N_5888,N_812,N_2132);
nor U5889 (N_5889,N_2857,N_4879);
and U5890 (N_5890,N_3860,N_105);
or U5891 (N_5891,N_4631,N_4092);
xnor U5892 (N_5892,N_4273,N_4812);
and U5893 (N_5893,N_4807,N_98);
nor U5894 (N_5894,N_3366,N_2553);
or U5895 (N_5895,N_847,N_1317);
xor U5896 (N_5896,N_1538,N_2198);
nor U5897 (N_5897,N_3463,N_685);
nand U5898 (N_5898,N_4595,N_2115);
nand U5899 (N_5899,N_262,N_275);
nand U5900 (N_5900,N_4413,N_1894);
xor U5901 (N_5901,N_2712,N_2085);
and U5902 (N_5902,N_2445,N_3354);
or U5903 (N_5903,N_391,N_4959);
or U5904 (N_5904,N_1855,N_4742);
and U5905 (N_5905,N_1362,N_2698);
or U5906 (N_5906,N_4623,N_4878);
or U5907 (N_5907,N_4442,N_1035);
nor U5908 (N_5908,N_4100,N_49);
and U5909 (N_5909,N_2835,N_3260);
and U5910 (N_5910,N_1202,N_3063);
nor U5911 (N_5911,N_2194,N_3092);
and U5912 (N_5912,N_3780,N_488);
or U5913 (N_5913,N_1401,N_4679);
or U5914 (N_5914,N_1742,N_2901);
or U5915 (N_5915,N_2155,N_4475);
xnor U5916 (N_5916,N_4882,N_3599);
xor U5917 (N_5917,N_1214,N_3430);
or U5918 (N_5918,N_45,N_4383);
nor U5919 (N_5919,N_820,N_4589);
and U5920 (N_5920,N_4392,N_2701);
xor U5921 (N_5921,N_1863,N_208);
nand U5922 (N_5922,N_2715,N_3554);
and U5923 (N_5923,N_2688,N_1747);
or U5924 (N_5924,N_1511,N_3475);
xnor U5925 (N_5925,N_282,N_1664);
nor U5926 (N_5926,N_4173,N_4602);
and U5927 (N_5927,N_3459,N_4833);
nor U5928 (N_5928,N_3169,N_3180);
and U5929 (N_5929,N_4915,N_4550);
nor U5930 (N_5930,N_2356,N_3010);
xnor U5931 (N_5931,N_2113,N_3909);
nand U5932 (N_5932,N_4110,N_2180);
nor U5933 (N_5933,N_118,N_385);
and U5934 (N_5934,N_1012,N_1748);
nand U5935 (N_5935,N_2836,N_1366);
and U5936 (N_5936,N_3068,N_3564);
nand U5937 (N_5937,N_4535,N_3211);
nand U5938 (N_5938,N_4464,N_3340);
xnor U5939 (N_5939,N_4664,N_2380);
and U5940 (N_5940,N_2195,N_2787);
and U5941 (N_5941,N_3697,N_2719);
and U5942 (N_5942,N_4831,N_4854);
nand U5943 (N_5943,N_2552,N_1170);
xnor U5944 (N_5944,N_1588,N_2144);
or U5945 (N_5945,N_4210,N_3258);
nor U5946 (N_5946,N_2314,N_3837);
or U5947 (N_5947,N_3038,N_4417);
and U5948 (N_5948,N_505,N_1526);
nand U5949 (N_5949,N_3408,N_3176);
nand U5950 (N_5950,N_3706,N_3355);
or U5951 (N_5951,N_946,N_1384);
and U5952 (N_5952,N_1332,N_1850);
nand U5953 (N_5953,N_4560,N_4091);
or U5954 (N_5954,N_878,N_2078);
nand U5955 (N_5955,N_12,N_3103);
and U5956 (N_5956,N_1770,N_787);
nor U5957 (N_5957,N_2776,N_2976);
nand U5958 (N_5958,N_4948,N_3949);
nor U5959 (N_5959,N_4491,N_2822);
xnor U5960 (N_5960,N_2875,N_4312);
nor U5961 (N_5961,N_1448,N_4372);
nand U5962 (N_5962,N_127,N_3643);
or U5963 (N_5963,N_2788,N_1015);
nor U5964 (N_5964,N_3581,N_2589);
and U5965 (N_5965,N_219,N_4723);
or U5966 (N_5966,N_4726,N_1417);
nand U5967 (N_5967,N_704,N_2494);
nor U5968 (N_5968,N_1922,N_709);
or U5969 (N_5969,N_1586,N_3280);
xor U5970 (N_5970,N_2242,N_3490);
nand U5971 (N_5971,N_4165,N_4172);
xnor U5972 (N_5972,N_710,N_2754);
and U5973 (N_5973,N_3179,N_1621);
nand U5974 (N_5974,N_3302,N_4891);
and U5975 (N_5975,N_3247,N_4506);
nand U5976 (N_5976,N_742,N_1666);
nand U5977 (N_5977,N_4156,N_2302);
nand U5978 (N_5978,N_2547,N_3737);
xnor U5979 (N_5979,N_297,N_4287);
xor U5980 (N_5980,N_387,N_3703);
xor U5981 (N_5981,N_1795,N_345);
nor U5982 (N_5982,N_161,N_246);
and U5983 (N_5983,N_851,N_1361);
and U5984 (N_5984,N_3775,N_4843);
nand U5985 (N_5985,N_4783,N_3036);
and U5986 (N_5986,N_3141,N_3023);
nand U5987 (N_5987,N_124,N_4697);
xor U5988 (N_5988,N_197,N_1297);
xnor U5989 (N_5989,N_398,N_1238);
nor U5990 (N_5990,N_1058,N_2350);
nor U5991 (N_5991,N_1257,N_840);
nand U5992 (N_5992,N_773,N_4135);
xor U5993 (N_5993,N_2154,N_4625);
and U5994 (N_5994,N_2422,N_719);
and U5995 (N_5995,N_2517,N_1582);
nor U5996 (N_5996,N_3724,N_255);
or U5997 (N_5997,N_1987,N_429);
nor U5998 (N_5998,N_2050,N_1052);
or U5999 (N_5999,N_741,N_4710);
xor U6000 (N_6000,N_2057,N_3867);
and U6001 (N_6001,N_843,N_4867);
or U6002 (N_6002,N_772,N_2447);
or U6003 (N_6003,N_3831,N_3191);
nor U6004 (N_6004,N_527,N_2964);
nor U6005 (N_6005,N_1974,N_397);
or U6006 (N_6006,N_1329,N_4767);
or U6007 (N_6007,N_2012,N_1074);
or U6008 (N_6008,N_4858,N_2855);
or U6009 (N_6009,N_4928,N_4305);
and U6010 (N_6010,N_2384,N_2239);
nand U6011 (N_6011,N_2287,N_3417);
nor U6012 (N_6012,N_1612,N_3954);
nand U6013 (N_6013,N_2970,N_1694);
and U6014 (N_6014,N_3122,N_4196);
or U6015 (N_6015,N_3745,N_4267);
xor U6016 (N_6016,N_4686,N_2294);
nand U6017 (N_6017,N_4471,N_176);
xnor U6018 (N_6018,N_427,N_3674);
nor U6019 (N_6019,N_4621,N_2250);
nor U6020 (N_6020,N_3660,N_3869);
and U6021 (N_6021,N_672,N_2820);
nand U6022 (N_6022,N_2304,N_2311);
and U6023 (N_6023,N_4049,N_506);
nor U6024 (N_6024,N_1353,N_739);
nor U6025 (N_6025,N_2513,N_1891);
nand U6026 (N_6026,N_4378,N_689);
nand U6027 (N_6027,N_1301,N_4157);
nand U6028 (N_6028,N_2460,N_323);
xor U6029 (N_6029,N_2274,N_4271);
nand U6030 (N_6030,N_1290,N_781);
nand U6031 (N_6031,N_1882,N_842);
xnor U6032 (N_6032,N_558,N_3305);
or U6033 (N_6033,N_4009,N_2896);
nand U6034 (N_6034,N_1003,N_4786);
nor U6035 (N_6035,N_473,N_1203);
and U6036 (N_6036,N_3172,N_4908);
and U6037 (N_6037,N_3091,N_3486);
or U6038 (N_6038,N_1416,N_1428);
and U6039 (N_6039,N_4556,N_4153);
or U6040 (N_6040,N_435,N_1983);
nor U6041 (N_6041,N_874,N_4842);
or U6042 (N_6042,N_2079,N_3107);
or U6043 (N_6043,N_4154,N_3649);
nand U6044 (N_6044,N_4708,N_3223);
and U6045 (N_6045,N_2395,N_2686);
and U6046 (N_6046,N_1263,N_3770);
nor U6047 (N_6047,N_1429,N_4370);
or U6048 (N_6048,N_2980,N_1841);
nand U6049 (N_6049,N_4498,N_652);
or U6050 (N_6050,N_3935,N_4278);
nand U6051 (N_6051,N_3578,N_1399);
nor U6052 (N_6052,N_2618,N_3291);
xnor U6053 (N_6053,N_4426,N_3871);
nor U6054 (N_6054,N_70,N_3605);
and U6055 (N_6055,N_888,N_2176);
nor U6056 (N_6056,N_244,N_73);
and U6057 (N_6057,N_4175,N_3587);
nor U6058 (N_6058,N_4971,N_3815);
nor U6059 (N_6059,N_274,N_716);
and U6060 (N_6060,N_2515,N_4852);
xor U6061 (N_6061,N_2188,N_819);
and U6062 (N_6062,N_420,N_1247);
or U6063 (N_6063,N_4326,N_1097);
or U6064 (N_6064,N_1103,N_3343);
nor U6065 (N_6065,N_1374,N_1321);
nor U6066 (N_6066,N_4364,N_1305);
and U6067 (N_6067,N_4131,N_2635);
or U6068 (N_6068,N_804,N_4330);
xnor U6069 (N_6069,N_1010,N_75);
nor U6070 (N_6070,N_3096,N_3462);
xor U6071 (N_6071,N_3439,N_4507);
nand U6072 (N_6072,N_729,N_1705);
and U6073 (N_6073,N_3266,N_2641);
xor U6074 (N_6074,N_577,N_3406);
nand U6075 (N_6075,N_2437,N_3553);
or U6076 (N_6076,N_3700,N_4007);
and U6077 (N_6077,N_4791,N_2335);
xnor U6078 (N_6078,N_2915,N_358);
nor U6079 (N_6079,N_4923,N_483);
and U6080 (N_6080,N_4639,N_1768);
nor U6081 (N_6081,N_4806,N_3704);
or U6082 (N_6082,N_4735,N_1712);
nor U6083 (N_6083,N_4682,N_3963);
nand U6084 (N_6084,N_3743,N_1411);
and U6085 (N_6085,N_4303,N_4753);
and U6086 (N_6086,N_2271,N_1524);
nor U6087 (N_6087,N_2882,N_3855);
and U6088 (N_6088,N_3197,N_2627);
nor U6089 (N_6089,N_760,N_605);
nor U6090 (N_6090,N_376,N_4616);
or U6091 (N_6091,N_2101,N_2229);
or U6092 (N_6092,N_961,N_2560);
xor U6093 (N_6093,N_3938,N_2264);
and U6094 (N_6094,N_4662,N_3292);
or U6095 (N_6095,N_728,N_40);
nand U6096 (N_6096,N_4641,N_2498);
nand U6097 (N_6097,N_1691,N_2709);
xnor U6098 (N_6098,N_1758,N_4906);
xor U6099 (N_6099,N_1552,N_1501);
and U6100 (N_6100,N_1336,N_1166);
nor U6101 (N_6101,N_4246,N_3231);
xor U6102 (N_6102,N_4986,N_1284);
and U6103 (N_6103,N_2433,N_1811);
nor U6104 (N_6104,N_4924,N_1979);
nand U6105 (N_6105,N_4740,N_307);
or U6106 (N_6106,N_1420,N_174);
xnor U6107 (N_6107,N_1642,N_3230);
or U6108 (N_6108,N_3611,N_285);
nor U6109 (N_6109,N_2100,N_3449);
or U6110 (N_6110,N_1966,N_600);
or U6111 (N_6111,N_3143,N_2732);
and U6112 (N_6112,N_1139,N_1746);
nor U6113 (N_6113,N_1196,N_4197);
and U6114 (N_6114,N_2818,N_121);
or U6115 (N_6115,N_3885,N_1809);
and U6116 (N_6116,N_586,N_1827);
and U6117 (N_6117,N_4586,N_1044);
nand U6118 (N_6118,N_2059,N_885);
nor U6119 (N_6119,N_1028,N_1451);
xor U6120 (N_6120,N_1412,N_4773);
nor U6121 (N_6121,N_3790,N_1604);
and U6122 (N_6122,N_3409,N_1036);
and U6123 (N_6123,N_4161,N_4544);
xor U6124 (N_6124,N_2245,N_2485);
nor U6125 (N_6125,N_1860,N_3773);
nor U6126 (N_6126,N_2863,N_4945);
or U6127 (N_6127,N_913,N_2020);
nor U6128 (N_6128,N_4642,N_2528);
nor U6129 (N_6129,N_4929,N_3811);
xnor U6130 (N_6130,N_2780,N_1856);
nor U6131 (N_6131,N_3645,N_390);
or U6132 (N_6132,N_1073,N_87);
and U6133 (N_6133,N_2762,N_3472);
and U6134 (N_6134,N_2421,N_2755);
nor U6135 (N_6135,N_4811,N_4292);
or U6136 (N_6136,N_360,N_1040);
and U6137 (N_6137,N_1560,N_2254);
nor U6138 (N_6138,N_3995,N_3200);
and U6139 (N_6139,N_2259,N_4139);
nand U6140 (N_6140,N_1600,N_9);
nor U6141 (N_6141,N_2507,N_4968);
and U6142 (N_6142,N_1523,N_3856);
nand U6143 (N_6143,N_2330,N_3375);
or U6144 (N_6144,N_4622,N_1502);
and U6145 (N_6145,N_4626,N_1934);
or U6146 (N_6146,N_4599,N_3126);
nor U6147 (N_6147,N_4572,N_1283);
nand U6148 (N_6148,N_1442,N_536);
nor U6149 (N_6149,N_1859,N_3715);
nand U6150 (N_6150,N_4401,N_1785);
nor U6151 (N_6151,N_3407,N_2730);
and U6152 (N_6152,N_1208,N_3181);
xor U6153 (N_6153,N_312,N_4769);
nand U6154 (N_6154,N_125,N_1192);
nand U6155 (N_6155,N_83,N_189);
nor U6156 (N_6156,N_867,N_4674);
nor U6157 (N_6157,N_731,N_1315);
or U6158 (N_6158,N_4898,N_469);
and U6159 (N_6159,N_2936,N_4789);
or U6160 (N_6160,N_3318,N_1414);
or U6161 (N_6161,N_3389,N_3269);
or U6162 (N_6162,N_3646,N_2187);
nand U6163 (N_6163,N_4050,N_987);
or U6164 (N_6164,N_184,N_257);
and U6165 (N_6165,N_3127,N_1268);
or U6166 (N_6166,N_4265,N_97);
and U6167 (N_6167,N_1968,N_617);
or U6168 (N_6168,N_4250,N_1144);
and U6169 (N_6169,N_3579,N_100);
and U6170 (N_6170,N_480,N_2593);
and U6171 (N_6171,N_3391,N_3400);
and U6172 (N_6172,N_4318,N_1657);
nand U6173 (N_6173,N_954,N_4438);
or U6174 (N_6174,N_892,N_4068);
nand U6175 (N_6175,N_3928,N_782);
and U6176 (N_6176,N_4646,N_2844);
nand U6177 (N_6177,N_4494,N_1122);
and U6178 (N_6178,N_3492,N_1619);
nand U6179 (N_6179,N_1037,N_3626);
xor U6180 (N_6180,N_784,N_377);
nand U6181 (N_6181,N_3261,N_562);
and U6182 (N_6182,N_456,N_4431);
nor U6183 (N_6183,N_3618,N_2234);
nand U6184 (N_6184,N_4704,N_2943);
and U6185 (N_6185,N_3218,N_2087);
and U6186 (N_6186,N_994,N_801);
or U6187 (N_6187,N_1760,N_440);
nor U6188 (N_6188,N_2056,N_1461);
xor U6189 (N_6189,N_2888,N_3808);
or U6190 (N_6190,N_1680,N_3043);
nand U6191 (N_6191,N_2297,N_375);
nand U6192 (N_6192,N_2531,N_1293);
nor U6193 (N_6193,N_3064,N_2610);
nand U6194 (N_6194,N_2957,N_2053);
nand U6195 (N_6195,N_4409,N_4984);
xor U6196 (N_6196,N_4778,N_366);
nor U6197 (N_6197,N_1156,N_2643);
nor U6198 (N_6198,N_99,N_1394);
or U6199 (N_6199,N_4160,N_2014);
xor U6200 (N_6200,N_732,N_167);
and U6201 (N_6201,N_2299,N_3098);
and U6202 (N_6202,N_78,N_475);
and U6203 (N_6203,N_4112,N_267);
or U6204 (N_6204,N_1493,N_2345);
and U6205 (N_6205,N_3923,N_2146);
and U6206 (N_6206,N_158,N_4242);
nand U6207 (N_6207,N_4897,N_1686);
nor U6208 (N_6208,N_2684,N_926);
and U6209 (N_6209,N_1544,N_2051);
and U6210 (N_6210,N_1450,N_3873);
and U6211 (N_6211,N_762,N_4543);
and U6212 (N_6212,N_519,N_201);
and U6213 (N_6213,N_3996,N_3190);
nor U6214 (N_6214,N_1014,N_2827);
nand U6215 (N_6215,N_4430,N_4633);
and U6216 (N_6216,N_4394,N_2741);
or U6217 (N_6217,N_1246,N_3993);
nand U6218 (N_6218,N_628,N_1984);
xor U6219 (N_6219,N_2673,N_2929);
or U6220 (N_6220,N_1051,N_3676);
nand U6221 (N_6221,N_4896,N_3547);
nand U6222 (N_6222,N_4300,N_839);
and U6223 (N_6223,N_3377,N_1369);
nand U6224 (N_6224,N_2182,N_4195);
nand U6225 (N_6225,N_1045,N_2909);
and U6226 (N_6226,N_1838,N_1441);
and U6227 (N_6227,N_3917,N_876);
or U6228 (N_6228,N_3604,N_3663);
nor U6229 (N_6229,N_3630,N_2444);
or U6230 (N_6230,N_1241,N_1881);
nand U6231 (N_6231,N_4432,N_2959);
nor U6232 (N_6232,N_3251,N_3065);
nand U6233 (N_6233,N_1397,N_4113);
xnor U6234 (N_6234,N_1753,N_3799);
nor U6235 (N_6235,N_3052,N_862);
or U6236 (N_6236,N_733,N_780);
and U6237 (N_6237,N_4497,N_4069);
nor U6238 (N_6238,N_2191,N_2177);
nor U6239 (N_6239,N_1825,N_343);
and U6240 (N_6240,N_4217,N_4731);
or U6241 (N_6241,N_3334,N_2293);
nor U6242 (N_6242,N_3137,N_1209);
or U6243 (N_6243,N_4205,N_459);
nor U6244 (N_6244,N_2905,N_1419);
nand U6245 (N_6245,N_1669,N_4630);
or U6246 (N_6246,N_686,N_1099);
nand U6247 (N_6247,N_1132,N_2984);
and U6248 (N_6248,N_4015,N_3268);
and U6249 (N_6249,N_4284,N_4081);
nor U6250 (N_6250,N_694,N_1639);
nand U6251 (N_6251,N_943,N_919);
nor U6252 (N_6252,N_2885,N_1529);
and U6253 (N_6253,N_4057,N_3344);
nor U6254 (N_6254,N_4295,N_1635);
or U6255 (N_6255,N_2562,N_3296);
or U6256 (N_6256,N_825,N_4729);
xor U6257 (N_6257,N_3642,N_767);
nand U6258 (N_6258,N_4374,N_1790);
nor U6259 (N_6259,N_3705,N_1506);
nand U6260 (N_6260,N_2475,N_4011);
or U6261 (N_6261,N_4884,N_4818);
and U6262 (N_6262,N_1818,N_4796);
or U6263 (N_6263,N_4121,N_3974);
nor U6264 (N_6264,N_868,N_676);
and U6265 (N_6265,N_4382,N_1439);
or U6266 (N_6266,N_1421,N_751);
or U6267 (N_6267,N_3159,N_2272);
nand U6268 (N_6268,N_1191,N_3276);
xnor U6269 (N_6269,N_3600,N_4018);
nor U6270 (N_6270,N_4428,N_2578);
or U6271 (N_6271,N_3278,N_3493);
nor U6272 (N_6272,N_2076,N_593);
nand U6273 (N_6273,N_4001,N_240);
and U6274 (N_6274,N_4349,N_2696);
nand U6275 (N_6275,N_4654,N_4105);
nand U6276 (N_6276,N_303,N_1254);
xor U6277 (N_6277,N_555,N_2756);
nor U6278 (N_6278,N_4194,N_3393);
or U6279 (N_6279,N_39,N_4321);
and U6280 (N_6280,N_2834,N_1224);
and U6281 (N_6281,N_1964,N_383);
nor U6282 (N_6282,N_4063,N_1636);
and U6283 (N_6283,N_3517,N_4874);
or U6284 (N_6284,N_927,N_882);
nand U6285 (N_6285,N_2096,N_4218);
or U6286 (N_6286,N_1865,N_1528);
and U6287 (N_6287,N_3541,N_1042);
xor U6288 (N_6288,N_808,N_3607);
nand U6289 (N_6289,N_2649,N_3351);
xnor U6290 (N_6290,N_4213,N_3555);
or U6291 (N_6291,N_743,N_2948);
nor U6292 (N_6292,N_2067,N_4334);
nand U6293 (N_6293,N_3196,N_561);
xor U6294 (N_6294,N_1085,N_4310);
xnor U6295 (N_6295,N_3742,N_4360);
nand U6296 (N_6296,N_3595,N_295);
xor U6297 (N_6297,N_1857,N_4705);
xnor U6298 (N_6298,N_1135,N_1433);
or U6299 (N_6299,N_2670,N_2292);
nand U6300 (N_6300,N_1852,N_332);
nand U6301 (N_6301,N_2376,N_2583);
nor U6302 (N_6302,N_1148,N_1668);
and U6303 (N_6303,N_2877,N_3987);
xnor U6304 (N_6304,N_3813,N_3741);
nor U6305 (N_6305,N_4917,N_3285);
nor U6306 (N_6306,N_854,N_77);
nand U6307 (N_6307,N_4826,N_649);
or U6308 (N_6308,N_3157,N_4712);
and U6309 (N_6309,N_4692,N_3058);
and U6310 (N_6310,N_521,N_3594);
nor U6311 (N_6311,N_129,N_3243);
xnor U6312 (N_6312,N_3907,N_4953);
and U6313 (N_6313,N_93,N_4203);
nor U6314 (N_6314,N_1962,N_1294);
nand U6315 (N_6315,N_489,N_2699);
nand U6316 (N_6316,N_3820,N_1453);
nor U6317 (N_6317,N_4365,N_1844);
nand U6318 (N_6318,N_976,N_4582);
nand U6319 (N_6319,N_2678,N_2646);
nor U6320 (N_6320,N_4256,N_3342);
nand U6321 (N_6321,N_846,N_1091);
nand U6322 (N_6322,N_2028,N_3937);
or U6323 (N_6323,N_1963,N_337);
and U6324 (N_6324,N_2026,N_4359);
nor U6325 (N_6325,N_4559,N_1456);
and U6326 (N_6326,N_2483,N_4927);
xor U6327 (N_6327,N_2270,N_2480);
xor U6328 (N_6328,N_1207,N_3148);
nand U6329 (N_6329,N_4233,N_844);
xor U6330 (N_6330,N_4176,N_4371);
and U6331 (N_6331,N_2671,N_3787);
and U6332 (N_6332,N_408,N_4191);
nand U6333 (N_6333,N_1998,N_3825);
and U6334 (N_6334,N_3687,N_1720);
xnor U6335 (N_6335,N_2336,N_3692);
nor U6336 (N_6336,N_2795,N_1116);
or U6337 (N_6337,N_1057,N_4738);
and U6338 (N_6338,N_4065,N_37);
nor U6339 (N_6339,N_3099,N_3237);
nor U6340 (N_6340,N_2435,N_2365);
nor U6341 (N_6341,N_3850,N_1292);
nand U6342 (N_6342,N_1585,N_4120);
nand U6343 (N_6343,N_4366,N_3460);
or U6344 (N_6344,N_1059,N_4424);
and U6345 (N_6345,N_149,N_4825);
nand U6346 (N_6346,N_3303,N_2279);
and U6347 (N_6347,N_4293,N_442);
or U6348 (N_6348,N_1822,N_2178);
or U6349 (N_6349,N_2114,N_2571);
and U6350 (N_6350,N_3527,N_786);
and U6351 (N_6351,N_1026,N_182);
and U6352 (N_6352,N_4619,N_4747);
nor U6353 (N_6353,N_2266,N_1492);
or U6354 (N_6354,N_939,N_1624);
xor U6355 (N_6355,N_2893,N_1554);
nor U6356 (N_6356,N_3778,N_196);
xnor U6357 (N_6357,N_974,N_91);
or U6358 (N_6358,N_2642,N_210);
nor U6359 (N_6359,N_1978,N_1081);
xnor U6360 (N_6360,N_2508,N_1190);
xnor U6361 (N_6361,N_4026,N_1654);
nand U6362 (N_6362,N_359,N_2942);
or U6363 (N_6363,N_289,N_2276);
nand U6364 (N_6364,N_2904,N_3385);
xor U6365 (N_6365,N_2591,N_2309);
or U6366 (N_6366,N_106,N_667);
xnor U6367 (N_6367,N_27,N_1183);
nand U6368 (N_6368,N_4728,N_180);
nand U6369 (N_6369,N_1061,N_2665);
nand U6370 (N_6370,N_4587,N_4570);
nand U6371 (N_6371,N_4073,N_2477);
nor U6372 (N_6372,N_4501,N_3980);
nor U6373 (N_6373,N_696,N_71);
and U6374 (N_6374,N_133,N_4914);
and U6375 (N_6375,N_893,N_730);
nand U6376 (N_6376,N_3721,N_3308);
and U6377 (N_6377,N_1622,N_2296);
nand U6378 (N_6378,N_1871,N_3843);
nor U6379 (N_6379,N_2468,N_4490);
and U6380 (N_6380,N_1237,N_1634);
and U6381 (N_6381,N_447,N_4030);
nor U6382 (N_6382,N_3879,N_1539);
nor U6383 (N_6383,N_1609,N_1115);
or U6384 (N_6384,N_722,N_1513);
nor U6385 (N_6385,N_3328,N_1778);
or U6386 (N_6386,N_3536,N_3095);
and U6387 (N_6387,N_3022,N_942);
xor U6388 (N_6388,N_1153,N_2938);
and U6389 (N_6389,N_3910,N_4974);
nor U6390 (N_6390,N_1434,N_1626);
nand U6391 (N_6391,N_53,N_4920);
nor U6392 (N_6392,N_4012,N_3479);
and U6393 (N_6393,N_2821,N_3655);
and U6394 (N_6394,N_433,N_1440);
or U6395 (N_6395,N_13,N_2894);
nand U6396 (N_6396,N_3988,N_1465);
xor U6397 (N_6397,N_4164,N_2524);
and U6398 (N_6398,N_3193,N_1848);
nand U6399 (N_6399,N_2802,N_3084);
nand U6400 (N_6400,N_4485,N_746);
nor U6401 (N_6401,N_4725,N_1899);
or U6402 (N_6402,N_2248,N_3976);
and U6403 (N_6403,N_1614,N_446);
nand U6404 (N_6404,N_2891,N_3812);
or U6405 (N_6405,N_4298,N_3740);
nor U6406 (N_6406,N_441,N_2718);
and U6407 (N_6407,N_3414,N_548);
nand U6408 (N_6408,N_8,N_637);
and U6409 (N_6409,N_1762,N_2700);
xor U6410 (N_6410,N_3306,N_1151);
nor U6411 (N_6411,N_415,N_1527);
or U6412 (N_6412,N_2360,N_4992);
nand U6413 (N_6413,N_86,N_1090);
nand U6414 (N_6414,N_3102,N_185);
and U6415 (N_6415,N_2207,N_3754);
nand U6416 (N_6416,N_2375,N_4700);
and U6417 (N_6417,N_1249,N_44);
nand U6418 (N_6418,N_3348,N_738);
nor U6419 (N_6419,N_4655,N_3399);
nand U6420 (N_6420,N_989,N_4410);
nor U6421 (N_6421,N_2257,N_3339);
or U6422 (N_6422,N_4212,N_4344);
and U6423 (N_6423,N_3749,N_4316);
nor U6424 (N_6424,N_2420,N_2606);
nand U6425 (N_6425,N_4226,N_1002);
and U6426 (N_6426,N_3982,N_2064);
and U6427 (N_6427,N_2737,N_2220);
or U6428 (N_6428,N_515,N_3313);
and U6429 (N_6429,N_3420,N_4542);
or U6430 (N_6430,N_1189,N_770);
nand U6431 (N_6431,N_2010,N_4396);
or U6432 (N_6432,N_4618,N_1432);
and U6433 (N_6433,N_4313,N_1929);
nand U6434 (N_6434,N_4037,N_4865);
and U6435 (N_6435,N_3832,N_4014);
xor U6436 (N_6436,N_4672,N_2414);
xnor U6437 (N_6437,N_1086,N_3257);
nand U6438 (N_6438,N_903,N_2920);
nand U6439 (N_6439,N_1531,N_4950);
and U6440 (N_6440,N_4988,N_154);
xor U6441 (N_6441,N_1266,N_1032);
nand U6442 (N_6442,N_4214,N_3055);
or U6443 (N_6443,N_4021,N_3615);
nor U6444 (N_6444,N_1400,N_1610);
xnor U6445 (N_6445,N_3386,N_3394);
and U6446 (N_6446,N_934,N_4320);
and U6447 (N_6447,N_1842,N_2840);
or U6448 (N_6448,N_3970,N_947);
nand U6449 (N_6449,N_4650,N_4768);
nand U6450 (N_6450,N_2383,N_3163);
nand U6451 (N_6451,N_2647,N_2651);
or U6452 (N_6452,N_434,N_2197);
nor U6453 (N_6453,N_4414,N_2841);
xnor U6454 (N_6454,N_2518,N_454);
or U6455 (N_6455,N_3789,N_4640);
and U6456 (N_6456,N_1495,N_402);
nor U6457 (N_6457,N_832,N_1480);
nor U6458 (N_6458,N_4573,N_3557);
nand U6459 (N_6459,N_2619,N_3925);
xor U6460 (N_6460,N_3067,N_4283);
nor U6461 (N_6461,N_2770,N_1941);
or U6462 (N_6462,N_1279,N_4963);
nand U6463 (N_6463,N_2320,N_657);
or U6464 (N_6464,N_708,N_3902);
and U6465 (N_6465,N_2978,N_115);
or U6466 (N_6466,N_2614,N_4286);
nor U6467 (N_6467,N_3863,N_721);
or U6468 (N_6468,N_4721,N_2919);
xnor U6469 (N_6469,N_1788,N_4956);
and U6470 (N_6470,N_1498,N_3213);
or U6471 (N_6471,N_108,N_636);
nand U6472 (N_6472,N_4976,N_4868);
nor U6473 (N_6473,N_57,N_3971);
nand U6474 (N_6474,N_909,N_2456);
or U6475 (N_6475,N_1377,N_1444);
nor U6476 (N_6476,N_4393,N_428);
or U6477 (N_6477,N_4319,N_3504);
nor U6478 (N_6478,N_1367,N_4148);
or U6479 (N_6479,N_2124,N_1630);
and U6480 (N_6480,N_479,N_4734);
nor U6481 (N_6481,N_2680,N_1104);
nand U6482 (N_6482,N_1233,N_1155);
and U6483 (N_6483,N_3989,N_1749);
nor U6484 (N_6484,N_4529,N_872);
or U6485 (N_6485,N_587,N_3133);
nor U6486 (N_6486,N_1299,N_2252);
nand U6487 (N_6487,N_4661,N_4045);
and U6488 (N_6488,N_663,N_317);
or U6489 (N_6489,N_3652,N_1376);
nand U6490 (N_6490,N_1,N_4533);
nand U6491 (N_6491,N_4547,N_2231);
nor U6492 (N_6492,N_3418,N_2086);
nand U6493 (N_6493,N_3432,N_920);
and U6494 (N_6494,N_1076,N_3933);
or U6495 (N_6495,N_4824,N_3085);
nor U6496 (N_6496,N_4268,N_638);
nor U6497 (N_6497,N_4558,N_1435);
nand U6498 (N_6498,N_2310,N_1695);
nor U6499 (N_6499,N_3173,N_4427);
or U6500 (N_6500,N_817,N_229);
or U6501 (N_6501,N_171,N_4143);
nor U6502 (N_6502,N_278,N_591);
nor U6503 (N_6503,N_1830,N_3317);
or U6504 (N_6504,N_457,N_1289);
xor U6505 (N_6505,N_3229,N_3034);
or U6506 (N_6506,N_3939,N_3168);
or U6507 (N_6507,N_674,N_1034);
and U6508 (N_6508,N_3694,N_1791);
and U6509 (N_6509,N_313,N_4047);
and U6510 (N_6510,N_2506,N_3881);
nor U6511 (N_6511,N_1252,N_2482);
xnor U6512 (N_6512,N_3468,N_2900);
nor U6513 (N_6513,N_4220,N_3336);
nor U6514 (N_6514,N_3376,N_4180);
nand U6515 (N_6515,N_2282,N_4216);
nor U6516 (N_6516,N_734,N_2917);
or U6517 (N_6517,N_4489,N_4206);
or U6518 (N_6518,N_3577,N_3513);
or U6519 (N_6519,N_2042,N_3464);
xnor U6520 (N_6520,N_2381,N_4000);
nor U6521 (N_6521,N_2260,N_4973);
and U6522 (N_6522,N_1161,N_3729);
or U6523 (N_6523,N_3214,N_1306);
nor U6524 (N_6524,N_286,N_3709);
nor U6525 (N_6525,N_4053,N_187);
nand U6526 (N_6526,N_4792,N_3932);
and U6527 (N_6527,N_2268,N_249);
nand U6528 (N_6528,N_753,N_4188);
and U6529 (N_6529,N_3060,N_2289);
or U6530 (N_6530,N_2743,N_1615);
xor U6531 (N_6531,N_170,N_554);
nor U6532 (N_6532,N_3195,N_2565);
nand U6533 (N_6533,N_2346,N_1897);
nand U6534 (N_6534,N_4757,N_4231);
and U6535 (N_6535,N_2009,N_4269);
nor U6536 (N_6536,N_4340,N_1125);
and U6537 (N_6537,N_2362,N_1212);
nor U6538 (N_6538,N_612,N_141);
nor U6539 (N_6539,N_4433,N_3371);
and U6540 (N_6540,N_935,N_3310);
nor U6541 (N_6541,N_10,N_1499);
xor U6542 (N_6542,N_136,N_4814);
nor U6543 (N_6543,N_4472,N_151);
or U6544 (N_6544,N_1961,N_384);
xnor U6545 (N_6545,N_985,N_3717);
and U6546 (N_6546,N_582,N_1618);
nor U6547 (N_6547,N_821,N_2205);
and U6548 (N_6548,N_4568,N_4615);
and U6549 (N_6549,N_644,N_1677);
or U6550 (N_6550,N_1083,N_4694);
nor U6551 (N_6551,N_4449,N_759);
nor U6552 (N_6552,N_4944,N_2216);
nand U6553 (N_6553,N_2809,N_765);
nand U6554 (N_6554,N_2521,N_294);
and U6555 (N_6555,N_534,N_1684);
nand U6556 (N_6556,N_232,N_2588);
or U6557 (N_6557,N_2963,N_1641);
and U6558 (N_6558,N_3828,N_3661);
nor U6559 (N_6559,N_1665,N_4075);
and U6560 (N_6560,N_2111,N_3733);
nor U6561 (N_6561,N_653,N_157);
and U6562 (N_6562,N_2739,N_890);
and U6563 (N_6563,N_1275,N_2071);
and U6564 (N_6564,N_1031,N_3606);
nor U6565 (N_6565,N_2659,N_3498);
and U6566 (N_6566,N_525,N_3078);
or U6567 (N_6567,N_607,N_4836);
nand U6568 (N_6568,N_2974,N_3483);
and U6569 (N_6569,N_2397,N_3277);
and U6570 (N_6570,N_2703,N_2968);
and U6571 (N_6571,N_3027,N_953);
and U6572 (N_6572,N_4942,N_986);
nand U6573 (N_6573,N_1650,N_4804);
xor U6574 (N_6574,N_3369,N_2838);
and U6575 (N_6575,N_2326,N_2217);
nand U6576 (N_6576,N_4707,N_3927);
nand U6577 (N_6577,N_357,N_3562);
xor U6578 (N_6578,N_1688,N_1230);
and U6579 (N_6579,N_1993,N_4142);
and U6580 (N_6580,N_3666,N_3934);
nor U6581 (N_6581,N_4876,N_3307);
nand U6582 (N_6582,N_1182,N_2449);
or U6583 (N_6583,N_3678,N_42);
xor U6584 (N_6584,N_3883,N_2973);
and U6585 (N_6585,N_2074,N_1514);
nand U6586 (N_6586,N_3245,N_3160);
or U6587 (N_6587,N_3722,N_2388);
nand U6588 (N_6588,N_271,N_1398);
or U6589 (N_6589,N_3322,N_4649);
and U6590 (N_6590,N_3853,N_2940);
xnor U6591 (N_6591,N_1373,N_4941);
or U6592 (N_6592,N_1005,N_988);
nor U6593 (N_6593,N_4810,N_3887);
nor U6594 (N_6594,N_362,N_1685);
nor U6595 (N_6595,N_3267,N_4822);
nand U6596 (N_6596,N_4670,N_823);
and U6597 (N_6597,N_367,N_123);
or U6598 (N_6598,N_3543,N_2752);
or U6599 (N_6599,N_2423,N_2241);
xor U6600 (N_6600,N_308,N_4448);
nor U6601 (N_6601,N_231,N_2373);
nand U6602 (N_6602,N_774,N_2728);
or U6603 (N_6603,N_4144,N_2986);
nor U6604 (N_6604,N_4743,N_1274);
and U6605 (N_6605,N_2186,N_315);
and U6606 (N_6606,N_2953,N_1152);
nand U6607 (N_6607,N_2374,N_3913);
nor U6608 (N_6608,N_2927,N_3079);
or U6609 (N_6609,N_224,N_2206);
or U6610 (N_6610,N_2765,N_2416);
nand U6611 (N_6611,N_2876,N_2131);
and U6612 (N_6612,N_218,N_2419);
xor U6613 (N_6613,N_4264,N_2491);
nor U6614 (N_6614,N_2987,N_1127);
nand U6615 (N_6615,N_4402,N_3941);
or U6616 (N_6616,N_4636,N_1172);
nand U6617 (N_6617,N_4932,N_322);
nor U6618 (N_6618,N_1784,N_4289);
or U6619 (N_6619,N_1396,N_3991);
nand U6620 (N_6620,N_340,N_4124);
and U6621 (N_6621,N_3563,N_3005);
and U6622 (N_6622,N_1718,N_1347);
nand U6623 (N_6623,N_54,N_69);
and U6624 (N_6624,N_3767,N_1121);
and U6625 (N_6625,N_1479,N_204);
nor U6626 (N_6626,N_3381,N_2634);
xnor U6627 (N_6627,N_3702,N_248);
or U6628 (N_6628,N_3494,N_4457);
and U6629 (N_6629,N_4097,N_2110);
nor U6630 (N_6630,N_2650,N_978);
nand U6631 (N_6631,N_3516,N_4554);
nor U6632 (N_6632,N_1154,N_3452);
or U6633 (N_6633,N_233,N_3405);
nand U6634 (N_6634,N_3030,N_4574);
nand U6635 (N_6635,N_2327,N_4949);
nor U6636 (N_6636,N_65,N_1210);
or U6637 (N_6637,N_4718,N_3640);
nand U6638 (N_6638,N_3592,N_228);
or U6639 (N_6639,N_1689,N_3613);
xor U6640 (N_6640,N_3151,N_1326);
and U6641 (N_6641,N_1169,N_1706);
or U6642 (N_6642,N_783,N_4555);
or U6643 (N_6643,N_3217,N_3603);
nand U6644 (N_6644,N_2249,N_4653);
nor U6645 (N_6645,N_4857,N_2958);
or U6646 (N_6646,N_2322,N_3428);
nand U6647 (N_6647,N_2579,N_3635);
or U6648 (N_6648,N_439,N_1660);
nor U6649 (N_6649,N_46,N_404);
xnor U6650 (N_6650,N_625,N_802);
and U6651 (N_6651,N_3166,N_2500);
nand U6652 (N_6652,N_2189,N_3940);
nor U6653 (N_6653,N_4055,N_3509);
and U6654 (N_6654,N_798,N_1267);
and U6655 (N_6655,N_2596,N_2621);
nor U6656 (N_6656,N_3786,N_1167);
or U6657 (N_6657,N_3998,N_930);
nand U6658 (N_6658,N_217,N_2179);
and U6659 (N_6659,N_4019,N_4597);
or U6660 (N_6660,N_549,N_2332);
nor U6661 (N_6661,N_3772,N_4952);
nor U6662 (N_6662,N_4683,N_951);
or U6663 (N_6663,N_2544,N_1242);
and U6664 (N_6664,N_4358,N_572);
or U6665 (N_6665,N_958,N_4461);
nor U6666 (N_6666,N_1165,N_4502);
xor U6667 (N_6667,N_3854,N_1972);
nor U6668 (N_6668,N_1924,N_533);
nand U6669 (N_6669,N_4864,N_1994);
nor U6670 (N_6670,N_4534,N_2142);
and U6671 (N_6671,N_4478,N_4270);
or U6672 (N_6672,N_3478,N_4101);
or U6673 (N_6673,N_1106,N_411);
xor U6674 (N_6674,N_4465,N_4185);
xor U6675 (N_6675,N_3835,N_2073);
nand U6676 (N_6676,N_2166,N_213);
nor U6677 (N_6677,N_330,N_960);
xnor U6678 (N_6678,N_4788,N_4186);
or U6679 (N_6679,N_3100,N_4518);
nor U6680 (N_6680,N_4787,N_396);
nand U6681 (N_6681,N_3727,N_1880);
or U6682 (N_6682,N_660,N_1815);
nor U6683 (N_6683,N_2775,N_2024);
nand U6684 (N_6684,N_671,N_2951);
nor U6685 (N_6685,N_1142,N_683);
nor U6686 (N_6686,N_4363,N_771);
nor U6687 (N_6687,N_3104,N_355);
nor U6688 (N_6688,N_3826,N_2960);
nand U6689 (N_6689,N_4419,N_2109);
or U6690 (N_6690,N_3357,N_2554);
and U6691 (N_6691,N_1174,N_1658);
nand U6692 (N_6692,N_2966,N_2222);
nor U6693 (N_6693,N_3759,N_3152);
nor U6694 (N_6694,N_4627,N_2536);
and U6695 (N_6695,N_432,N_34);
xor U6696 (N_6696,N_2476,N_2902);
nand U6697 (N_6697,N_2399,N_220);
or U6698 (N_6698,N_2158,N_2660);
nor U6699 (N_6699,N_944,N_925);
nor U6700 (N_6700,N_1608,N_2566);
nor U6701 (N_6701,N_3695,N_703);
xnor U6702 (N_6702,N_1046,N_1295);
and U6703 (N_6703,N_4744,N_1302);
or U6704 (N_6704,N_2464,N_4771);
or U6705 (N_6705,N_421,N_658);
and U6706 (N_6706,N_3284,N_4809);
nor U6707 (N_6707,N_1215,N_28);
and U6708 (N_6708,N_4830,N_4799);
or U6709 (N_6709,N_866,N_2956);
nand U6710 (N_6710,N_2934,N_4058);
nand U6711 (N_6711,N_4509,N_2555);
or U6712 (N_6712,N_3844,N_2657);
and U6713 (N_6713,N_2585,N_2269);
xor U6714 (N_6714,N_4936,N_4991);
or U6715 (N_6715,N_321,N_1123);
nor U6716 (N_6716,N_3827,N_3329);
or U6717 (N_6717,N_2587,N_2156);
or U6718 (N_6718,N_3436,N_655);
or U6719 (N_6719,N_293,N_4939);
nor U6720 (N_6720,N_2325,N_995);
and U6721 (N_6721,N_2063,N_2586);
or U6722 (N_6722,N_3264,N_604);
nand U6723 (N_6723,N_1281,N_4899);
nor U6724 (N_6724,N_1339,N_3731);
nand U6725 (N_6725,N_4198,N_2348);
nor U6726 (N_6726,N_1812,N_3699);
or U6727 (N_6727,N_1054,N_2406);
nor U6728 (N_6728,N_4062,N_3106);
nor U6729 (N_6729,N_1910,N_2440);
and U6730 (N_6730,N_3774,N_2431);
and U6731 (N_6731,N_2418,N_1500);
or U6732 (N_6732,N_2525,N_3713);
xnor U6733 (N_6733,N_1659,N_3482);
nand U6734 (N_6734,N_4311,N_4793);
nor U6735 (N_6735,N_3013,N_789);
nand U6736 (N_6736,N_406,N_31);
or U6737 (N_6737,N_4093,N_273);
or U6738 (N_6738,N_3207,N_3833);
xor U6739 (N_6739,N_494,N_331);
or U6740 (N_6740,N_4628,N_3446);
nand U6741 (N_6741,N_4921,N_2994);
xor U6742 (N_6742,N_3361,N_2316);
and U6743 (N_6743,N_2033,N_349);
nor U6744 (N_6744,N_1545,N_3144);
nor U6745 (N_6745,N_973,N_1113);
and U6746 (N_6746,N_2203,N_791);
and U6747 (N_6747,N_1474,N_1470);
nand U6748 (N_6748,N_1519,N_138);
nand U6749 (N_6749,N_831,N_353);
nor U6750 (N_6750,N_4229,N_2062);
and U6751 (N_6751,N_1890,N_2962);
nand U6752 (N_6752,N_4351,N_1426);
nor U6753 (N_6753,N_14,N_673);
or U6754 (N_6754,N_1638,N_4733);
and U6755 (N_6755,N_2810,N_4086);
or U6756 (N_6756,N_2192,N_4656);
and U6757 (N_6757,N_1415,N_883);
and U6758 (N_6758,N_4698,N_965);
nand U6759 (N_6759,N_3788,N_632);
nor U6760 (N_6760,N_1443,N_3899);
or U6761 (N_6761,N_2031,N_3545);
or U6762 (N_6762,N_3046,N_1218);
nor U6763 (N_6763,N_222,N_4104);
and U6764 (N_6764,N_1269,N_2461);
nor U6765 (N_6765,N_1251,N_3955);
nand U6766 (N_6766,N_1445,N_865);
and U6767 (N_6767,N_2941,N_553);
nor U6768 (N_6768,N_3273,N_4051);
nand U6769 (N_6769,N_1716,N_1147);
xor U6770 (N_6770,N_2196,N_4724);
and U6771 (N_6771,N_4972,N_1869);
and U6772 (N_6772,N_3026,N_2745);
nor U6773 (N_6773,N_1195,N_542);
nand U6774 (N_6774,N_570,N_3846);
nand U6775 (N_6775,N_3506,N_2022);
xor U6776 (N_6776,N_4727,N_1546);
nor U6777 (N_6777,N_1038,N_1438);
nand U6778 (N_6778,N_470,N_3623);
or U6779 (N_6779,N_1704,N_3782);
nand U6780 (N_6780,N_2224,N_35);
and U6781 (N_6781,N_2702,N_251);
nand U6782 (N_6782,N_3402,N_3132);
and U6783 (N_6783,N_3403,N_4893);
and U6784 (N_6784,N_4317,N_4181);
nor U6785 (N_6785,N_855,N_290);
or U6786 (N_6786,N_4479,N_1602);
nand U6787 (N_6787,N_477,N_3440);
nor U6788 (N_6788,N_4539,N_3135);
nand U6789 (N_6789,N_4463,N_528);
nor U6790 (N_6790,N_2396,N_4255);
nand U6791 (N_6791,N_2607,N_566);
and U6792 (N_6792,N_4583,N_3429);
or U6793 (N_6793,N_2281,N_659);
nor U6794 (N_6794,N_4447,N_4651);
nand U6795 (N_6795,N_4277,N_4064);
nor U6796 (N_6796,N_4166,N_3204);
and U6797 (N_6797,N_2520,N_1661);
xnor U6798 (N_6798,N_3920,N_4332);
nand U6799 (N_6799,N_2867,N_1835);
nand U6800 (N_6800,N_3425,N_2806);
and U6801 (N_6801,N_3314,N_1819);
xor U6802 (N_6802,N_4684,N_2466);
or U6803 (N_6803,N_2184,N_687);
nand U6804 (N_6804,N_4297,N_2313);
and U6805 (N_6805,N_1217,N_2127);
nand U6806 (N_6806,N_3156,N_1888);
and U6807 (N_6807,N_465,N_788);
nor U6808 (N_6808,N_601,N_2613);
nor U6809 (N_6809,N_1713,N_298);
nor U6810 (N_6810,N_1007,N_64);
nor U6811 (N_6811,N_2870,N_2007);
or U6812 (N_6812,N_1898,N_481);
nor U6813 (N_6813,N_2060,N_3093);
and U6814 (N_6814,N_4190,N_1889);
and U6815 (N_6815,N_2092,N_3);
nor U6816 (N_6816,N_993,N_578);
and U6817 (N_6817,N_4634,N_3380);
or U6818 (N_6818,N_2228,N_2658);
and U6819 (N_6819,N_3202,N_826);
xor U6820 (N_6820,N_445,N_2557);
nand U6821 (N_6821,N_3077,N_4258);
nand U6822 (N_6822,N_2772,N_2751);
nor U6823 (N_6823,N_4482,N_1895);
nor U6824 (N_6824,N_1970,N_3785);
nand U6825 (N_6825,N_3086,N_2721);
or U6826 (N_6826,N_2136,N_1379);
nand U6827 (N_6827,N_1952,N_3616);
and U6828 (N_6828,N_4681,N_2134);
nand U6829 (N_6829,N_4816,N_132);
nand U6830 (N_6830,N_2679,N_3321);
and U6831 (N_6831,N_4459,N_1937);
and U6832 (N_6832,N_413,N_4685);
nand U6833 (N_6833,N_4900,N_1989);
nor U6834 (N_6834,N_4117,N_2817);
or U6835 (N_6835,N_1780,N_2479);
and U6836 (N_6836,N_2538,N_2510);
and U6837 (N_6837,N_3999,N_3708);
and U6838 (N_6838,N_2267,N_272);
and U6839 (N_6839,N_969,N_4937);
xor U6840 (N_6840,N_1323,N_691);
or U6841 (N_6841,N_1980,N_2639);
xor U6842 (N_6842,N_4785,N_778);
and U6843 (N_6843,N_3139,N_814);
nor U6844 (N_6844,N_4089,N_476);
nand U6845 (N_6845,N_2597,N_266);
or U6846 (N_6846,N_254,N_4416);
or U6847 (N_6847,N_2558,N_3948);
and U6848 (N_6848,N_2595,N_1893);
and U6849 (N_6849,N_1616,N_3747);
or U6850 (N_6850,N_1316,N_693);
nor U6851 (N_6851,N_4361,N_3981);
or U6852 (N_6852,N_4990,N_2061);
nand U6853 (N_6853,N_256,N_4467);
xnor U6854 (N_6854,N_1380,N_1386);
nor U6855 (N_6855,N_1258,N_17);
or U6856 (N_6856,N_2159,N_1948);
and U6857 (N_6857,N_1004,N_3028);
nand U6858 (N_6858,N_2654,N_2367);
or U6859 (N_6859,N_1211,N_2128);
nor U6860 (N_6860,N_2599,N_1101);
or U6861 (N_6861,N_4673,N_3332);
and U6862 (N_6862,N_1418,N_2425);
nand U6863 (N_6863,N_1769,N_3598);
and U6864 (N_6864,N_2747,N_3845);
or U6865 (N_6865,N_410,N_4947);
or U6866 (N_6866,N_354,N_776);
nor U6867 (N_6867,N_444,N_2170);
nand U6868 (N_6868,N_209,N_2914);
nor U6869 (N_6869,N_1199,N_2767);
xnor U6870 (N_6870,N_226,N_305);
or U6871 (N_6871,N_466,N_1678);
and U6872 (N_6872,N_3566,N_3900);
and U6873 (N_6873,N_3210,N_1030);
nor U6874 (N_6874,N_316,N_4871);
nand U6875 (N_6875,N_3294,N_4548);
xor U6876 (N_6876,N_3189,N_2211);
or U6877 (N_6877,N_1967,N_4129);
or U6878 (N_6878,N_718,N_51);
and U6879 (N_6879,N_2286,N_2899);
or U6880 (N_6880,N_2652,N_645);
nor U6881 (N_6881,N_1719,N_3108);
and U6882 (N_6882,N_3584,N_1335);
nand U6883 (N_6883,N_3158,N_181);
or U6884 (N_6884,N_1969,N_2043);
xor U6885 (N_6885,N_1318,N_3882);
or U6886 (N_6886,N_1774,N_1272);
or U6887 (N_6887,N_4458,N_1733);
nand U6888 (N_6888,N_996,N_1064);
or U6889 (N_6889,N_1024,N_76);
xnor U6890 (N_6890,N_3382,N_3942);
or U6891 (N_6891,N_1951,N_1409);
and U6892 (N_6892,N_2075,N_3411);
nor U6893 (N_6893,N_381,N_2886);
or U6894 (N_6894,N_1149,N_3448);
or U6895 (N_6895,N_928,N_59);
and U6896 (N_6896,N_4149,N_4763);
nor U6897 (N_6897,N_4512,N_486);
nor U6898 (N_6898,N_4552,N_4832);
xnor U6899 (N_6899,N_3112,N_2471);
xor U6900 (N_6900,N_4244,N_1779);
and U6901 (N_6901,N_4338,N_692);
nand U6902 (N_6902,N_1221,N_1473);
xor U6903 (N_6903,N_589,N_4859);
and U6904 (N_6904,N_177,N_2704);
and U6905 (N_6905,N_2093,N_4193);
and U6906 (N_6906,N_2681,N_399);
nor U6907 (N_6907,N_4381,N_1547);
nand U6908 (N_6908,N_4999,N_1764);
and U6909 (N_6909,N_4083,N_580);
or U6910 (N_6910,N_1136,N_2164);
xnor U6911 (N_6911,N_4020,N_389);
and U6912 (N_6912,N_4617,N_3484);
or U6913 (N_6913,N_4964,N_4145);
nand U6914 (N_6914,N_4517,N_3575);
and U6915 (N_6915,N_2001,N_3781);
and U6916 (N_6916,N_4141,N_1933);
and U6917 (N_6917,N_564,N_3337);
nor U6918 (N_6918,N_3859,N_3994);
or U6919 (N_6919,N_4845,N_1935);
or U6920 (N_6920,N_264,N_400);
and U6921 (N_6921,N_2537,N_1950);
and U6922 (N_6922,N_724,N_4982);
and U6923 (N_6923,N_2212,N_2047);
or U6924 (N_6924,N_3803,N_837);
or U6925 (N_6925,N_227,N_2575);
nor U6926 (N_6926,N_2006,N_2106);
xnor U6927 (N_6927,N_20,N_4002);
nor U6928 (N_6928,N_509,N_1112);
nor U6929 (N_6929,N_4620,N_3228);
nand U6930 (N_6930,N_4336,N_4230);
nand U6931 (N_6931,N_140,N_2450);
nand U6932 (N_6932,N_1593,N_3219);
xor U6933 (N_6933,N_1096,N_2275);
or U6934 (N_6934,N_2551,N_3006);
xor U6935 (N_6935,N_1108,N_1601);
or U6936 (N_6936,N_1971,N_4079);
xnor U6937 (N_6937,N_1270,N_1351);
nand U6938 (N_6938,N_4561,N_1334);
nand U6939 (N_6939,N_3894,N_3795);
xor U6940 (N_6940,N_1562,N_4527);
xor U6941 (N_6941,N_2990,N_4094);
and U6942 (N_6942,N_2463,N_346);
nand U6943 (N_6943,N_4553,N_4888);
or U6944 (N_6944,N_215,N_2084);
or U6945 (N_6945,N_1826,N_3689);
or U6946 (N_6946,N_1878,N_1577);
nand U6947 (N_6947,N_3551,N_356);
and U6948 (N_6948,N_4033,N_301);
or U6949 (N_6949,N_3912,N_1067);
or U6950 (N_6950,N_2871,N_2713);
or U6951 (N_6951,N_302,N_3539);
nand U6952 (N_6952,N_4341,N_3631);
nor U6953 (N_6953,N_2070,N_2015);
or U6954 (N_6954,N_1973,N_3487);
nor U6955 (N_6955,N_1754,N_3051);
nand U6956 (N_6956,N_4962,N_4368);
or U6957 (N_6957,N_861,N_2214);
or U6958 (N_6958,N_382,N_1392);
nor U6959 (N_6959,N_2052,N_3840);
xnor U6960 (N_6960,N_4676,N_3960);
xnor U6961 (N_6961,N_606,N_2683);
nand U6962 (N_6962,N_3807,N_173);
and U6963 (N_6963,N_4848,N_4853);
xor U6964 (N_6964,N_2235,N_296);
nand U6965 (N_6965,N_3199,N_4687);
xnor U6966 (N_6966,N_1072,N_3235);
and U6967 (N_6967,N_3224,N_4837);
or U6968 (N_6968,N_2505,N_3901);
xnor U6969 (N_6969,N_983,N_4469);
or U6970 (N_6970,N_2139,N_1810);
and U6971 (N_6971,N_501,N_1388);
nor U6972 (N_6972,N_212,N_1915);
nand U6973 (N_6973,N_3438,N_2209);
and U6974 (N_6974,N_3447,N_1570);
nand U6975 (N_6975,N_3362,N_4350);
or U6976 (N_6976,N_1288,N_669);
or U6977 (N_6977,N_998,N_2038);
and U6978 (N_6978,N_1672,N_4404);
and U6979 (N_6979,N_3865,N_3003);
nand U6980 (N_6980,N_736,N_1488);
or U6981 (N_6981,N_3944,N_556);
nand U6982 (N_6982,N_3265,N_1789);
and U6983 (N_6983,N_679,N_2018);
nand U6984 (N_6984,N_1359,N_4500);
nand U6985 (N_6985,N_829,N_1699);
xor U6986 (N_6986,N_2949,N_1484);
xnor U6987 (N_6987,N_1912,N_3866);
and U6988 (N_6988,N_4224,N_1105);
nand U6989 (N_6989,N_4301,N_80);
nand U6990 (N_6990,N_3735,N_4114);
nor U6991 (N_6991,N_4957,N_419);
and U6992 (N_6992,N_4039,N_2856);
nor U6993 (N_6993,N_1278,N_4052);
xor U6994 (N_6994,N_2582,N_3171);
nand U6995 (N_6995,N_2509,N_2612);
nor U6996 (N_6996,N_1620,N_4462);
and U6997 (N_6997,N_2107,N_3891);
or U6998 (N_6998,N_1629,N_3801);
nand U6999 (N_6999,N_394,N_55);
nor U7000 (N_7000,N_2137,N_4127);
nand U7001 (N_7001,N_2140,N_260);
and U7002 (N_7002,N_4680,N_4715);
and U7003 (N_7003,N_1491,N_2965);
nor U7004 (N_7004,N_4671,N_4829);
and U7005 (N_7005,N_139,N_474);
and U7006 (N_7006,N_4790,N_2880);
nor U7007 (N_7007,N_3335,N_1497);
xnor U7008 (N_7008,N_2352,N_4577);
or U7009 (N_7009,N_1590,N_1477);
and U7010 (N_7010,N_2620,N_1342);
or U7011 (N_7011,N_3281,N_3401);
nor U7012 (N_7012,N_1874,N_4702);
or U7013 (N_7013,N_864,N_3893);
xnor U7014 (N_7014,N_3205,N_1884);
nor U7015 (N_7015,N_4329,N_775);
nand U7016 (N_7016,N_1625,N_2860);
or U7017 (N_7017,N_1875,N_5);
nor U7018 (N_7018,N_4777,N_3728);
nor U7019 (N_7019,N_3537,N_4140);
xor U7020 (N_7020,N_2526,N_56);
and U7021 (N_7021,N_2323,N_2489);
or U7022 (N_7022,N_484,N_1926);
and U7023 (N_7023,N_2354,N_4613);
or U7024 (N_7024,N_4451,N_1126);
and U7025 (N_7025,N_4911,N_2122);
xor U7026 (N_7026,N_1648,N_3719);
nand U7027 (N_7027,N_4912,N_3958);
xnor U7028 (N_7028,N_2785,N_3057);
or U7029 (N_7029,N_1364,N_58);
nor U7030 (N_7030,N_327,N_460);
nor U7031 (N_7031,N_1048,N_3986);
nand U7032 (N_7032,N_2408,N_3794);
and U7033 (N_7033,N_4815,N_1916);
nor U7034 (N_7034,N_409,N_4919);
and U7035 (N_7035,N_614,N_162);
and U7036 (N_7036,N_1494,N_1313);
nand U7037 (N_7037,N_4455,N_145);
or U7038 (N_7038,N_3461,N_1345);
and U7039 (N_7039,N_235,N_3188);
nand U7040 (N_7040,N_910,N_3911);
or U7041 (N_7041,N_203,N_4985);
nand U7042 (N_7042,N_598,N_3456);
and U7043 (N_7043,N_2102,N_1171);
nand U7044 (N_7044,N_2089,N_3326);
nand U7045 (N_7045,N_4541,N_3636);
or U7046 (N_7046,N_3842,N_4146);
nand U7047 (N_7047,N_4309,N_3134);
nor U7048 (N_7048,N_2947,N_3233);
nor U7049 (N_7049,N_3760,N_2262);
or U7050 (N_7050,N_3227,N_2773);
and U7051 (N_7051,N_1734,N_2989);
or U7052 (N_7052,N_4040,N_4440);
nand U7053 (N_7053,N_2305,N_2455);
nor U7054 (N_7054,N_2873,N_4207);
and U7055 (N_7055,N_3009,N_3783);
xnor U7056 (N_7056,N_2952,N_2039);
nor U7057 (N_7057,N_4085,N_2);
nand U7058 (N_7058,N_904,N_1100);
nand U7059 (N_7059,N_3324,N_797);
and U7060 (N_7060,N_959,N_1300);
or U7061 (N_7061,N_1427,N_1341);
nor U7062 (N_7062,N_4118,N_2866);
and U7063 (N_7063,N_3966,N_921);
xor U7064 (N_7064,N_1314,N_504);
nor U7065 (N_7065,N_4946,N_1995);
nor U7066 (N_7066,N_2637,N_3167);
and U7067 (N_7067,N_3720,N_2190);
xor U7068 (N_7068,N_2337,N_1020);
xor U7069 (N_7069,N_1489,N_2133);
xor U7070 (N_7070,N_2574,N_698);
nor U7071 (N_7071,N_4493,N_3262);
nand U7072 (N_7072,N_2999,N_259);
or U7073 (N_7073,N_3821,N_1986);
nand U7074 (N_7074,N_4201,N_94);
or U7075 (N_7075,N_1727,N_4955);
and U7076 (N_7076,N_1079,N_1250);
and U7077 (N_7077,N_1606,N_1589);
and U7078 (N_7078,N_1536,N_144);
and U7079 (N_7079,N_4996,N_3851);
nand U7080 (N_7080,N_3192,N_2771);
and U7081 (N_7081,N_3973,N_1892);
and U7082 (N_7082,N_4545,N_4099);
nor U7083 (N_7083,N_2983,N_4004);
nor U7084 (N_7084,N_2908,N_4168);
and U7085 (N_7085,N_1117,N_845);
xnor U7086 (N_7086,N_2412,N_4872);
nor U7087 (N_7087,N_887,N_748);
and U7088 (N_7088,N_405,N_2540);
and U7089 (N_7089,N_223,N_684);
nand U7090 (N_7090,N_4076,N_4397);
or U7091 (N_7091,N_2622,N_388);
nor U7092 (N_7092,N_929,N_3693);
nand U7093 (N_7093,N_970,N_1128);
or U7094 (N_7094,N_3320,N_1728);
nor U7095 (N_7095,N_3968,N_755);
nand U7096 (N_7096,N_523,N_792);
or U7097 (N_7097,N_2869,N_3481);
xor U7098 (N_7098,N_3041,N_2312);
nand U7099 (N_7099,N_2404,N_500);
xnor U7100 (N_7100,N_1087,N_3924);
xor U7101 (N_7101,N_4006,N_4978);
and U7102 (N_7102,N_1611,N_2379);
nor U7103 (N_7103,N_2331,N_4765);
nor U7104 (N_7104,N_1767,N_4566);
nor U7105 (N_7105,N_1308,N_4821);
or U7106 (N_7106,N_4564,N_4693);
or U7107 (N_7107,N_3323,N_3295);
nand U7108 (N_7108,N_761,N_306);
xor U7109 (N_7109,N_90,N_2868);
or U7110 (N_7110,N_4515,N_2664);
nor U7111 (N_7111,N_373,N_907);
nand U7112 (N_7112,N_3624,N_4399);
nor U7113 (N_7113,N_975,N_3384);
and U7114 (N_7114,N_2758,N_4405);
nor U7115 (N_7115,N_2432,N_931);
nand U7116 (N_7116,N_2748,N_1016);
or U7117 (N_7117,N_2842,N_836);
and U7118 (N_7118,N_4958,N_2761);
nand U7119 (N_7119,N_3542,N_635);
or U7120 (N_7120,N_1722,N_107);
xor U7121 (N_7121,N_48,N_3950);
xnor U7122 (N_7122,N_2792,N_1867);
nand U7123 (N_7123,N_966,N_1674);
xnor U7124 (N_7124,N_3686,N_3922);
nand U7125 (N_7125,N_2921,N_4044);
nor U7126 (N_7126,N_2161,N_1206);
and U7127 (N_7127,N_3398,N_1357);
nor U7128 (N_7128,N_3936,N_1829);
and U7129 (N_7129,N_3074,N_2910);
nand U7130 (N_7130,N_1184,N_4904);
nand U7131 (N_7131,N_1331,N_3347);
nand U7132 (N_7132,N_588,N_1387);
xnor U7133 (N_7133,N_4503,N_3967);
or U7134 (N_7134,N_61,N_371);
or U7135 (N_7135,N_2843,N_3510);
or U7136 (N_7136,N_512,N_702);
or U7137 (N_7137,N_4102,N_1006);
xnor U7138 (N_7138,N_221,N_3105);
and U7139 (N_7139,N_2256,N_4759);
or U7140 (N_7140,N_3017,N_2667);
or U7141 (N_7141,N_2933,N_2731);
or U7142 (N_7142,N_4354,N_1541);
nor U7143 (N_7143,N_2334,N_3488);
nand U7144 (N_7144,N_2714,N_4088);
or U7145 (N_7145,N_2576,N_43);
nand U7146 (N_7146,N_668,N_1702);
nand U7147 (N_7147,N_807,N_3520);
nand U7148 (N_7148,N_766,N_938);
and U7149 (N_7149,N_1873,N_166);
nand U7150 (N_7150,N_2441,N_2829);
nor U7151 (N_7151,N_4764,N_1793);
nor U7152 (N_7152,N_2233,N_2569);
or U7153 (N_7153,N_4537,N_697);
xnor U7154 (N_7154,N_3090,N_3061);
and U7155 (N_7155,N_2717,N_688);
xnor U7156 (N_7156,N_3413,N_2349);
nor U7157 (N_7157,N_2069,N_239);
or U7158 (N_7158,N_1063,N_3426);
and U7159 (N_7159,N_3049,N_3753);
and U7160 (N_7160,N_979,N_2845);
and U7161 (N_7161,N_2490,N_4048);
nand U7162 (N_7162,N_503,N_769);
and U7163 (N_7163,N_706,N_3797);
and U7164 (N_7164,N_1204,N_677);
and U7165 (N_7165,N_1471,N_1120);
and U7166 (N_7166,N_2391,N_763);
and U7167 (N_7167,N_4657,N_4720);
nor U7168 (N_7168,N_3083,N_3346);
nand U7169 (N_7169,N_1137,N_1923);
nor U7170 (N_7170,N_1235,N_1738);
xnor U7171 (N_7171,N_4158,N_1041);
nor U7172 (N_7172,N_314,N_3601);
and U7173 (N_7173,N_4403,N_1557);
nor U7174 (N_7174,N_1794,N_3961);
xor U7175 (N_7175,N_1522,N_3110);
nand U7176 (N_7176,N_2244,N_195);
nand U7177 (N_7177,N_4847,N_199);
nor U7178 (N_7178,N_4450,N_2825);
or U7179 (N_7179,N_3664,N_3075);
nor U7180 (N_7180,N_72,N_567);
nand U7181 (N_7181,N_1847,N_283);
xor U7182 (N_7182,N_2769,N_1255);
and U7183 (N_7183,N_3282,N_4179);
or U7184 (N_7184,N_2169,N_1584);
or U7185 (N_7185,N_1371,N_4488);
and U7186 (N_7186,N_2434,N_2174);
or U7187 (N_7187,N_2366,N_2889);
nand U7188 (N_7188,N_3628,N_3800);
xnor U7189 (N_7189,N_3272,N_4013);
and U7190 (N_7190,N_4109,N_1338);
nor U7191 (N_7191,N_4995,N_3316);
or U7192 (N_7192,N_2628,N_1311);
nor U7193 (N_7193,N_3593,N_3198);
and U7194 (N_7194,N_2118,N_2278);
and U7195 (N_7195,N_3427,N_2246);
or U7196 (N_7196,N_2872,N_4418);
or U7197 (N_7197,N_4983,N_4531);
and U7198 (N_7198,N_2644,N_744);
or U7199 (N_7199,N_117,N_2534);
nor U7200 (N_7200,N_4178,N_4998);
xnor U7201 (N_7201,N_3550,N_2165);
nor U7202 (N_7202,N_3029,N_3149);
nor U7203 (N_7203,N_2300,N_1049);
xor U7204 (N_7204,N_1069,N_202);
nand U7205 (N_7205,N_2095,N_2225);
nand U7206 (N_7206,N_569,N_3725);
nor U7207 (N_7207,N_1792,N_2098);
nand U7208 (N_7208,N_4997,N_3514);
nand U7209 (N_7209,N_4675,N_192);
and U7210 (N_7210,N_2103,N_1773);
and U7211 (N_7211,N_467,N_1055);
or U7212 (N_7212,N_4031,N_4385);
xor U7213 (N_7213,N_368,N_3007);
or U7214 (N_7214,N_2833,N_89);
nor U7215 (N_7215,N_1319,N_3412);
nor U7216 (N_7216,N_2852,N_4774);
nor U7217 (N_7217,N_4980,N_4192);
and U7218 (N_7218,N_2707,N_268);
and U7219 (N_7219,N_963,N_3572);
nand U7220 (N_7220,N_4395,N_1023);
nand U7221 (N_7221,N_1109,N_3502);
nand U7222 (N_7222,N_4989,N_1757);
and U7223 (N_7223,N_438,N_2768);
and U7224 (N_7224,N_1649,N_4580);
or U7225 (N_7225,N_3671,N_3304);
nand U7226 (N_7226,N_1907,N_2691);
xor U7227 (N_7227,N_4849,N_2800);
and U7228 (N_7228,N_2794,N_3665);
xor U7229 (N_7229,N_964,N_1820);
and U7230 (N_7230,N_3001,N_4605);
nand U7231 (N_7231,N_2119,N_3289);
xor U7232 (N_7232,N_2740,N_1687);
and U7233 (N_7233,N_3311,N_918);
nand U7234 (N_7234,N_3319,N_1751);
and U7235 (N_7235,N_3471,N_2682);
nor U7236 (N_7236,N_1800,N_4041);
nor U7237 (N_7237,N_4136,N_3508);
nor U7238 (N_7238,N_4182,N_3416);
or U7239 (N_7239,N_4443,N_4035);
or U7240 (N_7240,N_498,N_4750);
nand U7241 (N_7241,N_557,N_3531);
nand U7242 (N_7242,N_2796,N_1853);
nand U7243 (N_7243,N_3701,N_3714);
and U7244 (N_7244,N_3710,N_1071);
or U7245 (N_7245,N_2944,N_2329);
xor U7246 (N_7246,N_3802,N_3182);
and U7247 (N_7247,N_292,N_3990);
and U7248 (N_7248,N_4499,N_3004);
or U7249 (N_7249,N_999,N_491);
nand U7250 (N_7250,N_1486,N_3619);
or U7251 (N_7251,N_328,N_923);
nor U7252 (N_7252,N_4016,N_4391);
and U7253 (N_7253,N_4525,N_664);
nor U7254 (N_7254,N_2034,N_2430);
nor U7255 (N_7255,N_2993,N_2486);
nand U7256 (N_7256,N_1540,N_3422);
and U7257 (N_7257,N_284,N_2514);
or U7258 (N_7258,N_3568,N_24);
nor U7259 (N_7259,N_130,N_160);
or U7260 (N_7260,N_4594,N_2150);
nor U7261 (N_7261,N_2410,N_3072);
and U7262 (N_7262,N_1846,N_1330);
or U7263 (N_7263,N_2438,N_386);
and U7264 (N_7264,N_3876,N_622);
xor U7265 (N_7265,N_1236,N_3116);
xnor U7266 (N_7266,N_4645,N_1413);
nand U7267 (N_7267,N_4227,N_3610);
or U7268 (N_7268,N_1533,N_1627);
or U7269 (N_7269,N_4367,N_4398);
nor U7270 (N_7270,N_417,N_2757);
and U7271 (N_7271,N_351,N_3746);
and U7272 (N_7272,N_3045,N_3565);
or U7273 (N_7273,N_3716,N_4335);
and U7274 (N_7274,N_3008,N_3145);
or U7275 (N_7275,N_4199,N_378);
or U7276 (N_7276,N_2689,N_723);
or U7277 (N_7277,N_3796,N_2017);
and U7278 (N_7278,N_364,N_4237);
and U7279 (N_7279,N_982,N_4159);
or U7280 (N_7280,N_3637,N_2865);
nor U7281 (N_7281,N_3765,N_3586);
nand U7282 (N_7282,N_2413,N_4122);
or U7283 (N_7283,N_2631,N_3011);
or U7284 (N_7284,N_1363,N_418);
nand U7285 (N_7285,N_1693,N_2532);
or U7286 (N_7286,N_1019,N_2054);
or U7287 (N_7287,N_2950,N_3904);
and U7288 (N_7288,N_793,N_2969);
or U7289 (N_7289,N_2729,N_3561);
and U7290 (N_7290,N_1340,N_2879);
and U7291 (N_7291,N_493,N_1205);
nand U7292 (N_7292,N_18,N_1750);
or U7293 (N_7293,N_1765,N_2819);
nand U7294 (N_7294,N_3848,N_4183);
nor U7295 (N_7295,N_3349,N_1145);
and U7296 (N_7296,N_2130,N_1775);
xor U7297 (N_7297,N_2895,N_3529);
or U7298 (N_7298,N_3771,N_2598);
nand U7299 (N_7299,N_3730,N_981);
nor U7300 (N_7300,N_3076,N_850);
xor U7301 (N_7301,N_4328,N_1957);
and U7302 (N_7302,N_1743,N_1368);
and U7303 (N_7303,N_1824,N_3206);
xnor U7304 (N_7304,N_971,N_3524);
or U7305 (N_7305,N_1530,N_1739);
xor U7306 (N_7306,N_1475,N_2451);
or U7307 (N_7307,N_1490,N_451);
and U7308 (N_7308,N_610,N_3474);
or U7309 (N_7309,N_630,N_1988);
nand U7310 (N_7310,N_403,N_1548);
nor U7311 (N_7311,N_1178,N_1393);
and U7312 (N_7312,N_4261,N_547);
and U7313 (N_7313,N_102,N_4883);
nand U7314 (N_7314,N_1717,N_1927);
nor U7315 (N_7315,N_905,N_4805);
or U7316 (N_7316,N_1265,N_3688);
nand U7317 (N_7317,N_416,N_4758);
and U7318 (N_7318,N_1796,N_740);
or U7319 (N_7319,N_1287,N_4752);
nor U7320 (N_7320,N_3834,N_4025);
nand U7321 (N_7321,N_29,N_3685);
or U7322 (N_7322,N_329,N_4437);
and U7323 (N_7323,N_4719,N_4699);
nand U7324 (N_7324,N_2013,N_4669);
or U7325 (N_7325,N_1324,N_750);
or U7326 (N_7326,N_3241,N_3895);
or U7327 (N_7327,N_4355,N_3824);
and U7328 (N_7328,N_1454,N_253);
nor U7329 (N_7329,N_3511,N_3580);
xnor U7330 (N_7330,N_3293,N_4798);
nor U7331 (N_7331,N_3582,N_2625);
xor U7332 (N_7332,N_3779,N_1093);
nor U7333 (N_7333,N_2344,N_4379);
or U7334 (N_7334,N_4072,N_1089);
and U7335 (N_7335,N_3255,N_2439);
nor U7336 (N_7336,N_3784,N_1679);
nor U7337 (N_7337,N_737,N_3044);
or U7338 (N_7338,N_1173,N_4965);
nor U7339 (N_7339,N_3194,N_3039);
nand U7340 (N_7340,N_1303,N_1248);
nand U7341 (N_7341,N_656,N_2359);
or U7342 (N_7342,N_4887,N_1797);
nor U7343 (N_7343,N_4722,N_2632);
nor U7344 (N_7344,N_1571,N_4090);
nand U7345 (N_7345,N_4249,N_957);
nor U7346 (N_7346,N_2561,N_2088);
or U7347 (N_7347,N_4077,N_3491);
nor U7348 (N_7348,N_2290,N_1596);
nor U7349 (N_7349,N_1675,N_2470);
nand U7350 (N_7350,N_1662,N_3644);
nand U7351 (N_7351,N_4480,N_3419);
and U7352 (N_7352,N_4345,N_1193);
or U7353 (N_7353,N_3748,N_4606);
and U7354 (N_7354,N_1458,N_3442);
xor U7355 (N_7355,N_1180,N_2837);
and U7356 (N_7356,N_3125,N_26);
nor U7357 (N_7357,N_4632,N_2117);
nor U7358 (N_7358,N_717,N_1385);
nor U7359 (N_7359,N_4280,N_3249);
or U7360 (N_7360,N_1831,N_3177);
nor U7361 (N_7361,N_2669,N_95);
nand U7362 (N_7362,N_280,N_1870);
nand U7363 (N_7363,N_4754,N_516);
nor U7364 (N_7364,N_1227,N_2791);
and U7365 (N_7365,N_1578,N_916);
and U7366 (N_7366,N_3538,N_2798);
and U7367 (N_7367,N_3985,N_3668);
or U7368 (N_7368,N_2584,N_4347);
or U7369 (N_7369,N_715,N_1745);
nor U7370 (N_7370,N_4647,N_4614);
and U7371 (N_7371,N_4761,N_1655);
nor U7372 (N_7372,N_1390,N_997);
or U7373 (N_7373,N_3680,N_4126);
and U7374 (N_7374,N_1561,N_4775);
and U7375 (N_7375,N_1551,N_3215);
and U7376 (N_7376,N_1999,N_3549);
nand U7377 (N_7377,N_2333,N_1487);
and U7378 (N_7378,N_3962,N_830);
nand U7379 (N_7379,N_860,N_4302);
and U7380 (N_7380,N_3969,N_2782);
xor U7381 (N_7381,N_3415,N_3275);
nand U7382 (N_7382,N_1692,N_3625);
or U7383 (N_7383,N_2347,N_2777);
or U7384 (N_7384,N_4926,N_3535);
nor U7385 (N_7385,N_374,N_594);
or U7386 (N_7386,N_2002,N_1814);
or U7387 (N_7387,N_452,N_911);
nor U7388 (N_7388,N_2008,N_828);
xor U7389 (N_7389,N_3162,N_1163);
nor U7390 (N_7390,N_510,N_1469);
nand U7391 (N_7391,N_2992,N_2720);
or U7392 (N_7392,N_4067,N_875);
nor U7393 (N_7393,N_945,N_230);
and U7394 (N_7394,N_3288,N_3138);
nand U7395 (N_7395,N_1060,N_4665);
nand U7396 (N_7396,N_1447,N_4977);
or U7397 (N_7397,N_590,N_310);
or U7398 (N_7398,N_207,N_4889);
or U7399 (N_7399,N_2049,N_1949);
and U7400 (N_7400,N_342,N_3062);
nand U7401 (N_7401,N_3404,N_1094);
nor U7402 (N_7402,N_4322,N_1803);
nand U7403 (N_7403,N_3792,N_2458);
nand U7404 (N_7404,N_3519,N_2227);
and U7405 (N_7405,N_1711,N_4979);
nor U7406 (N_7406,N_790,N_2426);
nor U7407 (N_7407,N_2183,N_1707);
nor U7408 (N_7408,N_4098,N_900);
nand U7409 (N_7409,N_2797,N_146);
or U7410 (N_7410,N_3877,N_818);
nand U7411 (N_7411,N_4516,N_3540);
and U7412 (N_7412,N_4223,N_1936);
nand U7413 (N_7413,N_4406,N_4240);
nand U7414 (N_7414,N_4324,N_335);
and U7415 (N_7415,N_1521,N_779);
xor U7416 (N_7416,N_3670,N_4373);
nor U7417 (N_7417,N_3897,N_690);
or U7418 (N_7418,N_3059,N_725);
nor U7419 (N_7419,N_243,N_1309);
and U7420 (N_7420,N_4189,N_412);
nor U7421 (N_7421,N_2213,N_1652);
xnor U7422 (N_7422,N_2675,N_3119);
and U7423 (N_7423,N_2495,N_3259);
xnor U7424 (N_7424,N_3226,N_1772);
nor U7425 (N_7425,N_2723,N_1579);
nand U7426 (N_7426,N_615,N_165);
or U7427 (N_7427,N_277,N_3254);
nand U7428 (N_7428,N_3290,N_1365);
nor U7429 (N_7429,N_2890,N_3174);
nor U7430 (N_7430,N_1459,N_4549);
nand U7431 (N_7431,N_4781,N_2826);
or U7432 (N_7432,N_112,N_1220);
or U7433 (N_7433,N_3847,N_471);
nor U7434 (N_7434,N_2083,N_4875);
nand U7435 (N_7435,N_1761,N_3370);
nand U7436 (N_7436,N_119,N_3707);
and U7437 (N_7437,N_941,N_2488);
nor U7438 (N_7438,N_2023,N_1821);
xnor U7439 (N_7439,N_2368,N_1310);
and U7440 (N_7440,N_3818,N_3768);
and U7441 (N_7441,N_4935,N_3146);
and U7442 (N_7442,N_583,N_4346);
and U7443 (N_7443,N_1909,N_2208);
xor U7444 (N_7444,N_4901,N_2694);
nand U7445 (N_7445,N_1515,N_2029);
and U7446 (N_7446,N_3286,N_2502);
nor U7447 (N_7447,N_4204,N_1673);
nand U7448 (N_7448,N_2108,N_3392);
and U7449 (N_7449,N_1592,N_2535);
and U7450 (N_7450,N_2925,N_2832);
and U7451 (N_7451,N_3521,N_2750);
and U7452 (N_7452,N_1232,N_1200);
and U7453 (N_7453,N_1813,N_2030);
nand U7454 (N_7454,N_32,N_3298);
nand U7455 (N_7455,N_3764,N_4477);
and U7456 (N_7456,N_3608,N_4931);
xnor U7457 (N_7457,N_2530,N_2315);
and U7458 (N_7458,N_1572,N_3878);
xnor U7459 (N_7459,N_1741,N_4132);
xor U7460 (N_7460,N_3629,N_713);
nand U7461 (N_7461,N_1839,N_3496);
and U7462 (N_7462,N_1808,N_300);
nor U7463 (N_7463,N_3914,N_3242);
nand U7464 (N_7464,N_1201,N_2265);
and U7465 (N_7465,N_4128,N_4262);
xnor U7466 (N_7466,N_924,N_3115);
or U7467 (N_7467,N_4036,N_4435);
nand U7468 (N_7468,N_1231,N_3596);
or U7469 (N_7469,N_3457,N_4869);
or U7470 (N_7470,N_1965,N_4886);
nor U7471 (N_7471,N_4841,N_1607);
or U7472 (N_7472,N_339,N_2243);
nand U7473 (N_7473,N_2094,N_4412);
or U7474 (N_7474,N_1510,N_2911);
nor U7475 (N_7475,N_4637,N_4362);
nand U7476 (N_7476,N_1507,N_4741);
nor U7477 (N_7477,N_4624,N_2979);
or U7478 (N_7478,N_3359,N_1349);
or U7479 (N_7479,N_3576,N_3073);
nand U7480 (N_7480,N_3930,N_2705);
or U7481 (N_7481,N_1312,N_1564);
xnor U7482 (N_7482,N_1291,N_3094);
or U7483 (N_7483,N_3184,N_2629);
nand U7484 (N_7484,N_869,N_1485);
and U7485 (N_7485,N_395,N_2831);
nand U7486 (N_7486,N_2931,N_3591);
xnor U7487 (N_7487,N_4562,N_2288);
nand U7488 (N_7488,N_1900,N_4314);
or U7489 (N_7489,N_4943,N_1320);
nor U7490 (N_7490,N_216,N_2492);
and U7491 (N_7491,N_4910,N_63);
and U7492 (N_7492,N_3682,N_2781);
xnor U7493 (N_7493,N_4510,N_1226);
nor U7494 (N_7494,N_3465,N_318);
or U7495 (N_7495,N_1977,N_101);
nor U7496 (N_7496,N_2722,N_4263);
and U7497 (N_7497,N_4760,N_52);
or U7498 (N_7498,N_3534,N_1573);
and U7499 (N_7499,N_1017,N_4243);
or U7500 (N_7500,N_3676,N_4546);
nor U7501 (N_7501,N_2275,N_978);
nor U7502 (N_7502,N_798,N_2295);
nor U7503 (N_7503,N_2100,N_2595);
or U7504 (N_7504,N_202,N_921);
nor U7505 (N_7505,N_808,N_242);
nor U7506 (N_7506,N_2298,N_4446);
nand U7507 (N_7507,N_330,N_2113);
nor U7508 (N_7508,N_4126,N_4710);
or U7509 (N_7509,N_3946,N_1506);
nor U7510 (N_7510,N_3793,N_3056);
nor U7511 (N_7511,N_2825,N_973);
nor U7512 (N_7512,N_3156,N_2635);
xor U7513 (N_7513,N_4629,N_1719);
and U7514 (N_7514,N_634,N_1123);
nor U7515 (N_7515,N_1744,N_2524);
nor U7516 (N_7516,N_4715,N_3690);
nand U7517 (N_7517,N_1150,N_4803);
nor U7518 (N_7518,N_1387,N_2706);
nor U7519 (N_7519,N_809,N_3446);
nand U7520 (N_7520,N_2476,N_4446);
nand U7521 (N_7521,N_3079,N_4227);
and U7522 (N_7522,N_414,N_1436);
or U7523 (N_7523,N_4951,N_1137);
xor U7524 (N_7524,N_3326,N_4733);
and U7525 (N_7525,N_4705,N_1975);
nand U7526 (N_7526,N_4452,N_3973);
nand U7527 (N_7527,N_2065,N_1188);
or U7528 (N_7528,N_4278,N_4196);
or U7529 (N_7529,N_4814,N_4372);
or U7530 (N_7530,N_4808,N_2068);
and U7531 (N_7531,N_956,N_2112);
nand U7532 (N_7532,N_2449,N_184);
nand U7533 (N_7533,N_1527,N_4267);
and U7534 (N_7534,N_351,N_243);
nor U7535 (N_7535,N_1345,N_1693);
or U7536 (N_7536,N_675,N_4365);
nor U7537 (N_7537,N_3170,N_448);
nor U7538 (N_7538,N_4094,N_4327);
nand U7539 (N_7539,N_3024,N_3075);
or U7540 (N_7540,N_3923,N_3632);
xor U7541 (N_7541,N_3658,N_2313);
or U7542 (N_7542,N_2194,N_1500);
and U7543 (N_7543,N_1933,N_4511);
nor U7544 (N_7544,N_1928,N_2810);
and U7545 (N_7545,N_1303,N_4095);
and U7546 (N_7546,N_2432,N_2672);
nand U7547 (N_7547,N_4917,N_306);
nor U7548 (N_7548,N_648,N_100);
nor U7549 (N_7549,N_1984,N_4518);
and U7550 (N_7550,N_4676,N_1642);
nor U7551 (N_7551,N_799,N_3013);
xor U7552 (N_7552,N_1339,N_3525);
or U7553 (N_7553,N_2003,N_1384);
nand U7554 (N_7554,N_1931,N_2461);
nand U7555 (N_7555,N_4369,N_1917);
and U7556 (N_7556,N_1075,N_3822);
nor U7557 (N_7557,N_3294,N_1508);
or U7558 (N_7558,N_3631,N_3838);
and U7559 (N_7559,N_1374,N_1392);
nor U7560 (N_7560,N_203,N_1368);
nor U7561 (N_7561,N_2710,N_2103);
nor U7562 (N_7562,N_4767,N_1821);
or U7563 (N_7563,N_2547,N_2346);
and U7564 (N_7564,N_54,N_3594);
or U7565 (N_7565,N_2570,N_2382);
nor U7566 (N_7566,N_711,N_4802);
and U7567 (N_7567,N_2773,N_1716);
or U7568 (N_7568,N_2271,N_2881);
or U7569 (N_7569,N_2557,N_531);
nand U7570 (N_7570,N_183,N_3651);
and U7571 (N_7571,N_477,N_3263);
xnor U7572 (N_7572,N_3276,N_2998);
nand U7573 (N_7573,N_3952,N_1335);
nand U7574 (N_7574,N_4659,N_2551);
and U7575 (N_7575,N_1839,N_1080);
or U7576 (N_7576,N_573,N_3424);
nand U7577 (N_7577,N_2010,N_173);
or U7578 (N_7578,N_4307,N_3053);
nand U7579 (N_7579,N_4736,N_3347);
or U7580 (N_7580,N_3382,N_573);
or U7581 (N_7581,N_3649,N_4885);
nor U7582 (N_7582,N_2657,N_2767);
nand U7583 (N_7583,N_1342,N_3356);
nand U7584 (N_7584,N_2107,N_2862);
or U7585 (N_7585,N_3833,N_1909);
xnor U7586 (N_7586,N_3203,N_2238);
nor U7587 (N_7587,N_4263,N_4243);
and U7588 (N_7588,N_3345,N_288);
nand U7589 (N_7589,N_804,N_3521);
nand U7590 (N_7590,N_3486,N_1616);
nand U7591 (N_7591,N_174,N_2260);
and U7592 (N_7592,N_48,N_4781);
nor U7593 (N_7593,N_200,N_1722);
nor U7594 (N_7594,N_4616,N_4277);
nor U7595 (N_7595,N_1064,N_92);
nor U7596 (N_7596,N_2399,N_2548);
or U7597 (N_7597,N_1844,N_4039);
xnor U7598 (N_7598,N_2630,N_3837);
nor U7599 (N_7599,N_251,N_2415);
or U7600 (N_7600,N_3278,N_3414);
or U7601 (N_7601,N_4859,N_1290);
or U7602 (N_7602,N_2137,N_1306);
xnor U7603 (N_7603,N_1139,N_3255);
nand U7604 (N_7604,N_2725,N_122);
nand U7605 (N_7605,N_1070,N_4444);
or U7606 (N_7606,N_3085,N_1653);
nor U7607 (N_7607,N_2544,N_1159);
nor U7608 (N_7608,N_1355,N_3883);
or U7609 (N_7609,N_4981,N_3387);
nor U7610 (N_7610,N_4245,N_2141);
nand U7611 (N_7611,N_3055,N_2670);
and U7612 (N_7612,N_4278,N_2511);
and U7613 (N_7613,N_3110,N_1577);
nor U7614 (N_7614,N_3030,N_466);
nor U7615 (N_7615,N_3312,N_4362);
nor U7616 (N_7616,N_2642,N_4042);
nor U7617 (N_7617,N_2434,N_3170);
nand U7618 (N_7618,N_625,N_2205);
and U7619 (N_7619,N_4715,N_2721);
or U7620 (N_7620,N_1666,N_3923);
or U7621 (N_7621,N_993,N_2615);
nand U7622 (N_7622,N_1142,N_1930);
and U7623 (N_7623,N_1404,N_3192);
and U7624 (N_7624,N_840,N_4867);
nor U7625 (N_7625,N_3764,N_3853);
or U7626 (N_7626,N_1918,N_3918);
and U7627 (N_7627,N_3946,N_1079);
or U7628 (N_7628,N_880,N_1314);
nor U7629 (N_7629,N_2116,N_846);
nand U7630 (N_7630,N_2770,N_4174);
and U7631 (N_7631,N_3616,N_495);
nand U7632 (N_7632,N_3504,N_4331);
nand U7633 (N_7633,N_2735,N_1632);
nand U7634 (N_7634,N_1076,N_4727);
and U7635 (N_7635,N_946,N_3398);
and U7636 (N_7636,N_4452,N_2536);
nor U7637 (N_7637,N_4908,N_1566);
nor U7638 (N_7638,N_146,N_2022);
and U7639 (N_7639,N_4986,N_278);
nand U7640 (N_7640,N_3953,N_637);
and U7641 (N_7641,N_1170,N_1983);
or U7642 (N_7642,N_1670,N_3134);
and U7643 (N_7643,N_941,N_890);
or U7644 (N_7644,N_2948,N_1178);
nor U7645 (N_7645,N_79,N_1469);
or U7646 (N_7646,N_698,N_4608);
nor U7647 (N_7647,N_4649,N_4469);
nor U7648 (N_7648,N_4954,N_1718);
xor U7649 (N_7649,N_3054,N_3815);
nor U7650 (N_7650,N_708,N_4497);
or U7651 (N_7651,N_438,N_695);
nand U7652 (N_7652,N_2472,N_2145);
nand U7653 (N_7653,N_3175,N_862);
or U7654 (N_7654,N_4252,N_3682);
nand U7655 (N_7655,N_3016,N_4393);
nor U7656 (N_7656,N_1756,N_1920);
nor U7657 (N_7657,N_3466,N_4279);
nand U7658 (N_7658,N_47,N_542);
and U7659 (N_7659,N_3824,N_1782);
nor U7660 (N_7660,N_1493,N_4533);
nand U7661 (N_7661,N_3661,N_4531);
and U7662 (N_7662,N_3335,N_333);
nor U7663 (N_7663,N_3743,N_4639);
nand U7664 (N_7664,N_1417,N_4865);
xnor U7665 (N_7665,N_4315,N_1659);
or U7666 (N_7666,N_3807,N_4443);
nand U7667 (N_7667,N_3064,N_2429);
nand U7668 (N_7668,N_2531,N_34);
or U7669 (N_7669,N_3974,N_4916);
xnor U7670 (N_7670,N_1958,N_4918);
or U7671 (N_7671,N_1742,N_2226);
xor U7672 (N_7672,N_3141,N_4278);
nand U7673 (N_7673,N_3705,N_1737);
nor U7674 (N_7674,N_1304,N_4444);
or U7675 (N_7675,N_2784,N_2253);
xor U7676 (N_7676,N_388,N_3406);
or U7677 (N_7677,N_3476,N_284);
and U7678 (N_7678,N_2493,N_68);
or U7679 (N_7679,N_504,N_3972);
nor U7680 (N_7680,N_3644,N_2054);
and U7681 (N_7681,N_3367,N_1300);
nand U7682 (N_7682,N_3343,N_853);
and U7683 (N_7683,N_2801,N_2361);
xor U7684 (N_7684,N_2268,N_3592);
xor U7685 (N_7685,N_1156,N_214);
nor U7686 (N_7686,N_4918,N_2404);
nand U7687 (N_7687,N_3155,N_1748);
nor U7688 (N_7688,N_2988,N_2486);
or U7689 (N_7689,N_3483,N_567);
and U7690 (N_7690,N_2536,N_3755);
nand U7691 (N_7691,N_1010,N_1210);
nor U7692 (N_7692,N_43,N_4315);
nand U7693 (N_7693,N_124,N_1369);
or U7694 (N_7694,N_3186,N_4220);
nand U7695 (N_7695,N_899,N_767);
or U7696 (N_7696,N_3171,N_1297);
nor U7697 (N_7697,N_3130,N_1712);
nor U7698 (N_7698,N_3011,N_1583);
nand U7699 (N_7699,N_4257,N_4833);
nor U7700 (N_7700,N_2372,N_1634);
nand U7701 (N_7701,N_356,N_493);
nor U7702 (N_7702,N_818,N_2772);
nand U7703 (N_7703,N_2556,N_2060);
or U7704 (N_7704,N_2033,N_1648);
nor U7705 (N_7705,N_861,N_3633);
or U7706 (N_7706,N_4628,N_2235);
and U7707 (N_7707,N_4591,N_959);
xor U7708 (N_7708,N_59,N_1523);
nand U7709 (N_7709,N_28,N_3520);
or U7710 (N_7710,N_4160,N_3770);
and U7711 (N_7711,N_1900,N_2867);
nand U7712 (N_7712,N_3850,N_3460);
and U7713 (N_7713,N_3383,N_3784);
and U7714 (N_7714,N_3082,N_3203);
nand U7715 (N_7715,N_4631,N_2477);
or U7716 (N_7716,N_1261,N_4620);
nor U7717 (N_7717,N_4821,N_3039);
or U7718 (N_7718,N_2728,N_1338);
nor U7719 (N_7719,N_1837,N_4106);
or U7720 (N_7720,N_766,N_609);
nor U7721 (N_7721,N_839,N_736);
nor U7722 (N_7722,N_1778,N_850);
nand U7723 (N_7723,N_4446,N_1729);
xor U7724 (N_7724,N_886,N_1715);
nand U7725 (N_7725,N_3512,N_4850);
nand U7726 (N_7726,N_4994,N_2815);
nor U7727 (N_7727,N_538,N_4225);
and U7728 (N_7728,N_4465,N_1138);
xor U7729 (N_7729,N_593,N_417);
nor U7730 (N_7730,N_3875,N_1805);
xor U7731 (N_7731,N_2748,N_2846);
nand U7732 (N_7732,N_2927,N_1545);
nand U7733 (N_7733,N_3065,N_3688);
or U7734 (N_7734,N_3104,N_3307);
and U7735 (N_7735,N_2621,N_3159);
and U7736 (N_7736,N_583,N_4549);
or U7737 (N_7737,N_2757,N_1087);
and U7738 (N_7738,N_1293,N_4753);
xnor U7739 (N_7739,N_2277,N_3566);
or U7740 (N_7740,N_3070,N_729);
nand U7741 (N_7741,N_2287,N_4141);
nand U7742 (N_7742,N_1314,N_578);
or U7743 (N_7743,N_2450,N_665);
nand U7744 (N_7744,N_3757,N_2723);
and U7745 (N_7745,N_376,N_828);
or U7746 (N_7746,N_2738,N_2360);
xnor U7747 (N_7747,N_4277,N_3604);
or U7748 (N_7748,N_2504,N_4730);
or U7749 (N_7749,N_2274,N_714);
or U7750 (N_7750,N_3139,N_2705);
or U7751 (N_7751,N_1854,N_2217);
nand U7752 (N_7752,N_2454,N_1462);
nand U7753 (N_7753,N_102,N_4450);
nor U7754 (N_7754,N_2441,N_3988);
nand U7755 (N_7755,N_4859,N_1015);
xnor U7756 (N_7756,N_897,N_746);
or U7757 (N_7757,N_1432,N_1947);
and U7758 (N_7758,N_3504,N_3456);
xor U7759 (N_7759,N_1851,N_4115);
and U7760 (N_7760,N_1179,N_3051);
xnor U7761 (N_7761,N_662,N_92);
nand U7762 (N_7762,N_2871,N_373);
or U7763 (N_7763,N_2311,N_2667);
or U7764 (N_7764,N_4993,N_3811);
nor U7765 (N_7765,N_1713,N_2756);
and U7766 (N_7766,N_2639,N_1608);
nor U7767 (N_7767,N_1089,N_514);
or U7768 (N_7768,N_1451,N_3985);
xnor U7769 (N_7769,N_3877,N_582);
and U7770 (N_7770,N_2112,N_4916);
or U7771 (N_7771,N_1284,N_1212);
nand U7772 (N_7772,N_1181,N_4975);
nand U7773 (N_7773,N_2583,N_212);
and U7774 (N_7774,N_1576,N_3732);
and U7775 (N_7775,N_685,N_1731);
xor U7776 (N_7776,N_995,N_3695);
or U7777 (N_7777,N_3021,N_2400);
nor U7778 (N_7778,N_3481,N_1738);
nand U7779 (N_7779,N_850,N_584);
or U7780 (N_7780,N_2697,N_2756);
or U7781 (N_7781,N_2564,N_1157);
nand U7782 (N_7782,N_1914,N_71);
nand U7783 (N_7783,N_3973,N_1401);
nor U7784 (N_7784,N_633,N_25);
nand U7785 (N_7785,N_1833,N_1720);
and U7786 (N_7786,N_4147,N_304);
and U7787 (N_7787,N_4904,N_3833);
nor U7788 (N_7788,N_1027,N_4389);
nand U7789 (N_7789,N_1139,N_4337);
or U7790 (N_7790,N_4157,N_3178);
xnor U7791 (N_7791,N_37,N_2074);
nor U7792 (N_7792,N_1028,N_3189);
nor U7793 (N_7793,N_3622,N_4658);
or U7794 (N_7794,N_3545,N_1207);
nor U7795 (N_7795,N_1808,N_1610);
nand U7796 (N_7796,N_4916,N_2104);
and U7797 (N_7797,N_1118,N_4264);
nand U7798 (N_7798,N_4976,N_360);
nand U7799 (N_7799,N_3616,N_3178);
nor U7800 (N_7800,N_2947,N_2998);
nand U7801 (N_7801,N_2497,N_3597);
and U7802 (N_7802,N_2001,N_615);
xor U7803 (N_7803,N_2958,N_2112);
nand U7804 (N_7804,N_4588,N_3515);
xor U7805 (N_7805,N_4732,N_3077);
nor U7806 (N_7806,N_355,N_3346);
or U7807 (N_7807,N_2661,N_3959);
nand U7808 (N_7808,N_3508,N_3090);
nor U7809 (N_7809,N_1787,N_3968);
and U7810 (N_7810,N_2937,N_2068);
or U7811 (N_7811,N_2506,N_1528);
nor U7812 (N_7812,N_1134,N_408);
nor U7813 (N_7813,N_2237,N_3862);
nand U7814 (N_7814,N_71,N_466);
or U7815 (N_7815,N_2468,N_946);
nand U7816 (N_7816,N_488,N_3033);
or U7817 (N_7817,N_628,N_4526);
nand U7818 (N_7818,N_1635,N_4879);
or U7819 (N_7819,N_779,N_4178);
xnor U7820 (N_7820,N_3198,N_1345);
nand U7821 (N_7821,N_740,N_4138);
and U7822 (N_7822,N_2556,N_1627);
or U7823 (N_7823,N_2486,N_2842);
nand U7824 (N_7824,N_1575,N_2795);
and U7825 (N_7825,N_141,N_894);
or U7826 (N_7826,N_3520,N_3690);
nand U7827 (N_7827,N_1878,N_2230);
nand U7828 (N_7828,N_3972,N_1435);
nor U7829 (N_7829,N_3580,N_3013);
xnor U7830 (N_7830,N_2457,N_1425);
and U7831 (N_7831,N_3219,N_1054);
xnor U7832 (N_7832,N_3353,N_284);
nand U7833 (N_7833,N_1177,N_2754);
or U7834 (N_7834,N_1247,N_3081);
xor U7835 (N_7835,N_1407,N_2667);
nor U7836 (N_7836,N_2805,N_3955);
or U7837 (N_7837,N_414,N_1737);
nor U7838 (N_7838,N_2349,N_413);
nand U7839 (N_7839,N_4986,N_2069);
or U7840 (N_7840,N_2117,N_2087);
or U7841 (N_7841,N_3720,N_2768);
nor U7842 (N_7842,N_640,N_2302);
nor U7843 (N_7843,N_3186,N_3458);
xor U7844 (N_7844,N_690,N_4782);
nor U7845 (N_7845,N_431,N_3747);
xor U7846 (N_7846,N_923,N_4687);
nor U7847 (N_7847,N_2660,N_1130);
and U7848 (N_7848,N_1331,N_2603);
or U7849 (N_7849,N_1830,N_2175);
nor U7850 (N_7850,N_61,N_798);
xor U7851 (N_7851,N_4330,N_1458);
nor U7852 (N_7852,N_898,N_3235);
xnor U7853 (N_7853,N_4884,N_371);
or U7854 (N_7854,N_3603,N_2280);
nand U7855 (N_7855,N_4011,N_4977);
or U7856 (N_7856,N_4161,N_1573);
or U7857 (N_7857,N_3158,N_812);
and U7858 (N_7858,N_3468,N_1322);
nand U7859 (N_7859,N_3037,N_4980);
nand U7860 (N_7860,N_4011,N_3898);
nand U7861 (N_7861,N_729,N_3132);
nand U7862 (N_7862,N_4021,N_2480);
or U7863 (N_7863,N_1035,N_571);
nor U7864 (N_7864,N_115,N_119);
and U7865 (N_7865,N_2770,N_191);
or U7866 (N_7866,N_953,N_3046);
and U7867 (N_7867,N_1042,N_550);
nand U7868 (N_7868,N_3528,N_4804);
nand U7869 (N_7869,N_3400,N_1477);
nand U7870 (N_7870,N_4536,N_1254);
or U7871 (N_7871,N_530,N_2990);
xor U7872 (N_7872,N_3444,N_508);
nand U7873 (N_7873,N_56,N_2261);
and U7874 (N_7874,N_3781,N_3354);
nor U7875 (N_7875,N_2177,N_2099);
nand U7876 (N_7876,N_2164,N_2070);
and U7877 (N_7877,N_795,N_3036);
and U7878 (N_7878,N_4971,N_4208);
or U7879 (N_7879,N_584,N_3430);
nor U7880 (N_7880,N_626,N_4672);
or U7881 (N_7881,N_4367,N_331);
nand U7882 (N_7882,N_849,N_1479);
or U7883 (N_7883,N_4483,N_912);
nor U7884 (N_7884,N_265,N_3605);
nor U7885 (N_7885,N_2544,N_1278);
nand U7886 (N_7886,N_3097,N_3422);
nand U7887 (N_7887,N_1651,N_2958);
or U7888 (N_7888,N_3083,N_1724);
and U7889 (N_7889,N_133,N_530);
nor U7890 (N_7890,N_1786,N_2504);
nor U7891 (N_7891,N_2795,N_1260);
nor U7892 (N_7892,N_3013,N_812);
and U7893 (N_7893,N_59,N_1397);
nand U7894 (N_7894,N_34,N_2819);
nand U7895 (N_7895,N_1239,N_1925);
or U7896 (N_7896,N_1287,N_2110);
or U7897 (N_7897,N_1785,N_4909);
or U7898 (N_7898,N_1343,N_1362);
nor U7899 (N_7899,N_4606,N_444);
and U7900 (N_7900,N_551,N_3592);
xnor U7901 (N_7901,N_4454,N_351);
xor U7902 (N_7902,N_1256,N_516);
nand U7903 (N_7903,N_2409,N_844);
nor U7904 (N_7904,N_2883,N_3475);
nand U7905 (N_7905,N_3829,N_663);
and U7906 (N_7906,N_460,N_2574);
or U7907 (N_7907,N_1048,N_836);
xor U7908 (N_7908,N_3717,N_3952);
nand U7909 (N_7909,N_3366,N_4173);
or U7910 (N_7910,N_4257,N_2963);
and U7911 (N_7911,N_484,N_628);
nor U7912 (N_7912,N_1082,N_2692);
nand U7913 (N_7913,N_4130,N_1429);
nand U7914 (N_7914,N_2791,N_2361);
or U7915 (N_7915,N_838,N_3657);
and U7916 (N_7916,N_2359,N_484);
or U7917 (N_7917,N_1704,N_3584);
or U7918 (N_7918,N_4969,N_1095);
or U7919 (N_7919,N_311,N_2292);
nor U7920 (N_7920,N_2690,N_2693);
or U7921 (N_7921,N_2747,N_3407);
nor U7922 (N_7922,N_4100,N_3901);
or U7923 (N_7923,N_3701,N_4502);
nor U7924 (N_7924,N_4287,N_586);
xnor U7925 (N_7925,N_538,N_1297);
or U7926 (N_7926,N_1744,N_1594);
and U7927 (N_7927,N_2781,N_820);
nor U7928 (N_7928,N_2937,N_2728);
or U7929 (N_7929,N_4190,N_3386);
nor U7930 (N_7930,N_4586,N_3881);
and U7931 (N_7931,N_1503,N_835);
or U7932 (N_7932,N_354,N_2998);
or U7933 (N_7933,N_0,N_4710);
and U7934 (N_7934,N_4723,N_2205);
nor U7935 (N_7935,N_150,N_1377);
and U7936 (N_7936,N_383,N_110);
nand U7937 (N_7937,N_4970,N_4993);
xor U7938 (N_7938,N_3657,N_1801);
and U7939 (N_7939,N_4703,N_2966);
or U7940 (N_7940,N_871,N_2411);
or U7941 (N_7941,N_325,N_1218);
nor U7942 (N_7942,N_2770,N_748);
nand U7943 (N_7943,N_2028,N_1231);
nor U7944 (N_7944,N_4089,N_2008);
or U7945 (N_7945,N_3301,N_4005);
or U7946 (N_7946,N_1884,N_1766);
nor U7947 (N_7947,N_2630,N_2877);
nand U7948 (N_7948,N_3249,N_2816);
nand U7949 (N_7949,N_310,N_3688);
and U7950 (N_7950,N_36,N_3835);
nand U7951 (N_7951,N_4482,N_1573);
or U7952 (N_7952,N_3509,N_2266);
or U7953 (N_7953,N_1336,N_4393);
nand U7954 (N_7954,N_998,N_1992);
nand U7955 (N_7955,N_286,N_2672);
nand U7956 (N_7956,N_3216,N_868);
nor U7957 (N_7957,N_1201,N_3702);
and U7958 (N_7958,N_3964,N_1491);
or U7959 (N_7959,N_2471,N_4256);
nand U7960 (N_7960,N_3523,N_4431);
and U7961 (N_7961,N_48,N_1870);
nand U7962 (N_7962,N_2442,N_1102);
nor U7963 (N_7963,N_204,N_745);
nand U7964 (N_7964,N_1383,N_2936);
nor U7965 (N_7965,N_1365,N_1414);
or U7966 (N_7966,N_3275,N_1159);
nor U7967 (N_7967,N_2999,N_4181);
nand U7968 (N_7968,N_2088,N_4039);
and U7969 (N_7969,N_279,N_1965);
xor U7970 (N_7970,N_888,N_2366);
or U7971 (N_7971,N_3247,N_1923);
and U7972 (N_7972,N_1828,N_1452);
and U7973 (N_7973,N_3192,N_4391);
nand U7974 (N_7974,N_376,N_4761);
nor U7975 (N_7975,N_1140,N_1378);
xnor U7976 (N_7976,N_248,N_2044);
or U7977 (N_7977,N_1443,N_2138);
nand U7978 (N_7978,N_1028,N_4227);
nand U7979 (N_7979,N_1213,N_986);
and U7980 (N_7980,N_4139,N_452);
or U7981 (N_7981,N_3346,N_527);
nor U7982 (N_7982,N_788,N_127);
xnor U7983 (N_7983,N_4301,N_1092);
and U7984 (N_7984,N_2480,N_4384);
xor U7985 (N_7985,N_4082,N_1364);
or U7986 (N_7986,N_2057,N_4487);
nor U7987 (N_7987,N_1508,N_4198);
or U7988 (N_7988,N_3270,N_1329);
and U7989 (N_7989,N_1196,N_4493);
or U7990 (N_7990,N_2481,N_3378);
nor U7991 (N_7991,N_3186,N_1429);
and U7992 (N_7992,N_2207,N_652);
nor U7993 (N_7993,N_3238,N_2140);
nor U7994 (N_7994,N_2311,N_2809);
and U7995 (N_7995,N_3183,N_1755);
or U7996 (N_7996,N_1940,N_4967);
nor U7997 (N_7997,N_4813,N_4799);
nor U7998 (N_7998,N_1061,N_4737);
and U7999 (N_7999,N_3690,N_3419);
nand U8000 (N_8000,N_1423,N_3898);
and U8001 (N_8001,N_256,N_2535);
and U8002 (N_8002,N_2358,N_982);
nor U8003 (N_8003,N_740,N_59);
or U8004 (N_8004,N_1209,N_1067);
nand U8005 (N_8005,N_3781,N_1055);
and U8006 (N_8006,N_3128,N_2223);
and U8007 (N_8007,N_2961,N_3862);
and U8008 (N_8008,N_201,N_4910);
nor U8009 (N_8009,N_2504,N_1519);
nor U8010 (N_8010,N_2810,N_247);
nand U8011 (N_8011,N_2888,N_1760);
nand U8012 (N_8012,N_4444,N_4461);
nand U8013 (N_8013,N_4345,N_4118);
and U8014 (N_8014,N_3300,N_1552);
and U8015 (N_8015,N_2221,N_2416);
nor U8016 (N_8016,N_3482,N_3337);
and U8017 (N_8017,N_1792,N_3064);
nand U8018 (N_8018,N_525,N_761);
or U8019 (N_8019,N_1946,N_4190);
nor U8020 (N_8020,N_38,N_4668);
and U8021 (N_8021,N_3932,N_2690);
and U8022 (N_8022,N_2339,N_3644);
nand U8023 (N_8023,N_3952,N_317);
or U8024 (N_8024,N_1895,N_4141);
and U8025 (N_8025,N_2246,N_25);
nor U8026 (N_8026,N_4978,N_1059);
xor U8027 (N_8027,N_1956,N_2993);
nor U8028 (N_8028,N_2204,N_368);
and U8029 (N_8029,N_1160,N_3541);
and U8030 (N_8030,N_4832,N_2101);
and U8031 (N_8031,N_3228,N_344);
nor U8032 (N_8032,N_1936,N_2580);
or U8033 (N_8033,N_3320,N_3443);
nor U8034 (N_8034,N_135,N_3250);
nor U8035 (N_8035,N_1444,N_4680);
nand U8036 (N_8036,N_2276,N_4395);
or U8037 (N_8037,N_3883,N_4345);
nand U8038 (N_8038,N_2718,N_1662);
nand U8039 (N_8039,N_4104,N_2471);
nor U8040 (N_8040,N_1877,N_2983);
or U8041 (N_8041,N_3858,N_3354);
nand U8042 (N_8042,N_408,N_3319);
or U8043 (N_8043,N_1227,N_2775);
nand U8044 (N_8044,N_3270,N_686);
or U8045 (N_8045,N_2411,N_779);
or U8046 (N_8046,N_3840,N_3792);
xor U8047 (N_8047,N_4161,N_4024);
or U8048 (N_8048,N_758,N_4229);
nand U8049 (N_8049,N_188,N_1707);
or U8050 (N_8050,N_4731,N_1357);
and U8051 (N_8051,N_3922,N_2601);
nor U8052 (N_8052,N_2880,N_2409);
or U8053 (N_8053,N_4722,N_1760);
xor U8054 (N_8054,N_4662,N_3856);
nor U8055 (N_8055,N_2690,N_3779);
nor U8056 (N_8056,N_2987,N_3539);
nand U8057 (N_8057,N_4862,N_4547);
nor U8058 (N_8058,N_3261,N_3812);
or U8059 (N_8059,N_1163,N_830);
nor U8060 (N_8060,N_3271,N_2592);
nand U8061 (N_8061,N_1921,N_3877);
or U8062 (N_8062,N_3059,N_2711);
nor U8063 (N_8063,N_4755,N_1457);
nand U8064 (N_8064,N_144,N_2753);
nand U8065 (N_8065,N_174,N_1692);
xor U8066 (N_8066,N_536,N_137);
nand U8067 (N_8067,N_1632,N_4903);
xnor U8068 (N_8068,N_2949,N_387);
and U8069 (N_8069,N_3849,N_2423);
xnor U8070 (N_8070,N_4172,N_365);
nand U8071 (N_8071,N_4244,N_2620);
or U8072 (N_8072,N_4754,N_3774);
or U8073 (N_8073,N_2684,N_2755);
and U8074 (N_8074,N_2467,N_2403);
or U8075 (N_8075,N_4995,N_748);
and U8076 (N_8076,N_4495,N_600);
nor U8077 (N_8077,N_1739,N_3003);
nand U8078 (N_8078,N_1785,N_333);
nand U8079 (N_8079,N_104,N_1836);
nor U8080 (N_8080,N_3366,N_2001);
xor U8081 (N_8081,N_3379,N_624);
and U8082 (N_8082,N_3793,N_4160);
xnor U8083 (N_8083,N_660,N_892);
nand U8084 (N_8084,N_1590,N_1091);
nand U8085 (N_8085,N_2979,N_4981);
or U8086 (N_8086,N_1099,N_4981);
nand U8087 (N_8087,N_3040,N_3335);
nor U8088 (N_8088,N_1595,N_3990);
and U8089 (N_8089,N_2283,N_3702);
and U8090 (N_8090,N_1137,N_716);
or U8091 (N_8091,N_4131,N_4693);
or U8092 (N_8092,N_3785,N_3022);
nor U8093 (N_8093,N_964,N_4100);
or U8094 (N_8094,N_871,N_1069);
nor U8095 (N_8095,N_3352,N_695);
or U8096 (N_8096,N_3370,N_2670);
and U8097 (N_8097,N_4952,N_255);
nand U8098 (N_8098,N_2992,N_3686);
nand U8099 (N_8099,N_781,N_4056);
nand U8100 (N_8100,N_2836,N_1677);
nor U8101 (N_8101,N_1271,N_4917);
nand U8102 (N_8102,N_673,N_2175);
and U8103 (N_8103,N_1710,N_723);
xnor U8104 (N_8104,N_3669,N_353);
nand U8105 (N_8105,N_4722,N_4808);
and U8106 (N_8106,N_4185,N_1504);
and U8107 (N_8107,N_154,N_327);
xor U8108 (N_8108,N_3890,N_3017);
nor U8109 (N_8109,N_1201,N_2777);
and U8110 (N_8110,N_2174,N_838);
nor U8111 (N_8111,N_4669,N_1663);
or U8112 (N_8112,N_2380,N_3046);
nand U8113 (N_8113,N_3534,N_3398);
or U8114 (N_8114,N_3160,N_1770);
nand U8115 (N_8115,N_2532,N_3008);
or U8116 (N_8116,N_4076,N_2218);
xnor U8117 (N_8117,N_4006,N_1959);
nand U8118 (N_8118,N_4164,N_1940);
and U8119 (N_8119,N_3237,N_215);
nor U8120 (N_8120,N_2131,N_1472);
nor U8121 (N_8121,N_2909,N_3951);
or U8122 (N_8122,N_767,N_908);
nand U8123 (N_8123,N_4364,N_3383);
nor U8124 (N_8124,N_601,N_454);
xnor U8125 (N_8125,N_2424,N_2658);
xnor U8126 (N_8126,N_4308,N_3985);
xnor U8127 (N_8127,N_197,N_1101);
nor U8128 (N_8128,N_2708,N_4181);
nand U8129 (N_8129,N_4476,N_3998);
and U8130 (N_8130,N_2759,N_4212);
and U8131 (N_8131,N_356,N_1924);
nor U8132 (N_8132,N_3896,N_3531);
and U8133 (N_8133,N_171,N_3798);
nand U8134 (N_8134,N_4422,N_1169);
nand U8135 (N_8135,N_612,N_4309);
nor U8136 (N_8136,N_4461,N_1045);
or U8137 (N_8137,N_4135,N_4511);
and U8138 (N_8138,N_3001,N_1223);
or U8139 (N_8139,N_53,N_4750);
xor U8140 (N_8140,N_383,N_3229);
and U8141 (N_8141,N_547,N_4546);
or U8142 (N_8142,N_1423,N_1326);
nand U8143 (N_8143,N_4729,N_3989);
nor U8144 (N_8144,N_3612,N_610);
and U8145 (N_8145,N_2806,N_3256);
nand U8146 (N_8146,N_3081,N_2067);
and U8147 (N_8147,N_464,N_2709);
or U8148 (N_8148,N_4217,N_158);
or U8149 (N_8149,N_2640,N_1013);
and U8150 (N_8150,N_782,N_2469);
nor U8151 (N_8151,N_3246,N_4410);
and U8152 (N_8152,N_2946,N_3049);
or U8153 (N_8153,N_1061,N_4292);
nor U8154 (N_8154,N_2347,N_1378);
nor U8155 (N_8155,N_4740,N_3771);
and U8156 (N_8156,N_4796,N_4174);
or U8157 (N_8157,N_2501,N_1589);
or U8158 (N_8158,N_3231,N_728);
nor U8159 (N_8159,N_3972,N_3715);
xnor U8160 (N_8160,N_4371,N_2288);
nand U8161 (N_8161,N_4618,N_4755);
nor U8162 (N_8162,N_4547,N_3326);
nor U8163 (N_8163,N_1179,N_3324);
nor U8164 (N_8164,N_2557,N_1524);
nor U8165 (N_8165,N_118,N_1026);
and U8166 (N_8166,N_1359,N_2391);
nor U8167 (N_8167,N_1588,N_1035);
nand U8168 (N_8168,N_3309,N_908);
nor U8169 (N_8169,N_2036,N_2661);
or U8170 (N_8170,N_2072,N_2987);
nor U8171 (N_8171,N_4767,N_782);
or U8172 (N_8172,N_4236,N_4062);
nand U8173 (N_8173,N_1134,N_3737);
and U8174 (N_8174,N_4097,N_4886);
and U8175 (N_8175,N_584,N_166);
or U8176 (N_8176,N_3301,N_4504);
nor U8177 (N_8177,N_3601,N_618);
nand U8178 (N_8178,N_2187,N_3719);
nor U8179 (N_8179,N_27,N_3916);
nor U8180 (N_8180,N_2483,N_2215);
nand U8181 (N_8181,N_4747,N_2063);
and U8182 (N_8182,N_1984,N_606);
or U8183 (N_8183,N_1231,N_1690);
or U8184 (N_8184,N_3449,N_2162);
and U8185 (N_8185,N_671,N_1466);
or U8186 (N_8186,N_2786,N_1300);
nand U8187 (N_8187,N_4046,N_4770);
or U8188 (N_8188,N_2609,N_2499);
xor U8189 (N_8189,N_4570,N_4268);
or U8190 (N_8190,N_3085,N_3546);
nand U8191 (N_8191,N_2982,N_2977);
nor U8192 (N_8192,N_2069,N_2800);
or U8193 (N_8193,N_670,N_2191);
and U8194 (N_8194,N_2907,N_396);
or U8195 (N_8195,N_629,N_884);
xor U8196 (N_8196,N_2701,N_943);
nand U8197 (N_8197,N_748,N_4628);
nor U8198 (N_8198,N_1099,N_3455);
or U8199 (N_8199,N_323,N_4052);
xor U8200 (N_8200,N_363,N_2922);
or U8201 (N_8201,N_4555,N_4179);
and U8202 (N_8202,N_3827,N_3332);
xnor U8203 (N_8203,N_200,N_1713);
xnor U8204 (N_8204,N_4693,N_64);
nand U8205 (N_8205,N_3467,N_854);
or U8206 (N_8206,N_4395,N_4974);
and U8207 (N_8207,N_3115,N_4635);
and U8208 (N_8208,N_1487,N_3856);
xor U8209 (N_8209,N_971,N_4947);
or U8210 (N_8210,N_890,N_2306);
xnor U8211 (N_8211,N_2736,N_1028);
nor U8212 (N_8212,N_4286,N_3267);
or U8213 (N_8213,N_2710,N_2085);
nor U8214 (N_8214,N_4589,N_2065);
and U8215 (N_8215,N_3122,N_4727);
nor U8216 (N_8216,N_10,N_4775);
nor U8217 (N_8217,N_1499,N_1558);
nor U8218 (N_8218,N_3869,N_4032);
or U8219 (N_8219,N_534,N_934);
xor U8220 (N_8220,N_3686,N_3721);
nand U8221 (N_8221,N_1912,N_2211);
nand U8222 (N_8222,N_2550,N_1230);
and U8223 (N_8223,N_455,N_2703);
xor U8224 (N_8224,N_1106,N_1186);
nor U8225 (N_8225,N_716,N_4929);
and U8226 (N_8226,N_530,N_3223);
or U8227 (N_8227,N_2783,N_4264);
or U8228 (N_8228,N_3211,N_1097);
and U8229 (N_8229,N_1053,N_1750);
nand U8230 (N_8230,N_2482,N_1486);
nor U8231 (N_8231,N_1629,N_4043);
and U8232 (N_8232,N_783,N_4291);
and U8233 (N_8233,N_501,N_348);
or U8234 (N_8234,N_1276,N_902);
or U8235 (N_8235,N_3468,N_4080);
nand U8236 (N_8236,N_1790,N_1939);
nor U8237 (N_8237,N_3444,N_2371);
or U8238 (N_8238,N_701,N_1661);
and U8239 (N_8239,N_2995,N_3797);
nor U8240 (N_8240,N_1879,N_633);
and U8241 (N_8241,N_4616,N_3744);
or U8242 (N_8242,N_3655,N_3606);
nor U8243 (N_8243,N_3360,N_303);
xor U8244 (N_8244,N_1142,N_4172);
and U8245 (N_8245,N_2318,N_2365);
and U8246 (N_8246,N_2910,N_2296);
nor U8247 (N_8247,N_800,N_3728);
nor U8248 (N_8248,N_4939,N_450);
xor U8249 (N_8249,N_350,N_3590);
or U8250 (N_8250,N_4867,N_4999);
nor U8251 (N_8251,N_1032,N_2132);
and U8252 (N_8252,N_4778,N_2717);
and U8253 (N_8253,N_1916,N_1275);
nand U8254 (N_8254,N_671,N_550);
nor U8255 (N_8255,N_4351,N_1063);
and U8256 (N_8256,N_3406,N_1580);
nand U8257 (N_8257,N_4287,N_3323);
and U8258 (N_8258,N_3797,N_4065);
xnor U8259 (N_8259,N_2892,N_3262);
or U8260 (N_8260,N_3334,N_2687);
and U8261 (N_8261,N_3280,N_1956);
nand U8262 (N_8262,N_4254,N_4688);
nand U8263 (N_8263,N_3891,N_4826);
or U8264 (N_8264,N_4349,N_4556);
nand U8265 (N_8265,N_4678,N_1265);
nand U8266 (N_8266,N_1089,N_2606);
and U8267 (N_8267,N_579,N_3054);
or U8268 (N_8268,N_3899,N_2534);
nor U8269 (N_8269,N_1706,N_4813);
nor U8270 (N_8270,N_2542,N_3056);
nand U8271 (N_8271,N_2605,N_165);
nor U8272 (N_8272,N_4046,N_3724);
or U8273 (N_8273,N_1855,N_913);
nand U8274 (N_8274,N_4634,N_3857);
nor U8275 (N_8275,N_3016,N_2212);
or U8276 (N_8276,N_2042,N_327);
nand U8277 (N_8277,N_3114,N_1991);
nor U8278 (N_8278,N_3526,N_801);
and U8279 (N_8279,N_3426,N_4726);
xor U8280 (N_8280,N_954,N_4927);
nor U8281 (N_8281,N_629,N_3288);
nor U8282 (N_8282,N_1355,N_3083);
nor U8283 (N_8283,N_2797,N_731);
or U8284 (N_8284,N_163,N_1987);
and U8285 (N_8285,N_1020,N_3699);
and U8286 (N_8286,N_2323,N_1851);
nand U8287 (N_8287,N_1221,N_4446);
nand U8288 (N_8288,N_582,N_3797);
nor U8289 (N_8289,N_1898,N_277);
and U8290 (N_8290,N_2064,N_524);
nor U8291 (N_8291,N_1173,N_1547);
or U8292 (N_8292,N_1860,N_4194);
xor U8293 (N_8293,N_1197,N_3371);
xor U8294 (N_8294,N_851,N_4123);
and U8295 (N_8295,N_287,N_1744);
or U8296 (N_8296,N_2731,N_2512);
nand U8297 (N_8297,N_3731,N_2979);
and U8298 (N_8298,N_4676,N_804);
or U8299 (N_8299,N_1570,N_2642);
nor U8300 (N_8300,N_4280,N_2839);
or U8301 (N_8301,N_4855,N_3890);
nand U8302 (N_8302,N_977,N_4161);
xor U8303 (N_8303,N_3514,N_4221);
nand U8304 (N_8304,N_958,N_4071);
nand U8305 (N_8305,N_1199,N_3286);
xor U8306 (N_8306,N_2768,N_684);
nand U8307 (N_8307,N_1650,N_3254);
or U8308 (N_8308,N_4926,N_502);
xnor U8309 (N_8309,N_4419,N_3252);
and U8310 (N_8310,N_1692,N_4463);
nand U8311 (N_8311,N_4689,N_3881);
nand U8312 (N_8312,N_1469,N_4092);
nand U8313 (N_8313,N_1380,N_4665);
nand U8314 (N_8314,N_2186,N_270);
nor U8315 (N_8315,N_335,N_3213);
or U8316 (N_8316,N_4609,N_1770);
nor U8317 (N_8317,N_924,N_4943);
xor U8318 (N_8318,N_828,N_1822);
nor U8319 (N_8319,N_211,N_2156);
nand U8320 (N_8320,N_3480,N_4569);
xor U8321 (N_8321,N_4141,N_4670);
nand U8322 (N_8322,N_588,N_3460);
nand U8323 (N_8323,N_2072,N_4265);
nand U8324 (N_8324,N_2879,N_4278);
xnor U8325 (N_8325,N_2744,N_4110);
nor U8326 (N_8326,N_3248,N_2362);
or U8327 (N_8327,N_3947,N_2447);
xor U8328 (N_8328,N_547,N_1340);
and U8329 (N_8329,N_260,N_830);
or U8330 (N_8330,N_3989,N_3794);
and U8331 (N_8331,N_1344,N_1733);
or U8332 (N_8332,N_554,N_1794);
nor U8333 (N_8333,N_3619,N_1434);
nor U8334 (N_8334,N_674,N_2878);
and U8335 (N_8335,N_2030,N_1624);
xor U8336 (N_8336,N_1610,N_2845);
or U8337 (N_8337,N_2496,N_163);
nand U8338 (N_8338,N_1996,N_2903);
or U8339 (N_8339,N_2841,N_2842);
and U8340 (N_8340,N_4714,N_2275);
nor U8341 (N_8341,N_3849,N_3770);
nor U8342 (N_8342,N_501,N_3427);
nand U8343 (N_8343,N_1788,N_4808);
or U8344 (N_8344,N_4564,N_1155);
nand U8345 (N_8345,N_2460,N_2516);
nor U8346 (N_8346,N_1511,N_1975);
xnor U8347 (N_8347,N_4584,N_4665);
and U8348 (N_8348,N_3559,N_1482);
nor U8349 (N_8349,N_2852,N_4373);
nand U8350 (N_8350,N_550,N_3651);
nand U8351 (N_8351,N_4625,N_3364);
xnor U8352 (N_8352,N_3303,N_2034);
and U8353 (N_8353,N_4511,N_4123);
and U8354 (N_8354,N_1628,N_694);
and U8355 (N_8355,N_263,N_4640);
nand U8356 (N_8356,N_2699,N_1680);
nor U8357 (N_8357,N_2460,N_560);
nand U8358 (N_8358,N_3638,N_2340);
nor U8359 (N_8359,N_1306,N_1657);
nor U8360 (N_8360,N_4260,N_4506);
and U8361 (N_8361,N_16,N_1912);
or U8362 (N_8362,N_3762,N_3171);
or U8363 (N_8363,N_3960,N_3683);
or U8364 (N_8364,N_3818,N_3221);
or U8365 (N_8365,N_2060,N_4900);
nand U8366 (N_8366,N_1337,N_627);
nand U8367 (N_8367,N_4494,N_1636);
and U8368 (N_8368,N_3423,N_2511);
nand U8369 (N_8369,N_2450,N_2334);
xnor U8370 (N_8370,N_3001,N_3843);
or U8371 (N_8371,N_2160,N_959);
and U8372 (N_8372,N_3150,N_598);
nor U8373 (N_8373,N_1502,N_3100);
nor U8374 (N_8374,N_3644,N_3629);
or U8375 (N_8375,N_4710,N_926);
nor U8376 (N_8376,N_4303,N_115);
nand U8377 (N_8377,N_3815,N_3975);
nand U8378 (N_8378,N_2659,N_411);
and U8379 (N_8379,N_4910,N_865);
nor U8380 (N_8380,N_155,N_2575);
nand U8381 (N_8381,N_686,N_2959);
nor U8382 (N_8382,N_1750,N_1821);
nand U8383 (N_8383,N_1891,N_4100);
or U8384 (N_8384,N_2216,N_4189);
and U8385 (N_8385,N_1127,N_1914);
nand U8386 (N_8386,N_789,N_4115);
nand U8387 (N_8387,N_4579,N_2357);
or U8388 (N_8388,N_4321,N_2999);
or U8389 (N_8389,N_2160,N_4384);
nand U8390 (N_8390,N_2871,N_779);
nand U8391 (N_8391,N_1659,N_4095);
nor U8392 (N_8392,N_3199,N_4384);
or U8393 (N_8393,N_3900,N_290);
or U8394 (N_8394,N_1598,N_2689);
nand U8395 (N_8395,N_3522,N_1936);
xnor U8396 (N_8396,N_4275,N_4383);
nor U8397 (N_8397,N_2898,N_3026);
nand U8398 (N_8398,N_756,N_3985);
or U8399 (N_8399,N_4621,N_1157);
xnor U8400 (N_8400,N_3682,N_4397);
xor U8401 (N_8401,N_3011,N_3318);
nand U8402 (N_8402,N_3549,N_2792);
xor U8403 (N_8403,N_4549,N_1063);
xor U8404 (N_8404,N_4514,N_1622);
nor U8405 (N_8405,N_3634,N_704);
nand U8406 (N_8406,N_2290,N_262);
or U8407 (N_8407,N_4085,N_482);
nand U8408 (N_8408,N_3248,N_1066);
and U8409 (N_8409,N_950,N_3194);
nand U8410 (N_8410,N_4319,N_1964);
and U8411 (N_8411,N_4005,N_4066);
xor U8412 (N_8412,N_4985,N_3209);
and U8413 (N_8413,N_4590,N_3438);
and U8414 (N_8414,N_3413,N_1198);
nor U8415 (N_8415,N_3738,N_1373);
or U8416 (N_8416,N_1453,N_3767);
nand U8417 (N_8417,N_728,N_1692);
nor U8418 (N_8418,N_3106,N_2051);
or U8419 (N_8419,N_993,N_55);
xnor U8420 (N_8420,N_3998,N_3053);
nand U8421 (N_8421,N_3317,N_805);
nand U8422 (N_8422,N_1879,N_4750);
nand U8423 (N_8423,N_2136,N_913);
or U8424 (N_8424,N_2662,N_321);
or U8425 (N_8425,N_522,N_4276);
xor U8426 (N_8426,N_2155,N_411);
and U8427 (N_8427,N_3850,N_541);
or U8428 (N_8428,N_109,N_2373);
nand U8429 (N_8429,N_2602,N_591);
nand U8430 (N_8430,N_1641,N_2560);
nand U8431 (N_8431,N_2939,N_4416);
and U8432 (N_8432,N_3240,N_3969);
nor U8433 (N_8433,N_4211,N_2962);
nor U8434 (N_8434,N_3229,N_1897);
nand U8435 (N_8435,N_577,N_4728);
nor U8436 (N_8436,N_945,N_1204);
nor U8437 (N_8437,N_755,N_2370);
xnor U8438 (N_8438,N_1902,N_1248);
nand U8439 (N_8439,N_2707,N_2677);
or U8440 (N_8440,N_776,N_3325);
nor U8441 (N_8441,N_1443,N_2376);
and U8442 (N_8442,N_1921,N_1605);
or U8443 (N_8443,N_3035,N_3072);
xor U8444 (N_8444,N_3621,N_1722);
nand U8445 (N_8445,N_1342,N_3437);
nand U8446 (N_8446,N_1616,N_3932);
nor U8447 (N_8447,N_4552,N_1303);
nand U8448 (N_8448,N_993,N_3020);
nor U8449 (N_8449,N_3328,N_620);
nand U8450 (N_8450,N_1925,N_758);
nor U8451 (N_8451,N_4398,N_2365);
nor U8452 (N_8452,N_756,N_1453);
nand U8453 (N_8453,N_2081,N_4608);
and U8454 (N_8454,N_4938,N_4837);
xnor U8455 (N_8455,N_4040,N_3692);
or U8456 (N_8456,N_4368,N_1348);
or U8457 (N_8457,N_3023,N_4626);
and U8458 (N_8458,N_3220,N_4734);
xnor U8459 (N_8459,N_1204,N_4973);
or U8460 (N_8460,N_4754,N_4790);
nor U8461 (N_8461,N_1718,N_892);
nand U8462 (N_8462,N_1745,N_1070);
nand U8463 (N_8463,N_2035,N_2174);
or U8464 (N_8464,N_926,N_3490);
and U8465 (N_8465,N_2708,N_317);
nand U8466 (N_8466,N_3534,N_495);
nand U8467 (N_8467,N_279,N_2384);
or U8468 (N_8468,N_4263,N_435);
nor U8469 (N_8469,N_2302,N_4873);
or U8470 (N_8470,N_2267,N_2832);
nor U8471 (N_8471,N_2584,N_3880);
and U8472 (N_8472,N_2964,N_1243);
and U8473 (N_8473,N_3737,N_279);
nor U8474 (N_8474,N_2559,N_4091);
nand U8475 (N_8475,N_3916,N_3463);
xnor U8476 (N_8476,N_3884,N_164);
nand U8477 (N_8477,N_4057,N_1494);
nand U8478 (N_8478,N_1288,N_78);
or U8479 (N_8479,N_3088,N_1054);
nand U8480 (N_8480,N_3793,N_1972);
nor U8481 (N_8481,N_3436,N_3415);
xor U8482 (N_8482,N_1782,N_395);
nor U8483 (N_8483,N_4561,N_2250);
or U8484 (N_8484,N_300,N_2289);
nand U8485 (N_8485,N_656,N_3949);
nor U8486 (N_8486,N_271,N_2232);
nand U8487 (N_8487,N_4160,N_1744);
or U8488 (N_8488,N_1429,N_1396);
xnor U8489 (N_8489,N_3072,N_171);
and U8490 (N_8490,N_2713,N_363);
nand U8491 (N_8491,N_1088,N_4230);
and U8492 (N_8492,N_3181,N_191);
or U8493 (N_8493,N_423,N_4047);
xor U8494 (N_8494,N_4395,N_1025);
and U8495 (N_8495,N_4295,N_3020);
and U8496 (N_8496,N_3827,N_1609);
nor U8497 (N_8497,N_2526,N_902);
nand U8498 (N_8498,N_4647,N_1449);
or U8499 (N_8499,N_4668,N_447);
nor U8500 (N_8500,N_4826,N_2911);
or U8501 (N_8501,N_2901,N_4830);
nor U8502 (N_8502,N_2557,N_880);
nor U8503 (N_8503,N_618,N_2848);
xnor U8504 (N_8504,N_4709,N_797);
or U8505 (N_8505,N_909,N_2630);
nor U8506 (N_8506,N_70,N_3649);
xor U8507 (N_8507,N_1512,N_539);
or U8508 (N_8508,N_4975,N_2755);
nand U8509 (N_8509,N_3108,N_2797);
and U8510 (N_8510,N_3895,N_1575);
and U8511 (N_8511,N_130,N_3635);
xor U8512 (N_8512,N_4929,N_3903);
and U8513 (N_8513,N_918,N_3667);
nor U8514 (N_8514,N_3234,N_1790);
nand U8515 (N_8515,N_579,N_4836);
or U8516 (N_8516,N_4982,N_2029);
or U8517 (N_8517,N_524,N_4118);
nand U8518 (N_8518,N_2113,N_4719);
or U8519 (N_8519,N_4166,N_1102);
nor U8520 (N_8520,N_149,N_3545);
or U8521 (N_8521,N_3908,N_3909);
xor U8522 (N_8522,N_1117,N_4669);
or U8523 (N_8523,N_3906,N_1359);
nor U8524 (N_8524,N_2442,N_4869);
nand U8525 (N_8525,N_3688,N_3414);
or U8526 (N_8526,N_2461,N_3573);
or U8527 (N_8527,N_1298,N_1318);
or U8528 (N_8528,N_4413,N_2078);
nand U8529 (N_8529,N_529,N_2606);
xnor U8530 (N_8530,N_558,N_2009);
nand U8531 (N_8531,N_3630,N_945);
or U8532 (N_8532,N_2905,N_361);
and U8533 (N_8533,N_4446,N_3317);
or U8534 (N_8534,N_1005,N_880);
or U8535 (N_8535,N_4094,N_3292);
nor U8536 (N_8536,N_2654,N_3711);
or U8537 (N_8537,N_4049,N_4864);
nor U8538 (N_8538,N_3298,N_1842);
and U8539 (N_8539,N_3359,N_1310);
and U8540 (N_8540,N_795,N_4726);
nand U8541 (N_8541,N_2320,N_1766);
nand U8542 (N_8542,N_2926,N_220);
nor U8543 (N_8543,N_4866,N_4826);
nand U8544 (N_8544,N_766,N_3767);
nor U8545 (N_8545,N_499,N_686);
nor U8546 (N_8546,N_2614,N_802);
and U8547 (N_8547,N_184,N_3827);
nand U8548 (N_8548,N_3736,N_4275);
and U8549 (N_8549,N_4686,N_3896);
or U8550 (N_8550,N_1378,N_3283);
or U8551 (N_8551,N_412,N_3885);
nor U8552 (N_8552,N_2565,N_697);
or U8553 (N_8553,N_16,N_378);
nor U8554 (N_8554,N_2200,N_14);
and U8555 (N_8555,N_806,N_540);
or U8556 (N_8556,N_1333,N_526);
xor U8557 (N_8557,N_4608,N_2424);
or U8558 (N_8558,N_2135,N_2000);
nand U8559 (N_8559,N_321,N_2379);
and U8560 (N_8560,N_3968,N_2395);
nand U8561 (N_8561,N_534,N_4172);
nor U8562 (N_8562,N_3208,N_722);
nor U8563 (N_8563,N_1794,N_3154);
and U8564 (N_8564,N_4055,N_4814);
or U8565 (N_8565,N_791,N_3162);
nor U8566 (N_8566,N_3989,N_450);
nor U8567 (N_8567,N_2010,N_1765);
or U8568 (N_8568,N_102,N_1198);
or U8569 (N_8569,N_668,N_2493);
or U8570 (N_8570,N_2794,N_3812);
or U8571 (N_8571,N_899,N_4321);
nand U8572 (N_8572,N_2735,N_345);
and U8573 (N_8573,N_2608,N_2637);
nand U8574 (N_8574,N_4248,N_2799);
nor U8575 (N_8575,N_101,N_996);
and U8576 (N_8576,N_625,N_1114);
nor U8577 (N_8577,N_957,N_3705);
and U8578 (N_8578,N_3355,N_2107);
or U8579 (N_8579,N_3415,N_3797);
and U8580 (N_8580,N_3884,N_3217);
xnor U8581 (N_8581,N_266,N_1688);
nand U8582 (N_8582,N_2729,N_1537);
or U8583 (N_8583,N_486,N_2680);
nand U8584 (N_8584,N_3682,N_3519);
and U8585 (N_8585,N_1764,N_4079);
nand U8586 (N_8586,N_4644,N_3140);
or U8587 (N_8587,N_3083,N_1216);
nand U8588 (N_8588,N_4475,N_2834);
or U8589 (N_8589,N_255,N_440);
nand U8590 (N_8590,N_2816,N_4948);
or U8591 (N_8591,N_2534,N_590);
or U8592 (N_8592,N_3694,N_1261);
nor U8593 (N_8593,N_3616,N_615);
nand U8594 (N_8594,N_2112,N_1402);
or U8595 (N_8595,N_3828,N_2811);
and U8596 (N_8596,N_4800,N_3823);
nand U8597 (N_8597,N_354,N_3480);
nand U8598 (N_8598,N_3903,N_3954);
xor U8599 (N_8599,N_3797,N_711);
nand U8600 (N_8600,N_256,N_4851);
nand U8601 (N_8601,N_4902,N_657);
xnor U8602 (N_8602,N_1787,N_665);
nor U8603 (N_8603,N_3990,N_586);
xnor U8604 (N_8604,N_47,N_2157);
nand U8605 (N_8605,N_956,N_2808);
nand U8606 (N_8606,N_4586,N_4603);
and U8607 (N_8607,N_2440,N_1602);
and U8608 (N_8608,N_1253,N_3069);
xor U8609 (N_8609,N_1324,N_4904);
nand U8610 (N_8610,N_966,N_1947);
or U8611 (N_8611,N_987,N_4837);
or U8612 (N_8612,N_2657,N_1985);
nand U8613 (N_8613,N_1830,N_2165);
nand U8614 (N_8614,N_2651,N_373);
or U8615 (N_8615,N_4839,N_389);
and U8616 (N_8616,N_301,N_2092);
or U8617 (N_8617,N_797,N_1597);
and U8618 (N_8618,N_4285,N_1362);
or U8619 (N_8619,N_2858,N_304);
xnor U8620 (N_8620,N_2261,N_4112);
nand U8621 (N_8621,N_717,N_4818);
or U8622 (N_8622,N_4112,N_2162);
or U8623 (N_8623,N_3600,N_4391);
nor U8624 (N_8624,N_381,N_1986);
xor U8625 (N_8625,N_4011,N_342);
and U8626 (N_8626,N_460,N_101);
nor U8627 (N_8627,N_1464,N_3865);
nand U8628 (N_8628,N_4563,N_3860);
and U8629 (N_8629,N_4583,N_1378);
nand U8630 (N_8630,N_168,N_3172);
nor U8631 (N_8631,N_4207,N_3783);
nand U8632 (N_8632,N_159,N_4534);
nor U8633 (N_8633,N_896,N_1134);
nand U8634 (N_8634,N_3623,N_448);
nor U8635 (N_8635,N_827,N_1976);
nor U8636 (N_8636,N_2730,N_3439);
nand U8637 (N_8637,N_3866,N_2926);
nand U8638 (N_8638,N_2437,N_118);
and U8639 (N_8639,N_3418,N_4595);
nand U8640 (N_8640,N_4691,N_4608);
nand U8641 (N_8641,N_555,N_3177);
nand U8642 (N_8642,N_239,N_1680);
nor U8643 (N_8643,N_4932,N_2605);
xor U8644 (N_8644,N_2920,N_4771);
nor U8645 (N_8645,N_4417,N_2033);
or U8646 (N_8646,N_2339,N_4169);
or U8647 (N_8647,N_4741,N_3430);
and U8648 (N_8648,N_1754,N_4426);
nand U8649 (N_8649,N_2551,N_1433);
or U8650 (N_8650,N_4808,N_1015);
nand U8651 (N_8651,N_3774,N_2649);
and U8652 (N_8652,N_3129,N_1397);
or U8653 (N_8653,N_4294,N_2544);
or U8654 (N_8654,N_4805,N_1205);
nand U8655 (N_8655,N_353,N_4281);
or U8656 (N_8656,N_653,N_943);
and U8657 (N_8657,N_285,N_2013);
and U8658 (N_8658,N_4476,N_4396);
nand U8659 (N_8659,N_693,N_425);
or U8660 (N_8660,N_2856,N_4932);
nor U8661 (N_8661,N_2215,N_1831);
or U8662 (N_8662,N_853,N_3906);
nand U8663 (N_8663,N_649,N_2334);
and U8664 (N_8664,N_3896,N_1228);
or U8665 (N_8665,N_1718,N_3547);
and U8666 (N_8666,N_1408,N_3613);
and U8667 (N_8667,N_2822,N_3378);
nor U8668 (N_8668,N_2647,N_2891);
nand U8669 (N_8669,N_2407,N_2361);
nand U8670 (N_8670,N_146,N_1544);
and U8671 (N_8671,N_4193,N_3637);
xor U8672 (N_8672,N_1531,N_303);
and U8673 (N_8673,N_2206,N_2069);
xor U8674 (N_8674,N_4868,N_4025);
or U8675 (N_8675,N_3822,N_3610);
and U8676 (N_8676,N_2771,N_1683);
and U8677 (N_8677,N_101,N_2103);
and U8678 (N_8678,N_2546,N_1523);
and U8679 (N_8679,N_4635,N_307);
nor U8680 (N_8680,N_202,N_3070);
and U8681 (N_8681,N_2035,N_3996);
nand U8682 (N_8682,N_2413,N_889);
nor U8683 (N_8683,N_4463,N_3837);
nor U8684 (N_8684,N_2935,N_2640);
or U8685 (N_8685,N_3187,N_1128);
nor U8686 (N_8686,N_791,N_365);
and U8687 (N_8687,N_3177,N_2887);
nand U8688 (N_8688,N_62,N_2668);
and U8689 (N_8689,N_4920,N_1389);
nor U8690 (N_8690,N_4590,N_4505);
nor U8691 (N_8691,N_2727,N_3776);
and U8692 (N_8692,N_3849,N_3544);
nand U8693 (N_8693,N_1184,N_3489);
or U8694 (N_8694,N_3547,N_98);
nand U8695 (N_8695,N_329,N_1557);
or U8696 (N_8696,N_3171,N_27);
or U8697 (N_8697,N_1052,N_3910);
nand U8698 (N_8698,N_2963,N_4074);
nand U8699 (N_8699,N_1887,N_1586);
nor U8700 (N_8700,N_3798,N_1112);
nor U8701 (N_8701,N_3179,N_1980);
nand U8702 (N_8702,N_4078,N_211);
nor U8703 (N_8703,N_401,N_2885);
and U8704 (N_8704,N_3222,N_1597);
nor U8705 (N_8705,N_2957,N_1833);
or U8706 (N_8706,N_4763,N_3188);
xor U8707 (N_8707,N_4448,N_4713);
nand U8708 (N_8708,N_1324,N_118);
or U8709 (N_8709,N_3340,N_3180);
or U8710 (N_8710,N_2813,N_879);
nand U8711 (N_8711,N_2996,N_986);
nand U8712 (N_8712,N_3590,N_4689);
or U8713 (N_8713,N_1943,N_4060);
nand U8714 (N_8714,N_661,N_2103);
nor U8715 (N_8715,N_2929,N_3100);
nor U8716 (N_8716,N_4924,N_1757);
nand U8717 (N_8717,N_3363,N_2247);
nand U8718 (N_8718,N_1333,N_4305);
or U8719 (N_8719,N_436,N_2814);
nand U8720 (N_8720,N_2915,N_4924);
nor U8721 (N_8721,N_873,N_2538);
or U8722 (N_8722,N_888,N_1271);
nand U8723 (N_8723,N_4798,N_2804);
and U8724 (N_8724,N_2685,N_3131);
and U8725 (N_8725,N_4213,N_2771);
nand U8726 (N_8726,N_1000,N_377);
and U8727 (N_8727,N_370,N_4610);
or U8728 (N_8728,N_1615,N_303);
nor U8729 (N_8729,N_4987,N_4012);
nor U8730 (N_8730,N_28,N_939);
or U8731 (N_8731,N_2811,N_1179);
or U8732 (N_8732,N_1042,N_732);
and U8733 (N_8733,N_1868,N_2631);
and U8734 (N_8734,N_2257,N_1583);
nand U8735 (N_8735,N_4162,N_4203);
xor U8736 (N_8736,N_1095,N_1129);
and U8737 (N_8737,N_3236,N_4886);
nor U8738 (N_8738,N_1446,N_4931);
nand U8739 (N_8739,N_1933,N_2284);
nor U8740 (N_8740,N_1496,N_681);
or U8741 (N_8741,N_4399,N_4321);
nand U8742 (N_8742,N_3547,N_2131);
and U8743 (N_8743,N_3274,N_3338);
xnor U8744 (N_8744,N_377,N_3063);
and U8745 (N_8745,N_1158,N_1670);
nor U8746 (N_8746,N_1868,N_1375);
and U8747 (N_8747,N_4331,N_3513);
and U8748 (N_8748,N_2873,N_3918);
nor U8749 (N_8749,N_1856,N_2114);
nand U8750 (N_8750,N_3579,N_116);
nor U8751 (N_8751,N_2572,N_416);
nand U8752 (N_8752,N_2296,N_1916);
nor U8753 (N_8753,N_4073,N_3591);
xnor U8754 (N_8754,N_786,N_2254);
and U8755 (N_8755,N_4937,N_2093);
and U8756 (N_8756,N_739,N_906);
nand U8757 (N_8757,N_1003,N_2229);
or U8758 (N_8758,N_202,N_4061);
nor U8759 (N_8759,N_3023,N_3856);
and U8760 (N_8760,N_314,N_741);
or U8761 (N_8761,N_2390,N_798);
xnor U8762 (N_8762,N_2377,N_1713);
nand U8763 (N_8763,N_1660,N_817);
and U8764 (N_8764,N_2467,N_3217);
xor U8765 (N_8765,N_2058,N_527);
nand U8766 (N_8766,N_4578,N_2904);
nor U8767 (N_8767,N_2231,N_216);
nor U8768 (N_8768,N_39,N_986);
and U8769 (N_8769,N_4460,N_1402);
nor U8770 (N_8770,N_1198,N_3290);
nor U8771 (N_8771,N_1549,N_2492);
xnor U8772 (N_8772,N_554,N_1111);
xnor U8773 (N_8773,N_4093,N_1503);
nand U8774 (N_8774,N_2614,N_996);
xor U8775 (N_8775,N_2539,N_488);
xor U8776 (N_8776,N_1859,N_2689);
xnor U8777 (N_8777,N_4080,N_1305);
and U8778 (N_8778,N_4510,N_2629);
or U8779 (N_8779,N_3195,N_2372);
and U8780 (N_8780,N_4990,N_4276);
and U8781 (N_8781,N_2276,N_419);
nand U8782 (N_8782,N_3813,N_4140);
and U8783 (N_8783,N_4538,N_1690);
and U8784 (N_8784,N_4714,N_1910);
nand U8785 (N_8785,N_3976,N_1876);
xor U8786 (N_8786,N_2773,N_3771);
nand U8787 (N_8787,N_2568,N_2936);
and U8788 (N_8788,N_3167,N_3841);
nor U8789 (N_8789,N_3107,N_1147);
xnor U8790 (N_8790,N_3428,N_2432);
or U8791 (N_8791,N_214,N_3246);
nand U8792 (N_8792,N_404,N_3583);
or U8793 (N_8793,N_3386,N_622);
nor U8794 (N_8794,N_2891,N_3549);
nor U8795 (N_8795,N_539,N_407);
nor U8796 (N_8796,N_4046,N_1264);
or U8797 (N_8797,N_4971,N_4694);
nand U8798 (N_8798,N_2581,N_3188);
and U8799 (N_8799,N_1497,N_889);
xor U8800 (N_8800,N_3731,N_2633);
and U8801 (N_8801,N_4808,N_4735);
and U8802 (N_8802,N_3829,N_3955);
and U8803 (N_8803,N_1481,N_1176);
nand U8804 (N_8804,N_796,N_767);
and U8805 (N_8805,N_66,N_1693);
nand U8806 (N_8806,N_3256,N_3444);
and U8807 (N_8807,N_294,N_1116);
xnor U8808 (N_8808,N_1215,N_1751);
nand U8809 (N_8809,N_1660,N_805);
nor U8810 (N_8810,N_1985,N_1583);
nor U8811 (N_8811,N_3454,N_1515);
nand U8812 (N_8812,N_3749,N_233);
nand U8813 (N_8813,N_4086,N_3753);
and U8814 (N_8814,N_4405,N_3873);
and U8815 (N_8815,N_1733,N_1349);
and U8816 (N_8816,N_4297,N_4205);
or U8817 (N_8817,N_4212,N_4722);
and U8818 (N_8818,N_1868,N_3649);
nand U8819 (N_8819,N_3061,N_4665);
and U8820 (N_8820,N_2998,N_3232);
nor U8821 (N_8821,N_1662,N_1504);
nand U8822 (N_8822,N_983,N_2792);
nand U8823 (N_8823,N_4420,N_1738);
or U8824 (N_8824,N_3340,N_3668);
and U8825 (N_8825,N_62,N_4667);
or U8826 (N_8826,N_1264,N_1955);
or U8827 (N_8827,N_4277,N_4993);
nor U8828 (N_8828,N_1102,N_1071);
nor U8829 (N_8829,N_930,N_4145);
or U8830 (N_8830,N_1123,N_987);
or U8831 (N_8831,N_3440,N_3117);
nand U8832 (N_8832,N_2715,N_323);
and U8833 (N_8833,N_804,N_2864);
nand U8834 (N_8834,N_4317,N_2614);
xor U8835 (N_8835,N_4857,N_2178);
nor U8836 (N_8836,N_4338,N_4038);
and U8837 (N_8837,N_546,N_4536);
nand U8838 (N_8838,N_766,N_1624);
nor U8839 (N_8839,N_4458,N_1988);
or U8840 (N_8840,N_4782,N_94);
nor U8841 (N_8841,N_2729,N_870);
and U8842 (N_8842,N_318,N_33);
nand U8843 (N_8843,N_3040,N_4124);
nor U8844 (N_8844,N_255,N_2611);
or U8845 (N_8845,N_3163,N_2163);
nor U8846 (N_8846,N_459,N_4936);
nand U8847 (N_8847,N_3460,N_291);
nor U8848 (N_8848,N_1680,N_2230);
or U8849 (N_8849,N_792,N_381);
nand U8850 (N_8850,N_3539,N_2747);
nand U8851 (N_8851,N_401,N_4215);
and U8852 (N_8852,N_3415,N_1905);
nand U8853 (N_8853,N_1040,N_2862);
xnor U8854 (N_8854,N_464,N_244);
nand U8855 (N_8855,N_4722,N_2248);
nand U8856 (N_8856,N_2740,N_2520);
nand U8857 (N_8857,N_3829,N_963);
or U8858 (N_8858,N_783,N_4693);
and U8859 (N_8859,N_4714,N_941);
nand U8860 (N_8860,N_1417,N_4079);
or U8861 (N_8861,N_2068,N_1133);
or U8862 (N_8862,N_4626,N_3127);
xnor U8863 (N_8863,N_937,N_1236);
nor U8864 (N_8864,N_3320,N_4550);
nor U8865 (N_8865,N_150,N_549);
nand U8866 (N_8866,N_435,N_828);
nand U8867 (N_8867,N_420,N_1285);
xnor U8868 (N_8868,N_1309,N_1225);
and U8869 (N_8869,N_2806,N_595);
xnor U8870 (N_8870,N_3493,N_4854);
and U8871 (N_8871,N_4511,N_322);
or U8872 (N_8872,N_3222,N_1432);
and U8873 (N_8873,N_844,N_4447);
nand U8874 (N_8874,N_4940,N_438);
or U8875 (N_8875,N_1785,N_828);
or U8876 (N_8876,N_4946,N_1594);
nand U8877 (N_8877,N_4784,N_4785);
and U8878 (N_8878,N_1871,N_3475);
or U8879 (N_8879,N_4899,N_3383);
nor U8880 (N_8880,N_1310,N_783);
or U8881 (N_8881,N_3564,N_4871);
or U8882 (N_8882,N_926,N_1629);
xor U8883 (N_8883,N_4839,N_3668);
nand U8884 (N_8884,N_930,N_4230);
or U8885 (N_8885,N_3699,N_2816);
nor U8886 (N_8886,N_4503,N_2985);
nand U8887 (N_8887,N_428,N_4019);
and U8888 (N_8888,N_2045,N_4248);
nand U8889 (N_8889,N_3199,N_3183);
or U8890 (N_8890,N_126,N_271);
or U8891 (N_8891,N_1799,N_4426);
nand U8892 (N_8892,N_561,N_2870);
and U8893 (N_8893,N_513,N_42);
nand U8894 (N_8894,N_1163,N_4481);
nor U8895 (N_8895,N_3419,N_4814);
or U8896 (N_8896,N_763,N_2603);
nand U8897 (N_8897,N_1421,N_4017);
or U8898 (N_8898,N_4839,N_2794);
and U8899 (N_8899,N_897,N_145);
nand U8900 (N_8900,N_1826,N_137);
nand U8901 (N_8901,N_1204,N_4721);
and U8902 (N_8902,N_3533,N_4630);
and U8903 (N_8903,N_823,N_4554);
nand U8904 (N_8904,N_2318,N_2812);
or U8905 (N_8905,N_3343,N_671);
xnor U8906 (N_8906,N_543,N_4491);
nand U8907 (N_8907,N_4339,N_2533);
or U8908 (N_8908,N_1870,N_1061);
and U8909 (N_8909,N_1908,N_3105);
and U8910 (N_8910,N_515,N_1874);
or U8911 (N_8911,N_1973,N_592);
nand U8912 (N_8912,N_4206,N_2917);
nor U8913 (N_8913,N_3602,N_2580);
nand U8914 (N_8914,N_2963,N_4277);
or U8915 (N_8915,N_4519,N_228);
nand U8916 (N_8916,N_2620,N_1451);
and U8917 (N_8917,N_2588,N_3463);
xnor U8918 (N_8918,N_4571,N_3570);
nand U8919 (N_8919,N_2974,N_2828);
xnor U8920 (N_8920,N_2736,N_1916);
nand U8921 (N_8921,N_3595,N_2408);
or U8922 (N_8922,N_4089,N_2172);
nand U8923 (N_8923,N_3138,N_790);
and U8924 (N_8924,N_825,N_1886);
nor U8925 (N_8925,N_115,N_1859);
nor U8926 (N_8926,N_2234,N_2005);
nand U8927 (N_8927,N_4456,N_1429);
and U8928 (N_8928,N_4538,N_2786);
xnor U8929 (N_8929,N_887,N_2327);
or U8930 (N_8930,N_2829,N_1032);
xnor U8931 (N_8931,N_2187,N_4410);
nor U8932 (N_8932,N_2548,N_2210);
or U8933 (N_8933,N_1087,N_3753);
or U8934 (N_8934,N_4908,N_758);
and U8935 (N_8935,N_1727,N_3271);
nand U8936 (N_8936,N_3287,N_3413);
and U8937 (N_8937,N_3631,N_3241);
xor U8938 (N_8938,N_4539,N_3321);
nor U8939 (N_8939,N_2961,N_4488);
nor U8940 (N_8940,N_3555,N_3229);
nand U8941 (N_8941,N_512,N_1643);
and U8942 (N_8942,N_88,N_1386);
nor U8943 (N_8943,N_4248,N_3548);
or U8944 (N_8944,N_119,N_193);
nand U8945 (N_8945,N_876,N_2062);
xnor U8946 (N_8946,N_4681,N_1810);
nand U8947 (N_8947,N_3051,N_1492);
nand U8948 (N_8948,N_1140,N_4477);
or U8949 (N_8949,N_2570,N_4862);
or U8950 (N_8950,N_4109,N_3258);
and U8951 (N_8951,N_3772,N_2535);
nor U8952 (N_8952,N_1273,N_2593);
nor U8953 (N_8953,N_3331,N_3780);
nand U8954 (N_8954,N_2877,N_979);
nor U8955 (N_8955,N_1269,N_2220);
nor U8956 (N_8956,N_2694,N_337);
nand U8957 (N_8957,N_4315,N_4019);
xor U8958 (N_8958,N_4677,N_992);
nand U8959 (N_8959,N_1956,N_4649);
and U8960 (N_8960,N_2599,N_596);
nor U8961 (N_8961,N_1649,N_2840);
or U8962 (N_8962,N_421,N_3756);
nand U8963 (N_8963,N_1806,N_562);
nand U8964 (N_8964,N_3007,N_3334);
xnor U8965 (N_8965,N_2288,N_4038);
and U8966 (N_8966,N_1759,N_1395);
and U8967 (N_8967,N_4950,N_95);
xor U8968 (N_8968,N_1628,N_1092);
and U8969 (N_8969,N_1184,N_2904);
nand U8970 (N_8970,N_4402,N_118);
nor U8971 (N_8971,N_3923,N_3943);
or U8972 (N_8972,N_3667,N_4134);
nand U8973 (N_8973,N_507,N_2127);
nor U8974 (N_8974,N_3485,N_1055);
nor U8975 (N_8975,N_2835,N_4472);
nor U8976 (N_8976,N_316,N_2447);
nor U8977 (N_8977,N_4709,N_1120);
xor U8978 (N_8978,N_16,N_3306);
and U8979 (N_8979,N_4307,N_3355);
nand U8980 (N_8980,N_3680,N_1899);
or U8981 (N_8981,N_3370,N_2796);
nor U8982 (N_8982,N_3021,N_4925);
nand U8983 (N_8983,N_2178,N_3971);
nand U8984 (N_8984,N_3921,N_1950);
nor U8985 (N_8985,N_3492,N_4346);
nor U8986 (N_8986,N_184,N_1869);
and U8987 (N_8987,N_648,N_388);
and U8988 (N_8988,N_2786,N_1592);
or U8989 (N_8989,N_4322,N_2476);
nand U8990 (N_8990,N_342,N_2771);
nor U8991 (N_8991,N_3078,N_3812);
xnor U8992 (N_8992,N_4162,N_2681);
and U8993 (N_8993,N_1403,N_629);
and U8994 (N_8994,N_4860,N_4046);
nand U8995 (N_8995,N_137,N_3269);
nand U8996 (N_8996,N_1473,N_3165);
nor U8997 (N_8997,N_2270,N_82);
or U8998 (N_8998,N_3274,N_3635);
nand U8999 (N_8999,N_3503,N_497);
or U9000 (N_9000,N_2190,N_1473);
or U9001 (N_9001,N_3355,N_1961);
nor U9002 (N_9002,N_1158,N_4363);
nand U9003 (N_9003,N_4776,N_757);
nor U9004 (N_9004,N_3768,N_1322);
xor U9005 (N_9005,N_484,N_4288);
or U9006 (N_9006,N_3672,N_1229);
xnor U9007 (N_9007,N_3217,N_4836);
nor U9008 (N_9008,N_4159,N_3437);
nand U9009 (N_9009,N_968,N_4286);
nor U9010 (N_9010,N_4569,N_436);
nand U9011 (N_9011,N_821,N_928);
nand U9012 (N_9012,N_1113,N_1993);
nand U9013 (N_9013,N_3000,N_975);
nand U9014 (N_9014,N_3292,N_2068);
nand U9015 (N_9015,N_3574,N_1000);
nor U9016 (N_9016,N_3915,N_2595);
and U9017 (N_9017,N_3669,N_1147);
nor U9018 (N_9018,N_2463,N_335);
nand U9019 (N_9019,N_4691,N_706);
or U9020 (N_9020,N_3488,N_2078);
xor U9021 (N_9021,N_1250,N_1540);
nand U9022 (N_9022,N_3538,N_4712);
nand U9023 (N_9023,N_328,N_1415);
and U9024 (N_9024,N_246,N_2180);
nor U9025 (N_9025,N_155,N_4769);
nand U9026 (N_9026,N_4688,N_1489);
and U9027 (N_9027,N_3330,N_4989);
nor U9028 (N_9028,N_3416,N_998);
or U9029 (N_9029,N_345,N_2271);
nor U9030 (N_9030,N_147,N_2176);
and U9031 (N_9031,N_1712,N_1986);
or U9032 (N_9032,N_1239,N_3380);
nor U9033 (N_9033,N_4813,N_1954);
and U9034 (N_9034,N_2422,N_3004);
or U9035 (N_9035,N_3600,N_1528);
nand U9036 (N_9036,N_910,N_125);
or U9037 (N_9037,N_3152,N_3586);
nand U9038 (N_9038,N_1041,N_1537);
nor U9039 (N_9039,N_2461,N_3281);
nand U9040 (N_9040,N_4703,N_4949);
and U9041 (N_9041,N_1936,N_2321);
and U9042 (N_9042,N_4041,N_3927);
and U9043 (N_9043,N_4719,N_4863);
or U9044 (N_9044,N_1136,N_4161);
nor U9045 (N_9045,N_3610,N_2512);
or U9046 (N_9046,N_1636,N_24);
nor U9047 (N_9047,N_1623,N_2473);
nand U9048 (N_9048,N_878,N_4097);
or U9049 (N_9049,N_1325,N_1993);
nand U9050 (N_9050,N_957,N_1426);
or U9051 (N_9051,N_66,N_4683);
nand U9052 (N_9052,N_1425,N_2710);
or U9053 (N_9053,N_1941,N_949);
and U9054 (N_9054,N_410,N_3096);
and U9055 (N_9055,N_2675,N_1339);
nand U9056 (N_9056,N_2821,N_4556);
nand U9057 (N_9057,N_3627,N_4335);
and U9058 (N_9058,N_738,N_1821);
nor U9059 (N_9059,N_3932,N_3760);
xnor U9060 (N_9060,N_1010,N_1474);
or U9061 (N_9061,N_3613,N_4541);
or U9062 (N_9062,N_2542,N_3784);
xor U9063 (N_9063,N_3045,N_3663);
nor U9064 (N_9064,N_3869,N_290);
nand U9065 (N_9065,N_3068,N_4852);
and U9066 (N_9066,N_4217,N_2355);
nor U9067 (N_9067,N_4801,N_2035);
and U9068 (N_9068,N_3514,N_4448);
nand U9069 (N_9069,N_3954,N_1589);
or U9070 (N_9070,N_4702,N_2567);
xnor U9071 (N_9071,N_3259,N_2185);
xor U9072 (N_9072,N_4559,N_2315);
nor U9073 (N_9073,N_411,N_2698);
and U9074 (N_9074,N_192,N_2733);
nand U9075 (N_9075,N_1019,N_2610);
or U9076 (N_9076,N_4312,N_1553);
xnor U9077 (N_9077,N_2674,N_813);
nand U9078 (N_9078,N_441,N_1335);
nand U9079 (N_9079,N_3530,N_4482);
or U9080 (N_9080,N_3820,N_131);
nand U9081 (N_9081,N_3188,N_3382);
nor U9082 (N_9082,N_2132,N_4265);
xor U9083 (N_9083,N_3465,N_587);
or U9084 (N_9084,N_2414,N_4541);
nand U9085 (N_9085,N_637,N_2432);
or U9086 (N_9086,N_3582,N_1255);
or U9087 (N_9087,N_2621,N_1068);
nor U9088 (N_9088,N_87,N_3952);
and U9089 (N_9089,N_4440,N_1466);
and U9090 (N_9090,N_4108,N_1770);
nand U9091 (N_9091,N_2009,N_3278);
nand U9092 (N_9092,N_1273,N_683);
or U9093 (N_9093,N_3795,N_1996);
nor U9094 (N_9094,N_4669,N_2604);
or U9095 (N_9095,N_3627,N_1552);
nand U9096 (N_9096,N_712,N_1819);
and U9097 (N_9097,N_3880,N_4270);
or U9098 (N_9098,N_3614,N_1493);
nand U9099 (N_9099,N_3692,N_3778);
or U9100 (N_9100,N_3291,N_4896);
xor U9101 (N_9101,N_2766,N_1108);
and U9102 (N_9102,N_518,N_1359);
nor U9103 (N_9103,N_2574,N_3394);
nand U9104 (N_9104,N_2267,N_3498);
nor U9105 (N_9105,N_2794,N_2194);
nand U9106 (N_9106,N_2466,N_3503);
or U9107 (N_9107,N_917,N_2996);
nand U9108 (N_9108,N_1638,N_926);
and U9109 (N_9109,N_4536,N_3710);
or U9110 (N_9110,N_4011,N_4803);
or U9111 (N_9111,N_3332,N_4202);
and U9112 (N_9112,N_1646,N_26);
or U9113 (N_9113,N_929,N_2355);
nor U9114 (N_9114,N_537,N_2245);
or U9115 (N_9115,N_1363,N_4768);
or U9116 (N_9116,N_3220,N_4780);
xor U9117 (N_9117,N_831,N_2343);
and U9118 (N_9118,N_4269,N_1670);
and U9119 (N_9119,N_426,N_1389);
nor U9120 (N_9120,N_447,N_4843);
xor U9121 (N_9121,N_918,N_4344);
or U9122 (N_9122,N_4688,N_244);
or U9123 (N_9123,N_1413,N_2780);
nor U9124 (N_9124,N_1478,N_2075);
and U9125 (N_9125,N_428,N_4948);
nor U9126 (N_9126,N_3730,N_4506);
or U9127 (N_9127,N_1879,N_2806);
and U9128 (N_9128,N_3790,N_2249);
or U9129 (N_9129,N_2219,N_3186);
or U9130 (N_9130,N_2483,N_2327);
nor U9131 (N_9131,N_535,N_2565);
and U9132 (N_9132,N_1607,N_3251);
xnor U9133 (N_9133,N_2489,N_770);
xor U9134 (N_9134,N_2979,N_2669);
nand U9135 (N_9135,N_4861,N_2495);
nand U9136 (N_9136,N_2669,N_2076);
and U9137 (N_9137,N_739,N_2268);
and U9138 (N_9138,N_2649,N_720);
xor U9139 (N_9139,N_4716,N_2314);
or U9140 (N_9140,N_2654,N_4129);
or U9141 (N_9141,N_4274,N_4486);
or U9142 (N_9142,N_2690,N_974);
and U9143 (N_9143,N_403,N_3320);
xnor U9144 (N_9144,N_870,N_4250);
or U9145 (N_9145,N_600,N_1857);
xor U9146 (N_9146,N_3164,N_3805);
or U9147 (N_9147,N_2486,N_1739);
nor U9148 (N_9148,N_223,N_3641);
xor U9149 (N_9149,N_1386,N_1629);
and U9150 (N_9150,N_4935,N_2343);
xor U9151 (N_9151,N_4436,N_3156);
nor U9152 (N_9152,N_2006,N_3740);
and U9153 (N_9153,N_4712,N_517);
or U9154 (N_9154,N_4619,N_4407);
xnor U9155 (N_9155,N_727,N_3902);
nand U9156 (N_9156,N_1525,N_4693);
nor U9157 (N_9157,N_4355,N_2554);
nand U9158 (N_9158,N_457,N_3500);
and U9159 (N_9159,N_3439,N_2920);
or U9160 (N_9160,N_2153,N_4148);
or U9161 (N_9161,N_2979,N_2243);
or U9162 (N_9162,N_4719,N_2616);
or U9163 (N_9163,N_3870,N_2987);
nand U9164 (N_9164,N_4693,N_1103);
xnor U9165 (N_9165,N_4515,N_965);
nor U9166 (N_9166,N_2364,N_4181);
nand U9167 (N_9167,N_897,N_10);
or U9168 (N_9168,N_888,N_3835);
and U9169 (N_9169,N_2532,N_2143);
or U9170 (N_9170,N_841,N_743);
xnor U9171 (N_9171,N_105,N_4104);
and U9172 (N_9172,N_2301,N_2385);
nor U9173 (N_9173,N_1514,N_4842);
nand U9174 (N_9174,N_882,N_1658);
and U9175 (N_9175,N_897,N_682);
xnor U9176 (N_9176,N_2457,N_2065);
or U9177 (N_9177,N_197,N_2992);
and U9178 (N_9178,N_4119,N_4033);
and U9179 (N_9179,N_4362,N_3453);
or U9180 (N_9180,N_4398,N_3601);
or U9181 (N_9181,N_2204,N_1427);
or U9182 (N_9182,N_3281,N_3209);
nand U9183 (N_9183,N_2682,N_3554);
nand U9184 (N_9184,N_2795,N_4532);
or U9185 (N_9185,N_3121,N_3478);
xnor U9186 (N_9186,N_1851,N_4999);
or U9187 (N_9187,N_4569,N_3834);
and U9188 (N_9188,N_4138,N_2586);
nor U9189 (N_9189,N_2156,N_1760);
xnor U9190 (N_9190,N_1175,N_3092);
xnor U9191 (N_9191,N_2639,N_2820);
nand U9192 (N_9192,N_4179,N_2735);
nand U9193 (N_9193,N_2800,N_832);
and U9194 (N_9194,N_289,N_1220);
nand U9195 (N_9195,N_3062,N_2585);
xor U9196 (N_9196,N_2291,N_3795);
and U9197 (N_9197,N_124,N_2108);
and U9198 (N_9198,N_3891,N_1635);
and U9199 (N_9199,N_2597,N_4251);
and U9200 (N_9200,N_3230,N_2654);
and U9201 (N_9201,N_814,N_2798);
and U9202 (N_9202,N_1865,N_1179);
and U9203 (N_9203,N_631,N_3061);
and U9204 (N_9204,N_3635,N_3932);
nand U9205 (N_9205,N_4420,N_3979);
nor U9206 (N_9206,N_4063,N_2536);
nor U9207 (N_9207,N_4822,N_3212);
and U9208 (N_9208,N_1782,N_866);
nand U9209 (N_9209,N_3348,N_3781);
xor U9210 (N_9210,N_173,N_3210);
xor U9211 (N_9211,N_4396,N_2747);
or U9212 (N_9212,N_3648,N_3582);
and U9213 (N_9213,N_3016,N_1734);
or U9214 (N_9214,N_1395,N_4179);
nor U9215 (N_9215,N_1834,N_46);
nor U9216 (N_9216,N_3686,N_805);
nand U9217 (N_9217,N_655,N_2237);
nand U9218 (N_9218,N_397,N_4594);
nand U9219 (N_9219,N_3284,N_2420);
xnor U9220 (N_9220,N_4933,N_697);
or U9221 (N_9221,N_3764,N_1695);
xnor U9222 (N_9222,N_1765,N_1454);
or U9223 (N_9223,N_2524,N_812);
and U9224 (N_9224,N_891,N_1582);
and U9225 (N_9225,N_4167,N_4113);
or U9226 (N_9226,N_710,N_2758);
and U9227 (N_9227,N_3605,N_2808);
or U9228 (N_9228,N_2969,N_3339);
xor U9229 (N_9229,N_3797,N_4531);
and U9230 (N_9230,N_1470,N_1714);
and U9231 (N_9231,N_3994,N_4407);
or U9232 (N_9232,N_1123,N_2883);
nand U9233 (N_9233,N_1352,N_1946);
nor U9234 (N_9234,N_522,N_2372);
or U9235 (N_9235,N_3662,N_4678);
or U9236 (N_9236,N_1130,N_3741);
nand U9237 (N_9237,N_4792,N_4082);
nand U9238 (N_9238,N_395,N_3816);
nand U9239 (N_9239,N_4555,N_890);
and U9240 (N_9240,N_4454,N_4940);
nor U9241 (N_9241,N_4730,N_501);
and U9242 (N_9242,N_2213,N_1470);
nor U9243 (N_9243,N_2313,N_2031);
or U9244 (N_9244,N_591,N_837);
or U9245 (N_9245,N_1060,N_2845);
and U9246 (N_9246,N_4200,N_137);
nand U9247 (N_9247,N_3634,N_4355);
nand U9248 (N_9248,N_1859,N_3836);
xnor U9249 (N_9249,N_2651,N_2190);
and U9250 (N_9250,N_588,N_1099);
nor U9251 (N_9251,N_2117,N_571);
or U9252 (N_9252,N_3198,N_416);
xnor U9253 (N_9253,N_2443,N_3944);
nand U9254 (N_9254,N_3395,N_4461);
nor U9255 (N_9255,N_140,N_2756);
nand U9256 (N_9256,N_2161,N_84);
or U9257 (N_9257,N_4748,N_2931);
and U9258 (N_9258,N_2740,N_2824);
nand U9259 (N_9259,N_2217,N_4873);
nand U9260 (N_9260,N_2307,N_4426);
nor U9261 (N_9261,N_3741,N_1481);
xor U9262 (N_9262,N_1507,N_3306);
nand U9263 (N_9263,N_621,N_1081);
and U9264 (N_9264,N_3931,N_4395);
nand U9265 (N_9265,N_1984,N_199);
or U9266 (N_9266,N_3867,N_3815);
nor U9267 (N_9267,N_3417,N_968);
xor U9268 (N_9268,N_2845,N_4621);
nand U9269 (N_9269,N_3966,N_1682);
nand U9270 (N_9270,N_1513,N_1816);
and U9271 (N_9271,N_2696,N_492);
and U9272 (N_9272,N_4477,N_4297);
nand U9273 (N_9273,N_3486,N_220);
nand U9274 (N_9274,N_3535,N_3098);
nand U9275 (N_9275,N_4440,N_981);
and U9276 (N_9276,N_4669,N_1293);
nor U9277 (N_9277,N_2991,N_4911);
or U9278 (N_9278,N_4351,N_2111);
nor U9279 (N_9279,N_4235,N_1538);
nor U9280 (N_9280,N_4702,N_4914);
or U9281 (N_9281,N_4533,N_4377);
and U9282 (N_9282,N_4737,N_4055);
and U9283 (N_9283,N_2067,N_3626);
nand U9284 (N_9284,N_4164,N_4700);
or U9285 (N_9285,N_3413,N_4519);
or U9286 (N_9286,N_2357,N_1799);
nand U9287 (N_9287,N_2456,N_1401);
nand U9288 (N_9288,N_2424,N_1027);
and U9289 (N_9289,N_407,N_1600);
xnor U9290 (N_9290,N_3499,N_2295);
and U9291 (N_9291,N_3633,N_4600);
xor U9292 (N_9292,N_914,N_3212);
nand U9293 (N_9293,N_760,N_4747);
nand U9294 (N_9294,N_4783,N_2715);
xor U9295 (N_9295,N_691,N_2013);
nand U9296 (N_9296,N_2464,N_3524);
or U9297 (N_9297,N_4432,N_2405);
or U9298 (N_9298,N_3270,N_4081);
nor U9299 (N_9299,N_2159,N_426);
and U9300 (N_9300,N_1466,N_1069);
nand U9301 (N_9301,N_1837,N_3327);
xor U9302 (N_9302,N_3464,N_2747);
xor U9303 (N_9303,N_1058,N_2045);
nor U9304 (N_9304,N_1990,N_2355);
and U9305 (N_9305,N_4625,N_2822);
and U9306 (N_9306,N_3947,N_4571);
or U9307 (N_9307,N_3284,N_517);
xnor U9308 (N_9308,N_477,N_1289);
and U9309 (N_9309,N_3172,N_2421);
and U9310 (N_9310,N_4920,N_4377);
and U9311 (N_9311,N_66,N_370);
and U9312 (N_9312,N_395,N_2229);
and U9313 (N_9313,N_1816,N_1265);
nand U9314 (N_9314,N_4545,N_3112);
nand U9315 (N_9315,N_2898,N_2514);
nor U9316 (N_9316,N_4844,N_4873);
or U9317 (N_9317,N_2337,N_1420);
nand U9318 (N_9318,N_673,N_4958);
and U9319 (N_9319,N_2818,N_1639);
or U9320 (N_9320,N_4460,N_2548);
nor U9321 (N_9321,N_4193,N_2425);
nor U9322 (N_9322,N_3305,N_3105);
nand U9323 (N_9323,N_395,N_4032);
or U9324 (N_9324,N_3526,N_1848);
or U9325 (N_9325,N_505,N_3299);
or U9326 (N_9326,N_2301,N_261);
nor U9327 (N_9327,N_1142,N_1308);
and U9328 (N_9328,N_2709,N_1949);
nor U9329 (N_9329,N_190,N_1997);
xnor U9330 (N_9330,N_1062,N_3704);
and U9331 (N_9331,N_79,N_459);
or U9332 (N_9332,N_2158,N_3502);
and U9333 (N_9333,N_4060,N_2674);
xor U9334 (N_9334,N_4753,N_3391);
and U9335 (N_9335,N_1838,N_2797);
or U9336 (N_9336,N_1051,N_3585);
or U9337 (N_9337,N_806,N_2054);
and U9338 (N_9338,N_2617,N_1205);
or U9339 (N_9339,N_1330,N_424);
and U9340 (N_9340,N_2772,N_1055);
nand U9341 (N_9341,N_391,N_1920);
and U9342 (N_9342,N_3834,N_4952);
and U9343 (N_9343,N_2445,N_3060);
or U9344 (N_9344,N_1407,N_4259);
and U9345 (N_9345,N_4336,N_1585);
nor U9346 (N_9346,N_975,N_2188);
or U9347 (N_9347,N_735,N_813);
xor U9348 (N_9348,N_2391,N_3292);
nor U9349 (N_9349,N_4839,N_4005);
nor U9350 (N_9350,N_4899,N_3851);
nor U9351 (N_9351,N_1106,N_3615);
or U9352 (N_9352,N_3957,N_3708);
and U9353 (N_9353,N_1833,N_300);
or U9354 (N_9354,N_3119,N_4286);
xor U9355 (N_9355,N_850,N_3791);
xor U9356 (N_9356,N_2734,N_947);
and U9357 (N_9357,N_3808,N_1581);
or U9358 (N_9358,N_3746,N_3204);
nor U9359 (N_9359,N_1427,N_2783);
or U9360 (N_9360,N_3557,N_1014);
xor U9361 (N_9361,N_1390,N_443);
and U9362 (N_9362,N_1404,N_2799);
and U9363 (N_9363,N_1261,N_2308);
and U9364 (N_9364,N_4491,N_4652);
and U9365 (N_9365,N_3700,N_2792);
nor U9366 (N_9366,N_2656,N_2017);
nand U9367 (N_9367,N_2249,N_2362);
and U9368 (N_9368,N_195,N_4169);
nand U9369 (N_9369,N_2506,N_617);
nand U9370 (N_9370,N_2737,N_4880);
nor U9371 (N_9371,N_2170,N_2255);
nand U9372 (N_9372,N_2373,N_1861);
nor U9373 (N_9373,N_2822,N_1260);
or U9374 (N_9374,N_61,N_3222);
nand U9375 (N_9375,N_2769,N_2514);
nor U9376 (N_9376,N_3299,N_2880);
or U9377 (N_9377,N_3288,N_1974);
and U9378 (N_9378,N_4722,N_3559);
nor U9379 (N_9379,N_3361,N_4072);
nor U9380 (N_9380,N_2700,N_1161);
nand U9381 (N_9381,N_2953,N_1223);
and U9382 (N_9382,N_3810,N_3633);
and U9383 (N_9383,N_2202,N_433);
nand U9384 (N_9384,N_4812,N_734);
and U9385 (N_9385,N_3269,N_341);
and U9386 (N_9386,N_3291,N_1841);
and U9387 (N_9387,N_791,N_3305);
and U9388 (N_9388,N_1516,N_4568);
or U9389 (N_9389,N_963,N_3758);
nand U9390 (N_9390,N_3318,N_1665);
and U9391 (N_9391,N_3771,N_3111);
nand U9392 (N_9392,N_2884,N_3677);
nand U9393 (N_9393,N_1964,N_4998);
or U9394 (N_9394,N_417,N_2301);
nor U9395 (N_9395,N_70,N_3629);
or U9396 (N_9396,N_3110,N_4058);
and U9397 (N_9397,N_2187,N_364);
or U9398 (N_9398,N_4579,N_773);
nand U9399 (N_9399,N_1426,N_4529);
nand U9400 (N_9400,N_2764,N_1382);
or U9401 (N_9401,N_525,N_3316);
nor U9402 (N_9402,N_1744,N_1788);
and U9403 (N_9403,N_275,N_805);
xor U9404 (N_9404,N_468,N_69);
xnor U9405 (N_9405,N_717,N_3565);
nand U9406 (N_9406,N_2745,N_1422);
or U9407 (N_9407,N_2044,N_808);
xnor U9408 (N_9408,N_4073,N_4037);
nand U9409 (N_9409,N_3568,N_101);
nor U9410 (N_9410,N_4774,N_3772);
xnor U9411 (N_9411,N_2453,N_1648);
nor U9412 (N_9412,N_722,N_658);
nor U9413 (N_9413,N_2254,N_2015);
or U9414 (N_9414,N_1410,N_3704);
xnor U9415 (N_9415,N_2466,N_1858);
nand U9416 (N_9416,N_1050,N_3178);
nand U9417 (N_9417,N_4897,N_3948);
or U9418 (N_9418,N_3832,N_623);
and U9419 (N_9419,N_4945,N_4088);
and U9420 (N_9420,N_3603,N_2544);
xor U9421 (N_9421,N_29,N_2965);
and U9422 (N_9422,N_104,N_4430);
nand U9423 (N_9423,N_3303,N_20);
xnor U9424 (N_9424,N_3466,N_438);
and U9425 (N_9425,N_3045,N_1958);
nor U9426 (N_9426,N_3357,N_449);
or U9427 (N_9427,N_4540,N_3141);
nand U9428 (N_9428,N_2130,N_3209);
xnor U9429 (N_9429,N_1964,N_2255);
nand U9430 (N_9430,N_3084,N_94);
nor U9431 (N_9431,N_4655,N_550);
or U9432 (N_9432,N_3095,N_3804);
nand U9433 (N_9433,N_4715,N_2485);
and U9434 (N_9434,N_4152,N_3694);
nand U9435 (N_9435,N_2241,N_3198);
nand U9436 (N_9436,N_3497,N_3460);
nand U9437 (N_9437,N_925,N_1753);
and U9438 (N_9438,N_1515,N_3375);
or U9439 (N_9439,N_228,N_908);
or U9440 (N_9440,N_1592,N_4007);
nor U9441 (N_9441,N_3302,N_4505);
nand U9442 (N_9442,N_1650,N_2848);
or U9443 (N_9443,N_3557,N_832);
and U9444 (N_9444,N_3988,N_3888);
or U9445 (N_9445,N_4678,N_4243);
nor U9446 (N_9446,N_748,N_2359);
and U9447 (N_9447,N_4414,N_2894);
or U9448 (N_9448,N_749,N_4299);
nand U9449 (N_9449,N_2298,N_479);
and U9450 (N_9450,N_2826,N_1672);
or U9451 (N_9451,N_1270,N_1683);
nor U9452 (N_9452,N_2949,N_612);
nand U9453 (N_9453,N_3444,N_1690);
and U9454 (N_9454,N_715,N_3671);
nand U9455 (N_9455,N_347,N_1789);
nor U9456 (N_9456,N_1659,N_4963);
nand U9457 (N_9457,N_3407,N_3457);
and U9458 (N_9458,N_1433,N_3693);
or U9459 (N_9459,N_1611,N_1068);
nor U9460 (N_9460,N_2178,N_327);
nand U9461 (N_9461,N_3881,N_2194);
nand U9462 (N_9462,N_4437,N_2783);
nor U9463 (N_9463,N_4864,N_4598);
and U9464 (N_9464,N_3172,N_2043);
nor U9465 (N_9465,N_3906,N_1545);
nand U9466 (N_9466,N_175,N_1636);
nand U9467 (N_9467,N_476,N_3669);
nor U9468 (N_9468,N_651,N_725);
and U9469 (N_9469,N_543,N_3158);
nor U9470 (N_9470,N_163,N_4249);
nor U9471 (N_9471,N_947,N_1513);
nand U9472 (N_9472,N_4629,N_58);
or U9473 (N_9473,N_1262,N_4875);
nor U9474 (N_9474,N_3952,N_675);
or U9475 (N_9475,N_4711,N_2073);
or U9476 (N_9476,N_3561,N_1781);
and U9477 (N_9477,N_2898,N_4228);
and U9478 (N_9478,N_2369,N_2243);
nor U9479 (N_9479,N_1337,N_3230);
or U9480 (N_9480,N_2195,N_3489);
and U9481 (N_9481,N_319,N_1556);
nor U9482 (N_9482,N_1340,N_4639);
nor U9483 (N_9483,N_4565,N_1550);
and U9484 (N_9484,N_1307,N_3853);
nor U9485 (N_9485,N_698,N_4644);
and U9486 (N_9486,N_4922,N_2051);
nand U9487 (N_9487,N_4454,N_4515);
nor U9488 (N_9488,N_3369,N_3878);
xnor U9489 (N_9489,N_567,N_1543);
nand U9490 (N_9490,N_2481,N_2649);
nor U9491 (N_9491,N_147,N_2439);
nand U9492 (N_9492,N_121,N_1410);
and U9493 (N_9493,N_1770,N_748);
xor U9494 (N_9494,N_3071,N_1086);
nor U9495 (N_9495,N_669,N_1938);
nor U9496 (N_9496,N_4807,N_1904);
nor U9497 (N_9497,N_1171,N_570);
or U9498 (N_9498,N_4529,N_3189);
or U9499 (N_9499,N_4096,N_2107);
or U9500 (N_9500,N_322,N_4106);
nor U9501 (N_9501,N_1786,N_3743);
nor U9502 (N_9502,N_16,N_2371);
nand U9503 (N_9503,N_3232,N_4587);
and U9504 (N_9504,N_1522,N_3624);
nand U9505 (N_9505,N_2113,N_3179);
nand U9506 (N_9506,N_2268,N_3542);
nor U9507 (N_9507,N_4871,N_3203);
or U9508 (N_9508,N_4076,N_3442);
nor U9509 (N_9509,N_3855,N_598);
nor U9510 (N_9510,N_3195,N_2409);
or U9511 (N_9511,N_4234,N_3200);
and U9512 (N_9512,N_3089,N_4211);
nand U9513 (N_9513,N_666,N_939);
or U9514 (N_9514,N_4467,N_2303);
nand U9515 (N_9515,N_1151,N_4431);
or U9516 (N_9516,N_1120,N_3613);
nand U9517 (N_9517,N_1165,N_1116);
xor U9518 (N_9518,N_207,N_4329);
and U9519 (N_9519,N_1940,N_801);
nor U9520 (N_9520,N_4455,N_122);
or U9521 (N_9521,N_2666,N_3318);
nand U9522 (N_9522,N_3997,N_2332);
and U9523 (N_9523,N_3291,N_4695);
xnor U9524 (N_9524,N_653,N_1632);
nand U9525 (N_9525,N_4109,N_4695);
or U9526 (N_9526,N_4563,N_1613);
or U9527 (N_9527,N_4953,N_1770);
nor U9528 (N_9528,N_1133,N_1432);
nor U9529 (N_9529,N_846,N_762);
or U9530 (N_9530,N_2464,N_4528);
nor U9531 (N_9531,N_2320,N_4625);
nand U9532 (N_9532,N_4343,N_4719);
and U9533 (N_9533,N_2824,N_94);
and U9534 (N_9534,N_3259,N_3056);
nand U9535 (N_9535,N_3821,N_1854);
or U9536 (N_9536,N_3246,N_1217);
nand U9537 (N_9537,N_2244,N_2883);
or U9538 (N_9538,N_1649,N_2951);
and U9539 (N_9539,N_58,N_2013);
nor U9540 (N_9540,N_4629,N_3479);
or U9541 (N_9541,N_199,N_4261);
or U9542 (N_9542,N_4681,N_3696);
xnor U9543 (N_9543,N_4239,N_4957);
nor U9544 (N_9544,N_2262,N_3732);
and U9545 (N_9545,N_3407,N_2457);
or U9546 (N_9546,N_1219,N_520);
or U9547 (N_9547,N_4830,N_452);
and U9548 (N_9548,N_2424,N_4428);
or U9549 (N_9549,N_972,N_1280);
and U9550 (N_9550,N_286,N_2600);
and U9551 (N_9551,N_989,N_3263);
nor U9552 (N_9552,N_3526,N_2055);
and U9553 (N_9553,N_1036,N_4353);
nand U9554 (N_9554,N_3860,N_2971);
xnor U9555 (N_9555,N_4516,N_2620);
and U9556 (N_9556,N_295,N_407);
xor U9557 (N_9557,N_843,N_1813);
or U9558 (N_9558,N_1952,N_2794);
nand U9559 (N_9559,N_1300,N_3151);
nand U9560 (N_9560,N_4863,N_172);
nand U9561 (N_9561,N_178,N_1830);
nand U9562 (N_9562,N_4096,N_4994);
nor U9563 (N_9563,N_550,N_1095);
and U9564 (N_9564,N_624,N_1951);
and U9565 (N_9565,N_4857,N_1007);
and U9566 (N_9566,N_401,N_3333);
nor U9567 (N_9567,N_1843,N_691);
nand U9568 (N_9568,N_4183,N_780);
nor U9569 (N_9569,N_1565,N_3635);
nand U9570 (N_9570,N_4179,N_4183);
or U9571 (N_9571,N_760,N_435);
nor U9572 (N_9572,N_1827,N_2711);
nor U9573 (N_9573,N_1467,N_1443);
and U9574 (N_9574,N_2554,N_1911);
nor U9575 (N_9575,N_3460,N_4881);
nor U9576 (N_9576,N_3149,N_4520);
nand U9577 (N_9577,N_4844,N_3510);
nand U9578 (N_9578,N_3974,N_3080);
xor U9579 (N_9579,N_3355,N_3608);
or U9580 (N_9580,N_798,N_2061);
nor U9581 (N_9581,N_3668,N_808);
nor U9582 (N_9582,N_2944,N_2338);
xor U9583 (N_9583,N_4137,N_464);
or U9584 (N_9584,N_4139,N_3575);
xnor U9585 (N_9585,N_3883,N_2045);
or U9586 (N_9586,N_4834,N_4457);
nor U9587 (N_9587,N_1151,N_1996);
and U9588 (N_9588,N_4516,N_2509);
nor U9589 (N_9589,N_3085,N_4045);
and U9590 (N_9590,N_4382,N_4924);
nor U9591 (N_9591,N_2359,N_4400);
nor U9592 (N_9592,N_1597,N_3339);
nor U9593 (N_9593,N_4123,N_1669);
nand U9594 (N_9594,N_4141,N_2133);
nor U9595 (N_9595,N_3675,N_2544);
nand U9596 (N_9596,N_42,N_4455);
and U9597 (N_9597,N_2671,N_2104);
or U9598 (N_9598,N_2681,N_3919);
nor U9599 (N_9599,N_4245,N_1207);
nor U9600 (N_9600,N_3903,N_4410);
xnor U9601 (N_9601,N_2087,N_3591);
xor U9602 (N_9602,N_3257,N_342);
xor U9603 (N_9603,N_2345,N_1774);
nand U9604 (N_9604,N_3704,N_438);
nor U9605 (N_9605,N_4761,N_1360);
nor U9606 (N_9606,N_212,N_4812);
xor U9607 (N_9607,N_1916,N_1308);
nand U9608 (N_9608,N_4640,N_4936);
xor U9609 (N_9609,N_3475,N_1276);
nand U9610 (N_9610,N_2283,N_1230);
nor U9611 (N_9611,N_575,N_3617);
and U9612 (N_9612,N_299,N_887);
nand U9613 (N_9613,N_4422,N_1801);
and U9614 (N_9614,N_1404,N_2884);
or U9615 (N_9615,N_3983,N_4557);
nand U9616 (N_9616,N_4178,N_2);
nand U9617 (N_9617,N_755,N_1414);
xnor U9618 (N_9618,N_779,N_2483);
xor U9619 (N_9619,N_2982,N_3880);
nand U9620 (N_9620,N_1284,N_4901);
nand U9621 (N_9621,N_85,N_1835);
or U9622 (N_9622,N_4970,N_4603);
nor U9623 (N_9623,N_3642,N_4854);
and U9624 (N_9624,N_1280,N_4419);
xor U9625 (N_9625,N_4243,N_3174);
nor U9626 (N_9626,N_3875,N_4599);
nor U9627 (N_9627,N_2137,N_3557);
and U9628 (N_9628,N_3301,N_943);
and U9629 (N_9629,N_2214,N_2360);
and U9630 (N_9630,N_1488,N_4748);
or U9631 (N_9631,N_4465,N_452);
or U9632 (N_9632,N_198,N_4567);
and U9633 (N_9633,N_2200,N_1415);
or U9634 (N_9634,N_3971,N_1903);
and U9635 (N_9635,N_948,N_4117);
xor U9636 (N_9636,N_2799,N_1736);
nand U9637 (N_9637,N_2965,N_2408);
nand U9638 (N_9638,N_4968,N_3657);
nor U9639 (N_9639,N_4773,N_552);
nand U9640 (N_9640,N_1008,N_1237);
and U9641 (N_9641,N_894,N_1754);
nor U9642 (N_9642,N_1034,N_2505);
xor U9643 (N_9643,N_4436,N_4802);
or U9644 (N_9644,N_3902,N_4653);
xor U9645 (N_9645,N_2446,N_394);
or U9646 (N_9646,N_3822,N_991);
nor U9647 (N_9647,N_776,N_4538);
and U9648 (N_9648,N_545,N_1453);
or U9649 (N_9649,N_4659,N_2044);
nor U9650 (N_9650,N_3241,N_2076);
nand U9651 (N_9651,N_3587,N_609);
nand U9652 (N_9652,N_3201,N_3494);
or U9653 (N_9653,N_3317,N_3997);
and U9654 (N_9654,N_4887,N_4727);
nor U9655 (N_9655,N_506,N_1505);
and U9656 (N_9656,N_313,N_3969);
nor U9657 (N_9657,N_967,N_3974);
or U9658 (N_9658,N_4470,N_3534);
or U9659 (N_9659,N_1192,N_1585);
or U9660 (N_9660,N_4625,N_245);
and U9661 (N_9661,N_3959,N_1353);
nand U9662 (N_9662,N_961,N_3335);
nor U9663 (N_9663,N_2902,N_2887);
and U9664 (N_9664,N_1349,N_1958);
or U9665 (N_9665,N_4007,N_102);
nor U9666 (N_9666,N_3077,N_3361);
xor U9667 (N_9667,N_2722,N_2979);
or U9668 (N_9668,N_822,N_2182);
nor U9669 (N_9669,N_2411,N_4167);
or U9670 (N_9670,N_2869,N_8);
or U9671 (N_9671,N_3880,N_669);
nand U9672 (N_9672,N_3776,N_3625);
and U9673 (N_9673,N_323,N_3145);
or U9674 (N_9674,N_1222,N_58);
and U9675 (N_9675,N_1881,N_1964);
nand U9676 (N_9676,N_4811,N_2205);
nand U9677 (N_9677,N_3712,N_3398);
nor U9678 (N_9678,N_1015,N_4238);
and U9679 (N_9679,N_2913,N_2409);
and U9680 (N_9680,N_213,N_1850);
and U9681 (N_9681,N_2642,N_4453);
or U9682 (N_9682,N_4242,N_1564);
or U9683 (N_9683,N_3392,N_2274);
nand U9684 (N_9684,N_3951,N_1463);
and U9685 (N_9685,N_2134,N_4273);
nand U9686 (N_9686,N_2241,N_243);
nand U9687 (N_9687,N_3333,N_1316);
nand U9688 (N_9688,N_1238,N_3918);
and U9689 (N_9689,N_783,N_2715);
nand U9690 (N_9690,N_1712,N_2777);
nor U9691 (N_9691,N_3559,N_4230);
xor U9692 (N_9692,N_3106,N_331);
nor U9693 (N_9693,N_4332,N_2826);
or U9694 (N_9694,N_1677,N_4206);
nand U9695 (N_9695,N_2596,N_1778);
and U9696 (N_9696,N_963,N_2812);
or U9697 (N_9697,N_61,N_2555);
and U9698 (N_9698,N_1457,N_4739);
nor U9699 (N_9699,N_97,N_3385);
nand U9700 (N_9700,N_3577,N_220);
nand U9701 (N_9701,N_3362,N_3101);
nor U9702 (N_9702,N_4859,N_393);
nand U9703 (N_9703,N_1145,N_283);
nand U9704 (N_9704,N_3611,N_958);
or U9705 (N_9705,N_2423,N_1656);
nand U9706 (N_9706,N_170,N_338);
xnor U9707 (N_9707,N_4620,N_4965);
or U9708 (N_9708,N_4289,N_4084);
or U9709 (N_9709,N_4837,N_901);
nand U9710 (N_9710,N_4476,N_1012);
xnor U9711 (N_9711,N_2857,N_2376);
nor U9712 (N_9712,N_13,N_3506);
nor U9713 (N_9713,N_3546,N_199);
or U9714 (N_9714,N_3885,N_4294);
and U9715 (N_9715,N_389,N_59);
nor U9716 (N_9716,N_243,N_997);
or U9717 (N_9717,N_3170,N_1955);
xor U9718 (N_9718,N_2597,N_4137);
xnor U9719 (N_9719,N_992,N_807);
nor U9720 (N_9720,N_2263,N_924);
and U9721 (N_9721,N_3644,N_3774);
nand U9722 (N_9722,N_205,N_1676);
nand U9723 (N_9723,N_402,N_3330);
or U9724 (N_9724,N_3912,N_3246);
nor U9725 (N_9725,N_3118,N_4815);
nor U9726 (N_9726,N_604,N_2705);
xnor U9727 (N_9727,N_2219,N_4548);
xnor U9728 (N_9728,N_2598,N_4367);
nor U9729 (N_9729,N_2477,N_1552);
xor U9730 (N_9730,N_3606,N_3061);
nand U9731 (N_9731,N_2617,N_2573);
and U9732 (N_9732,N_3558,N_250);
or U9733 (N_9733,N_4065,N_1316);
nand U9734 (N_9734,N_4248,N_3204);
or U9735 (N_9735,N_4467,N_4176);
nand U9736 (N_9736,N_1358,N_2413);
or U9737 (N_9737,N_4222,N_2794);
nor U9738 (N_9738,N_4155,N_4938);
nand U9739 (N_9739,N_3015,N_3232);
and U9740 (N_9740,N_4024,N_2227);
nand U9741 (N_9741,N_2742,N_94);
nor U9742 (N_9742,N_4235,N_4806);
xor U9743 (N_9743,N_2501,N_35);
or U9744 (N_9744,N_3083,N_110);
or U9745 (N_9745,N_2427,N_3776);
xor U9746 (N_9746,N_182,N_174);
nor U9747 (N_9747,N_1037,N_2220);
nand U9748 (N_9748,N_2288,N_3686);
or U9749 (N_9749,N_3855,N_2510);
or U9750 (N_9750,N_2679,N_2558);
nor U9751 (N_9751,N_4226,N_210);
and U9752 (N_9752,N_3805,N_3890);
nor U9753 (N_9753,N_1413,N_1843);
nand U9754 (N_9754,N_2094,N_535);
nand U9755 (N_9755,N_2473,N_4391);
nor U9756 (N_9756,N_795,N_2260);
nor U9757 (N_9757,N_3583,N_420);
nand U9758 (N_9758,N_2697,N_4203);
and U9759 (N_9759,N_4129,N_3046);
or U9760 (N_9760,N_1987,N_4128);
and U9761 (N_9761,N_1504,N_3871);
nand U9762 (N_9762,N_2803,N_2999);
nand U9763 (N_9763,N_4716,N_119);
or U9764 (N_9764,N_2575,N_1821);
and U9765 (N_9765,N_382,N_1213);
and U9766 (N_9766,N_3061,N_590);
nor U9767 (N_9767,N_4164,N_2185);
or U9768 (N_9768,N_3181,N_4622);
nand U9769 (N_9769,N_4364,N_4695);
or U9770 (N_9770,N_4135,N_1675);
or U9771 (N_9771,N_3682,N_2309);
xnor U9772 (N_9772,N_1202,N_2559);
nor U9773 (N_9773,N_660,N_1334);
nor U9774 (N_9774,N_1944,N_2780);
nor U9775 (N_9775,N_4269,N_4992);
nand U9776 (N_9776,N_101,N_4706);
and U9777 (N_9777,N_2466,N_3929);
or U9778 (N_9778,N_1793,N_1886);
nand U9779 (N_9779,N_4614,N_1861);
xor U9780 (N_9780,N_2396,N_4012);
or U9781 (N_9781,N_1843,N_977);
or U9782 (N_9782,N_546,N_2877);
xor U9783 (N_9783,N_2594,N_4234);
and U9784 (N_9784,N_4548,N_3388);
xnor U9785 (N_9785,N_4691,N_2946);
nand U9786 (N_9786,N_3717,N_4072);
or U9787 (N_9787,N_2928,N_4275);
nand U9788 (N_9788,N_3059,N_3246);
xor U9789 (N_9789,N_754,N_2142);
nand U9790 (N_9790,N_2461,N_3279);
nor U9791 (N_9791,N_3268,N_59);
and U9792 (N_9792,N_4991,N_4519);
nand U9793 (N_9793,N_1907,N_4980);
or U9794 (N_9794,N_4637,N_161);
xor U9795 (N_9795,N_2699,N_1627);
or U9796 (N_9796,N_636,N_82);
xnor U9797 (N_9797,N_1707,N_68);
nor U9798 (N_9798,N_2864,N_2265);
and U9799 (N_9799,N_895,N_533);
or U9800 (N_9800,N_2099,N_998);
nor U9801 (N_9801,N_2723,N_1936);
and U9802 (N_9802,N_4294,N_4286);
xnor U9803 (N_9803,N_3077,N_1903);
or U9804 (N_9804,N_4256,N_1349);
nor U9805 (N_9805,N_4159,N_4847);
nand U9806 (N_9806,N_1250,N_3744);
or U9807 (N_9807,N_352,N_1525);
nand U9808 (N_9808,N_2384,N_3004);
nand U9809 (N_9809,N_4758,N_3993);
nor U9810 (N_9810,N_3796,N_3727);
nor U9811 (N_9811,N_4378,N_3189);
or U9812 (N_9812,N_3695,N_3775);
and U9813 (N_9813,N_1655,N_2353);
nor U9814 (N_9814,N_4652,N_2259);
and U9815 (N_9815,N_3294,N_3067);
and U9816 (N_9816,N_2023,N_1493);
and U9817 (N_9817,N_4803,N_2198);
nand U9818 (N_9818,N_4337,N_4996);
or U9819 (N_9819,N_326,N_718);
nand U9820 (N_9820,N_1292,N_1011);
or U9821 (N_9821,N_2764,N_1639);
and U9822 (N_9822,N_4813,N_1869);
nand U9823 (N_9823,N_2458,N_186);
nor U9824 (N_9824,N_2981,N_4671);
and U9825 (N_9825,N_1043,N_2837);
and U9826 (N_9826,N_336,N_2050);
and U9827 (N_9827,N_4944,N_3221);
or U9828 (N_9828,N_1604,N_3658);
nor U9829 (N_9829,N_3824,N_987);
or U9830 (N_9830,N_1662,N_585);
nor U9831 (N_9831,N_2886,N_4727);
xnor U9832 (N_9832,N_648,N_3392);
and U9833 (N_9833,N_3713,N_3993);
nand U9834 (N_9834,N_1130,N_4597);
xnor U9835 (N_9835,N_4805,N_4367);
nand U9836 (N_9836,N_3463,N_121);
xnor U9837 (N_9837,N_1919,N_453);
nand U9838 (N_9838,N_4427,N_4500);
or U9839 (N_9839,N_4914,N_1088);
nand U9840 (N_9840,N_101,N_2823);
and U9841 (N_9841,N_134,N_4097);
xnor U9842 (N_9842,N_4028,N_3129);
or U9843 (N_9843,N_2306,N_4460);
and U9844 (N_9844,N_106,N_2022);
nand U9845 (N_9845,N_4167,N_1055);
nor U9846 (N_9846,N_1364,N_1854);
nor U9847 (N_9847,N_1237,N_1848);
and U9848 (N_9848,N_2657,N_436);
or U9849 (N_9849,N_2657,N_2888);
nand U9850 (N_9850,N_3558,N_4133);
or U9851 (N_9851,N_2160,N_3706);
and U9852 (N_9852,N_316,N_2713);
or U9853 (N_9853,N_715,N_1734);
xnor U9854 (N_9854,N_3686,N_1625);
or U9855 (N_9855,N_2523,N_3593);
xnor U9856 (N_9856,N_971,N_1019);
nor U9857 (N_9857,N_3234,N_4654);
xor U9858 (N_9858,N_459,N_1607);
xnor U9859 (N_9859,N_1320,N_581);
nand U9860 (N_9860,N_1682,N_2682);
nand U9861 (N_9861,N_2473,N_4414);
nand U9862 (N_9862,N_3230,N_3763);
xnor U9863 (N_9863,N_1477,N_951);
nand U9864 (N_9864,N_1330,N_1045);
and U9865 (N_9865,N_789,N_4029);
or U9866 (N_9866,N_3756,N_4767);
or U9867 (N_9867,N_2950,N_1099);
nor U9868 (N_9868,N_1860,N_3936);
or U9869 (N_9869,N_1831,N_1590);
and U9870 (N_9870,N_1008,N_2280);
nand U9871 (N_9871,N_1268,N_2588);
or U9872 (N_9872,N_4624,N_1604);
xor U9873 (N_9873,N_3564,N_1414);
nor U9874 (N_9874,N_2933,N_3190);
and U9875 (N_9875,N_742,N_4530);
xnor U9876 (N_9876,N_1764,N_3447);
nor U9877 (N_9877,N_2322,N_4684);
xnor U9878 (N_9878,N_2595,N_4358);
or U9879 (N_9879,N_4062,N_3512);
nand U9880 (N_9880,N_224,N_4737);
or U9881 (N_9881,N_2376,N_4834);
nand U9882 (N_9882,N_215,N_450);
nor U9883 (N_9883,N_3351,N_995);
nor U9884 (N_9884,N_1436,N_1683);
and U9885 (N_9885,N_454,N_1451);
and U9886 (N_9886,N_335,N_1420);
nor U9887 (N_9887,N_2376,N_4393);
or U9888 (N_9888,N_2406,N_2793);
and U9889 (N_9889,N_3212,N_3526);
or U9890 (N_9890,N_310,N_4344);
nor U9891 (N_9891,N_3353,N_2422);
nand U9892 (N_9892,N_1170,N_3904);
nand U9893 (N_9893,N_1875,N_2730);
nor U9894 (N_9894,N_3124,N_2320);
or U9895 (N_9895,N_2768,N_3079);
nand U9896 (N_9896,N_265,N_3081);
nand U9897 (N_9897,N_4520,N_1201);
or U9898 (N_9898,N_2245,N_1336);
nand U9899 (N_9899,N_3043,N_259);
and U9900 (N_9900,N_2891,N_3497);
and U9901 (N_9901,N_4090,N_2593);
or U9902 (N_9902,N_79,N_3889);
and U9903 (N_9903,N_161,N_4651);
nor U9904 (N_9904,N_3059,N_363);
nand U9905 (N_9905,N_1978,N_2583);
nand U9906 (N_9906,N_1211,N_3788);
nand U9907 (N_9907,N_1059,N_2969);
nand U9908 (N_9908,N_2307,N_3470);
nor U9909 (N_9909,N_4069,N_4508);
and U9910 (N_9910,N_2656,N_2436);
xnor U9911 (N_9911,N_1022,N_1079);
nor U9912 (N_9912,N_1381,N_1494);
or U9913 (N_9913,N_4478,N_3460);
nand U9914 (N_9914,N_4873,N_2223);
and U9915 (N_9915,N_1648,N_510);
nor U9916 (N_9916,N_3547,N_1015);
and U9917 (N_9917,N_2851,N_2123);
nand U9918 (N_9918,N_1127,N_2927);
or U9919 (N_9919,N_1208,N_1182);
and U9920 (N_9920,N_397,N_600);
nand U9921 (N_9921,N_1337,N_1620);
nand U9922 (N_9922,N_1022,N_318);
or U9923 (N_9923,N_1994,N_80);
or U9924 (N_9924,N_4113,N_2386);
nand U9925 (N_9925,N_2457,N_2962);
nor U9926 (N_9926,N_1816,N_4993);
or U9927 (N_9927,N_3818,N_495);
nand U9928 (N_9928,N_2561,N_22);
or U9929 (N_9929,N_1088,N_1542);
and U9930 (N_9930,N_3916,N_4012);
nor U9931 (N_9931,N_67,N_268);
nor U9932 (N_9932,N_1277,N_534);
xor U9933 (N_9933,N_725,N_394);
and U9934 (N_9934,N_3633,N_2542);
nand U9935 (N_9935,N_752,N_941);
and U9936 (N_9936,N_4376,N_795);
and U9937 (N_9937,N_890,N_4820);
nor U9938 (N_9938,N_573,N_672);
nand U9939 (N_9939,N_2626,N_3044);
xor U9940 (N_9940,N_906,N_2332);
nor U9941 (N_9941,N_3977,N_2859);
or U9942 (N_9942,N_4486,N_437);
nand U9943 (N_9943,N_3710,N_1658);
nand U9944 (N_9944,N_3284,N_939);
nand U9945 (N_9945,N_4937,N_3245);
nor U9946 (N_9946,N_4778,N_416);
nand U9947 (N_9947,N_2588,N_2944);
nor U9948 (N_9948,N_1061,N_451);
or U9949 (N_9949,N_2880,N_2670);
xnor U9950 (N_9950,N_4112,N_4646);
nor U9951 (N_9951,N_215,N_2854);
nor U9952 (N_9952,N_3888,N_4452);
and U9953 (N_9953,N_966,N_3931);
nor U9954 (N_9954,N_3870,N_4184);
nand U9955 (N_9955,N_1619,N_2117);
or U9956 (N_9956,N_2352,N_2614);
and U9957 (N_9957,N_4743,N_1824);
and U9958 (N_9958,N_3207,N_2605);
xor U9959 (N_9959,N_1407,N_638);
and U9960 (N_9960,N_1851,N_2168);
and U9961 (N_9961,N_2693,N_1355);
nor U9962 (N_9962,N_4417,N_4193);
or U9963 (N_9963,N_4485,N_3324);
nand U9964 (N_9964,N_4013,N_64);
and U9965 (N_9965,N_3057,N_3028);
nor U9966 (N_9966,N_2312,N_2254);
nor U9967 (N_9967,N_2834,N_4609);
xnor U9968 (N_9968,N_3793,N_360);
and U9969 (N_9969,N_3773,N_3006);
nor U9970 (N_9970,N_3156,N_2179);
nor U9971 (N_9971,N_4944,N_2587);
and U9972 (N_9972,N_2332,N_4275);
nor U9973 (N_9973,N_680,N_798);
nor U9974 (N_9974,N_3456,N_2235);
nor U9975 (N_9975,N_1009,N_4941);
or U9976 (N_9976,N_3951,N_4260);
nor U9977 (N_9977,N_3490,N_4785);
nand U9978 (N_9978,N_4203,N_1007);
and U9979 (N_9979,N_2927,N_1839);
or U9980 (N_9980,N_4776,N_3947);
nor U9981 (N_9981,N_1057,N_1052);
and U9982 (N_9982,N_4659,N_4573);
and U9983 (N_9983,N_798,N_2018);
nor U9984 (N_9984,N_2060,N_3091);
nand U9985 (N_9985,N_2016,N_4780);
nor U9986 (N_9986,N_2126,N_1373);
xnor U9987 (N_9987,N_2970,N_1727);
or U9988 (N_9988,N_4889,N_1478);
or U9989 (N_9989,N_1462,N_1012);
nand U9990 (N_9990,N_2339,N_4736);
and U9991 (N_9991,N_1994,N_967);
xor U9992 (N_9992,N_4940,N_2628);
and U9993 (N_9993,N_4433,N_3288);
and U9994 (N_9994,N_2624,N_4038);
nand U9995 (N_9995,N_1731,N_772);
nand U9996 (N_9996,N_412,N_1152);
nor U9997 (N_9997,N_1906,N_2485);
nand U9998 (N_9998,N_3301,N_1383);
nor U9999 (N_9999,N_3603,N_3129);
or U10000 (N_10000,N_9535,N_8487);
nor U10001 (N_10001,N_6996,N_9124);
nand U10002 (N_10002,N_8670,N_6404);
nand U10003 (N_10003,N_8240,N_6283);
nand U10004 (N_10004,N_6538,N_8692);
nor U10005 (N_10005,N_7071,N_6450);
nand U10006 (N_10006,N_9242,N_6650);
nand U10007 (N_10007,N_6934,N_6354);
and U10008 (N_10008,N_7616,N_8470);
and U10009 (N_10009,N_6006,N_8511);
and U10010 (N_10010,N_8996,N_7620);
and U10011 (N_10011,N_6328,N_9008);
or U10012 (N_10012,N_9639,N_9072);
or U10013 (N_10013,N_5046,N_5634);
xor U10014 (N_10014,N_9963,N_5495);
xor U10015 (N_10015,N_9017,N_5534);
and U10016 (N_10016,N_9144,N_6360);
and U10017 (N_10017,N_6737,N_7497);
nand U10018 (N_10018,N_5474,N_8598);
and U10019 (N_10019,N_8795,N_8853);
or U10020 (N_10020,N_5759,N_5785);
or U10021 (N_10021,N_7574,N_9723);
and U10022 (N_10022,N_6466,N_8662);
or U10023 (N_10023,N_5226,N_6147);
or U10024 (N_10024,N_6408,N_7954);
and U10025 (N_10025,N_9633,N_6436);
or U10026 (N_10026,N_7807,N_6540);
xor U10027 (N_10027,N_8407,N_6107);
nor U10028 (N_10028,N_5960,N_7244);
xnor U10029 (N_10029,N_8351,N_5408);
nor U10030 (N_10030,N_9977,N_6595);
or U10031 (N_10031,N_6598,N_5137);
or U10032 (N_10032,N_6614,N_7710);
nor U10033 (N_10033,N_6253,N_8397);
or U10034 (N_10034,N_8141,N_7337);
xor U10035 (N_10035,N_7908,N_9239);
or U10036 (N_10036,N_5524,N_9672);
nand U10037 (N_10037,N_9437,N_5669);
nand U10038 (N_10038,N_6684,N_9048);
nor U10039 (N_10039,N_8816,N_7619);
nand U10040 (N_10040,N_7602,N_8556);
and U10041 (N_10041,N_6805,N_6723);
nand U10042 (N_10042,N_8786,N_6722);
and U10043 (N_10043,N_6263,N_6523);
nand U10044 (N_10044,N_7783,N_6639);
and U10045 (N_10045,N_7320,N_5754);
or U10046 (N_10046,N_8994,N_7522);
or U10047 (N_10047,N_9755,N_9809);
and U10048 (N_10048,N_6551,N_7315);
or U10049 (N_10049,N_5141,N_9818);
nor U10050 (N_10050,N_6447,N_7463);
or U10051 (N_10051,N_5951,N_7462);
xnor U10052 (N_10052,N_8384,N_9976);
nor U10053 (N_10053,N_8251,N_9935);
and U10054 (N_10054,N_9308,N_5172);
nor U10055 (N_10055,N_7998,N_8650);
nor U10056 (N_10056,N_6034,N_8291);
and U10057 (N_10057,N_8239,N_6882);
nand U10058 (N_10058,N_8716,N_6660);
and U10059 (N_10059,N_5442,N_9363);
nand U10060 (N_10060,N_9073,N_7832);
and U10061 (N_10061,N_7525,N_6988);
or U10062 (N_10062,N_8526,N_7495);
xnor U10063 (N_10063,N_5385,N_9270);
nor U10064 (N_10064,N_5610,N_8329);
nand U10065 (N_10065,N_8707,N_9855);
xor U10066 (N_10066,N_6385,N_6790);
and U10067 (N_10067,N_6745,N_6346);
or U10068 (N_10068,N_7514,N_8117);
nor U10069 (N_10069,N_5433,N_8159);
nand U10070 (N_10070,N_9047,N_5290);
and U10071 (N_10071,N_6195,N_8867);
xnor U10072 (N_10072,N_8602,N_9225);
xor U10073 (N_10073,N_6806,N_7855);
nor U10074 (N_10074,N_5393,N_5917);
and U10075 (N_10075,N_9329,N_9177);
nor U10076 (N_10076,N_5642,N_7909);
and U10077 (N_10077,N_7284,N_9952);
nor U10078 (N_10078,N_9813,N_9282);
xnor U10079 (N_10079,N_7453,N_5996);
nor U10080 (N_10080,N_6956,N_7851);
and U10081 (N_10081,N_7032,N_6871);
and U10082 (N_10082,N_7267,N_6089);
nor U10083 (N_10083,N_6141,N_6571);
and U10084 (N_10084,N_8821,N_8633);
and U10085 (N_10085,N_8922,N_5804);
nand U10086 (N_10086,N_9160,N_6331);
or U10087 (N_10087,N_8366,N_5438);
nor U10088 (N_10088,N_9769,N_9758);
nor U10089 (N_10089,N_6101,N_6087);
nand U10090 (N_10090,N_9369,N_6062);
or U10091 (N_10091,N_9076,N_6705);
nand U10092 (N_10092,N_8225,N_7650);
nor U10093 (N_10093,N_9942,N_9186);
nor U10094 (N_10094,N_5021,N_8903);
and U10095 (N_10095,N_8464,N_7962);
and U10096 (N_10096,N_9461,N_8262);
xnor U10097 (N_10097,N_7104,N_9792);
nor U10098 (N_10098,N_6116,N_9722);
nor U10099 (N_10099,N_9805,N_5125);
nand U10100 (N_10100,N_9812,N_9284);
nand U10101 (N_10101,N_5116,N_7377);
nand U10102 (N_10102,N_9417,N_6434);
or U10103 (N_10103,N_6130,N_5163);
and U10104 (N_10104,N_6809,N_7044);
or U10105 (N_10105,N_5915,N_5028);
and U10106 (N_10106,N_9362,N_5449);
nand U10107 (N_10107,N_7404,N_7075);
and U10108 (N_10108,N_9463,N_5631);
or U10109 (N_10109,N_5587,N_5364);
nand U10110 (N_10110,N_9014,N_6597);
nand U10111 (N_10111,N_7774,N_6319);
or U10112 (N_10112,N_6405,N_9286);
nor U10113 (N_10113,N_7705,N_9745);
nor U10114 (N_10114,N_8241,N_8886);
nor U10115 (N_10115,N_5373,N_7393);
nand U10116 (N_10116,N_7974,N_8899);
and U10117 (N_10117,N_8749,N_8451);
nor U10118 (N_10118,N_8669,N_6248);
or U10119 (N_10119,N_5292,N_9896);
nor U10120 (N_10120,N_8847,N_8720);
nand U10121 (N_10121,N_5686,N_7116);
and U10122 (N_10122,N_6740,N_8590);
nor U10123 (N_10123,N_7970,N_6202);
and U10124 (N_10124,N_9243,N_5151);
xor U10125 (N_10125,N_5242,N_8076);
or U10126 (N_10126,N_7333,N_9569);
or U10127 (N_10127,N_6798,N_8544);
nor U10128 (N_10128,N_9193,N_6841);
nand U10129 (N_10129,N_9836,N_9474);
or U10130 (N_10130,N_8188,N_5263);
nor U10131 (N_10131,N_6568,N_6171);
or U10132 (N_10132,N_7049,N_6341);
or U10133 (N_10133,N_7652,N_8691);
nor U10134 (N_10134,N_7670,N_9978);
and U10135 (N_10135,N_9589,N_8815);
nor U10136 (N_10136,N_5530,N_7613);
or U10137 (N_10137,N_9106,N_8110);
and U10138 (N_10138,N_9638,N_8017);
nor U10139 (N_10139,N_8713,N_6640);
nor U10140 (N_10140,N_8671,N_9222);
nor U10141 (N_10141,N_5112,N_9546);
xor U10142 (N_10142,N_8194,N_6449);
and U10143 (N_10143,N_9167,N_7510);
nor U10144 (N_10144,N_5856,N_9399);
nor U10145 (N_10145,N_6863,N_9786);
nand U10146 (N_10146,N_9148,N_8873);
xor U10147 (N_10147,N_7504,N_8489);
nand U10148 (N_10148,N_9534,N_8756);
nand U10149 (N_10149,N_8212,N_9772);
nand U10150 (N_10150,N_9069,N_5439);
or U10151 (N_10151,N_8521,N_5714);
nand U10152 (N_10152,N_7224,N_5051);
and U10153 (N_10153,N_5467,N_7070);
nand U10154 (N_10154,N_8626,N_7081);
or U10155 (N_10155,N_8991,N_5562);
nor U10156 (N_10156,N_6410,N_7371);
nor U10157 (N_10157,N_8325,N_7185);
and U10158 (N_10158,N_9176,N_8642);
nor U10159 (N_10159,N_8485,N_5415);
nor U10160 (N_10160,N_7667,N_9957);
xnor U10161 (N_10161,N_7438,N_5710);
nor U10162 (N_10162,N_5690,N_8610);
nand U10163 (N_10163,N_5480,N_9760);
or U10164 (N_10164,N_6463,N_8297);
xnor U10165 (N_10165,N_8981,N_8810);
nand U10166 (N_10166,N_7280,N_6300);
nand U10167 (N_10167,N_8379,N_7260);
nand U10168 (N_10168,N_7669,N_7999);
nor U10169 (N_10169,N_8805,N_5810);
nand U10170 (N_10170,N_7595,N_7300);
nand U10171 (N_10171,N_6743,N_7556);
nand U10172 (N_10172,N_7996,N_5875);
nor U10173 (N_10173,N_6496,N_8014);
or U10174 (N_10174,N_5428,N_9274);
nor U10175 (N_10175,N_9512,N_6681);
and U10176 (N_10176,N_8295,N_7328);
xnor U10177 (N_10177,N_7390,N_5411);
nand U10178 (N_10178,N_7584,N_9765);
nor U10179 (N_10179,N_7323,N_7858);
xor U10180 (N_10180,N_5831,N_7961);
nand U10181 (N_10181,N_6854,N_8580);
and U10182 (N_10182,N_8798,N_5413);
or U10183 (N_10183,N_5236,N_6898);
nor U10184 (N_10184,N_7831,N_8646);
or U10185 (N_10185,N_9783,N_9257);
and U10186 (N_10186,N_9366,N_6083);
and U10187 (N_10187,N_6995,N_5152);
xnor U10188 (N_10188,N_9502,N_9273);
nor U10189 (N_10189,N_9340,N_8841);
nor U10190 (N_10190,N_7155,N_5945);
and U10191 (N_10191,N_8656,N_8394);
or U10192 (N_10192,N_9246,N_6005);
nand U10193 (N_10193,N_5414,N_6622);
nand U10194 (N_10194,N_6528,N_5320);
or U10195 (N_10195,N_9892,N_6268);
and U10196 (N_10196,N_6509,N_6605);
and U10197 (N_10197,N_9307,N_6702);
nor U10198 (N_10198,N_6813,N_9599);
and U10199 (N_10199,N_7102,N_5515);
and U10200 (N_10200,N_6741,N_8595);
nand U10201 (N_10201,N_8863,N_7364);
xnor U10202 (N_10202,N_5463,N_9424);
and U10203 (N_10203,N_6292,N_9198);
and U10204 (N_10204,N_7158,N_7217);
nor U10205 (N_10205,N_5266,N_6656);
nor U10206 (N_10206,N_5384,N_6693);
nand U10207 (N_10207,N_8211,N_9305);
nor U10208 (N_10208,N_9192,N_6137);
nor U10209 (N_10209,N_5532,N_9622);
nor U10210 (N_10210,N_5342,N_8307);
nor U10211 (N_10211,N_9635,N_8686);
nor U10212 (N_10212,N_6356,N_8573);
nand U10213 (N_10213,N_9734,N_9318);
nor U10214 (N_10214,N_5916,N_8699);
and U10215 (N_10215,N_5312,N_5942);
or U10216 (N_10216,N_9782,N_8173);
or U10217 (N_10217,N_5221,N_5429);
and U10218 (N_10218,N_7615,N_6688);
and U10219 (N_10219,N_6288,N_9968);
nor U10220 (N_10220,N_5963,N_8750);
and U10221 (N_10221,N_5982,N_5579);
nand U10222 (N_10222,N_9372,N_6383);
nor U10223 (N_10223,N_7310,N_5258);
nor U10224 (N_10224,N_9597,N_5636);
nor U10225 (N_10225,N_8653,N_7451);
and U10226 (N_10226,N_9762,N_7901);
nor U10227 (N_10227,N_9398,N_5023);
nor U10228 (N_10228,N_8500,N_5874);
and U10229 (N_10229,N_8389,N_7589);
or U10230 (N_10230,N_9278,N_6920);
and U10231 (N_10231,N_6669,N_8907);
or U10232 (N_10232,N_9007,N_5217);
nand U10233 (N_10233,N_6054,N_5984);
nand U10234 (N_10234,N_5869,N_5732);
nand U10235 (N_10235,N_9841,N_5847);
nor U10236 (N_10236,N_8091,N_7985);
nor U10237 (N_10237,N_7922,N_7604);
or U10238 (N_10238,N_9481,N_5854);
nand U10239 (N_10239,N_5542,N_6227);
or U10240 (N_10240,N_9736,N_6550);
nor U10241 (N_10241,N_5735,N_8917);
xnor U10242 (N_10242,N_6767,N_7027);
and U10243 (N_10243,N_5435,N_6964);
nor U10244 (N_10244,N_8914,N_8119);
or U10245 (N_10245,N_7663,N_5593);
or U10246 (N_10246,N_6269,N_8254);
xor U10247 (N_10247,N_8049,N_8918);
or U10248 (N_10248,N_5314,N_7618);
and U10249 (N_10249,N_7289,N_6063);
or U10250 (N_10250,N_8261,N_8850);
and U10251 (N_10251,N_8731,N_7428);
or U10252 (N_10252,N_9970,N_9272);
or U10253 (N_10253,N_7129,N_6162);
and U10254 (N_10254,N_6224,N_6439);
nor U10255 (N_10255,N_9563,N_5144);
and U10256 (N_10256,N_8746,N_9334);
xor U10257 (N_10257,N_6877,N_8054);
or U10258 (N_10258,N_5693,N_6541);
nand U10259 (N_10259,N_5048,N_9729);
and U10260 (N_10260,N_9676,N_8469);
and U10261 (N_10261,N_5793,N_5424);
nor U10262 (N_10262,N_6843,N_5671);
or U10263 (N_10263,N_7416,N_8507);
nand U10264 (N_10264,N_5138,N_6186);
or U10265 (N_10265,N_7824,N_7009);
or U10266 (N_10266,N_5155,N_7761);
or U10267 (N_10267,N_5621,N_7542);
nor U10268 (N_10268,N_8024,N_5889);
nor U10269 (N_10269,N_9031,N_9728);
nor U10270 (N_10270,N_6233,N_6500);
nor U10271 (N_10271,N_8553,N_5126);
nand U10272 (N_10272,N_7162,N_6768);
nor U10273 (N_10273,N_9063,N_9617);
and U10274 (N_10274,N_8986,N_8101);
xor U10275 (N_10275,N_6714,N_8620);
and U10276 (N_10276,N_5904,N_7876);
and U10277 (N_10277,N_8979,N_9229);
or U10278 (N_10278,N_9907,N_9315);
or U10279 (N_10279,N_6475,N_9687);
nor U10280 (N_10280,N_7329,N_6651);
nand U10281 (N_10281,N_8066,N_7225);
and U10282 (N_10282,N_8475,N_5811);
nor U10283 (N_10283,N_7527,N_7380);
xnor U10284 (N_10284,N_5676,N_8523);
or U10285 (N_10285,N_8356,N_5601);
or U10286 (N_10286,N_6816,N_5719);
nand U10287 (N_10287,N_5822,N_9263);
nor U10288 (N_10288,N_7738,N_5727);
xnor U10289 (N_10289,N_9157,N_7771);
and U10290 (N_10290,N_8121,N_5997);
and U10291 (N_10291,N_8326,N_8210);
nor U10292 (N_10292,N_8622,N_7157);
nand U10293 (N_10293,N_9411,N_7294);
nor U10294 (N_10294,N_5476,N_6978);
and U10295 (N_10295,N_9804,N_5571);
or U10296 (N_10296,N_5279,N_5723);
nor U10297 (N_10297,N_6844,N_6867);
nand U10298 (N_10298,N_5131,N_8327);
or U10299 (N_10299,N_8369,N_9297);
or U10300 (N_10300,N_9798,N_6349);
nand U10301 (N_10301,N_9650,N_7696);
and U10302 (N_10302,N_9886,N_7817);
nand U10303 (N_10303,N_7742,N_8216);
or U10304 (N_10304,N_9560,N_7021);
nand U10305 (N_10305,N_8037,N_5655);
nand U10306 (N_10306,N_9109,N_5472);
or U10307 (N_10307,N_6774,N_6144);
nor U10308 (N_10308,N_5849,N_5733);
nand U10309 (N_10309,N_6869,N_7422);
or U10310 (N_10310,N_5128,N_5801);
nor U10311 (N_10311,N_5012,N_5936);
nor U10312 (N_10312,N_7821,N_8365);
or U10313 (N_10313,N_6044,N_6191);
or U10314 (N_10314,N_9238,N_6691);
and U10315 (N_10315,N_7064,N_7906);
nor U10316 (N_10316,N_9834,N_9483);
xor U10317 (N_10317,N_9686,N_5296);
or U10318 (N_10318,N_6909,N_6853);
nand U10319 (N_10319,N_5341,N_6378);
xnor U10320 (N_10320,N_5972,N_6462);
or U10321 (N_10321,N_5285,N_5444);
and U10322 (N_10322,N_5157,N_5086);
or U10323 (N_10323,N_5005,N_8231);
and U10324 (N_10324,N_8951,N_7701);
xor U10325 (N_10325,N_6223,N_5232);
or U10326 (N_10326,N_6336,N_6673);
nand U10327 (N_10327,N_6464,N_5335);
nand U10328 (N_10328,N_9982,N_7854);
or U10329 (N_10329,N_7773,N_8934);
or U10330 (N_10330,N_7234,N_6471);
or U10331 (N_10331,N_9613,N_7309);
or U10332 (N_10332,N_7077,N_9923);
nor U10333 (N_10333,N_6226,N_9390);
or U10334 (N_10334,N_6015,N_6317);
nand U10335 (N_10335,N_8882,N_7779);
nand U10336 (N_10336,N_8399,N_7391);
or U10337 (N_10337,N_8811,N_8198);
nand U10338 (N_10338,N_5955,N_5127);
nor U10339 (N_10339,N_9585,N_6197);
or U10340 (N_10340,N_6470,N_5797);
or U10341 (N_10341,N_6947,N_9895);
or U10342 (N_10342,N_7412,N_9394);
xor U10343 (N_10343,N_6819,N_7426);
nor U10344 (N_10344,N_9831,N_7699);
nor U10345 (N_10345,N_6583,N_6071);
or U10346 (N_10346,N_9423,N_9071);
xor U10347 (N_10347,N_8808,N_5036);
or U10348 (N_10348,N_5598,N_5886);
and U10349 (N_10349,N_7690,N_5700);
and U10350 (N_10350,N_8782,N_8519);
and U10351 (N_10351,N_6661,N_9256);
xnor U10352 (N_10352,N_5615,N_8911);
and U10353 (N_10353,N_7100,N_8709);
nor U10354 (N_10354,N_9756,N_8904);
nor U10355 (N_10355,N_5452,N_5612);
nand U10356 (N_10356,N_9688,N_5469);
nor U10357 (N_10357,N_8495,N_8280);
xor U10358 (N_10358,N_7760,N_7111);
or U10359 (N_10359,N_6393,N_7512);
and U10360 (N_10360,N_8547,N_8134);
xor U10361 (N_10361,N_9467,N_6807);
or U10362 (N_10362,N_6779,N_5145);
nand U10363 (N_10363,N_5677,N_5164);
nand U10364 (N_10364,N_6310,N_6706);
nor U10365 (N_10365,N_8617,N_5349);
nand U10366 (N_10366,N_7809,N_8276);
nand U10367 (N_10367,N_7836,N_7033);
or U10368 (N_10368,N_7557,N_8813);
nor U10369 (N_10369,N_8288,N_6563);
xor U10370 (N_10370,N_8830,N_9517);
xor U10371 (N_10371,N_8582,N_5441);
nand U10372 (N_10372,N_6753,N_5479);
or U10373 (N_10373,N_5362,N_9086);
nand U10374 (N_10374,N_9924,N_6746);
or U10375 (N_10375,N_9010,N_5839);
nor U10376 (N_10376,N_7857,N_9494);
nand U10377 (N_10377,N_5715,N_9727);
or U10378 (N_10378,N_6339,N_9107);
or U10379 (N_10379,N_8565,N_7754);
xor U10380 (N_10380,N_9887,N_7379);
nand U10381 (N_10381,N_8828,N_5771);
and U10382 (N_10382,N_8203,N_8467);
and U10383 (N_10383,N_7258,N_7538);
nor U10384 (N_10384,N_9861,N_5999);
nand U10385 (N_10385,N_8688,N_5691);
nor U10386 (N_10386,N_6106,N_9099);
nand U10387 (N_10387,N_5460,N_6763);
nand U10388 (N_10388,N_8406,N_5873);
or U10389 (N_10389,N_9021,N_6771);
nor U10390 (N_10390,N_5037,N_5319);
and U10391 (N_10391,N_6537,N_8310);
nand U10392 (N_10392,N_7312,N_9678);
or U10393 (N_10393,N_7537,N_7934);
nand U10394 (N_10394,N_6432,N_9004);
nand U10395 (N_10395,N_8160,N_9025);
nor U10396 (N_10396,N_9104,N_5506);
and U10397 (N_10397,N_9506,N_9095);
nand U10398 (N_10398,N_8456,N_9060);
or U10399 (N_10399,N_7656,N_8800);
xor U10400 (N_10400,N_6874,N_5851);
or U10401 (N_10401,N_9379,N_6053);
nor U10402 (N_10402,N_7240,N_9605);
or U10403 (N_10403,N_7108,N_9511);
nand U10404 (N_10404,N_5981,N_9466);
or U10405 (N_10405,N_5248,N_5775);
or U10406 (N_10406,N_6736,N_9888);
and U10407 (N_10407,N_9715,N_9878);
nor U10408 (N_10408,N_7283,N_9002);
nand U10409 (N_10409,N_6367,N_7725);
nand U10410 (N_10410,N_9735,N_6321);
nand U10411 (N_10411,N_6007,N_9930);
and U10412 (N_10412,N_9959,N_7372);
and U10413 (N_10413,N_6517,N_8877);
nand U10414 (N_10414,N_8158,N_8906);
nand U10415 (N_10415,N_6648,N_8170);
and U10416 (N_10416,N_9139,N_5074);
nor U10417 (N_10417,N_9138,N_5153);
and U10418 (N_10418,N_6817,N_5979);
nand U10419 (N_10419,N_9279,N_6014);
or U10420 (N_10420,N_7113,N_5149);
xor U10421 (N_10421,N_5751,N_8884);
nor U10422 (N_10422,N_7849,N_6369);
and U10423 (N_10423,N_5203,N_9983);
and U10424 (N_10424,N_9022,N_9870);
nand U10425 (N_10425,N_6050,N_7219);
or U10426 (N_10426,N_8010,N_8417);
nand U10427 (N_10427,N_8734,N_5573);
and U10428 (N_10428,N_5956,N_8084);
nand U10429 (N_10429,N_8772,N_6780);
nor U10430 (N_10430,N_8320,N_8107);
nor U10431 (N_10431,N_7061,N_8197);
xnor U10432 (N_10432,N_8775,N_9460);
and U10433 (N_10433,N_9480,N_9752);
nor U10434 (N_10434,N_6849,N_6951);
nand U10435 (N_10435,N_6894,N_7264);
and U10436 (N_10436,N_5055,N_5702);
and U10437 (N_10437,N_7282,N_8287);
or U10438 (N_10438,N_7846,N_9524);
and U10439 (N_10439,N_9995,N_8442);
nor U10440 (N_10440,N_8564,N_8583);
and U10441 (N_10441,N_6564,N_7782);
xor U10442 (N_10442,N_9355,N_5599);
nor U10443 (N_10443,N_7415,N_5905);
nor U10444 (N_10444,N_5918,N_9941);
and U10445 (N_10445,N_6976,N_8094);
nor U10446 (N_10446,N_8232,N_9053);
or U10447 (N_10447,N_6121,N_9425);
or U10448 (N_10448,N_8074,N_7532);
or U10449 (N_10449,N_7753,N_7420);
or U10450 (N_10450,N_5376,N_8586);
and U10451 (N_10451,N_5744,N_7327);
nor U10452 (N_10452,N_7570,N_8001);
nand U10453 (N_10453,N_7878,N_5070);
or U10454 (N_10454,N_8997,N_9578);
and U10455 (N_10455,N_7127,N_9570);
nand U10456 (N_10456,N_7356,N_6052);
or U10457 (N_10457,N_8779,N_7603);
nand U10458 (N_10458,N_8787,N_6018);
nand U10459 (N_10459,N_7401,N_6670);
or U10460 (N_10460,N_7900,N_7581);
nand U10461 (N_10461,N_7866,N_5208);
nor U10462 (N_10462,N_7547,N_5019);
nor U10463 (N_10463,N_7548,N_6212);
nand U10464 (N_10464,N_8560,N_9051);
nor U10465 (N_10465,N_6739,N_9026);
nand U10466 (N_10466,N_8948,N_6940);
nor U10467 (N_10467,N_9544,N_5846);
and U10468 (N_10468,N_6299,N_7124);
nand U10469 (N_10469,N_5786,N_9264);
or U10470 (N_10470,N_5344,N_7055);
and U10471 (N_10471,N_7718,N_5422);
nand U10472 (N_10472,N_6151,N_6388);
nand U10473 (N_10473,N_5239,N_9190);
nor U10474 (N_10474,N_7659,N_6896);
nand U10475 (N_10475,N_5018,N_8625);
nand U10476 (N_10476,N_5196,N_5374);
xor U10477 (N_10477,N_6266,N_8140);
nor U10478 (N_10478,N_9259,N_9169);
nor U10479 (N_10479,N_7160,N_7069);
nor U10480 (N_10480,N_8100,N_7918);
or U10481 (N_10481,N_9434,N_9636);
xnor U10482 (N_10482,N_9822,N_9491);
and U10483 (N_10483,N_8163,N_5641);
nand U10484 (N_10484,N_5106,N_8898);
nand U10485 (N_10485,N_9652,N_7957);
nand U10486 (N_10486,N_6423,N_5082);
or U10487 (N_10487,N_7795,N_7191);
nand U10488 (N_10488,N_7423,N_5400);
or U10489 (N_10489,N_7091,N_7638);
or U10490 (N_10490,N_7879,N_5377);
nand U10491 (N_10491,N_8661,N_5567);
nor U10492 (N_10492,N_6267,N_8226);
or U10493 (N_10493,N_9405,N_6036);
or U10494 (N_10494,N_7230,N_9960);
xnor U10495 (N_10495,N_5517,N_5174);
nand U10496 (N_10496,N_7881,N_6396);
nand U10497 (N_10497,N_5678,N_8176);
and U10498 (N_10498,N_6984,N_6347);
or U10499 (N_10499,N_7730,N_5586);
nand U10500 (N_10500,N_7509,N_7344);
nor U10501 (N_10501,N_9777,N_7727);
nand U10502 (N_10502,N_9821,N_5866);
nor U10503 (N_10503,N_8569,N_8184);
nand U10504 (N_10504,N_7079,N_9328);
nand U10505 (N_10505,N_7822,N_7402);
nor U10506 (N_10506,N_7458,N_6971);
nand U10507 (N_10507,N_8488,N_9179);
or U10508 (N_10508,N_9174,N_6389);
and U10509 (N_10509,N_5765,N_7776);
nor U10510 (N_10510,N_7014,N_5156);
or U10511 (N_10511,N_9431,N_9972);
xor U10512 (N_10512,N_6842,N_5205);
nand U10513 (N_10513,N_7357,N_9630);
nand U10514 (N_10514,N_8436,N_7790);
xor U10515 (N_10515,N_9248,N_5329);
or U10516 (N_10516,N_9839,N_9219);
nand U10517 (N_10517,N_5522,N_8302);
nor U10518 (N_10518,N_7456,N_6770);
and U10519 (N_10519,N_5766,N_6507);
and U10520 (N_10520,N_5398,N_7942);
or U10521 (N_10521,N_7814,N_9943);
and U10522 (N_10522,N_9247,N_7500);
nor U10523 (N_10523,N_9317,N_6987);
nor U10524 (N_10524,N_5520,N_8415);
xor U10525 (N_10525,N_7259,N_7958);
and U10526 (N_10526,N_8529,N_8153);
nor U10527 (N_10527,N_6038,N_7653);
and U10528 (N_10528,N_7484,N_8777);
nor U10529 (N_10529,N_6980,N_6282);
and U10530 (N_10530,N_8640,N_9851);
or U10531 (N_10531,N_9620,N_6552);
xnor U10532 (N_10532,N_8073,N_6272);
nand U10533 (N_10533,N_9367,N_8584);
nor U10534 (N_10534,N_8512,N_9649);
and U10535 (N_10535,N_9429,N_8978);
and U10536 (N_10536,N_6917,N_8304);
or U10537 (N_10537,N_6277,N_5173);
or U10538 (N_10538,N_5574,N_6683);
nand U10539 (N_10539,N_6658,N_7980);
or U10540 (N_10540,N_7012,N_5122);
nand U10541 (N_10541,N_9513,N_5421);
nand U10542 (N_10542,N_6031,N_5338);
nand U10543 (N_10543,N_6295,N_7048);
and U10544 (N_10544,N_9486,N_7593);
xnor U10545 (N_10545,N_6060,N_7916);
and U10546 (N_10546,N_5741,N_8860);
and U10547 (N_10547,N_8908,N_7915);
and U10548 (N_10548,N_7103,N_7599);
or U10549 (N_10549,N_8732,N_6484);
xor U10550 (N_10550,N_6324,N_7350);
nand U10551 (N_10551,N_5355,N_8059);
nand U10552 (N_10552,N_7627,N_7549);
xnor U10553 (N_10553,N_7982,N_5670);
and U10554 (N_10554,N_6792,N_7200);
nor U10555 (N_10555,N_7744,N_8657);
or U10556 (N_10556,N_6264,N_7206);
nand U10557 (N_10557,N_5666,N_6219);
and U10558 (N_10558,N_8545,N_5454);
and U10559 (N_10559,N_8318,N_6503);
nand U10560 (N_10560,N_8090,N_5576);
nor U10561 (N_10561,N_5406,N_5526);
nor U10562 (N_10562,N_9226,N_8829);
nor U10563 (N_10563,N_5059,N_9303);
nor U10564 (N_10564,N_7955,N_9114);
or U10565 (N_10565,N_8289,N_7953);
or U10566 (N_10566,N_7023,N_8892);
xnor U10567 (N_10567,N_9890,N_8422);
or U10568 (N_10568,N_8315,N_6677);
xnor U10569 (N_10569,N_8792,N_8615);
and U10570 (N_10570,N_5729,N_5638);
or U10571 (N_10571,N_5013,N_6667);
nor U10572 (N_10572,N_5124,N_6865);
or U10573 (N_10573,N_5644,N_5381);
and U10574 (N_10574,N_8537,N_9116);
and U10575 (N_10575,N_7554,N_7439);
or U10576 (N_10576,N_8483,N_6124);
nor U10577 (N_10577,N_8002,N_9852);
nor U10578 (N_10578,N_6961,N_7037);
xor U10579 (N_10579,N_7662,N_7810);
and U10580 (N_10580,N_7898,N_5931);
and U10581 (N_10581,N_5633,N_6533);
nor U10582 (N_10582,N_5011,N_5519);
or U10583 (N_10583,N_8046,N_6316);
xnor U10584 (N_10584,N_9515,N_5078);
nand U10585 (N_10585,N_8614,N_6919);
nor U10586 (N_10586,N_8207,N_8865);
and U10587 (N_10587,N_5412,N_9146);
or U10588 (N_10588,N_8826,N_6453);
and U10589 (N_10589,N_9862,N_8683);
nor U10590 (N_10590,N_8592,N_7746);
nand U10591 (N_10591,N_8740,N_5301);
or U10592 (N_10592,N_9265,N_6883);
and U10593 (N_10593,N_6353,N_6590);
and U10594 (N_10594,N_6315,N_6111);
nand U10595 (N_10595,N_9564,N_8803);
xnor U10596 (N_10596,N_6625,N_9224);
or U10597 (N_10597,N_7010,N_5547);
and U10598 (N_10598,N_9213,N_8956);
or U10599 (N_10599,N_9766,N_5003);
and U10600 (N_10600,N_5632,N_9078);
nand U10601 (N_10601,N_5749,N_7640);
nand U10602 (N_10602,N_7226,N_7747);
nor U10603 (N_10603,N_9612,N_7411);
nand U10604 (N_10604,N_5933,N_5318);
xnor U10605 (N_10605,N_8600,N_6698);
or U10606 (N_10606,N_5966,N_5752);
or U10607 (N_10607,N_9457,N_8837);
nor U10608 (N_10608,N_8502,N_6442);
nand U10609 (N_10609,N_9731,N_8844);
nand U10610 (N_10610,N_7311,N_7201);
or U10611 (N_10611,N_9497,N_6562);
xor U10612 (N_10612,N_6884,N_9689);
and U10613 (N_10613,N_5625,N_9435);
nand U10614 (N_10614,N_6398,N_6900);
xor U10615 (N_10615,N_6072,N_9062);
xor U10616 (N_10616,N_9269,N_9925);
nand U10617 (N_10617,N_6446,N_6855);
or U10618 (N_10618,N_7261,N_8578);
nor U10619 (N_10619,N_5483,N_6886);
nor U10620 (N_10620,N_5274,N_5343);
nor U10621 (N_10621,N_9127,N_8839);
and U10622 (N_10622,N_8196,N_7764);
nor U10623 (N_10623,N_5551,N_7455);
nor U10624 (N_10624,N_9093,N_6003);
and U10625 (N_10625,N_8542,N_8714);
or U10626 (N_10626,N_8999,N_5323);
nand U10627 (N_10627,N_8319,N_5927);
xor U10628 (N_10628,N_9126,N_6543);
nand U10629 (N_10629,N_8687,N_8630);
xnor U10630 (N_10630,N_6218,N_6561);
and U10631 (N_10631,N_5720,N_8257);
nand U10632 (N_10632,N_5473,N_8995);
or U10633 (N_10633,N_5100,N_8838);
nand U10634 (N_10634,N_9671,N_9388);
or U10635 (N_10635,N_7852,N_8452);
and U10636 (N_10636,N_5947,N_9281);
and U10637 (N_10637,N_5178,N_6472);
nor U10638 (N_10638,N_9651,N_9920);
or U10639 (N_10639,N_8175,N_5548);
and U10640 (N_10640,N_7122,N_9298);
or U10641 (N_10641,N_9921,N_5685);
and U10642 (N_10642,N_5095,N_8277);
nand U10643 (N_10643,N_5553,N_7285);
nand U10644 (N_10644,N_7053,N_7834);
or U10645 (N_10645,N_8114,N_9295);
xor U10646 (N_10646,N_5139,N_7435);
nand U10647 (N_10647,N_8344,N_6857);
nor U10648 (N_10648,N_9313,N_9207);
xnor U10649 (N_10649,N_9801,N_6033);
nand U10650 (N_10650,N_9879,N_5523);
or U10651 (N_10651,N_8386,N_5140);
and U10652 (N_10652,N_9714,N_6856);
nor U10653 (N_10653,N_5024,N_7178);
nor U10654 (N_10654,N_7301,N_9212);
or U10655 (N_10655,N_8797,N_5605);
nor U10656 (N_10656,N_5660,N_5731);
nor U10657 (N_10657,N_8199,N_9568);
nor U10658 (N_10658,N_5629,N_9045);
xnor U10659 (N_10659,N_8631,N_9111);
and U10660 (N_10660,N_9618,N_8796);
nor U10661 (N_10661,N_7241,N_6904);
nor U10662 (N_10662,N_5289,N_8174);
nand U10663 (N_10663,N_9449,N_8424);
nor U10664 (N_10664,N_5465,N_5351);
or U10665 (N_10665,N_7273,N_7352);
and U10666 (N_10666,N_6615,N_7485);
nor U10667 (N_10667,N_5025,N_7332);
nand U10668 (N_10668,N_9302,N_8658);
and U10669 (N_10669,N_9900,N_6024);
nand U10670 (N_10670,N_8784,N_8987);
nor U10671 (N_10671,N_8942,N_9747);
xor U10672 (N_10672,N_5975,N_6664);
or U10673 (N_10673,N_9365,N_6707);
and U10674 (N_10674,N_9200,N_6414);
nand U10675 (N_10675,N_7735,N_6603);
xor U10676 (N_10676,N_6482,N_5147);
nor U10677 (N_10677,N_6214,N_5973);
or U10678 (N_10678,N_8361,N_7349);
nor U10679 (N_10679,N_8028,N_5697);
or U10680 (N_10680,N_8887,N_5109);
or U10681 (N_10681,N_6427,N_5707);
nor U10682 (N_10682,N_7437,N_8753);
nand U10683 (N_10683,N_9726,N_9899);
nor U10684 (N_10684,N_5782,N_5045);
or U10685 (N_10685,N_5658,N_6502);
nor U10686 (N_10686,N_9971,N_5410);
nor U10687 (N_10687,N_5093,N_9529);
and U10688 (N_10688,N_8285,N_8763);
or U10689 (N_10689,N_8020,N_9287);
or U10690 (N_10690,N_7762,N_5698);
and U10691 (N_10691,N_7691,N_9386);
nor U10692 (N_10692,N_8460,N_9871);
and U10693 (N_10693,N_8780,N_8179);
nand U10694 (N_10694,N_5992,N_6686);
and U10695 (N_10695,N_7678,N_9335);
or U10696 (N_10696,N_9271,N_9973);
and U10697 (N_10697,N_6008,N_6302);
nand U10698 (N_10698,N_9946,N_8928);
and U10699 (N_10699,N_9012,N_5663);
and U10700 (N_10700,N_8127,N_6177);
nor U10701 (N_10701,N_9950,N_6772);
nand U10702 (N_10702,N_8855,N_8738);
nor U10703 (N_10703,N_6818,N_5284);
nor U10704 (N_10704,N_8336,N_9038);
or U10705 (N_10705,N_6252,N_7741);
and U10706 (N_10706,N_7316,N_7794);
nand U10707 (N_10707,N_6993,N_8312);
or U10708 (N_10708,N_9903,N_9280);
xnor U10709 (N_10709,N_7511,N_6397);
xor U10710 (N_10710,N_9667,N_9050);
nor U10711 (N_10711,N_6709,N_5608);
nand U10712 (N_10712,N_7843,N_7502);
or U10713 (N_10713,N_6574,N_9759);
or U10714 (N_10714,N_9416,N_8003);
and U10715 (N_10715,N_6512,N_8668);
nor U10716 (N_10716,N_7739,N_5777);
nor U10717 (N_10717,N_5769,N_8354);
nand U10718 (N_10718,N_5737,N_7304);
and U10719 (N_10719,N_9566,N_8353);
nor U10720 (N_10720,N_9347,N_9754);
and U10721 (N_10721,N_5635,N_7360);
and U10722 (N_10722,N_5651,N_6019);
and U10723 (N_10723,N_8804,N_7400);
and U10724 (N_10724,N_6099,N_9277);
nor U10725 (N_10725,N_8413,N_5878);
nor U10726 (N_10726,N_5119,N_7567);
nor U10727 (N_10727,N_7923,N_9947);
nand U10728 (N_10728,N_7136,N_8205);
nor U10729 (N_10729,N_8936,N_5647);
nand U10730 (N_10730,N_8168,N_6433);
nor U10731 (N_10731,N_7016,N_5993);
and U10732 (N_10732,N_6327,N_7789);
xor U10733 (N_10733,N_5107,N_7378);
and U10734 (N_10734,N_6326,N_5330);
or U10735 (N_10735,N_9865,N_6260);
nand U10736 (N_10736,N_5742,N_7383);
or U10737 (N_10737,N_7193,N_5383);
or U10738 (N_10738,N_9509,N_9586);
nand U10739 (N_10739,N_6148,N_8181);
or U10740 (N_10740,N_8696,N_9316);
and U10741 (N_10741,N_9110,N_7221);
nor U10742 (N_10742,N_9955,N_5768);
nor U10743 (N_10743,N_8377,N_8984);
nor U10744 (N_10744,N_6235,N_6174);
and U10745 (N_10745,N_5481,N_5930);
nand U10746 (N_10746,N_8149,N_9985);
or U10747 (N_10747,N_9697,N_6308);
nand U10748 (N_10748,N_8375,N_5272);
nor U10749 (N_10749,N_5630,N_6998);
and U10750 (N_10750,N_9717,N_6905);
nor U10751 (N_10751,N_9135,N_8596);
and U10752 (N_10752,N_7068,N_7288);
nand U10753 (N_10753,N_9969,N_6037);
nand U10754 (N_10754,N_5921,N_6558);
nand U10755 (N_10755,N_8895,N_5876);
nor U10756 (N_10756,N_5260,N_6628);
nand U10757 (N_10757,N_9709,N_6426);
xor U10758 (N_10758,N_9507,N_9013);
nand U10759 (N_10759,N_6955,N_6152);
or U10760 (N_10760,N_6110,N_5105);
xnor U10761 (N_10761,N_6468,N_8405);
nand U10762 (N_10762,N_5004,N_9237);
or U10763 (N_10763,N_8388,N_5937);
xor U10764 (N_10764,N_9409,N_6135);
nor U10765 (N_10765,N_7395,N_6333);
nor U10766 (N_10766,N_6733,N_7138);
and U10767 (N_10767,N_7913,N_6196);
or U10768 (N_10768,N_9656,N_5543);
nand U10769 (N_10769,N_9774,N_7476);
or U10770 (N_10770,N_8684,N_6285);
nor U10771 (N_10771,N_6198,N_9223);
xnor U10772 (N_10772,N_6584,N_9090);
nor U10773 (N_10773,N_6560,N_7719);
nor U10774 (N_10774,N_6029,N_9575);
nor U10775 (N_10775,N_5038,N_6636);
and U10776 (N_10776,N_6279,N_7173);
or U10777 (N_10777,N_6764,N_8982);
or U10778 (N_10778,N_9376,N_9859);
and U10779 (N_10779,N_6572,N_5595);
or U10780 (N_10780,N_7305,N_8439);
nor U10781 (N_10781,N_9962,N_9825);
nand U10782 (N_10782,N_6073,N_6754);
and U10783 (N_10783,N_5561,N_9323);
and U10784 (N_10784,N_5695,N_5368);
or U10785 (N_10785,N_5814,N_6322);
nand U10786 (N_10786,N_9289,N_7978);
nor U10787 (N_10787,N_7180,N_8157);
or U10788 (N_10788,N_8098,N_9419);
nor U10789 (N_10789,N_7891,N_6513);
and U10790 (N_10790,N_6644,N_8881);
or U10791 (N_10791,N_6589,N_7209);
nand U10792 (N_10792,N_7013,N_9356);
and U10793 (N_10793,N_6424,N_5504);
nor U10794 (N_10794,N_6160,N_9220);
or U10795 (N_10795,N_9360,N_5322);
xor U10796 (N_10796,N_9125,N_6192);
or U10797 (N_10797,N_5389,N_6695);
nand U10798 (N_10798,N_6997,N_6609);
and U10799 (N_10799,N_6417,N_6352);
and U10800 (N_10800,N_9603,N_6088);
nor U10801 (N_10801,N_6362,N_7099);
nor U10802 (N_10802,N_9954,N_6910);
nand U10803 (N_10803,N_7755,N_6678);
and U10804 (N_10804,N_8165,N_9454);
nand U10805 (N_10805,N_7561,N_7635);
and U10806 (N_10806,N_9520,N_5783);
nand U10807 (N_10807,N_7363,N_5711);
nor U10808 (N_10808,N_8806,N_5867);
or U10809 (N_10809,N_9301,N_7591);
and U10810 (N_10810,N_6963,N_7058);
and U10811 (N_10811,N_7712,N_6112);
and U10812 (N_10812,N_5827,N_5002);
or U10813 (N_10813,N_9310,N_6936);
or U10814 (N_10814,N_5577,N_7944);
nor U10815 (N_10815,N_6897,N_6422);
nor U10816 (N_10816,N_7279,N_6619);
or U10817 (N_10817,N_7022,N_5948);
and U10818 (N_10818,N_7680,N_9456);
and U10819 (N_10819,N_7706,N_8131);
and U10820 (N_10820,N_9746,N_7336);
nor U10821 (N_10821,N_5175,N_7269);
or U10822 (N_10822,N_9961,N_6815);
or U10823 (N_10823,N_7644,N_8445);
and U10824 (N_10824,N_8644,N_7681);
xnor U10825 (N_10825,N_7346,N_9040);
or U10826 (N_10826,N_7247,N_9931);
nor U10827 (N_10827,N_7249,N_5132);
xor U10828 (N_10828,N_9155,N_5363);
or U10829 (N_10829,N_6585,N_7085);
xnor U10830 (N_10830,N_5249,N_6504);
nor U10831 (N_10831,N_5764,N_7535);
and U10832 (N_10832,N_7171,N_8478);
and U10833 (N_10833,N_8778,N_5090);
or U10834 (N_10834,N_6068,N_8929);
nor U10835 (N_10835,N_8209,N_5807);
and U10836 (N_10836,N_8659,N_5667);
nor U10837 (N_10837,N_5108,N_5626);
nand U10838 (N_10838,N_6486,N_6962);
and U10839 (N_10839,N_6945,N_7417);
and U10840 (N_10840,N_5297,N_7883);
nor U10841 (N_10841,N_5150,N_5808);
nand U10842 (N_10842,N_5578,N_8585);
nor U10843 (N_10843,N_5559,N_6912);
nand U10844 (N_10844,N_9387,N_8023);
nand U10845 (N_10845,N_7271,N_7490);
and U10846 (N_10846,N_8463,N_6967);
nand U10847 (N_10847,N_6136,N_6337);
or U10848 (N_10848,N_8450,N_6076);
nand U10849 (N_10849,N_5825,N_8941);
nand U10850 (N_10850,N_7494,N_7317);
nand U10851 (N_10851,N_5081,N_5405);
nand U10852 (N_10852,N_9091,N_6173);
or U10853 (N_10853,N_9665,N_5896);
nor U10854 (N_10854,N_5016,N_6359);
nand U10855 (N_10855,N_9391,N_8700);
nor U10856 (N_10856,N_9402,N_6114);
and U10857 (N_10857,N_7086,N_9082);
nand U10858 (N_10858,N_5853,N_7819);
nor U10859 (N_10859,N_9791,N_8154);
xnor U10860 (N_10860,N_5757,N_6168);
or U10861 (N_10861,N_9645,N_9132);
xnor U10862 (N_10862,N_8710,N_6665);
or U10863 (N_10863,N_5763,N_6401);
nand U10864 (N_10864,N_8970,N_6781);
nand U10865 (N_10865,N_9351,N_6529);
or U10866 (N_10866,N_8359,N_7036);
and U10867 (N_10867,N_7496,N_9100);
nand U10868 (N_10868,N_8429,N_9221);
nand U10869 (N_10869,N_8067,N_6932);
nor U10870 (N_10870,N_5282,N_8723);
or U10871 (N_10871,N_8482,N_5919);
nor U10872 (N_10872,N_5471,N_8089);
nand U10873 (N_10873,N_5954,N_6974);
xnor U10874 (N_10874,N_9232,N_5380);
or U10875 (N_10875,N_6635,N_6125);
xor U10876 (N_10876,N_9011,N_5193);
nand U10877 (N_10877,N_8966,N_7028);
or U10878 (N_10878,N_8649,N_9680);
nor U10879 (N_10879,N_6935,N_5588);
nor U10880 (N_10880,N_8789,N_5397);
and U10881 (N_10881,N_5220,N_7833);
nand U10882 (N_10882,N_9594,N_5842);
or U10883 (N_10883,N_8263,N_6965);
and U10884 (N_10884,N_9115,N_7894);
nand U10885 (N_10885,N_5549,N_7633);
and U10886 (N_10886,N_6251,N_9661);
and U10887 (N_10887,N_9545,N_7050);
xor U10888 (N_10888,N_8739,N_6626);
or U10889 (N_10889,N_6836,N_6246);
nor U10890 (N_10890,N_9181,N_6244);
or U10891 (N_10891,N_8831,N_8449);
or U10892 (N_10892,N_9572,N_8550);
nor U10893 (N_10893,N_5505,N_5110);
nand U10894 (N_10894,N_6042,N_6445);
nor U10895 (N_10895,N_5557,N_9796);
nand U10896 (N_10896,N_9556,N_7207);
nand U10897 (N_10897,N_5830,N_8299);
xnor U10898 (N_10898,N_7418,N_7179);
nor U10899 (N_10899,N_8949,N_7528);
or U10900 (N_10900,N_8599,N_8607);
or U10901 (N_10901,N_6991,N_7339);
or U10902 (N_10902,N_7105,N_6773);
and U10903 (N_10903,N_5664,N_8817);
and U10904 (N_10904,N_9856,N_6576);
nand U10905 (N_10905,N_7609,N_9685);
nand U10906 (N_10906,N_8697,N_6056);
nor U10907 (N_10907,N_8932,N_7558);
nor U10908 (N_10908,N_9487,N_8541);
nor U10909 (N_10909,N_8543,N_9994);
nand U10910 (N_10910,N_8430,N_5787);
or U10911 (N_10911,N_7592,N_5231);
nor U10912 (N_10912,N_8264,N_5353);
or U10913 (N_10913,N_8132,N_7150);
nand U10914 (N_10914,N_7523,N_7868);
xnor U10915 (N_10915,N_9833,N_6966);
and U10916 (N_10916,N_8448,N_9787);
nand U10917 (N_10917,N_6649,N_9690);
or U10918 (N_10918,N_9346,N_8678);
or U10919 (N_10919,N_5895,N_5591);
or U10920 (N_10920,N_6575,N_7612);
nand U10921 (N_10921,N_9342,N_7856);
nor U10922 (N_10922,N_9602,N_6096);
or U10923 (N_10923,N_6657,N_6140);
and U10924 (N_10924,N_8051,N_6075);
nand U10925 (N_10925,N_5071,N_7479);
nand U10926 (N_10926,N_5219,N_5171);
or U10927 (N_10927,N_9185,N_9552);
nor U10928 (N_10928,N_8548,N_5427);
and U10929 (N_10929,N_9702,N_9514);
nand U10930 (N_10930,N_9761,N_7467);
nor U10931 (N_10931,N_8705,N_5462);
nor U10932 (N_10932,N_8546,N_7607);
nor U10933 (N_10933,N_6613,N_9421);
nor U10934 (N_10934,N_9085,N_6802);
and U10935 (N_10935,N_7869,N_5458);
or U10936 (N_10936,N_6364,N_5030);
nor U10937 (N_10937,N_5327,N_6030);
nand U10938 (N_10938,N_9075,N_9205);
nor U10939 (N_10939,N_7223,N_7787);
nand U10940 (N_10940,N_8491,N_9571);
and U10941 (N_10941,N_8516,N_5350);
nor U10942 (N_10942,N_9614,N_7231);
xnor U10943 (N_10943,N_9129,N_7433);
xnor U10944 (N_10944,N_7236,N_7469);
and U10945 (N_10945,N_9118,N_7679);
and U10946 (N_10946,N_8619,N_7011);
or U10947 (N_10947,N_9142,N_6289);
nand U10948 (N_10948,N_9767,N_7194);
nand U10949 (N_10949,N_6931,N_6163);
and U10950 (N_10950,N_8983,N_7732);
and U10951 (N_10951,N_6633,N_5494);
xor U10952 (N_10952,N_5583,N_6495);
or U10953 (N_10953,N_7893,N_5080);
and U10954 (N_10954,N_9197,N_6986);
xnor U10955 (N_10955,N_7096,N_6851);
xor U10956 (N_10956,N_6420,N_9361);
nand U10957 (N_10957,N_8474,N_6641);
and U10958 (N_10958,N_9321,N_5325);
nor U10959 (N_10959,N_9530,N_7060);
or U10960 (N_10960,N_7564,N_9949);
nand U10961 (N_10961,N_8317,N_6825);
or U10962 (N_10962,N_7666,N_9776);
or U10963 (N_10963,N_7563,N_9385);
and U10964 (N_10964,N_9465,N_6494);
and U10965 (N_10965,N_6047,N_7109);
or U10966 (N_10966,N_9744,N_7107);
nor U10967 (N_10967,N_7098,N_7183);
and U10968 (N_10968,N_6234,N_6200);
and U10969 (N_10969,N_6866,N_5228);
nor U10970 (N_10970,N_6146,N_7386);
nand U10971 (N_10971,N_8637,N_6437);
nand U10972 (N_10972,N_5304,N_6017);
nand U10973 (N_10973,N_7097,N_7345);
nor U10974 (N_10974,N_5006,N_9311);
or U10975 (N_10975,N_6777,N_5146);
xor U10976 (N_10976,N_5316,N_8189);
nor U10977 (N_10977,N_7263,N_6654);
or U10978 (N_10978,N_7376,N_8824);
nor U10979 (N_10979,N_6026,N_9240);
and U10980 (N_10980,N_7624,N_5008);
nand U10981 (N_10981,N_8677,N_5202);
nand U10982 (N_10982,N_7526,N_6176);
and U10983 (N_10983,N_8403,N_8222);
nor U10984 (N_10984,N_6663,N_6715);
xnor U10985 (N_10985,N_7948,N_5790);
and U10986 (N_10986,N_5114,N_5035);
and U10987 (N_10987,N_8969,N_8760);
nor U10988 (N_10988,N_7292,N_6758);
and U10989 (N_10989,N_8080,N_9842);
nor U10990 (N_10990,N_5540,N_7015);
nor U10991 (N_10991,N_9217,N_9909);
or U10992 (N_10992,N_5944,N_9133);
or U10993 (N_10993,N_5470,N_8755);
and U10994 (N_10994,N_8115,N_5340);
or U10995 (N_10995,N_8193,N_6992);
nand U10996 (N_10996,N_8284,N_7228);
or U10997 (N_10997,N_8331,N_9793);
or U10998 (N_10998,N_7248,N_6880);
nand U10999 (N_10999,N_9348,N_6386);
and U11000 (N_11000,N_8950,N_9079);
and U11001 (N_11001,N_9934,N_9912);
nor U11002 (N_11002,N_6216,N_8048);
or U11003 (N_11003,N_7335,N_5659);
nor U11004 (N_11004,N_9166,N_8426);
nand U11005 (N_11005,N_8864,N_8878);
and U11006 (N_11006,N_5267,N_9393);
and U11007 (N_11007,N_6201,N_5204);
nor U11008 (N_11008,N_7862,N_8082);
or U11009 (N_11009,N_5773,N_6793);
nor U11010 (N_11010,N_9415,N_7562);
and U11011 (N_11011,N_7665,N_5058);
or U11012 (N_11012,N_8171,N_6444);
xor U11013 (N_11013,N_5692,N_8725);
nor U11014 (N_11014,N_5277,N_6703);
and U11015 (N_11015,N_6942,N_6493);
nand U11016 (N_11016,N_9732,N_8639);
nand U11017 (N_11017,N_9574,N_8694);
or U11018 (N_11018,N_7368,N_7214);
nand U11019 (N_11019,N_7002,N_5426);
xnor U11020 (N_11020,N_6452,N_9150);
or U11021 (N_11021,N_9108,N_9666);
and U11022 (N_11022,N_5064,N_9202);
and U11023 (N_11023,N_7749,N_5333);
nand U11024 (N_11024,N_8202,N_7134);
and U11025 (N_11025,N_6236,N_7343);
xnor U11026 (N_11026,N_5501,N_6810);
and U11027 (N_11027,N_5020,N_5716);
nand U11028 (N_11028,N_7413,N_5478);
nand U11029 (N_11029,N_5556,N_9283);
nand U11030 (N_11030,N_7427,N_9945);
nor U11031 (N_11031,N_8019,N_9642);
or U11032 (N_11032,N_7979,N_5166);
nor U11033 (N_11033,N_5726,N_7559);
and U11034 (N_11034,N_8433,N_7290);
nor U11035 (N_11035,N_6968,N_5154);
or U11036 (N_11036,N_6366,N_6858);
nor U11037 (N_11037,N_7019,N_8757);
nor U11038 (N_11038,N_6184,N_6286);
or U11039 (N_11039,N_9832,N_9214);
nor U11040 (N_11040,N_8745,N_7275);
or U11041 (N_11041,N_8105,N_5718);
and U11042 (N_11042,N_5420,N_5117);
xor U11043 (N_11043,N_9608,N_8957);
nor U11044 (N_11044,N_6127,N_7245);
or U11045 (N_11045,N_7188,N_5740);
and U11046 (N_11046,N_6981,N_9668);
and U11047 (N_11047,N_8588,N_9953);
nor U11048 (N_11048,N_6717,N_9991);
nor U11049 (N_11049,N_9795,N_5934);
nor U11050 (N_11050,N_9576,N_5665);
or U11051 (N_11051,N_6161,N_8258);
nor U11052 (N_11052,N_6632,N_8192);
nand U11053 (N_11053,N_8961,N_6610);
xor U11054 (N_11054,N_7367,N_7566);
or U11055 (N_11055,N_6608,N_9503);
nor U11056 (N_11056,N_8027,N_7142);
nand U11057 (N_11057,N_9654,N_8385);
nand U11058 (N_11058,N_6012,N_7572);
nand U11059 (N_11059,N_9854,N_8102);
nor U11060 (N_11060,N_6539,N_8221);
and U11061 (N_11061,N_6238,N_5396);
or U11062 (N_11062,N_9001,N_7634);
nand U11063 (N_11063,N_5067,N_9990);
and U11064 (N_11064,N_8279,N_6631);
nand U11065 (N_11065,N_9849,N_6418);
or U11066 (N_11066,N_8910,N_5360);
nor U11067 (N_11067,N_9306,N_5802);
nand U11068 (N_11068,N_8292,N_8651);
nand U11069 (N_11069,N_6207,N_9857);
or U11070 (N_11070,N_7174,N_9737);
nand U11071 (N_11071,N_9884,N_7932);
or U11072 (N_11072,N_9646,N_7850);
and U11073 (N_11073,N_9543,N_7521);
nand U11074 (N_11074,N_5053,N_9655);
xor U11075 (N_11075,N_8747,N_7059);
and U11076 (N_11076,N_9596,N_6342);
and U11077 (N_11077,N_6875,N_5815);
nand U11078 (N_11078,N_9748,N_7605);
and U11079 (N_11079,N_6392,N_8471);
and U11080 (N_11080,N_5857,N_7394);
or U11081 (N_11081,N_8728,N_9784);
and U11082 (N_11082,N_7806,N_5872);
or U11083 (N_11083,N_7610,N_5967);
and U11084 (N_11084,N_6188,N_8065);
or U11085 (N_11085,N_5541,N_5084);
nor U11086 (N_11086,N_5165,N_7095);
and U11087 (N_11087,N_7639,N_6953);
nor U11088 (N_11088,N_7531,N_8842);
or U11089 (N_11089,N_7823,N_7674);
or U11090 (N_11090,N_8256,N_9610);
nor U11091 (N_11091,N_7066,N_9395);
xor U11092 (N_11092,N_8660,N_6642);
nand U11093 (N_11093,N_6973,N_7151);
or U11094 (N_11094,N_5366,N_5345);
xor U11095 (N_11095,N_7046,N_9288);
and U11096 (N_11096,N_9341,N_6428);
nor U11097 (N_11097,N_7205,N_5841);
or U11098 (N_11098,N_6311,N_6274);
or U11099 (N_11099,N_5238,N_8562);
and U11100 (N_11100,N_6915,N_9527);
nor U11101 (N_11101,N_9476,N_7373);
or U11102 (N_11102,N_7076,N_5762);
and U11103 (N_11103,N_5240,N_8920);
or U11104 (N_11104,N_9339,N_8085);
and U11105 (N_11105,N_9951,N_6730);
or U11106 (N_11106,N_7268,N_5871);
xor U11107 (N_11107,N_6400,N_7074);
nand U11108 (N_11108,N_6149,N_9300);
nor U11109 (N_11109,N_8876,N_5168);
nor U11110 (N_11110,N_6542,N_7990);
xnor U11111 (N_11111,N_5218,N_5015);
and U11112 (N_11112,N_9615,N_7154);
nor U11113 (N_11113,N_5498,N_9848);
nand U11114 (N_11114,N_7257,N_8937);
and U11115 (N_11115,N_8574,N_9218);
and U11116 (N_11116,N_8015,N_5445);
or U11117 (N_11117,N_8593,N_7553);
nand U11118 (N_11118,N_5708,N_5184);
nand U11119 (N_11119,N_9718,N_9810);
or U11120 (N_11120,N_5352,N_7130);
nand U11121 (N_11121,N_8333,N_5791);
nor U11122 (N_11122,N_6674,N_8985);
or U11123 (N_11123,N_9915,N_7169);
nor U11124 (N_11124,N_7251,N_5315);
nor U11125 (N_11125,N_7131,N_9253);
and U11126 (N_11126,N_5684,N_7969);
nand U11127 (N_11127,N_8306,N_7161);
or U11128 (N_11128,N_7892,N_6505);
nor U11129 (N_11129,N_6830,N_9080);
and U11130 (N_11130,N_9713,N_8390);
or U11131 (N_11131,N_6199,N_7927);
and U11132 (N_11132,N_6926,N_5281);
nor U11133 (N_11133,N_5159,N_8311);
and U11134 (N_11134,N_7964,N_7025);
nand U11135 (N_11135,N_9525,N_9916);
nand U11136 (N_11136,N_7321,N_9098);
nor U11137 (N_11137,N_7370,N_5336);
and U11138 (N_11138,N_8524,N_8224);
xnor U11139 (N_11139,N_8809,N_5034);
nor U11140 (N_11140,N_6895,N_8167);
nand U11141 (N_11141,N_7303,N_9522);
nand U11142 (N_11142,N_5390,N_5694);
nand U11143 (N_11143,N_9840,N_7084);
nand U11144 (N_11144,N_8195,N_8352);
xnor U11145 (N_11145,N_7041,N_8802);
and U11146 (N_11146,N_5600,N_7544);
or U11147 (N_11147,N_8416,N_6850);
and U11148 (N_11148,N_9658,N_9432);
nand U11149 (N_11149,N_8822,N_5858);
or U11150 (N_11150,N_5487,N_6845);
nor U11151 (N_11151,N_9781,N_6181);
nand U11152 (N_11152,N_9860,N_8974);
or U11153 (N_11153,N_9471,N_7585);
xnor U11154 (N_11154,N_6097,N_8177);
nor U11155 (N_11155,N_7630,N_7202);
or U11156 (N_11156,N_7092,N_6501);
nand U11157 (N_11157,N_5946,N_6690);
and U11158 (N_11158,N_5291,N_6259);
xnor U11159 (N_11159,N_7796,N_5772);
or U11160 (N_11160,N_6175,N_9975);
nor U11161 (N_11161,N_5488,N_7880);
nand U11162 (N_11162,N_6335,N_5833);
nand U11163 (N_11163,N_9882,N_7873);
and U11164 (N_11164,N_6179,N_6721);
and U11165 (N_11165,N_9549,N_8618);
nor U11166 (N_11166,N_6172,N_7459);
nand U11167 (N_11167,N_6402,N_7752);
nor U11168 (N_11168,N_9988,N_9797);
nand U11169 (N_11169,N_7056,N_6368);
nor U11170 (N_11170,N_9473,N_8616);
and U11171 (N_11171,N_7030,N_7682);
or U11172 (N_11172,N_8253,N_8963);
or U11173 (N_11173,N_8421,N_7430);
and U11174 (N_11174,N_6421,N_6049);
nor U11175 (N_11175,N_9230,N_8807);
nor U11176 (N_11176,N_9326,N_8298);
nand U11177 (N_11177,N_8566,N_7723);
nand U11178 (N_11178,N_5868,N_6384);
nand U11179 (N_11179,N_5091,N_6989);
or U11180 (N_11180,N_5932,N_6629);
or U11181 (N_11181,N_7128,N_6022);
or U11182 (N_11182,N_8013,N_7444);
and U11183 (N_11183,N_6602,N_5348);
xor U11184 (N_11184,N_7992,N_6776);
and U11185 (N_11185,N_7265,N_5950);
nand U11186 (N_11186,N_8825,N_9984);
or U11187 (N_11187,N_6524,N_6169);
or U11188 (N_11188,N_6580,N_5820);
nor U11189 (N_11189,N_7460,N_7334);
nand U11190 (N_11190,N_7448,N_7658);
and U11191 (N_11191,N_7905,N_7195);
and U11192 (N_11192,N_7676,N_9554);
or U11193 (N_11193,N_7687,N_5459);
nand U11194 (N_11194,N_7587,N_9033);
or U11195 (N_11195,N_9538,N_6985);
nand U11196 (N_11196,N_8034,N_9030);
xor U11197 (N_11197,N_5940,N_7307);
nand U11198 (N_11198,N_6783,N_9948);
nor U11199 (N_11199,N_6206,N_6257);
xor U11200 (N_11200,N_9980,N_7407);
or U11201 (N_11201,N_5717,N_5294);
and U11202 (N_11202,N_9939,N_7825);
xor U11203 (N_11203,N_6954,N_6567);
or U11204 (N_11204,N_9122,N_6262);
nor U11205 (N_11205,N_8693,N_9662);
nor U11206 (N_11206,N_7874,N_8721);
nor U11207 (N_11207,N_6078,N_6194);
or U11208 (N_11208,N_8695,N_9331);
nor U11209 (N_11209,N_5645,N_8959);
or U11210 (N_11210,N_6086,N_7326);
or U11211 (N_11211,N_9493,N_9875);
nand U11212 (N_11212,N_8420,N_6275);
nand U11213 (N_11213,N_7828,N_9336);
xnor U11214 (N_11214,N_6429,N_8321);
and U11215 (N_11215,N_5040,N_9712);
and U11216 (N_11216,N_8381,N_8376);
nand U11217 (N_11217,N_7034,N_5130);
or U11218 (N_11218,N_5356,N_5531);
nand U11219 (N_11219,N_9249,N_7778);
or U11220 (N_11220,N_6687,N_5186);
or U11221 (N_11221,N_8689,N_8058);
and U11222 (N_11222,N_5076,N_5379);
nand U11223 (N_11223,N_5622,N_7067);
xnor U11224 (N_11224,N_7904,N_6645);
xnor U11225 (N_11225,N_9806,N_7483);
xnor U11226 (N_11226,N_8303,N_9187);
and U11227 (N_11227,N_7487,N_9944);
nor U11228 (N_11228,N_9101,N_7000);
nand U11229 (N_11229,N_6180,N_6240);
and U11230 (N_11230,N_8236,N_6153);
nand U11231 (N_11231,N_5183,N_8230);
nand U11232 (N_11232,N_8552,N_6438);
nand U11233 (N_11233,N_9105,N_5295);
nor U11234 (N_11234,N_7181,N_8664);
nor U11235 (N_11235,N_7888,N_9640);
and U11236 (N_11236,N_7374,N_7579);
nand U11237 (N_11237,N_7818,N_7262);
nor U11238 (N_11238,N_7914,N_5899);
nor U11239 (N_11239,N_8587,N_7457);
and U11240 (N_11240,N_5957,N_5836);
nand U11241 (N_11241,N_5923,N_8145);
nor U11242 (N_11242,N_9629,N_5305);
and U11243 (N_11243,N_8849,N_9845);
nand U11244 (N_11244,N_9404,N_8672);
and U11245 (N_11245,N_7756,N_8190);
and U11246 (N_11246,N_9422,N_5900);
or U11247 (N_11247,N_8801,N_7441);
nor U11248 (N_11248,N_9508,N_6911);
nor U11249 (N_11249,N_9450,N_6228);
and U11250 (N_11250,N_7399,N_6872);
nor U11251 (N_11251,N_8061,N_7470);
nand U11252 (N_11252,N_7938,N_6557);
nor U11253 (N_11253,N_7534,N_7791);
nor U11254 (N_11254,N_7645,N_9414);
or U11255 (N_11255,N_9235,N_7765);
nor U11256 (N_11256,N_8355,N_5998);
nor U11257 (N_11257,N_8378,N_6510);
and U11258 (N_11258,N_8611,N_5903);
nand U11259 (N_11259,N_8056,N_5796);
nand U11260 (N_11260,N_5280,N_6247);
or U11261 (N_11261,N_7045,N_8229);
and U11262 (N_11262,N_9262,N_8836);
or U11263 (N_11263,N_7031,N_6659);
or U11264 (N_11264,N_5566,N_7446);
nor U11265 (N_11265,N_7695,N_6860);
or U11266 (N_11266,N_8510,N_7550);
nor U11267 (N_11267,N_7902,N_5436);
or U11268 (N_11268,N_5758,N_5209);
or U11269 (N_11269,N_5550,N_9710);
xnor U11270 (N_11270,N_9019,N_7235);
and U11271 (N_11271,N_9338,N_7295);
and U11272 (N_11272,N_8924,N_8086);
and U11273 (N_11273,N_6312,N_9140);
nand U11274 (N_11274,N_6838,N_9309);
and U11275 (N_11275,N_6109,N_5594);
nor U11276 (N_11276,N_6716,N_9170);
nor U11277 (N_11277,N_9261,N_9817);
nand U11278 (N_11278,N_5275,N_6531);
nand U11279 (N_11279,N_6010,N_9590);
xnor U11280 (N_11280,N_7940,N_9227);
or U11281 (N_11281,N_8508,N_8832);
xor U11282 (N_11282,N_7939,N_8976);
or U11283 (N_11283,N_8539,N_5042);
and U11284 (N_11284,N_8237,N_9433);
and U11285 (N_11285,N_7903,N_9028);
and U11286 (N_11286,N_8125,N_7541);
or U11287 (N_11287,N_6646,N_8708);
nor U11288 (N_11288,N_9864,N_6000);
and U11289 (N_11289,N_8477,N_7946);
nor U11290 (N_11290,N_8185,N_5450);
and U11291 (N_11291,N_9490,N_8868);
nand U11292 (N_11292,N_7657,N_9067);
or U11293 (N_11293,N_8282,N_7125);
and U11294 (N_11294,N_9657,N_7683);
nor U11295 (N_11295,N_9438,N_8766);
nor U11296 (N_11296,N_6193,N_5883);
nand U11297 (N_11297,N_6028,N_9757);
xnor U11298 (N_11298,N_8070,N_9228);
nor U11299 (N_11299,N_6506,N_9659);
nand U11300 (N_11300,N_8742,N_5029);
nand U11301 (N_11301,N_7536,N_7298);
xnor U11302 (N_11302,N_7227,N_9631);
xor U11303 (N_11303,N_5104,N_5845);
nor U11304 (N_11304,N_5910,N_9163);
nor U11305 (N_11305,N_9441,N_7065);
or U11306 (N_11306,N_5617,N_7675);
nand U11307 (N_11307,N_6488,N_6903);
nor U11308 (N_11308,N_9183,N_8113);
or U11309 (N_11309,N_8634,N_5987);
or U11310 (N_11310,N_6448,N_5674);
nand U11311 (N_11311,N_8217,N_7114);
nand U11312 (N_11312,N_8492,N_8041);
or U11313 (N_11313,N_6611,N_5800);
and U11314 (N_11314,N_7991,N_7689);
nor U11315 (N_11315,N_7966,N_5492);
nor U11316 (N_11316,N_7007,N_8988);
and U11317 (N_11317,N_5191,N_9137);
or U11318 (N_11318,N_5499,N_7697);
or U11319 (N_11319,N_7668,N_9141);
nand U11320 (N_11320,N_5404,N_5437);
nor U11321 (N_11321,N_5861,N_7529);
or U11322 (N_11322,N_8818,N_6318);
nor U11323 (N_11323,N_5721,N_9055);
nand U11324 (N_11324,N_9134,N_6868);
or U11325 (N_11325,N_6726,N_5824);
xnor U11326 (N_11326,N_5654,N_6620);
nand U11327 (N_11327,N_6803,N_7786);
nand U11328 (N_11328,N_8129,N_7425);
xor U11329 (N_11329,N_5358,N_5185);
nor U11330 (N_11330,N_8719,N_6225);
and U11331 (N_11331,N_8635,N_8520);
xnor U11332 (N_11332,N_9052,N_9216);
and U11333 (N_11333,N_8912,N_8440);
nand U11334 (N_11334,N_9208,N_5293);
nand U11335 (N_11335,N_9462,N_5813);
nor U11336 (N_11336,N_7196,N_7421);
or U11337 (N_11337,N_5888,N_8402);
nor U11338 (N_11338,N_5848,N_6074);
and U11339 (N_11339,N_8427,N_6786);
nor U11340 (N_11340,N_6332,N_6638);
or U11341 (N_11341,N_5563,N_5809);
nor U11342 (N_11342,N_8923,N_8033);
nor U11343 (N_11343,N_7005,N_9092);
nor U11344 (N_11344,N_6081,N_5092);
or U11345 (N_11345,N_5781,N_5098);
and U11346 (N_11346,N_9940,N_8880);
or U11347 (N_11347,N_6554,N_6828);
or U11348 (N_11348,N_6839,N_9151);
nand U11349 (N_11349,N_7975,N_5544);
and U11350 (N_11350,N_5497,N_9046);
nor U11351 (N_11351,N_6380,N_6406);
xnor U11352 (N_11352,N_8896,N_6041);
and U11353 (N_11353,N_6891,N_5941);
and U11354 (N_11354,N_7976,N_5224);
and U11355 (N_11355,N_9986,N_5978);
and U11356 (N_11356,N_5525,N_8111);
nor U11357 (N_11357,N_9070,N_8459);
or U11358 (N_11358,N_5986,N_6467);
and U11359 (N_11359,N_7919,N_8243);
nand U11360 (N_11360,N_6515,N_8479);
nor U11361 (N_11361,N_6616,N_5898);
nor U11362 (N_11362,N_7445,N_9350);
nor U11363 (N_11363,N_9407,N_7583);
or U11364 (N_11364,N_6727,N_8095);
nor U11365 (N_11365,N_6889,N_6412);
and U11366 (N_11366,N_8118,N_7164);
nand U11367 (N_11367,N_9917,N_7815);
or U11368 (N_11368,N_5672,N_5170);
xnor U11369 (N_11369,N_5652,N_8846);
nor U11370 (N_11370,N_7864,N_5734);
nand U11371 (N_11371,N_5065,N_5197);
nand U11372 (N_11372,N_7801,N_8517);
nor U11373 (N_11373,N_9725,N_5965);
nand U11374 (N_11374,N_5509,N_7018);
and U11375 (N_11375,N_7361,N_6742);
nand U11376 (N_11376,N_7884,N_7763);
and U11377 (N_11377,N_5257,N_5306);
nor U11378 (N_11378,N_5417,N_8137);
xnor U11379 (N_11379,N_8208,N_8045);
nand U11380 (N_11380,N_5795,N_8083);
and U11381 (N_11381,N_5361,N_9704);
or U11382 (N_11382,N_9445,N_9236);
xnor U11383 (N_11383,N_6065,N_8497);
nor U11384 (N_11384,N_6549,N_9863);
nand U11385 (N_11385,N_5736,N_9412);
or U11386 (N_11386,N_7491,N_5088);
nor U11387 (N_11387,N_6307,N_8206);
nand U11388 (N_11388,N_6759,N_7552);
nor U11389 (N_11389,N_9064,N_8011);
nor U11390 (N_11390,N_9172,N_7140);
nand U11391 (N_11391,N_6837,N_5066);
xnor U11392 (N_11392,N_6928,N_9794);
nor U11393 (N_11393,N_9993,N_8555);
and U11394 (N_11394,N_9866,N_8947);
nor U11395 (N_11395,N_5099,N_6519);
nand U11396 (N_11396,N_5214,N_8676);
nor U11397 (N_11397,N_9904,N_8255);
or U11398 (N_11398,N_7351,N_7925);
nand U11399 (N_11399,N_6313,N_5970);
xnor U11400 (N_11400,N_8641,N_7686);
and U11401 (N_11401,N_5639,N_9799);
or U11402 (N_11402,N_5653,N_9703);
nand U11403 (N_11403,N_6165,N_7988);
xor U11404 (N_11404,N_5068,N_6832);
nor U11405 (N_11405,N_5935,N_9452);
or U11406 (N_11406,N_7039,N_7943);
nor U11407 (N_11407,N_8706,N_7837);
nor U11408 (N_11408,N_9158,N_6306);
nand U11409 (N_11409,N_6516,N_5158);
or U11410 (N_11410,N_7119,N_5288);
nand U11411 (N_11411,N_9641,N_5527);
nor U11412 (N_11412,N_9898,N_7643);
nor U11413 (N_11413,N_9999,N_8161);
or U11414 (N_11414,N_5334,N_9624);
nand U11415 (N_11415,N_9083,N_9189);
and U11416 (N_11416,N_8055,N_6958);
or U11417 (N_11417,N_8271,N_8341);
or U11418 (N_11418,N_8252,N_5994);
xor U11419 (N_11419,N_6355,N_5057);
and U11420 (N_11420,N_9057,N_6697);
nor U11421 (N_11421,N_9319,N_9770);
nor U11422 (N_11422,N_6565,N_7911);
and U11423 (N_11423,N_6834,N_8260);
or U11424 (N_11424,N_7115,N_8730);
and U11425 (N_11425,N_8717,N_6011);
nor U11426 (N_11426,N_5760,N_8410);
nor U11427 (N_11427,N_7410,N_6440);
or U11428 (N_11428,N_5262,N_7802);
nand U11429 (N_11429,N_8357,N_9632);
or U11430 (N_11430,N_5565,N_5195);
nor U11431 (N_11431,N_5007,N_7871);
or U11432 (N_11432,N_5256,N_5924);
nor U11433 (N_11433,N_8265,N_5774);
nor U11434 (N_11434,N_5378,N_8833);
or U11435 (N_11435,N_6278,N_8428);
nor U11436 (N_11436,N_7865,N_7348);
xnor U11437 (N_11437,N_9811,N_8638);
nor U11438 (N_11438,N_7576,N_5864);
and U11439 (N_11439,N_6077,N_6846);
xor U11440 (N_11440,N_6004,N_6652);
xor U11441 (N_11441,N_6334,N_9084);
or U11442 (N_11442,N_6351,N_5443);
or U11443 (N_11443,N_9785,N_8346);
nand U11444 (N_11444,N_7887,N_8843);
nor U11445 (N_11445,N_9830,N_5575);
xnor U11446 (N_11446,N_9039,N_9088);
nor U11447 (N_11447,N_6164,N_7848);
or U11448 (N_11448,N_5706,N_8939);
and U11449 (N_11449,N_8538,N_9152);
nand U11450 (N_11450,N_8109,N_7518);
or U11451 (N_11451,N_9906,N_5837);
nand U11452 (N_11452,N_8438,N_8628);
or U11453 (N_11453,N_8169,N_9173);
xnor U11454 (N_11454,N_8558,N_7406);
and U11455 (N_11455,N_9358,N_8645);
or U11456 (N_11456,N_6887,N_6689);
and U11457 (N_11457,N_5120,N_7928);
and U11458 (N_11458,N_8971,N_5235);
or U11459 (N_11459,N_5902,N_7646);
and U11460 (N_11460,N_9565,N_5298);
and U11461 (N_11461,N_6593,N_6949);
and U11462 (N_11462,N_5959,N_5269);
or U11463 (N_11463,N_8458,N_8313);
nor U11464 (N_11464,N_8363,N_8901);
or U11465 (N_11465,N_5958,N_7960);
nor U11466 (N_11466,N_8123,N_9472);
nand U11467 (N_11467,N_5724,N_8627);
xnor U11468 (N_11468,N_9061,N_5096);
and U11469 (N_11469,N_7842,N_9579);
and U11470 (N_11470,N_8768,N_9911);
nor U11471 (N_11471,N_7973,N_5371);
nand U11472 (N_11472,N_7641,N_8248);
nand U11473 (N_11473,N_5369,N_5806);
and U11474 (N_11474,N_7147,N_9332);
and U11475 (N_11475,N_7688,N_5753);
nand U11476 (N_11476,N_6765,N_7703);
nor U11477 (N_11477,N_7745,N_9724);
or U11478 (N_11478,N_5237,N_8680);
or U11479 (N_11479,N_7724,N_6747);
nor U11480 (N_11480,N_6245,N_7748);
and U11481 (N_11481,N_8581,N_8530);
nor U11482 (N_11482,N_8466,N_5991);
nor U11483 (N_11483,N_7578,N_7052);
or U11484 (N_11484,N_5788,N_7001);
and U11485 (N_11485,N_6769,N_9255);
nand U11486 (N_11486,N_7208,N_8905);
or U11487 (N_11487,N_6600,N_5200);
or U11488 (N_11488,N_7358,N_7896);
nor U11489 (N_11489,N_5988,N_5590);
nor U11490 (N_11490,N_7573,N_5585);
nor U11491 (N_11491,N_8952,N_6941);
or U11492 (N_11492,N_9820,N_9501);
or U11493 (N_11493,N_8769,N_7993);
xor U11494 (N_11494,N_9451,N_8493);
nor U11495 (N_11495,N_6215,N_7861);
and U11496 (N_11496,N_6243,N_7062);
nor U11497 (N_11497,N_9381,N_6023);
nor U11498 (N_11498,N_9042,N_6290);
nor U11499 (N_11499,N_7281,N_5816);
nand U11500 (N_11500,N_5079,N_9653);
nor U11501 (N_11501,N_9584,N_9698);
and U11502 (N_11502,N_8242,N_6425);
nor U11503 (N_11503,N_8432,N_8874);
or U11504 (N_11504,N_9516,N_7388);
nand U11505 (N_11505,N_5276,N_7211);
nand U11506 (N_11506,N_9320,N_9059);
nor U11507 (N_11507,N_9029,N_6592);
nor U11508 (N_11508,N_5464,N_7355);
nand U11509 (N_11509,N_9044,N_7040);
and U11510 (N_11510,N_7721,N_5961);
nand U11511 (N_11511,N_7726,N_9739);
nor U11512 (N_11512,N_8057,N_7568);
and U11513 (N_11513,N_6933,N_9479);
nor U11514 (N_11514,N_5083,N_8891);
nand U11515 (N_11515,N_5382,N_6925);
nor U11516 (N_11516,N_6411,N_5246);
nor U11517 (N_11517,N_7473,N_6990);
nand U11518 (N_11518,N_8278,N_7729);
nand U11519 (N_11519,N_6242,N_8106);
or U11520 (N_11520,N_7621,N_9562);
nand U11521 (N_11521,N_6885,N_8794);
and U11522 (N_11522,N_8525,N_5689);
and U11523 (N_11523,N_9582,N_5346);
and U11524 (N_11524,N_5014,N_5882);
xnor U11525 (N_11525,N_7397,N_6273);
nand U11526 (N_11526,N_5060,N_6117);
xor U11527 (N_11527,N_8322,N_5703);
nand U11528 (N_11528,N_7515,N_9588);
nor U11529 (N_11529,N_8834,N_8945);
and U11530 (N_11530,N_9162,N_5143);
and U11531 (N_11531,N_9673,N_6893);
nor U11532 (N_11532,N_6708,N_5311);
nor U11533 (N_11533,N_9669,N_8093);
nand U11534 (N_11534,N_6607,N_6182);
nand U11535 (N_11535,N_5728,N_5976);
or U11536 (N_11536,N_8736,N_9542);
or U11537 (N_11537,N_7799,N_5877);
nor U11538 (N_11538,N_8401,N_8561);
nor U11539 (N_11539,N_6924,N_8266);
or U11540 (N_11540,N_7935,N_5118);
and U11541 (N_11541,N_8162,N_6757);
nand U11542 (N_11542,N_7608,N_9835);
nor U11543 (N_11543,N_7051,N_7442);
nand U11544 (N_11544,N_5624,N_5243);
nor U11545 (N_11545,N_9478,N_6864);
and U11546 (N_11546,N_8752,N_6100);
nand U11547 (N_11547,N_9815,N_9677);
or U11548 (N_11548,N_6634,N_5033);
nand U11549 (N_11549,N_5409,N_7210);
nor U11550 (N_11550,N_6525,N_5767);
nand U11551 (N_11551,N_9807,N_8540);
nor U11552 (N_11552,N_7910,N_7365);
nor U11553 (N_11553,N_6901,N_9410);
nand U11554 (N_11554,N_5572,N_5681);
and U11555 (N_11555,N_6020,N_9378);
or U11556 (N_11556,N_7189,N_9905);
nand U11557 (N_11557,N_5511,N_9936);
nand U11558 (N_11558,N_5798,N_9191);
or U11559 (N_11559,N_8393,N_8182);
and U11560 (N_11560,N_7078,N_5039);
nand U11561 (N_11561,N_9477,N_8349);
xnor U11562 (N_11562,N_6485,N_8549);
nor U11563 (N_11563,N_8409,N_5687);
or U11564 (N_11564,N_7297,N_5913);
nor U11565 (N_11565,N_7213,N_5701);
or U11566 (N_11566,N_8305,N_5049);
or U11567 (N_11567,N_5401,N_8854);
or U11568 (N_11568,N_6637,N_7499);
and U11569 (N_11569,N_8654,N_8135);
and U11570 (N_11570,N_7387,N_9094);
nor U11571 (N_11571,N_8219,N_7308);
nor U11572 (N_11572,N_6133,N_6469);
nor U11573 (N_11573,N_5456,N_8776);
nand U11574 (N_11574,N_6403,N_6498);
and U11575 (N_11575,N_8472,N_8770);
or U11576 (N_11576,N_7443,N_9648);
or U11577 (N_11577,N_6013,N_7492);
xnor U11578 (N_11578,N_5210,N_7728);
nand U11579 (N_11579,N_9550,N_9660);
and U11580 (N_11580,N_8496,N_8441);
nand U11581 (N_11581,N_7839,N_6205);
and U11582 (N_11582,N_6916,N_6085);
xor U11583 (N_11583,N_5347,N_7813);
nand U11584 (N_11584,N_5198,N_8018);
or U11585 (N_11585,N_9204,N_6025);
nor U11586 (N_11586,N_9359,N_6876);
and U11587 (N_11587,N_9926,N_8215);
nor U11588 (N_11588,N_8044,N_9113);
nor U11589 (N_11589,N_9136,N_7933);
nand U11590 (N_11590,N_8751,N_5880);
nand U11591 (N_11591,N_5448,N_6581);
nand U11592 (N_11592,N_6979,N_7877);
nor U11593 (N_11593,N_8958,N_6454);
or U11594 (N_11594,N_7477,N_7146);
or U11595 (N_11595,N_8006,N_5475);
nand U11596 (N_11596,N_7080,N_6118);
nand U11597 (N_11597,N_8761,N_8727);
nand U11598 (N_11598,N_6569,N_5709);
xor U11599 (N_11599,N_7713,N_5604);
or U11600 (N_11600,N_9519,N_5968);
and U11601 (N_11601,N_7432,N_5225);
nor U11602 (N_11602,N_5286,N_6413);
or U11603 (N_11603,N_7968,N_8883);
nor U11604 (N_11604,N_7218,N_7986);
nor U11605 (N_11605,N_7575,N_6643);
and U11606 (N_11606,N_7751,N_5502);
nor U11607 (N_11607,N_5643,N_7590);
nand U11608 (N_11608,N_9741,N_5597);
nor U11609 (N_11609,N_9475,N_9488);
nor U11610 (N_11610,N_8454,N_9000);
or U11611 (N_11611,N_8373,N_6929);
xor U11612 (N_11612,N_7588,N_6157);
nor U11613 (N_11613,N_9296,N_5077);
or U11614 (N_11614,N_7889,N_6343);
or U11615 (N_11615,N_7921,N_7121);
or U11616 (N_11616,N_5490,N_6699);
and U11617 (N_11617,N_9123,N_5251);
nor U11618 (N_11618,N_8380,N_5317);
nand U11619 (N_11619,N_7929,N_8534);
or U11620 (N_11620,N_7003,N_9682);
or U11621 (N_11621,N_8116,N_8314);
or U11622 (N_11622,N_8869,N_6596);
nor U11623 (N_11623,N_8146,N_5179);
or U11624 (N_11624,N_6079,N_6069);
nor U11625 (N_11625,N_8238,N_7577);
xor U11626 (N_11626,N_8704,N_7389);
and U11627 (N_11627,N_8990,N_6451);
nor U11628 (N_11628,N_9600,N_7949);
nor U11629 (N_11629,N_8345,N_8589);
or U11630 (N_11630,N_8533,N_5552);
nor U11631 (N_11631,N_9324,N_7083);
nor U11632 (N_11632,N_8935,N_9428);
or U11633 (N_11633,N_8682,N_8133);
and U11634 (N_11634,N_6878,N_7094);
nand U11635 (N_11635,N_9068,N_8214);
and U11636 (N_11636,N_5969,N_7937);
xnor U11637 (N_11637,N_8063,N_9380);
or U11638 (N_11638,N_8940,N_8575);
and U11639 (N_11639,N_7772,N_7447);
or U11640 (N_11640,N_8960,N_8690);
and U11641 (N_11641,N_8673,N_9749);
and U11642 (N_11642,N_5233,N_7829);
nand U11643 (N_11643,N_5089,N_8712);
or U11644 (N_11644,N_6514,N_6760);
xnor U11645 (N_11645,N_6178,N_5730);
or U11646 (N_11646,N_5780,N_6108);
and U11647 (N_11647,N_5909,N_8476);
and U11648 (N_11648,N_9164,N_5539);
or U11649 (N_11649,N_9368,N_8667);
and U11650 (N_11650,N_9981,N_5162);
xor U11651 (N_11651,N_7278,N_7685);
nor U11652 (N_11652,N_6329,N_8663);
or U11653 (N_11653,N_6797,N_9149);
nor U11654 (N_11654,N_6092,N_6831);
or U11655 (N_11655,N_6982,N_7628);
xnor U11656 (N_11656,N_7565,N_9773);
nor U11657 (N_11657,N_5241,N_9621);
and U11658 (N_11658,N_8754,N_7651);
nor U11659 (N_11659,N_9382,N_8000);
or U11660 (N_11660,N_8840,N_8425);
nor U11661 (N_11661,N_7947,N_8603);
and U11662 (N_11662,N_9097,N_7461);
nor U11663 (N_11663,N_5799,N_5115);
nand U11664 (N_11664,N_9587,N_7715);
or U11665 (N_11665,N_5995,N_8308);
nor U11666 (N_11666,N_8835,N_9541);
and U11667 (N_11667,N_5339,N_7471);
or U11668 (N_11668,N_5953,N_8200);
nand U11669 (N_11669,N_7704,N_6021);
and U11670 (N_11670,N_6294,N_9468);
xor U11671 (N_11671,N_5949,N_8374);
nor U11672 (N_11672,N_5628,N_9814);
or U11673 (N_11673,N_7601,N_7734);
or U11674 (N_11674,N_5589,N_6419);
nor U11675 (N_11675,N_7770,N_9234);
or U11676 (N_11676,N_9958,N_7853);
nand U11677 (N_11677,N_6375,N_8953);
nand U11678 (N_11678,N_9683,N_9345);
nand U11679 (N_11679,N_6586,N_5230);
and U11680 (N_11680,N_6799,N_6009);
xor U11681 (N_11681,N_6710,N_9701);
nand U11682 (N_11682,N_6822,N_6606);
xor U11683 (N_11683,N_8791,N_9066);
nand U11684 (N_11684,N_5989,N_6477);
or U11685 (N_11685,N_9156,N_5746);
and U11686 (N_11686,N_6304,N_9553);
nand U11687 (N_11687,N_8269,N_7101);
or U11688 (N_11688,N_9771,N_8178);
nand U11689 (N_11689,N_7580,N_9577);
nor U11690 (N_11690,N_7369,N_5656);
nor U11691 (N_11691,N_5485,N_5592);
nand U11692 (N_11692,N_9089,N_8652);
nand U11693 (N_11693,N_8703,N_7493);
or U11694 (N_11694,N_8120,N_8060);
xnor U11695 (N_11695,N_6051,N_8722);
or U11696 (N_11696,N_7629,N_6712);
xnor U11697 (N_11697,N_8931,N_5865);
and U11698 (N_11698,N_9913,N_6788);
and U11699 (N_11699,N_9455,N_6859);
nor U11700 (N_11700,N_9396,N_5250);
or U11701 (N_11701,N_5085,N_9919);
or U11702 (N_11702,N_5662,N_7649);
nand U11703 (N_11703,N_8733,N_7941);
nor U11704 (N_11704,N_5000,N_9159);
or U11705 (N_11705,N_9215,N_9974);
and U11706 (N_11706,N_9023,N_9838);
nor U11707 (N_11707,N_9790,N_9180);
xnor U11708 (N_11708,N_6261,N_8698);
nor U11709 (N_11709,N_5570,N_8819);
nand U11710 (N_11710,N_9005,N_5177);
or U11711 (N_11711,N_8062,N_8005);
and U11712 (N_11712,N_9171,N_5500);
and U11713 (N_11713,N_8316,N_5245);
xnor U11714 (N_11714,N_6399,N_8972);
nor U11715 (N_11715,N_6094,N_5713);
and U11716 (N_11716,N_6918,N_8396);
or U11717 (N_11717,N_9037,N_5657);
nand U11718 (N_11718,N_9850,N_7047);
or U11719 (N_11719,N_6061,N_8324);
xnor U11720 (N_11720,N_7145,N_8234);
or U11721 (N_11721,N_7698,N_9206);
nand U11722 (N_11722,N_5770,N_9231);
or U11723 (N_11723,N_8612,N_6254);
and U11724 (N_11724,N_7981,N_6134);
or U11725 (N_11725,N_5722,N_5897);
and U11726 (N_11726,N_8035,N_6119);
nor U11727 (N_11727,N_8281,N_5136);
or U11728 (N_11728,N_7431,N_9868);
xnor U11729 (N_11729,N_7232,N_8715);
nand U11730 (N_11730,N_7930,N_6796);
and U11731 (N_11731,N_7072,N_6719);
nor U11732 (N_11732,N_7717,N_7498);
or U11733 (N_11733,N_9357,N_7555);
xnor U11734 (N_11734,N_7716,N_7543);
and U11735 (N_11735,N_9161,N_7454);
nand U11736 (N_11736,N_9964,N_6271);
or U11737 (N_11737,N_8328,N_8075);
or U11738 (N_11738,N_6139,N_9750);
nand U11739 (N_11739,N_9561,N_9742);
or U11740 (N_11740,N_7952,N_9738);
xnor U11741 (N_11741,N_8038,N_8097);
or U11742 (N_11742,N_6662,N_8139);
nand U11743 (N_11743,N_9408,N_9663);
nand U11744 (N_11744,N_9370,N_5097);
and U11745 (N_11745,N_9178,N_8933);
nand U11746 (N_11746,N_6145,N_9009);
or U11747 (N_11747,N_6210,N_5069);
and U11748 (N_11748,N_8187,N_6511);
or U11749 (N_11749,N_6409,N_8437);
xor U11750 (N_11750,N_7168,N_6888);
or U11751 (N_11751,N_7750,N_5188);
nor U11752 (N_11752,N_6579,N_5564);
or U11753 (N_11753,N_7381,N_9015);
nand U11754 (N_11754,N_5794,N_9276);
or U11755 (N_11755,N_6761,N_6520);
and U11756 (N_11756,N_5812,N_7781);
and U11757 (N_11757,N_7405,N_9967);
nand U11758 (N_11758,N_8632,N_8743);
and U11759 (N_11759,N_9716,N_9006);
nor U11760 (N_11760,N_7501,N_5894);
xnor U11761 (N_11761,N_9389,N_8515);
nor U11762 (N_11762,N_7042,N_5054);
nor U11763 (N_11763,N_8138,N_8773);
or U11764 (N_11764,N_5860,N_7392);
or U11765 (N_11765,N_7475,N_8943);
nor U11766 (N_11766,N_8342,N_9492);
or U11767 (N_11767,N_8604,N_9691);
or U11768 (N_11768,N_8096,N_5213);
or U11769 (N_11769,N_9293,N_6546);
xor U11770 (N_11770,N_5252,N_6296);
and U11771 (N_11771,N_7872,N_8201);
xor U11772 (N_11772,N_6381,N_7586);
or U11773 (N_11773,N_8514,N_8431);
nand U11774 (N_11774,N_9364,N_8340);
nand U11775 (N_11775,N_6458,N_7186);
xnor U11776 (N_11776,N_7330,N_9692);
nand U11777 (N_11777,N_6762,N_7474);
and U11778 (N_11778,N_7520,N_6208);
nor U11779 (N_11779,N_9880,N_5254);
nor U11780 (N_11780,N_9383,N_5546);
nand U11781 (N_11781,N_9555,N_7338);
or U11782 (N_11782,N_8391,N_5890);
or U11783 (N_11783,N_6751,N_7384);
nor U11784 (N_11784,N_8827,N_5466);
and U11785 (N_11785,N_8748,N_7505);
nand U11786 (N_11786,N_8909,N_7648);
and U11787 (N_11787,N_5834,N_9872);
xnor U11788 (N_11788,N_7424,N_7664);
xnor U11789 (N_11789,N_9131,N_9285);
nand U11790 (N_11790,N_5392,N_5938);
or U11791 (N_11791,N_6655,N_9203);
nor U11792 (N_11792,N_5425,N_7684);
xor U11793 (N_11793,N_7239,N_9020);
nand U11794 (N_11794,N_8498,N_7302);
nand U11795 (N_11795,N_9675,N_9877);
or U11796 (N_11796,N_8504,N_5568);
nor U11797 (N_11797,N_7216,N_5750);
nand U11798 (N_11798,N_6131,N_9598);
nor U11799 (N_11799,N_7306,N_7780);
or U11800 (N_11800,N_9819,N_6132);
and U11801 (N_11801,N_8759,N_9557);
nand U11802 (N_11802,N_8364,N_9401);
nand U11803 (N_11803,N_9439,N_8362);
or U11804 (N_11804,N_6090,N_9484);
nor U11805 (N_11805,N_9165,N_8370);
nor U11806 (N_11806,N_9540,N_6474);
nor U11807 (N_11807,N_6457,N_7983);
and U11808 (N_11808,N_6497,N_7073);
nand U11809 (N_11809,N_6701,N_6820);
or U11810 (N_11810,N_8025,N_5367);
or U11811 (N_11811,N_7163,N_7184);
and U11812 (N_11812,N_5535,N_7875);
nor U11813 (N_11813,N_7702,N_8400);
xor U11814 (N_11814,N_5661,N_5440);
nor U11815 (N_11815,N_7816,N_6594);
nand U11816 (N_11816,N_9120,N_6058);
nor U11817 (N_11817,N_5859,N_7945);
and U11818 (N_11818,N_8790,N_5920);
nand U11819 (N_11819,N_5637,N_7785);
nand U11820 (N_11820,N_8398,N_5222);
nand U11821 (N_11821,N_5370,N_9867);
nor U11822 (N_11822,N_7758,N_7215);
or U11823 (N_11823,N_7847,N_8367);
nor U11824 (N_11824,N_6416,N_8079);
nand U11825 (N_11825,N_7385,N_6833);
nor U11826 (N_11826,N_5063,N_6480);
or U11827 (N_11827,N_6158,N_7560);
nand U11828 (N_11828,N_9041,N_8665);
nor U11829 (N_11829,N_8885,N_5255);
or U11830 (N_11830,N_7143,N_6994);
and U11831 (N_11831,N_6624,N_8522);
nor U11832 (N_11832,N_9374,N_9526);
nand U11833 (N_11833,N_5850,N_7141);
and U11834 (N_11834,N_5418,N_5453);
or U11835 (N_11835,N_5623,N_8039);
xnor U11836 (N_11836,N_6694,N_5649);
and U11837 (N_11837,N_5614,N_8047);
nand U11838 (N_11838,N_9444,N_7478);
xor U11839 (N_11839,N_6728,N_6983);
and U11840 (N_11840,N_7995,N_7117);
and U11841 (N_11841,N_7313,N_6478);
and U11842 (N_11842,N_9979,N_8605);
nand U11843 (N_11843,N_5926,N_6229);
xnor U11844 (N_11844,N_9349,N_7614);
nor U11845 (N_11845,N_6155,N_6879);
and U11846 (N_11846,N_8980,N_7325);
and U11847 (N_11847,N_9392,N_7434);
nor U11848 (N_11848,N_6104,N_7931);
or U11849 (N_11849,N_5962,N_6039);
and U11850 (N_11850,N_6032,N_8126);
nor U11851 (N_11851,N_9330,N_8103);
and U11852 (N_11852,N_9016,N_6491);
nor U11853 (N_11853,N_7331,N_6345);
xor U11854 (N_11854,N_8501,N_8858);
and U11855 (N_11855,N_9824,N_8016);
or U11856 (N_11856,N_5047,N_7845);
or U11857 (N_11857,N_9996,N_9081);
xor U11858 (N_11858,N_6435,N_8172);
nand U11859 (N_11859,N_9436,N_8513);
or U11860 (N_11860,N_9510,N_9252);
nand U11861 (N_11861,N_9504,N_6826);
or U11862 (N_11862,N_8233,N_8629);
nand U11863 (N_11863,N_9902,N_6755);
nand U11864 (N_11864,N_5738,N_8793);
nand U11865 (N_11865,N_6305,N_5914);
or U11866 (N_11866,N_9453,N_8259);
nor U11867 (N_11867,N_5190,N_7353);
and U11868 (N_11868,N_9266,N_6142);
or U11869 (N_11869,N_8468,N_9403);
nand U11870 (N_11870,N_6170,N_5818);
nand U11871 (N_11871,N_9694,N_6340);
and U11872 (N_11872,N_8764,N_8267);
xnor U11873 (N_11873,N_8571,N_7449);
nor U11874 (N_11874,N_7743,N_7530);
nor U11875 (N_11875,N_9290,N_6946);
or U11876 (N_11876,N_6122,N_6829);
or U11877 (N_11877,N_7830,N_8335);
and U11878 (N_11878,N_8551,N_8897);
or U11879 (N_11879,N_7123,N_9117);
nand U11880 (N_11880,N_6704,N_6187);
xor U11881 (N_11881,N_5922,N_8967);
and U11882 (N_11882,N_5508,N_6927);
nor U11883 (N_11883,N_9637,N_7252);
nor U11884 (N_11884,N_9294,N_6363);
xor U11885 (N_11885,N_8785,N_5283);
xor U11886 (N_11886,N_7693,N_7625);
nand U11887 (N_11887,N_7606,N_7167);
or U11888 (N_11888,N_8486,N_9209);
xor U11889 (N_11889,N_5180,N_6394);
nand U11890 (N_11890,N_6952,N_8228);
nor U11891 (N_11891,N_5518,N_7250);
and U11892 (N_11892,N_8052,N_6756);
or U11893 (N_11893,N_6521,N_9499);
nand U11894 (N_11894,N_6407,N_8128);
nand U11895 (N_11895,N_7804,N_5832);
nand U11896 (N_11896,N_5503,N_6067);
nand U11897 (N_11897,N_9580,N_6323);
and U11898 (N_11898,N_5619,N_7617);
nor U11899 (N_11899,N_8915,N_7488);
nor U11900 (N_11900,N_5022,N_8494);
or U11901 (N_11901,N_8334,N_7314);
nand U11902 (N_11902,N_7967,N_7882);
nand U11903 (N_11903,N_9827,N_8418);
nand U11904 (N_11904,N_9885,N_7768);
nor U11905 (N_11905,N_7222,N_5817);
nand U11906 (N_11906,N_5977,N_8601);
nand U11907 (N_11907,N_6348,N_5884);
nor U11908 (N_11908,N_5216,N_8412);
or U11909 (N_11909,N_8666,N_5688);
xor U11910 (N_11910,N_8332,N_8247);
and U11911 (N_11911,N_6873,N_5881);
nor U11912 (N_11912,N_5537,N_6057);
nor U11913 (N_11913,N_7533,N_6870);
nand U11914 (N_11914,N_6824,N_7546);
and U11915 (N_11915,N_6487,N_5271);
or U11916 (N_11916,N_5273,N_7740);
and U11917 (N_11917,N_8050,N_9847);
and U11918 (N_11918,N_5602,N_6526);
nand U11919 (N_11919,N_5265,N_7596);
or U11920 (N_11920,N_5789,N_6696);
and U11921 (N_11921,N_9420,N_8527);
and U11922 (N_11922,N_6016,N_8820);
nor U11923 (N_11923,N_5223,N_6371);
nand U11924 (N_11924,N_9446,N_9458);
xnor U11925 (N_11925,N_7984,N_6766);
or U11926 (N_11926,N_5227,N_5673);
and U11927 (N_11927,N_8888,N_8223);
or U11928 (N_11928,N_6959,N_7255);
or U11929 (N_11929,N_7242,N_8029);
or U11930 (N_11930,N_8636,N_8621);
and U11931 (N_11931,N_7172,N_9426);
nand U11932 (N_11932,N_8735,N_9883);
or U11933 (N_11933,N_6621,N_7382);
nor U11934 (N_11934,N_6204,N_9375);
and U11935 (N_11935,N_9837,N_5943);
and U11936 (N_11936,N_9711,N_7912);
and U11937 (N_11937,N_9928,N_9377);
nor U11938 (N_11938,N_8347,N_6752);
nand U11939 (N_11939,N_6361,N_5061);
and U11940 (N_11940,N_8900,N_7340);
xor U11941 (N_11941,N_6821,N_7276);
xor U11942 (N_11942,N_6250,N_5402);
nand U11943 (N_11943,N_8609,N_5187);
xnor U11944 (N_11944,N_8088,N_6782);
or U11945 (N_11945,N_9333,N_6545);
or U11946 (N_11946,N_9573,N_5313);
nand U11947 (N_11947,N_8962,N_5699);
xor U11948 (N_11948,N_6914,N_9643);
xnor U11949 (N_11949,N_7835,N_5416);
and U11950 (N_11950,N_8447,N_5001);
nor U11951 (N_11951,N_5761,N_7506);
nand U11952 (N_11952,N_5133,N_5983);
nor U11953 (N_11953,N_9299,N_6902);
nor U11954 (N_11954,N_5419,N_7182);
nor U11955 (N_11955,N_7788,N_7636);
nor U11956 (N_11956,N_5805,N_8998);
or U11957 (N_11957,N_6297,N_7956);
nor U11958 (N_11958,N_5516,N_9548);
and U11959 (N_11959,N_7840,N_6103);
nor U11960 (N_11960,N_7708,N_5554);
or U11961 (N_11961,N_5640,N_8408);
xor U11962 (N_11962,N_8729,N_8358);
or U11963 (N_11963,N_9168,N_6668);
nand U11964 (N_11964,N_5971,N_5247);
and U11965 (N_11965,N_7212,N_8275);
nand U11966 (N_11966,N_9074,N_5705);
and U11967 (N_11967,N_7897,N_8294);
xnor U11968 (N_11968,N_7190,N_5359);
and U11969 (N_11969,N_5891,N_8563);
nor U11970 (N_11970,N_7486,N_5182);
or U11971 (N_11971,N_6732,N_8213);
or U11972 (N_11972,N_7197,N_9354);
and U11973 (N_11973,N_5451,N_7647);
nand U11974 (N_11974,N_5974,N_7632);
nand U11975 (N_11975,N_9768,N_8092);
nand U11976 (N_11976,N_8147,N_9337);
nor U11977 (N_11977,N_9464,N_9829);
or U11978 (N_11978,N_9459,N_6748);
nand U11979 (N_11979,N_6231,N_8300);
nand U11980 (N_11980,N_7057,N_5569);
xor U11981 (N_11981,N_6365,N_7132);
nand U11982 (N_11982,N_6692,N_6476);
nand U11983 (N_11983,N_5489,N_8444);
and U11984 (N_11984,N_5264,N_6150);
nor U11985 (N_11985,N_7731,N_5952);
nor U11986 (N_11986,N_6679,N_7489);
nand U11987 (N_11987,N_9740,N_5032);
nor U11988 (N_11988,N_5009,N_7767);
and U11989 (N_11989,N_8220,N_6814);
nand U11990 (N_11990,N_8004,N_9693);
or U11991 (N_11991,N_8343,N_5094);
or U11992 (N_11992,N_6577,N_9371);
xnor U11993 (N_11993,N_5161,N_9616);
nand U11994 (N_11994,N_8143,N_7156);
nor U11995 (N_11995,N_9537,N_6492);
nand U11996 (N_11996,N_6280,N_5244);
and U11997 (N_11997,N_9720,N_7137);
nand U11998 (N_11998,N_5457,N_5461);
or U11999 (N_11999,N_5725,N_8112);
nand U12000 (N_12000,N_9992,N_6922);
nand U12001 (N_12001,N_8330,N_9027);
and U12002 (N_12002,N_5212,N_5062);
nand U12003 (N_12003,N_5925,N_5648);
and U12004 (N_12004,N_6325,N_8296);
or U12005 (N_12005,N_9966,N_7811);
nand U12006 (N_12006,N_9495,N_7165);
or U12007 (N_12007,N_7229,N_6113);
or U12008 (N_12008,N_9893,N_7797);
nor U12009 (N_12009,N_6738,N_6080);
nor U12010 (N_12010,N_6518,N_8350);
and U12011 (N_12011,N_8465,N_9684);
and U12012 (N_12012,N_9254,N_5618);
or U12013 (N_12013,N_5496,N_7318);
nand U12014 (N_12014,N_8455,N_7220);
and U12015 (N_12015,N_5027,N_6735);
and U12016 (N_12016,N_7238,N_5980);
nand U12017 (N_12017,N_6553,N_7472);
xnor U12018 (N_12018,N_7524,N_6675);
nand U12019 (N_12019,N_9314,N_6350);
or U12020 (N_12020,N_5668,N_6098);
nand U12021 (N_12021,N_6848,N_7513);
and U12022 (N_12022,N_7660,N_6921);
xor U12023 (N_12023,N_7299,N_6599);
nor U12024 (N_12024,N_5844,N_8509);
or U12025 (N_12025,N_8009,N_7977);
and U12026 (N_12026,N_5447,N_7826);
nor U12027 (N_12027,N_8531,N_5056);
or U12028 (N_12028,N_5743,N_6330);
nor U12029 (N_12029,N_5041,N_8919);
and U12030 (N_12030,N_5331,N_6734);
nand U12031 (N_12031,N_6618,N_5430);
or U12032 (N_12032,N_5375,N_9593);
nor U12033 (N_12033,N_6156,N_7482);
nor U12034 (N_12034,N_5512,N_7722);
nor U12035 (N_12035,N_5609,N_5606);
nand U12036 (N_12036,N_5778,N_9130);
or U12037 (N_12037,N_7692,N_9505);
and U12038 (N_12038,N_5075,N_6082);
or U12039 (N_12039,N_5332,N_8186);
or U12040 (N_12040,N_8623,N_6374);
xnor U12041 (N_12041,N_8872,N_9922);
nor U12042 (N_12042,N_5507,N_8913);
nand U12043 (N_12043,N_5354,N_6489);
and U12044 (N_12044,N_7203,N_6185);
and U12045 (N_12045,N_9003,N_8674);
nand U12046 (N_12046,N_9018,N_7139);
nand U12047 (N_12047,N_6239,N_9681);
nand U12048 (N_12048,N_7798,N_8104);
xor U12049 (N_12049,N_9035,N_7926);
and U12050 (N_12050,N_5555,N_7187);
nand U12051 (N_12051,N_8925,N_9427);
and U12052 (N_12052,N_7611,N_7466);
or U12053 (N_12053,N_5581,N_8250);
and U12054 (N_12054,N_8702,N_6685);
xor U12055 (N_12055,N_6791,N_6483);
nor U12056 (N_12056,N_9844,N_8227);
nor U12057 (N_12057,N_6977,N_7106);
or U12058 (N_12058,N_6459,N_6907);
nand U12059 (N_12059,N_8042,N_9874);
nand U12060 (N_12060,N_6129,N_5268);
and U12061 (N_12061,N_6627,N_6490);
and U12062 (N_12062,N_6167,N_6718);
and U12063 (N_12063,N_6301,N_9043);
or U12064 (N_12064,N_6823,N_8480);
nor U12065 (N_12065,N_8286,N_9989);
or U12066 (N_12066,N_8462,N_8711);
nor U12067 (N_12067,N_6680,N_9733);
and U12068 (N_12068,N_9551,N_7516);
and U12069 (N_12069,N_9894,N_9721);
xnor U12070 (N_12070,N_5779,N_8767);
and U12071 (N_12071,N_6303,N_6102);
and U12072 (N_12072,N_9592,N_9440);
or U12073 (N_12073,N_5803,N_6530);
and U12074 (N_12074,N_6249,N_6258);
nand U12075 (N_12075,N_8557,N_9998);
nand U12076 (N_12076,N_5199,N_5840);
and U12077 (N_12077,N_7020,N_6209);
and U12078 (N_12078,N_7733,N_9927);
nand U12079 (N_12079,N_5747,N_6281);
nand U12080 (N_12080,N_7920,N_7112);
nand U12081 (N_12081,N_9112,N_5835);
nor U12082 (N_12082,N_7808,N_9199);
nor U12083 (N_12083,N_6430,N_5113);
nand U12084 (N_12084,N_7503,N_9559);
xnor U12085 (N_12085,N_7569,N_9153);
nor U12086 (N_12086,N_6372,N_9780);
nand U12087 (N_12087,N_8927,N_5852);
or U12088 (N_12088,N_8031,N_6623);
and U12089 (N_12089,N_8862,N_6725);
nand U12090 (N_12090,N_6536,N_6314);
and U12091 (N_12091,N_6913,N_5309);
xnor U12092 (N_12092,N_9823,N_7766);
nand U12093 (N_12093,N_9344,N_5189);
xor U12094 (N_12094,N_6544,N_6800);
nand U12095 (N_12095,N_7237,N_6944);
and U12096 (N_12096,N_5885,N_8902);
nand U12097 (N_12097,N_8930,N_8142);
or U12098 (N_12098,N_5253,N_9627);
nor U12099 (N_12099,N_6055,N_6159);
nand U12100 (N_12100,N_8473,N_9145);
nand U12101 (N_12101,N_7820,N_5324);
or U12102 (N_12102,N_7166,N_7175);
or U12103 (N_12103,N_7296,N_7480);
nand U12104 (N_12104,N_8007,N_5407);
and U12105 (N_12105,N_8151,N_7950);
nor U12106 (N_12106,N_9956,N_8893);
nand U12107 (N_12107,N_6811,N_7917);
or U12108 (N_12108,N_8099,N_6128);
nand U12109 (N_12109,N_6027,N_8506);
and U12110 (N_12110,N_5031,N_8762);
nand U12111 (N_12111,N_7737,N_9442);
nor U12112 (N_12112,N_5101,N_6861);
nor U12113 (N_12113,N_7863,N_5682);
and U12114 (N_12114,N_6559,N_7707);
or U12115 (N_12115,N_5434,N_7465);
nor U12116 (N_12116,N_9327,N_9184);
nor U12117 (N_12117,N_9611,N_5259);
nor U12118 (N_12118,N_8890,N_8180);
or U12119 (N_12119,N_8643,N_8781);
and U12120 (N_12120,N_8273,N_7319);
nor U12121 (N_12121,N_6975,N_5229);
nor U12122 (N_12122,N_8164,N_5423);
nand U12123 (N_12123,N_5603,N_9581);
and U12124 (N_12124,N_7429,N_9626);
and U12125 (N_12125,N_9121,N_9194);
nor U12126 (N_12126,N_6604,N_7409);
and U12127 (N_12127,N_6555,N_7192);
and U12128 (N_12128,N_7159,N_8944);
or U12129 (N_12129,N_7700,N_5533);
nor U12130 (N_12130,N_6969,N_8124);
or U12131 (N_12131,N_7093,N_6284);
nor U12132 (N_12132,N_9719,N_7270);
or U12133 (N_12133,N_5300,N_5142);
nor U12134 (N_12134,N_5821,N_7170);
or U12135 (N_12135,N_5395,N_8387);
nand U12136 (N_12136,N_6091,N_7626);
nand U12137 (N_12137,N_8946,N_6890);
or U12138 (N_12138,N_7256,N_7342);
nor U12139 (N_12139,N_9523,N_6256);
or U12140 (N_12140,N_5862,N_9536);
or U12141 (N_12141,N_7594,N_5169);
nor U12142 (N_12142,N_7885,N_7793);
or U12143 (N_12143,N_6035,N_8150);
or U12144 (N_12144,N_6731,N_9604);
or U12145 (N_12145,N_7951,N_6309);
and U12146 (N_12146,N_9103,N_7890);
nor U12147 (N_12147,N_7038,N_9292);
nor U12148 (N_12148,N_7063,N_8993);
xor U12149 (N_12149,N_5308,N_6217);
nand U12150 (N_12150,N_8481,N_7396);
or U12151 (N_12151,N_9250,N_7354);
and U12152 (N_12152,N_7545,N_5906);
nand U12153 (N_12153,N_8348,N_7359);
xor U12154 (N_12154,N_6230,N_9901);
nor U12155 (N_12155,N_7481,N_5582);
or U12156 (N_12156,N_9803,N_6666);
nor U12157 (N_12157,N_9034,N_9670);
nor U12158 (N_12158,N_6906,N_7812);
or U12159 (N_12159,N_8072,N_6950);
xnor U12160 (N_12160,N_5912,N_7895);
and U12161 (N_12161,N_7860,N_9397);
or U12162 (N_12162,N_6255,N_8528);
nand U12163 (N_12163,N_7540,N_9664);
nand U12164 (N_12164,N_8268,N_7769);
or U12165 (N_12165,N_9547,N_7971);
xnor U12166 (N_12166,N_7452,N_8624);
and U12167 (N_12167,N_6789,N_9595);
and U12168 (N_12168,N_8423,N_6784);
nor U12169 (N_12169,N_5514,N_8021);
nor U12170 (N_12170,N_7997,N_7133);
nand U12171 (N_12171,N_8576,N_7720);
or U12172 (N_12172,N_9533,N_6938);
or U12173 (N_12173,N_5887,N_7694);
xnor U12174 (N_12174,N_5863,N_6183);
and U12175 (N_12175,N_7341,N_6221);
nand U12176 (N_12176,N_8737,N_6370);
nor U12177 (N_12177,N_6431,N_6460);
nand U12178 (N_12178,N_8871,N_6220);
nand U12179 (N_12179,N_5111,N_8283);
xnor U12180 (N_12180,N_6972,N_6892);
nor U12181 (N_12181,N_9869,N_5528);
and U12182 (N_12182,N_7120,N_6923);
nor U12183 (N_12183,N_9816,N_9609);
nand U12184 (N_12184,N_9619,N_9910);
nor U12185 (N_12185,N_6508,N_9775);
nand U12186 (N_12186,N_9897,N_8414);
xor U12187 (N_12187,N_7654,N_8068);
and U12188 (N_12188,N_7987,N_8274);
or U12189 (N_12189,N_7403,N_9753);
nand U12190 (N_12190,N_9188,N_8204);
nand U12191 (N_12191,N_6154,N_9211);
nand U12192 (N_12192,N_7266,N_5929);
nand U12193 (N_12193,N_8964,N_6241);
or U12194 (N_12194,N_5696,N_7870);
nor U12195 (N_12195,N_9413,N_8857);
xnor U12196 (N_12196,N_7287,N_7398);
and U12197 (N_12197,N_7026,N_8490);
and U12198 (N_12198,N_9908,N_8536);
and U12199 (N_12199,N_5121,N_6443);
xor U12200 (N_12200,N_8532,N_9102);
nor U12201 (N_12201,N_9373,N_5287);
nor U12202 (N_12202,N_8744,N_7899);
nand U12203 (N_12203,N_6166,N_7254);
nand U12204 (N_12204,N_7004,N_7087);
nor U12205 (N_12205,N_6048,N_9077);
and U12206 (N_12206,N_8799,N_9500);
nand U12207 (N_12207,N_6588,N_7082);
or U12208 (N_12208,N_6320,N_7324);
nor U12209 (N_12209,N_5675,N_8435);
and U12210 (N_12210,N_5129,N_6391);
or U12211 (N_12211,N_7859,N_9708);
nor U12212 (N_12212,N_7736,N_9965);
and U12213 (N_12213,N_6043,N_6729);
nand U12214 (N_12214,N_6338,N_8606);
or U12215 (N_12215,N_7246,N_7408);
nand U12216 (N_12216,N_6002,N_5620);
xor U12217 (N_12217,N_7637,N_8446);
nor U12218 (N_12218,N_6120,N_9623);
nand U12219 (N_12219,N_6908,N_8783);
nand U12220 (N_12220,N_8765,N_8916);
nand U12221 (N_12221,N_6948,N_5679);
xor U12222 (N_12222,N_8989,N_5321);
xor U12223 (N_12223,N_9628,N_6570);
or U12224 (N_12224,N_5491,N_8064);
nand U12225 (N_12225,N_7965,N_5357);
and U12226 (N_12226,N_8675,N_7805);
and U12227 (N_12227,N_5302,N_5855);
or U12228 (N_12228,N_9937,N_7152);
and U12229 (N_12229,N_5307,N_7243);
and U12230 (N_12230,N_8036,N_6461);
nand U12231 (N_12231,N_9418,N_5613);
or U12232 (N_12232,N_9531,N_8613);
nor U12233 (N_12233,N_8681,N_8655);
nand U12234 (N_12234,N_6787,N_8301);
nand U12235 (N_12235,N_9933,N_9128);
nor U12236 (N_12236,N_7775,N_5683);
or U12237 (N_12237,N_6801,N_5206);
or U12238 (N_12238,N_9674,N_6724);
or U12239 (N_12239,N_6095,N_8337);
and U12240 (N_12240,N_6203,N_8647);
nor U12241 (N_12241,N_5536,N_9601);
or U12242 (N_12242,N_9096,N_6287);
or U12243 (N_12243,N_7366,N_9469);
or U12244 (N_12244,N_8108,N_5484);
nand U12245 (N_12245,N_9304,N_9521);
nand U12246 (N_12246,N_5477,N_9567);
or U12247 (N_12247,N_8568,N_8249);
and U12248 (N_12248,N_7035,N_5826);
and U12249 (N_12249,N_6999,N_6040);
nand U12250 (N_12250,N_7204,N_7972);
nor U12251 (N_12251,N_5337,N_9932);
or U12252 (N_12252,N_5299,N_6379);
nand U12253 (N_12253,N_8270,N_6601);
or U12254 (N_12254,N_8290,N_7088);
and U12255 (N_12255,N_8148,N_5403);
nor U12256 (N_12256,N_5148,N_6582);
nand U12257 (N_12257,N_8992,N_7907);
or U12258 (N_12258,N_7110,N_5310);
xor U12259 (N_12259,N_6358,N_7024);
nand U12260 (N_12260,N_9322,N_6456);
nor U12261 (N_12261,N_9430,N_8371);
xnor U12262 (N_12262,N_6591,N_7959);
nor U12263 (N_12263,N_5455,N_5160);
or U12264 (N_12264,N_7714,N_8577);
nor U12265 (N_12265,N_6881,N_6617);
nor U12266 (N_12266,N_9258,N_5792);
nand U12267 (N_12267,N_7043,N_8724);
or U12268 (N_12268,N_7253,N_6547);
nor U12269 (N_12269,N_7029,N_8973);
nand U12270 (N_12270,N_6344,N_7844);
or U12271 (N_12271,N_6847,N_7440);
nand U12272 (N_12272,N_8726,N_5391);
nand U12273 (N_12273,N_8218,N_6778);
nand U12274 (N_12274,N_9210,N_6293);
and U12275 (N_12275,N_8894,N_9802);
or U12276 (N_12276,N_8597,N_5611);
nor U12277 (N_12277,N_6373,N_5893);
or U12278 (N_12278,N_9764,N_9591);
and U12279 (N_12279,N_9789,N_7272);
or U12280 (N_12280,N_8866,N_6143);
and U12281 (N_12281,N_5964,N_5167);
xnor U12282 (N_12282,N_8823,N_6064);
or U12283 (N_12283,N_9447,N_6794);
and U12284 (N_12284,N_7551,N_8032);
nor U12285 (N_12285,N_8372,N_6291);
nand U12286 (N_12286,N_9778,N_5102);
or U12287 (N_12287,N_9929,N_8443);
xor U12288 (N_12288,N_5870,N_6532);
and U12289 (N_12289,N_7655,N_8030);
nor U12290 (N_12290,N_6573,N_9699);
or U12291 (N_12291,N_5755,N_7838);
nor U12292 (N_12292,N_7963,N_5560);
or U12293 (N_12293,N_8183,N_6578);
or U12294 (N_12294,N_9241,N_8851);
or U12295 (N_12295,N_6084,N_7582);
nand U12296 (N_12296,N_5627,N_9914);
nand U12297 (N_12297,N_8339,N_5843);
or U12298 (N_12298,N_7286,N_6970);
nor U12299 (N_12299,N_7757,N_8087);
nor U12300 (N_12300,N_6059,N_6522);
or U12301 (N_12301,N_5739,N_8954);
nand U12302 (N_12302,N_9201,N_6105);
nand U12303 (N_12303,N_8591,N_5493);
nor U12304 (N_12304,N_7661,N_5194);
nand U12305 (N_12305,N_6115,N_8293);
and U12306 (N_12306,N_9743,N_7464);
and U12307 (N_12307,N_8081,N_8246);
nand U12308 (N_12308,N_5828,N_9539);
nand U12309 (N_12309,N_9143,N_8968);
and U12310 (N_12310,N_5486,N_9245);
nor U12311 (N_12311,N_9343,N_7118);
or U12312 (N_12312,N_9606,N_5823);
and U12313 (N_12313,N_7800,N_5134);
nor U12314 (N_12314,N_7508,N_6527);
or U12315 (N_12315,N_7792,N_8559);
nand U12316 (N_12316,N_8130,N_9751);
nor U12317 (N_12317,N_5748,N_7827);
nand U12318 (N_12318,N_8648,N_9625);
or U12319 (N_12319,N_5072,N_7233);
nand U12320 (N_12320,N_8043,N_7671);
or U12321 (N_12321,N_7199,N_5545);
nor U12322 (N_12322,N_9800,N_5704);
xnor U12323 (N_12323,N_9291,N_8848);
and U12324 (N_12324,N_6566,N_5901);
or U12325 (N_12325,N_9119,N_6265);
and U12326 (N_12326,N_7149,N_8572);
nand U12327 (N_12327,N_5026,N_9583);
or U12328 (N_12328,N_9482,N_9485);
or U12329 (N_12329,N_8022,N_6070);
nor U12330 (N_12330,N_8053,N_6237);
or U12331 (N_12331,N_9448,N_6808);
or U12332 (N_12332,N_6276,N_5607);
or U12333 (N_12333,N_8771,N_6672);
and U12334 (N_12334,N_9779,N_8156);
nand U12335 (N_12335,N_6852,N_8554);
nand U12336 (N_12336,N_9881,N_9873);
or U12337 (N_12337,N_6189,N_8419);
nand U12338 (N_12338,N_9705,N_9808);
nand U12339 (N_12339,N_6465,N_8008);
nand U12340 (N_12340,N_8812,N_8975);
nand U12341 (N_12341,N_8879,N_7867);
and U12342 (N_12342,N_6298,N_5270);
and U12343 (N_12343,N_8535,N_6387);
or U12344 (N_12344,N_7571,N_8758);
nor U12345 (N_12345,N_5365,N_7803);
nand U12346 (N_12346,N_9644,N_9696);
and U12347 (N_12347,N_8685,N_8567);
or U12348 (N_12348,N_6376,N_8404);
and U12349 (N_12349,N_7090,N_8718);
or U12350 (N_12350,N_7277,N_8012);
and U12351 (N_12351,N_9087,N_9558);
nor U12352 (N_12352,N_7507,N_7622);
or U12353 (N_12353,N_5558,N_7008);
nand U12354 (N_12354,N_8856,N_5431);
nor U12355 (N_12355,N_7144,N_8040);
nand U12356 (N_12356,N_8814,N_7176);
nand U12357 (N_12357,N_5192,N_8461);
nand U12358 (N_12358,N_5372,N_5073);
xor U12359 (N_12359,N_5176,N_8338);
nand U12360 (N_12360,N_5234,N_6232);
nor U12361 (N_12361,N_5646,N_6957);
and U12362 (N_12362,N_9275,N_9828);
nand U12363 (N_12363,N_9997,N_5446);
or U12364 (N_12364,N_6548,N_9470);
and U12365 (N_12365,N_9175,N_5215);
or U12366 (N_12366,N_8191,N_9607);
and U12367 (N_12367,N_8503,N_7711);
nor U12368 (N_12368,N_9532,N_5911);
nor U12369 (N_12369,N_9918,N_8938);
nor U12370 (N_12370,N_8155,N_8368);
nand U12371 (N_12371,N_6395,N_9496);
nor U12372 (N_12372,N_6930,N_7322);
nor U12373 (N_12373,N_5650,N_5580);
nor U12374 (N_12374,N_5510,N_5017);
nand U12375 (N_12375,N_6647,N_9058);
or U12376 (N_12376,N_6804,N_8309);
nand U12377 (N_12377,N_8955,N_7539);
or U12378 (N_12378,N_5261,N_6840);
nor U12379 (N_12379,N_6862,N_8859);
xnor U12380 (N_12380,N_5278,N_8499);
or U12381 (N_12381,N_8360,N_6556);
and U12382 (N_12382,N_8395,N_8383);
or U12383 (N_12383,N_7597,N_6899);
xnor U12384 (N_12384,N_9707,N_8579);
nor U12385 (N_12385,N_8977,N_9700);
or U12386 (N_12386,N_9846,N_7006);
nor U12387 (N_12387,N_8788,N_6377);
xnor U12388 (N_12388,N_5990,N_5838);
nor U12389 (N_12389,N_8852,N_9036);
xor U12390 (N_12390,N_6479,N_6835);
and U12391 (N_12391,N_8244,N_9889);
and U12392 (N_12392,N_8608,N_7054);
nor U12393 (N_12393,N_9196,N_5211);
nor U12394 (N_12394,N_6676,N_6700);
and U12395 (N_12395,N_9244,N_7841);
or U12396 (N_12396,N_5207,N_7672);
or U12397 (N_12397,N_7450,N_5482);
nand U12398 (N_12398,N_6713,N_7924);
or U12399 (N_12399,N_8457,N_8122);
and U12400 (N_12400,N_8077,N_7419);
or U12401 (N_12401,N_5985,N_6211);
xnor U12402 (N_12402,N_6711,N_7274);
or U12403 (N_12403,N_5908,N_6775);
or U12404 (N_12404,N_7623,N_7598);
xnor U12405 (N_12405,N_9400,N_7936);
or U12406 (N_12406,N_8136,N_8774);
or U12407 (N_12407,N_5529,N_8069);
nor U12408 (N_12408,N_5521,N_5928);
nand U12409 (N_12409,N_6682,N_8144);
and U12410 (N_12410,N_9443,N_9891);
nand U12411 (N_12411,N_6943,N_9065);
and U12412 (N_12412,N_9325,N_6749);
nor U12413 (N_12413,N_5712,N_9987);
nand U12414 (N_12414,N_6812,N_8382);
or U12415 (N_12415,N_7362,N_9489);
or U12416 (N_12416,N_8570,N_8453);
nor U12417 (N_12417,N_6357,N_9267);
nand U12418 (N_12418,N_8870,N_8272);
nor U12419 (N_12419,N_9260,N_5399);
nand U12420 (N_12420,N_5596,N_6123);
nor U12421 (N_12421,N_5052,N_6093);
xnor U12422 (N_12422,N_6939,N_6382);
nand U12423 (N_12423,N_8875,N_5044);
or U12424 (N_12424,N_7089,N_9049);
or U12425 (N_12425,N_7375,N_6455);
nand U12426 (N_12426,N_9182,N_6001);
nor U12427 (N_12427,N_5892,N_9195);
and U12428 (N_12428,N_7517,N_9054);
or U12429 (N_12429,N_7600,N_6653);
and U12430 (N_12430,N_6415,N_8071);
and U12431 (N_12431,N_7135,N_6960);
nor U12432 (N_12432,N_9938,N_7709);
or U12433 (N_12433,N_7642,N_9826);
or U12434 (N_12434,N_5745,N_8518);
nor U12435 (N_12435,N_9352,N_9647);
nand U12436 (N_12436,N_8411,N_8434);
nand U12437 (N_12437,N_5468,N_5135);
and U12438 (N_12438,N_5394,N_5616);
xnor U12439 (N_12439,N_5303,N_6046);
nor U12440 (N_12440,N_7886,N_8392);
and U12441 (N_12441,N_5513,N_9498);
and U12442 (N_12442,N_7989,N_7017);
nand U12443 (N_12443,N_6744,N_5201);
and U12444 (N_12444,N_5680,N_8921);
or U12445 (N_12445,N_5907,N_8741);
nand U12446 (N_12446,N_5181,N_6390);
nand U12447 (N_12447,N_9518,N_6499);
or U12448 (N_12448,N_6222,N_6270);
nor U12449 (N_12449,N_7436,N_7148);
and U12450 (N_12450,N_8594,N_9763);
or U12451 (N_12451,N_6750,N_6671);
and U12452 (N_12452,N_8026,N_8965);
and U12453 (N_12453,N_9024,N_8078);
nand U12454 (N_12454,N_6630,N_9695);
or U12455 (N_12455,N_9312,N_6473);
xor U12456 (N_12456,N_5756,N_6720);
and U12457 (N_12457,N_7291,N_8889);
or U12458 (N_12458,N_5123,N_7519);
nand U12459 (N_12459,N_8926,N_5784);
and U12460 (N_12460,N_5087,N_6126);
and U12461 (N_12461,N_9853,N_7153);
or U12462 (N_12462,N_9788,N_9843);
nor U12463 (N_12463,N_8679,N_8484);
nand U12464 (N_12464,N_5819,N_7784);
xnor U12465 (N_12465,N_6587,N_7293);
nand U12466 (N_12466,N_7631,N_6937);
xnor U12467 (N_12467,N_9528,N_9154);
nand U12468 (N_12468,N_5050,N_6534);
nor U12469 (N_12469,N_9268,N_7177);
and U12470 (N_12470,N_6190,N_5776);
and U12471 (N_12471,N_8323,N_7673);
nor U12472 (N_12472,N_6785,N_9032);
or U12473 (N_12473,N_9730,N_5939);
nor U12474 (N_12474,N_9233,N_7777);
and U12475 (N_12475,N_5010,N_5388);
nor U12476 (N_12476,N_6066,N_7759);
nor U12477 (N_12477,N_5432,N_6213);
or U12478 (N_12478,N_6612,N_8152);
xnor U12479 (N_12479,N_9706,N_9876);
xor U12480 (N_12480,N_7347,N_6795);
or U12481 (N_12481,N_6827,N_7994);
nor U12482 (N_12482,N_7198,N_9353);
and U12483 (N_12483,N_5584,N_5326);
or U12484 (N_12484,N_5043,N_9634);
and U12485 (N_12485,N_5538,N_5387);
or U12486 (N_12486,N_5103,N_9858);
or U12487 (N_12487,N_6441,N_6045);
or U12488 (N_12488,N_5328,N_5879);
or U12489 (N_12489,N_9251,N_8505);
and U12490 (N_12490,N_8235,N_8245);
xor U12491 (N_12491,N_5386,N_8845);
xor U12492 (N_12492,N_8166,N_8861);
xor U12493 (N_12493,N_7677,N_9406);
and U12494 (N_12494,N_7414,N_6535);
and U12495 (N_12495,N_9679,N_8701);
and U12496 (N_12496,N_5829,N_7126);
nand U12497 (N_12497,N_9056,N_6481);
and U12498 (N_12498,N_6138,N_7468);
nand U12499 (N_12499,N_9147,N_9384);
nor U12500 (N_12500,N_6694,N_6200);
nor U12501 (N_12501,N_8227,N_7322);
nor U12502 (N_12502,N_8543,N_6796);
nor U12503 (N_12503,N_5726,N_5152);
or U12504 (N_12504,N_6036,N_7627);
and U12505 (N_12505,N_5134,N_6116);
nor U12506 (N_12506,N_8335,N_9105);
nor U12507 (N_12507,N_7564,N_5179);
nand U12508 (N_12508,N_9370,N_9123);
nor U12509 (N_12509,N_8838,N_8707);
xnor U12510 (N_12510,N_8447,N_5193);
and U12511 (N_12511,N_6807,N_5842);
and U12512 (N_12512,N_8969,N_8640);
and U12513 (N_12513,N_5627,N_7658);
or U12514 (N_12514,N_7074,N_7299);
and U12515 (N_12515,N_9893,N_5681);
nand U12516 (N_12516,N_9163,N_6218);
nor U12517 (N_12517,N_5841,N_8426);
and U12518 (N_12518,N_8936,N_7329);
or U12519 (N_12519,N_8548,N_9314);
nor U12520 (N_12520,N_8159,N_5873);
and U12521 (N_12521,N_8743,N_5019);
xor U12522 (N_12522,N_5043,N_5917);
and U12523 (N_12523,N_6933,N_7737);
xnor U12524 (N_12524,N_8140,N_9606);
and U12525 (N_12525,N_6782,N_8696);
xnor U12526 (N_12526,N_7152,N_9289);
and U12527 (N_12527,N_5844,N_5320);
nand U12528 (N_12528,N_9750,N_9929);
and U12529 (N_12529,N_5456,N_5027);
nor U12530 (N_12530,N_7374,N_7251);
or U12531 (N_12531,N_6043,N_5149);
nor U12532 (N_12532,N_5328,N_5005);
or U12533 (N_12533,N_5428,N_7287);
and U12534 (N_12534,N_7745,N_8240);
nor U12535 (N_12535,N_8506,N_6977);
nand U12536 (N_12536,N_5799,N_6492);
or U12537 (N_12537,N_6596,N_9524);
nand U12538 (N_12538,N_9721,N_6741);
or U12539 (N_12539,N_5301,N_8878);
xor U12540 (N_12540,N_6521,N_9041);
and U12541 (N_12541,N_9090,N_7893);
xnor U12542 (N_12542,N_9207,N_7496);
or U12543 (N_12543,N_5589,N_8336);
and U12544 (N_12544,N_7656,N_8602);
or U12545 (N_12545,N_9360,N_8343);
nor U12546 (N_12546,N_9206,N_5338);
nor U12547 (N_12547,N_8654,N_9247);
nand U12548 (N_12548,N_6518,N_6378);
or U12549 (N_12549,N_8712,N_7083);
or U12550 (N_12550,N_5801,N_8670);
or U12551 (N_12551,N_6540,N_8214);
and U12552 (N_12552,N_5443,N_6404);
and U12553 (N_12553,N_6065,N_7239);
nor U12554 (N_12554,N_9295,N_9762);
nor U12555 (N_12555,N_8728,N_7656);
and U12556 (N_12556,N_8988,N_8701);
or U12557 (N_12557,N_9413,N_8834);
and U12558 (N_12558,N_8770,N_6217);
nand U12559 (N_12559,N_6727,N_7451);
and U12560 (N_12560,N_9452,N_7662);
nand U12561 (N_12561,N_7508,N_5698);
or U12562 (N_12562,N_9514,N_9415);
nand U12563 (N_12563,N_7119,N_7248);
and U12564 (N_12564,N_9061,N_7777);
and U12565 (N_12565,N_8532,N_9885);
or U12566 (N_12566,N_8402,N_9862);
or U12567 (N_12567,N_8048,N_5953);
nor U12568 (N_12568,N_7422,N_6698);
nor U12569 (N_12569,N_7563,N_8277);
xnor U12570 (N_12570,N_9582,N_5812);
or U12571 (N_12571,N_7403,N_7883);
nand U12572 (N_12572,N_9190,N_6587);
xnor U12573 (N_12573,N_6650,N_9628);
nand U12574 (N_12574,N_9876,N_9065);
or U12575 (N_12575,N_7938,N_6726);
nor U12576 (N_12576,N_7409,N_7351);
nand U12577 (N_12577,N_5756,N_5556);
or U12578 (N_12578,N_9058,N_7883);
nor U12579 (N_12579,N_5400,N_7931);
xnor U12580 (N_12580,N_6601,N_8756);
xor U12581 (N_12581,N_6564,N_9464);
and U12582 (N_12582,N_5999,N_6521);
or U12583 (N_12583,N_6621,N_5957);
nor U12584 (N_12584,N_7233,N_8702);
or U12585 (N_12585,N_8690,N_5841);
and U12586 (N_12586,N_9883,N_8326);
nand U12587 (N_12587,N_8493,N_9240);
and U12588 (N_12588,N_5686,N_7933);
nor U12589 (N_12589,N_8064,N_9542);
nand U12590 (N_12590,N_9043,N_7266);
nor U12591 (N_12591,N_7661,N_6096);
and U12592 (N_12592,N_5606,N_8457);
or U12593 (N_12593,N_7514,N_5385);
or U12594 (N_12594,N_5364,N_6260);
nand U12595 (N_12595,N_7925,N_6624);
nand U12596 (N_12596,N_9018,N_7279);
or U12597 (N_12597,N_6047,N_8927);
nor U12598 (N_12598,N_5829,N_5421);
or U12599 (N_12599,N_8974,N_5020);
or U12600 (N_12600,N_6498,N_5523);
xnor U12601 (N_12601,N_6969,N_8307);
and U12602 (N_12602,N_8601,N_9276);
nor U12603 (N_12603,N_8496,N_7745);
nand U12604 (N_12604,N_7126,N_8730);
or U12605 (N_12605,N_5745,N_5466);
nor U12606 (N_12606,N_8621,N_9821);
or U12607 (N_12607,N_5533,N_7320);
or U12608 (N_12608,N_9175,N_6793);
nor U12609 (N_12609,N_9429,N_6258);
nor U12610 (N_12610,N_5727,N_8614);
or U12611 (N_12611,N_5398,N_9559);
or U12612 (N_12612,N_6259,N_6675);
or U12613 (N_12613,N_7442,N_6649);
xnor U12614 (N_12614,N_9009,N_8632);
nor U12615 (N_12615,N_6303,N_5312);
nand U12616 (N_12616,N_6418,N_9848);
or U12617 (N_12617,N_6882,N_9121);
xor U12618 (N_12618,N_7530,N_7697);
or U12619 (N_12619,N_6269,N_6929);
or U12620 (N_12620,N_6759,N_7051);
nor U12621 (N_12621,N_5466,N_8532);
nand U12622 (N_12622,N_5910,N_8020);
and U12623 (N_12623,N_7120,N_6256);
and U12624 (N_12624,N_7566,N_9012);
xnor U12625 (N_12625,N_5513,N_8123);
nand U12626 (N_12626,N_5827,N_7370);
nor U12627 (N_12627,N_9258,N_9225);
or U12628 (N_12628,N_9517,N_7246);
nor U12629 (N_12629,N_9529,N_5259);
nand U12630 (N_12630,N_8450,N_5077);
or U12631 (N_12631,N_5007,N_9595);
nand U12632 (N_12632,N_6801,N_9681);
and U12633 (N_12633,N_5572,N_7421);
nor U12634 (N_12634,N_8497,N_5290);
or U12635 (N_12635,N_7033,N_6436);
xnor U12636 (N_12636,N_5271,N_5736);
nor U12637 (N_12637,N_8484,N_9344);
and U12638 (N_12638,N_8287,N_7355);
nand U12639 (N_12639,N_6384,N_5099);
or U12640 (N_12640,N_5428,N_9913);
nand U12641 (N_12641,N_7804,N_9084);
nand U12642 (N_12642,N_6764,N_7613);
nand U12643 (N_12643,N_8800,N_7758);
and U12644 (N_12644,N_6046,N_7433);
nor U12645 (N_12645,N_7049,N_5502);
nand U12646 (N_12646,N_5598,N_6665);
nand U12647 (N_12647,N_6734,N_6380);
nor U12648 (N_12648,N_7546,N_6122);
xnor U12649 (N_12649,N_6861,N_5558);
xnor U12650 (N_12650,N_8192,N_7709);
or U12651 (N_12651,N_9384,N_9325);
or U12652 (N_12652,N_8612,N_8825);
or U12653 (N_12653,N_8598,N_7303);
or U12654 (N_12654,N_9834,N_5261);
nand U12655 (N_12655,N_9055,N_6066);
and U12656 (N_12656,N_6834,N_9560);
xnor U12657 (N_12657,N_8418,N_5904);
nand U12658 (N_12658,N_9002,N_7321);
nand U12659 (N_12659,N_7812,N_5494);
or U12660 (N_12660,N_5551,N_6281);
nor U12661 (N_12661,N_8473,N_7317);
and U12662 (N_12662,N_7715,N_9671);
and U12663 (N_12663,N_5226,N_5159);
xor U12664 (N_12664,N_5661,N_6236);
xnor U12665 (N_12665,N_9199,N_8432);
and U12666 (N_12666,N_5244,N_6886);
nand U12667 (N_12667,N_6003,N_8143);
and U12668 (N_12668,N_9619,N_5895);
nand U12669 (N_12669,N_5845,N_7579);
or U12670 (N_12670,N_7579,N_9544);
nand U12671 (N_12671,N_6052,N_5372);
or U12672 (N_12672,N_7673,N_6646);
nand U12673 (N_12673,N_7114,N_7448);
nand U12674 (N_12674,N_6964,N_7248);
or U12675 (N_12675,N_5034,N_6813);
nand U12676 (N_12676,N_9331,N_7343);
or U12677 (N_12677,N_6689,N_5878);
nand U12678 (N_12678,N_8088,N_5941);
and U12679 (N_12679,N_8990,N_9693);
nor U12680 (N_12680,N_7812,N_5968);
nand U12681 (N_12681,N_8610,N_5926);
and U12682 (N_12682,N_7544,N_6259);
and U12683 (N_12683,N_5272,N_5346);
or U12684 (N_12684,N_7310,N_7426);
nor U12685 (N_12685,N_8885,N_7590);
nor U12686 (N_12686,N_9386,N_9717);
nand U12687 (N_12687,N_9105,N_5392);
nand U12688 (N_12688,N_8948,N_9050);
and U12689 (N_12689,N_5859,N_5984);
nor U12690 (N_12690,N_7032,N_5481);
xnor U12691 (N_12691,N_9570,N_5541);
nand U12692 (N_12692,N_5411,N_7807);
or U12693 (N_12693,N_7396,N_7135);
xor U12694 (N_12694,N_8726,N_5784);
nor U12695 (N_12695,N_7946,N_6664);
xor U12696 (N_12696,N_5395,N_9425);
nor U12697 (N_12697,N_7453,N_5393);
or U12698 (N_12698,N_7263,N_7726);
and U12699 (N_12699,N_9770,N_9134);
nand U12700 (N_12700,N_5937,N_5245);
xor U12701 (N_12701,N_5191,N_5149);
nor U12702 (N_12702,N_9921,N_7718);
nor U12703 (N_12703,N_9091,N_5707);
or U12704 (N_12704,N_9932,N_5512);
nand U12705 (N_12705,N_6246,N_8123);
xor U12706 (N_12706,N_7718,N_9619);
nor U12707 (N_12707,N_5078,N_5561);
and U12708 (N_12708,N_5804,N_6085);
nor U12709 (N_12709,N_8121,N_7529);
nand U12710 (N_12710,N_6991,N_6115);
nor U12711 (N_12711,N_6539,N_5491);
nor U12712 (N_12712,N_6812,N_5237);
or U12713 (N_12713,N_6437,N_7635);
and U12714 (N_12714,N_6253,N_9702);
or U12715 (N_12715,N_7637,N_9255);
and U12716 (N_12716,N_9754,N_5995);
and U12717 (N_12717,N_8460,N_7874);
nand U12718 (N_12718,N_7145,N_6101);
and U12719 (N_12719,N_5765,N_7464);
nand U12720 (N_12720,N_6680,N_7683);
nor U12721 (N_12721,N_7889,N_7888);
nor U12722 (N_12722,N_6235,N_9267);
nor U12723 (N_12723,N_9788,N_8546);
or U12724 (N_12724,N_6698,N_8718);
or U12725 (N_12725,N_5373,N_6438);
nor U12726 (N_12726,N_9845,N_5332);
and U12727 (N_12727,N_9223,N_5941);
nor U12728 (N_12728,N_7673,N_9049);
nand U12729 (N_12729,N_5986,N_7691);
nor U12730 (N_12730,N_6217,N_9099);
nor U12731 (N_12731,N_9411,N_5627);
or U12732 (N_12732,N_5575,N_5096);
or U12733 (N_12733,N_8935,N_7930);
or U12734 (N_12734,N_6650,N_7013);
and U12735 (N_12735,N_5386,N_9634);
and U12736 (N_12736,N_6544,N_6402);
nand U12737 (N_12737,N_7326,N_5899);
nand U12738 (N_12738,N_8066,N_8170);
nand U12739 (N_12739,N_5673,N_9199);
nor U12740 (N_12740,N_6898,N_6161);
nor U12741 (N_12741,N_7241,N_8354);
nor U12742 (N_12742,N_7943,N_5755);
nor U12743 (N_12743,N_7666,N_6432);
and U12744 (N_12744,N_9932,N_9083);
nor U12745 (N_12745,N_9447,N_7513);
or U12746 (N_12746,N_8454,N_9396);
and U12747 (N_12747,N_8452,N_8441);
nor U12748 (N_12748,N_7808,N_9484);
or U12749 (N_12749,N_5931,N_8443);
xnor U12750 (N_12750,N_6905,N_9908);
or U12751 (N_12751,N_9273,N_9535);
nor U12752 (N_12752,N_9384,N_8911);
and U12753 (N_12753,N_9357,N_5539);
nand U12754 (N_12754,N_7705,N_7337);
nand U12755 (N_12755,N_9084,N_5206);
nor U12756 (N_12756,N_7116,N_7768);
nor U12757 (N_12757,N_5723,N_8874);
nand U12758 (N_12758,N_7390,N_8009);
nor U12759 (N_12759,N_5881,N_8611);
nand U12760 (N_12760,N_5948,N_7197);
nand U12761 (N_12761,N_6149,N_7103);
and U12762 (N_12762,N_5450,N_5435);
and U12763 (N_12763,N_7122,N_8267);
nor U12764 (N_12764,N_9186,N_5538);
nor U12765 (N_12765,N_8603,N_5023);
or U12766 (N_12766,N_6804,N_5680);
nand U12767 (N_12767,N_5430,N_5201);
or U12768 (N_12768,N_8275,N_5756);
or U12769 (N_12769,N_8454,N_7128);
nand U12770 (N_12770,N_7809,N_6470);
nor U12771 (N_12771,N_7586,N_9472);
or U12772 (N_12772,N_5064,N_9046);
or U12773 (N_12773,N_6156,N_9779);
xor U12774 (N_12774,N_9658,N_6313);
or U12775 (N_12775,N_9252,N_5550);
nand U12776 (N_12776,N_8794,N_7721);
nor U12777 (N_12777,N_8012,N_6582);
nor U12778 (N_12778,N_6854,N_7121);
nand U12779 (N_12779,N_9877,N_5385);
nor U12780 (N_12780,N_5106,N_9279);
and U12781 (N_12781,N_7253,N_8708);
xor U12782 (N_12782,N_7603,N_7578);
xor U12783 (N_12783,N_9806,N_7325);
or U12784 (N_12784,N_5374,N_6591);
nor U12785 (N_12785,N_9118,N_5499);
or U12786 (N_12786,N_7481,N_9441);
or U12787 (N_12787,N_5635,N_7469);
or U12788 (N_12788,N_8185,N_5223);
nand U12789 (N_12789,N_7051,N_6785);
nor U12790 (N_12790,N_7695,N_5918);
or U12791 (N_12791,N_5013,N_7829);
nor U12792 (N_12792,N_6124,N_8688);
or U12793 (N_12793,N_9042,N_7486);
nor U12794 (N_12794,N_6475,N_9699);
or U12795 (N_12795,N_8287,N_9866);
nand U12796 (N_12796,N_8981,N_8505);
or U12797 (N_12797,N_6888,N_7434);
nor U12798 (N_12798,N_6020,N_5243);
nor U12799 (N_12799,N_6350,N_6794);
or U12800 (N_12800,N_8825,N_6947);
nor U12801 (N_12801,N_9988,N_6558);
and U12802 (N_12802,N_9227,N_9607);
or U12803 (N_12803,N_5977,N_8714);
nor U12804 (N_12804,N_6913,N_5367);
nand U12805 (N_12805,N_9761,N_6036);
nand U12806 (N_12806,N_7788,N_8553);
nor U12807 (N_12807,N_6002,N_7999);
and U12808 (N_12808,N_5649,N_7022);
nor U12809 (N_12809,N_9209,N_6476);
or U12810 (N_12810,N_6848,N_5817);
or U12811 (N_12811,N_8849,N_9929);
nor U12812 (N_12812,N_7948,N_5196);
nor U12813 (N_12813,N_9908,N_6418);
or U12814 (N_12814,N_6523,N_7673);
and U12815 (N_12815,N_5669,N_8009);
or U12816 (N_12816,N_9480,N_8041);
nor U12817 (N_12817,N_8001,N_8529);
nor U12818 (N_12818,N_9274,N_6213);
nor U12819 (N_12819,N_7548,N_8793);
nor U12820 (N_12820,N_6404,N_6684);
nor U12821 (N_12821,N_6861,N_9434);
nand U12822 (N_12822,N_6239,N_5052);
xnor U12823 (N_12823,N_5225,N_8178);
nand U12824 (N_12824,N_5981,N_6814);
or U12825 (N_12825,N_5974,N_7517);
xor U12826 (N_12826,N_7050,N_9232);
and U12827 (N_12827,N_5665,N_5239);
nand U12828 (N_12828,N_9155,N_9305);
xor U12829 (N_12829,N_5435,N_5818);
and U12830 (N_12830,N_5429,N_6143);
and U12831 (N_12831,N_5080,N_7658);
xor U12832 (N_12832,N_8553,N_9750);
and U12833 (N_12833,N_9485,N_5486);
nand U12834 (N_12834,N_6581,N_6126);
and U12835 (N_12835,N_7899,N_9708);
nor U12836 (N_12836,N_5404,N_6421);
nand U12837 (N_12837,N_8221,N_5071);
or U12838 (N_12838,N_7791,N_8161);
and U12839 (N_12839,N_6931,N_6173);
or U12840 (N_12840,N_8119,N_5627);
nand U12841 (N_12841,N_9266,N_5096);
nor U12842 (N_12842,N_5202,N_6471);
nor U12843 (N_12843,N_5985,N_7774);
nand U12844 (N_12844,N_8321,N_7023);
or U12845 (N_12845,N_8287,N_8451);
or U12846 (N_12846,N_9941,N_7780);
and U12847 (N_12847,N_8494,N_9015);
nor U12848 (N_12848,N_6994,N_8542);
or U12849 (N_12849,N_6768,N_9359);
xor U12850 (N_12850,N_7280,N_9971);
and U12851 (N_12851,N_9203,N_5576);
or U12852 (N_12852,N_5515,N_5815);
xnor U12853 (N_12853,N_9760,N_7901);
or U12854 (N_12854,N_6082,N_8204);
and U12855 (N_12855,N_6335,N_6836);
nor U12856 (N_12856,N_6583,N_9537);
nor U12857 (N_12857,N_5301,N_6055);
and U12858 (N_12858,N_9853,N_7137);
and U12859 (N_12859,N_7572,N_7706);
nand U12860 (N_12860,N_5717,N_5070);
xor U12861 (N_12861,N_7503,N_8057);
nand U12862 (N_12862,N_7331,N_5184);
nor U12863 (N_12863,N_8100,N_7893);
and U12864 (N_12864,N_6933,N_6726);
and U12865 (N_12865,N_5678,N_6045);
or U12866 (N_12866,N_5525,N_9067);
nand U12867 (N_12867,N_6275,N_5371);
nor U12868 (N_12868,N_5291,N_6206);
nor U12869 (N_12869,N_9424,N_8615);
nor U12870 (N_12870,N_5581,N_6167);
nor U12871 (N_12871,N_8647,N_6026);
nor U12872 (N_12872,N_7727,N_7089);
and U12873 (N_12873,N_9684,N_5091);
xor U12874 (N_12874,N_8719,N_9715);
xor U12875 (N_12875,N_8730,N_5187);
and U12876 (N_12876,N_8003,N_5622);
or U12877 (N_12877,N_8492,N_9343);
and U12878 (N_12878,N_6878,N_9343);
or U12879 (N_12879,N_5278,N_9973);
or U12880 (N_12880,N_8024,N_8077);
and U12881 (N_12881,N_9483,N_5008);
nor U12882 (N_12882,N_6571,N_9969);
nand U12883 (N_12883,N_9059,N_8930);
nand U12884 (N_12884,N_7985,N_8627);
and U12885 (N_12885,N_8725,N_8643);
or U12886 (N_12886,N_8821,N_9551);
nor U12887 (N_12887,N_5705,N_6474);
nor U12888 (N_12888,N_6127,N_8523);
or U12889 (N_12889,N_8348,N_7785);
xor U12890 (N_12890,N_7281,N_7943);
xor U12891 (N_12891,N_6917,N_9163);
and U12892 (N_12892,N_7093,N_6976);
nor U12893 (N_12893,N_9520,N_8566);
nor U12894 (N_12894,N_6188,N_5760);
xor U12895 (N_12895,N_9332,N_9231);
and U12896 (N_12896,N_6644,N_6297);
or U12897 (N_12897,N_9174,N_8461);
nor U12898 (N_12898,N_5232,N_6983);
nor U12899 (N_12899,N_8821,N_9396);
nor U12900 (N_12900,N_8136,N_7825);
or U12901 (N_12901,N_8620,N_5505);
xnor U12902 (N_12902,N_8830,N_6194);
or U12903 (N_12903,N_6875,N_5264);
nor U12904 (N_12904,N_7978,N_7913);
and U12905 (N_12905,N_5742,N_5952);
or U12906 (N_12906,N_7169,N_9189);
nor U12907 (N_12907,N_7453,N_9870);
or U12908 (N_12908,N_8824,N_5672);
nor U12909 (N_12909,N_8843,N_9279);
nand U12910 (N_12910,N_9214,N_8738);
or U12911 (N_12911,N_8083,N_9182);
nor U12912 (N_12912,N_7621,N_8433);
and U12913 (N_12913,N_9421,N_9610);
nand U12914 (N_12914,N_9932,N_9092);
nand U12915 (N_12915,N_5587,N_5267);
or U12916 (N_12916,N_7127,N_7541);
nand U12917 (N_12917,N_7851,N_9570);
or U12918 (N_12918,N_9231,N_7184);
nor U12919 (N_12919,N_8427,N_6562);
nor U12920 (N_12920,N_7788,N_5273);
and U12921 (N_12921,N_6821,N_5539);
nor U12922 (N_12922,N_9367,N_7765);
nor U12923 (N_12923,N_9601,N_6837);
nor U12924 (N_12924,N_7554,N_9428);
or U12925 (N_12925,N_7094,N_9629);
nor U12926 (N_12926,N_6473,N_9690);
nand U12927 (N_12927,N_6295,N_6451);
xnor U12928 (N_12928,N_9345,N_8167);
nand U12929 (N_12929,N_6417,N_8644);
or U12930 (N_12930,N_7720,N_7208);
xnor U12931 (N_12931,N_6340,N_5690);
nor U12932 (N_12932,N_8379,N_9854);
nand U12933 (N_12933,N_8979,N_7948);
nand U12934 (N_12934,N_6770,N_9989);
or U12935 (N_12935,N_7130,N_7893);
or U12936 (N_12936,N_6510,N_9438);
nand U12937 (N_12937,N_9793,N_6767);
nor U12938 (N_12938,N_5360,N_5528);
nand U12939 (N_12939,N_9126,N_8263);
nor U12940 (N_12940,N_5486,N_6051);
and U12941 (N_12941,N_9534,N_7794);
and U12942 (N_12942,N_7539,N_7816);
and U12943 (N_12943,N_8097,N_7855);
nor U12944 (N_12944,N_8039,N_5660);
nand U12945 (N_12945,N_8821,N_9339);
nor U12946 (N_12946,N_9026,N_9627);
nand U12947 (N_12947,N_9871,N_8754);
and U12948 (N_12948,N_5972,N_9374);
and U12949 (N_12949,N_9234,N_7317);
and U12950 (N_12950,N_9874,N_7988);
and U12951 (N_12951,N_7630,N_7727);
and U12952 (N_12952,N_8793,N_5456);
and U12953 (N_12953,N_8882,N_9755);
xor U12954 (N_12954,N_7757,N_8427);
nand U12955 (N_12955,N_5520,N_7242);
nand U12956 (N_12956,N_9208,N_9264);
nor U12957 (N_12957,N_5074,N_7364);
nand U12958 (N_12958,N_8774,N_6690);
nor U12959 (N_12959,N_5542,N_9083);
nor U12960 (N_12960,N_8466,N_8707);
nand U12961 (N_12961,N_9763,N_8546);
and U12962 (N_12962,N_6297,N_6107);
or U12963 (N_12963,N_8894,N_6799);
nor U12964 (N_12964,N_9058,N_7128);
nand U12965 (N_12965,N_5890,N_8153);
and U12966 (N_12966,N_7931,N_9667);
nor U12967 (N_12967,N_9344,N_9508);
or U12968 (N_12968,N_8334,N_7708);
xnor U12969 (N_12969,N_6244,N_9049);
nor U12970 (N_12970,N_7852,N_7191);
nand U12971 (N_12971,N_8424,N_9725);
nor U12972 (N_12972,N_9959,N_7522);
and U12973 (N_12973,N_7124,N_5074);
xor U12974 (N_12974,N_6081,N_6375);
and U12975 (N_12975,N_8708,N_6248);
or U12976 (N_12976,N_6708,N_6877);
nor U12977 (N_12977,N_7356,N_9732);
or U12978 (N_12978,N_8498,N_6021);
xnor U12979 (N_12979,N_8590,N_9192);
or U12980 (N_12980,N_6061,N_5499);
and U12981 (N_12981,N_9870,N_7478);
nor U12982 (N_12982,N_8494,N_5958);
and U12983 (N_12983,N_5681,N_6379);
and U12984 (N_12984,N_9043,N_9890);
nor U12985 (N_12985,N_7173,N_5027);
and U12986 (N_12986,N_8827,N_8085);
and U12987 (N_12987,N_7414,N_9132);
nand U12988 (N_12988,N_9876,N_5262);
and U12989 (N_12989,N_6585,N_6118);
and U12990 (N_12990,N_9928,N_8004);
nor U12991 (N_12991,N_8041,N_7367);
nand U12992 (N_12992,N_7800,N_8690);
xor U12993 (N_12993,N_8806,N_5440);
and U12994 (N_12994,N_7218,N_6280);
nand U12995 (N_12995,N_9579,N_5607);
xnor U12996 (N_12996,N_7452,N_9400);
or U12997 (N_12997,N_9913,N_9270);
or U12998 (N_12998,N_8517,N_5367);
nand U12999 (N_12999,N_8571,N_9339);
or U13000 (N_13000,N_6802,N_9009);
nor U13001 (N_13001,N_6688,N_8825);
nand U13002 (N_13002,N_5638,N_8569);
nor U13003 (N_13003,N_9574,N_5329);
nor U13004 (N_13004,N_9437,N_9854);
nand U13005 (N_13005,N_5368,N_6164);
or U13006 (N_13006,N_7721,N_8433);
nor U13007 (N_13007,N_9106,N_5691);
or U13008 (N_13008,N_6237,N_9965);
nor U13009 (N_13009,N_7988,N_6011);
nand U13010 (N_13010,N_5875,N_8023);
and U13011 (N_13011,N_5450,N_7903);
and U13012 (N_13012,N_6732,N_5381);
and U13013 (N_13013,N_5656,N_8107);
or U13014 (N_13014,N_5052,N_5377);
nand U13015 (N_13015,N_5154,N_6146);
and U13016 (N_13016,N_6947,N_6545);
or U13017 (N_13017,N_9343,N_6276);
nor U13018 (N_13018,N_7653,N_9679);
nor U13019 (N_13019,N_7820,N_9152);
or U13020 (N_13020,N_7987,N_6938);
nor U13021 (N_13021,N_7340,N_9754);
nand U13022 (N_13022,N_5630,N_6460);
and U13023 (N_13023,N_8257,N_9032);
nor U13024 (N_13024,N_9273,N_6807);
nor U13025 (N_13025,N_7179,N_8783);
and U13026 (N_13026,N_5945,N_7769);
nand U13027 (N_13027,N_8249,N_8910);
or U13028 (N_13028,N_9208,N_7128);
and U13029 (N_13029,N_5245,N_6808);
and U13030 (N_13030,N_8565,N_5549);
or U13031 (N_13031,N_6609,N_6378);
nand U13032 (N_13032,N_7244,N_5388);
xnor U13033 (N_13033,N_8755,N_8922);
nor U13034 (N_13034,N_7615,N_9469);
or U13035 (N_13035,N_5547,N_9558);
nor U13036 (N_13036,N_5463,N_9414);
xor U13037 (N_13037,N_7350,N_9691);
nand U13038 (N_13038,N_7742,N_5671);
nand U13039 (N_13039,N_6871,N_7444);
nor U13040 (N_13040,N_5940,N_5419);
and U13041 (N_13041,N_9011,N_7357);
nor U13042 (N_13042,N_8058,N_8686);
xnor U13043 (N_13043,N_6073,N_9648);
nand U13044 (N_13044,N_8003,N_8080);
or U13045 (N_13045,N_5259,N_5219);
and U13046 (N_13046,N_8462,N_7818);
nor U13047 (N_13047,N_6921,N_8921);
or U13048 (N_13048,N_8482,N_7001);
and U13049 (N_13049,N_7178,N_6885);
or U13050 (N_13050,N_7369,N_7552);
or U13051 (N_13051,N_8213,N_7956);
nor U13052 (N_13052,N_7865,N_6782);
nor U13053 (N_13053,N_8019,N_5461);
xor U13054 (N_13054,N_8223,N_8573);
nor U13055 (N_13055,N_6659,N_5886);
nand U13056 (N_13056,N_9631,N_5838);
and U13057 (N_13057,N_8217,N_5520);
or U13058 (N_13058,N_5622,N_8239);
or U13059 (N_13059,N_8192,N_7269);
xnor U13060 (N_13060,N_7534,N_7347);
nor U13061 (N_13061,N_8317,N_8478);
nand U13062 (N_13062,N_9486,N_8178);
xor U13063 (N_13063,N_6979,N_7439);
or U13064 (N_13064,N_6465,N_7411);
and U13065 (N_13065,N_5736,N_7178);
nor U13066 (N_13066,N_9332,N_5861);
nor U13067 (N_13067,N_5110,N_7639);
nand U13068 (N_13068,N_6778,N_5219);
nand U13069 (N_13069,N_8136,N_6958);
nand U13070 (N_13070,N_9158,N_8088);
and U13071 (N_13071,N_6267,N_8381);
and U13072 (N_13072,N_6324,N_9502);
and U13073 (N_13073,N_7552,N_9730);
nand U13074 (N_13074,N_8821,N_6455);
nor U13075 (N_13075,N_8727,N_7358);
or U13076 (N_13076,N_7404,N_9236);
or U13077 (N_13077,N_6645,N_5143);
nand U13078 (N_13078,N_7668,N_7576);
nand U13079 (N_13079,N_6963,N_5449);
and U13080 (N_13080,N_8196,N_6028);
xor U13081 (N_13081,N_9134,N_9029);
or U13082 (N_13082,N_5948,N_5875);
and U13083 (N_13083,N_9772,N_9880);
and U13084 (N_13084,N_8767,N_9277);
nor U13085 (N_13085,N_6284,N_5354);
and U13086 (N_13086,N_7164,N_5086);
nand U13087 (N_13087,N_7374,N_5017);
nand U13088 (N_13088,N_6255,N_9954);
nor U13089 (N_13089,N_6096,N_6913);
nor U13090 (N_13090,N_6221,N_5560);
nand U13091 (N_13091,N_9696,N_8152);
nor U13092 (N_13092,N_6545,N_6387);
and U13093 (N_13093,N_9513,N_5383);
or U13094 (N_13094,N_9881,N_8280);
nor U13095 (N_13095,N_8752,N_8985);
nor U13096 (N_13096,N_7363,N_8973);
or U13097 (N_13097,N_6245,N_9216);
nand U13098 (N_13098,N_5435,N_8157);
or U13099 (N_13099,N_9750,N_8518);
nor U13100 (N_13100,N_6023,N_8655);
or U13101 (N_13101,N_7994,N_9358);
and U13102 (N_13102,N_6673,N_6283);
and U13103 (N_13103,N_6608,N_9482);
nor U13104 (N_13104,N_8074,N_6387);
or U13105 (N_13105,N_6763,N_6044);
or U13106 (N_13106,N_9496,N_8965);
nand U13107 (N_13107,N_5096,N_6181);
or U13108 (N_13108,N_8937,N_8822);
xor U13109 (N_13109,N_9681,N_8950);
xnor U13110 (N_13110,N_6363,N_6550);
and U13111 (N_13111,N_5707,N_9677);
or U13112 (N_13112,N_7860,N_9002);
or U13113 (N_13113,N_8668,N_6753);
and U13114 (N_13114,N_6919,N_5071);
nand U13115 (N_13115,N_7137,N_8810);
xnor U13116 (N_13116,N_6120,N_6613);
or U13117 (N_13117,N_8190,N_6770);
nor U13118 (N_13118,N_9393,N_6850);
and U13119 (N_13119,N_5765,N_5584);
nor U13120 (N_13120,N_8494,N_8216);
or U13121 (N_13121,N_6166,N_7568);
nor U13122 (N_13122,N_7012,N_9683);
and U13123 (N_13123,N_5535,N_8353);
nor U13124 (N_13124,N_9212,N_6530);
and U13125 (N_13125,N_8814,N_7797);
nor U13126 (N_13126,N_7532,N_6725);
nand U13127 (N_13127,N_8814,N_9518);
nand U13128 (N_13128,N_7479,N_8077);
nor U13129 (N_13129,N_5112,N_6972);
and U13130 (N_13130,N_6641,N_8943);
nor U13131 (N_13131,N_8914,N_6929);
nand U13132 (N_13132,N_5036,N_7869);
nor U13133 (N_13133,N_7886,N_9858);
or U13134 (N_13134,N_9999,N_7518);
xor U13135 (N_13135,N_6360,N_6327);
and U13136 (N_13136,N_5828,N_6935);
and U13137 (N_13137,N_9769,N_7012);
or U13138 (N_13138,N_9762,N_8151);
or U13139 (N_13139,N_8921,N_9783);
nand U13140 (N_13140,N_7461,N_7068);
or U13141 (N_13141,N_8246,N_7210);
nor U13142 (N_13142,N_5470,N_5528);
xnor U13143 (N_13143,N_7288,N_6984);
nor U13144 (N_13144,N_8189,N_7902);
or U13145 (N_13145,N_6329,N_6053);
nor U13146 (N_13146,N_8003,N_7291);
or U13147 (N_13147,N_6531,N_8421);
xnor U13148 (N_13148,N_5862,N_6847);
nor U13149 (N_13149,N_8099,N_8432);
or U13150 (N_13150,N_5731,N_7659);
nand U13151 (N_13151,N_5364,N_9920);
or U13152 (N_13152,N_8916,N_5738);
or U13153 (N_13153,N_9969,N_8641);
nor U13154 (N_13154,N_9830,N_6253);
xnor U13155 (N_13155,N_6105,N_7243);
or U13156 (N_13156,N_9564,N_7484);
and U13157 (N_13157,N_5897,N_5600);
or U13158 (N_13158,N_6006,N_5299);
nand U13159 (N_13159,N_5980,N_8197);
or U13160 (N_13160,N_5747,N_7667);
nand U13161 (N_13161,N_7426,N_6928);
xnor U13162 (N_13162,N_6067,N_8316);
or U13163 (N_13163,N_6754,N_7226);
nor U13164 (N_13164,N_8038,N_7427);
xnor U13165 (N_13165,N_7296,N_6331);
nand U13166 (N_13166,N_8130,N_5364);
nand U13167 (N_13167,N_7720,N_5376);
or U13168 (N_13168,N_8236,N_5705);
nand U13169 (N_13169,N_9586,N_8070);
nand U13170 (N_13170,N_8405,N_8982);
nor U13171 (N_13171,N_8301,N_6888);
or U13172 (N_13172,N_9637,N_9524);
nor U13173 (N_13173,N_5254,N_6236);
and U13174 (N_13174,N_8937,N_9402);
nand U13175 (N_13175,N_8807,N_6773);
and U13176 (N_13176,N_5411,N_6551);
or U13177 (N_13177,N_8651,N_5138);
nand U13178 (N_13178,N_7477,N_6021);
or U13179 (N_13179,N_7247,N_9801);
nand U13180 (N_13180,N_5121,N_7552);
or U13181 (N_13181,N_6111,N_9342);
and U13182 (N_13182,N_9740,N_8412);
nor U13183 (N_13183,N_5028,N_6897);
or U13184 (N_13184,N_9143,N_8844);
nor U13185 (N_13185,N_7569,N_8486);
nand U13186 (N_13186,N_6865,N_9028);
xnor U13187 (N_13187,N_8221,N_9697);
or U13188 (N_13188,N_8284,N_6446);
xor U13189 (N_13189,N_5210,N_7529);
or U13190 (N_13190,N_7193,N_9309);
xor U13191 (N_13191,N_5898,N_6443);
or U13192 (N_13192,N_5708,N_5131);
nand U13193 (N_13193,N_6956,N_9030);
or U13194 (N_13194,N_5473,N_5066);
or U13195 (N_13195,N_9114,N_7070);
and U13196 (N_13196,N_8441,N_9264);
and U13197 (N_13197,N_8813,N_5700);
and U13198 (N_13198,N_6987,N_7902);
xnor U13199 (N_13199,N_6589,N_6976);
nor U13200 (N_13200,N_9233,N_5530);
and U13201 (N_13201,N_7413,N_9161);
nand U13202 (N_13202,N_9018,N_5214);
and U13203 (N_13203,N_8335,N_6500);
or U13204 (N_13204,N_9229,N_8779);
nand U13205 (N_13205,N_6586,N_5491);
and U13206 (N_13206,N_5692,N_5463);
and U13207 (N_13207,N_5484,N_8771);
and U13208 (N_13208,N_7732,N_8290);
or U13209 (N_13209,N_8798,N_6417);
nor U13210 (N_13210,N_9864,N_7759);
or U13211 (N_13211,N_9896,N_6545);
nand U13212 (N_13212,N_8925,N_8681);
nand U13213 (N_13213,N_8971,N_5843);
or U13214 (N_13214,N_8651,N_6262);
nand U13215 (N_13215,N_9988,N_8701);
or U13216 (N_13216,N_5978,N_8366);
xor U13217 (N_13217,N_5999,N_5645);
and U13218 (N_13218,N_6326,N_8024);
nand U13219 (N_13219,N_9949,N_6551);
and U13220 (N_13220,N_5849,N_7164);
or U13221 (N_13221,N_6504,N_9100);
or U13222 (N_13222,N_9566,N_7154);
nor U13223 (N_13223,N_8444,N_7881);
or U13224 (N_13224,N_7483,N_8274);
xor U13225 (N_13225,N_9088,N_6893);
or U13226 (N_13226,N_6755,N_9356);
or U13227 (N_13227,N_7250,N_6504);
nor U13228 (N_13228,N_7573,N_6452);
nor U13229 (N_13229,N_9952,N_8395);
and U13230 (N_13230,N_8274,N_9374);
nor U13231 (N_13231,N_5038,N_9887);
nor U13232 (N_13232,N_7360,N_9690);
nor U13233 (N_13233,N_5456,N_5428);
or U13234 (N_13234,N_5956,N_8284);
nor U13235 (N_13235,N_9684,N_9163);
xnor U13236 (N_13236,N_6399,N_5929);
or U13237 (N_13237,N_5780,N_6885);
xnor U13238 (N_13238,N_7902,N_9936);
and U13239 (N_13239,N_6955,N_8342);
and U13240 (N_13240,N_6674,N_9647);
nand U13241 (N_13241,N_9392,N_9051);
and U13242 (N_13242,N_9461,N_6918);
xor U13243 (N_13243,N_8448,N_5126);
nand U13244 (N_13244,N_7879,N_6780);
nor U13245 (N_13245,N_7973,N_7813);
nor U13246 (N_13246,N_7243,N_9233);
or U13247 (N_13247,N_8329,N_7984);
nor U13248 (N_13248,N_7893,N_6891);
or U13249 (N_13249,N_7894,N_7717);
and U13250 (N_13250,N_7444,N_8942);
or U13251 (N_13251,N_5465,N_6015);
and U13252 (N_13252,N_9454,N_7524);
nor U13253 (N_13253,N_7015,N_8163);
and U13254 (N_13254,N_9181,N_7227);
and U13255 (N_13255,N_9356,N_9785);
nor U13256 (N_13256,N_6412,N_8312);
nor U13257 (N_13257,N_6779,N_9011);
and U13258 (N_13258,N_6697,N_7263);
nor U13259 (N_13259,N_5095,N_5594);
or U13260 (N_13260,N_6813,N_9426);
or U13261 (N_13261,N_8128,N_5742);
or U13262 (N_13262,N_8896,N_7669);
and U13263 (N_13263,N_5874,N_8473);
nand U13264 (N_13264,N_8239,N_6367);
and U13265 (N_13265,N_7605,N_9112);
nand U13266 (N_13266,N_7463,N_5448);
nor U13267 (N_13267,N_8193,N_8898);
or U13268 (N_13268,N_6532,N_6857);
nand U13269 (N_13269,N_5361,N_9301);
nand U13270 (N_13270,N_9554,N_9940);
xor U13271 (N_13271,N_6663,N_5899);
nor U13272 (N_13272,N_7996,N_7690);
nor U13273 (N_13273,N_8455,N_6201);
and U13274 (N_13274,N_5106,N_7051);
nor U13275 (N_13275,N_7471,N_8978);
and U13276 (N_13276,N_8031,N_9673);
nor U13277 (N_13277,N_8536,N_8162);
nand U13278 (N_13278,N_5236,N_7928);
nor U13279 (N_13279,N_9106,N_5588);
or U13280 (N_13280,N_6042,N_9763);
or U13281 (N_13281,N_7785,N_5067);
nand U13282 (N_13282,N_9555,N_9432);
or U13283 (N_13283,N_6805,N_7720);
nand U13284 (N_13284,N_9723,N_7307);
nand U13285 (N_13285,N_5758,N_9313);
nand U13286 (N_13286,N_5354,N_7035);
and U13287 (N_13287,N_6725,N_9599);
nand U13288 (N_13288,N_8911,N_7367);
nor U13289 (N_13289,N_6655,N_9040);
and U13290 (N_13290,N_8163,N_7550);
xnor U13291 (N_13291,N_5678,N_6063);
or U13292 (N_13292,N_9123,N_9295);
nor U13293 (N_13293,N_5376,N_6415);
or U13294 (N_13294,N_8589,N_6220);
or U13295 (N_13295,N_8867,N_8093);
nand U13296 (N_13296,N_6536,N_5977);
nor U13297 (N_13297,N_8966,N_9432);
or U13298 (N_13298,N_5433,N_9384);
nand U13299 (N_13299,N_7387,N_7806);
nand U13300 (N_13300,N_7870,N_5087);
xor U13301 (N_13301,N_8094,N_6563);
nand U13302 (N_13302,N_5266,N_7851);
and U13303 (N_13303,N_5678,N_5301);
nand U13304 (N_13304,N_7091,N_7665);
and U13305 (N_13305,N_5171,N_8091);
nand U13306 (N_13306,N_7776,N_6765);
or U13307 (N_13307,N_8411,N_7682);
nand U13308 (N_13308,N_7083,N_7156);
nor U13309 (N_13309,N_7256,N_5638);
xnor U13310 (N_13310,N_7789,N_6916);
or U13311 (N_13311,N_9091,N_5480);
nor U13312 (N_13312,N_9309,N_6585);
nor U13313 (N_13313,N_6540,N_5153);
nand U13314 (N_13314,N_6069,N_5446);
and U13315 (N_13315,N_6797,N_6193);
or U13316 (N_13316,N_9081,N_8449);
or U13317 (N_13317,N_8143,N_5072);
nand U13318 (N_13318,N_9646,N_5613);
nor U13319 (N_13319,N_9979,N_8223);
and U13320 (N_13320,N_7026,N_7656);
and U13321 (N_13321,N_8063,N_6921);
xnor U13322 (N_13322,N_6639,N_8444);
nand U13323 (N_13323,N_7309,N_7431);
nor U13324 (N_13324,N_5545,N_9068);
or U13325 (N_13325,N_7943,N_8346);
xor U13326 (N_13326,N_6006,N_5710);
or U13327 (N_13327,N_6083,N_8531);
nor U13328 (N_13328,N_7687,N_5983);
xor U13329 (N_13329,N_9292,N_6915);
and U13330 (N_13330,N_7826,N_9111);
and U13331 (N_13331,N_6478,N_8978);
nor U13332 (N_13332,N_8707,N_8580);
and U13333 (N_13333,N_6258,N_9539);
nor U13334 (N_13334,N_6354,N_9453);
nor U13335 (N_13335,N_8211,N_8367);
and U13336 (N_13336,N_9307,N_7048);
or U13337 (N_13337,N_8348,N_7076);
or U13338 (N_13338,N_9567,N_5850);
nor U13339 (N_13339,N_8194,N_6388);
nor U13340 (N_13340,N_8204,N_6066);
and U13341 (N_13341,N_8072,N_7463);
or U13342 (N_13342,N_5141,N_7418);
nor U13343 (N_13343,N_8216,N_8185);
and U13344 (N_13344,N_8051,N_7877);
or U13345 (N_13345,N_9424,N_7335);
nor U13346 (N_13346,N_6481,N_5537);
or U13347 (N_13347,N_6219,N_6070);
and U13348 (N_13348,N_8548,N_5082);
nor U13349 (N_13349,N_6548,N_9945);
nor U13350 (N_13350,N_9546,N_5864);
nor U13351 (N_13351,N_9086,N_9242);
nand U13352 (N_13352,N_6590,N_8324);
nor U13353 (N_13353,N_6724,N_7543);
or U13354 (N_13354,N_5746,N_7287);
or U13355 (N_13355,N_8084,N_6538);
nor U13356 (N_13356,N_9191,N_5339);
nor U13357 (N_13357,N_6795,N_6290);
nand U13358 (N_13358,N_8308,N_7305);
and U13359 (N_13359,N_9407,N_5312);
and U13360 (N_13360,N_5396,N_8013);
nor U13361 (N_13361,N_6886,N_9680);
or U13362 (N_13362,N_9513,N_7024);
nand U13363 (N_13363,N_6337,N_5234);
and U13364 (N_13364,N_6210,N_6164);
xnor U13365 (N_13365,N_7277,N_8599);
nor U13366 (N_13366,N_5501,N_6992);
nand U13367 (N_13367,N_7251,N_9588);
xor U13368 (N_13368,N_7292,N_7332);
nor U13369 (N_13369,N_8457,N_7492);
and U13370 (N_13370,N_8822,N_7334);
xor U13371 (N_13371,N_5986,N_8167);
and U13372 (N_13372,N_6794,N_6831);
and U13373 (N_13373,N_7758,N_8308);
and U13374 (N_13374,N_5710,N_9615);
or U13375 (N_13375,N_7400,N_5139);
xor U13376 (N_13376,N_5449,N_9382);
or U13377 (N_13377,N_7207,N_9774);
or U13378 (N_13378,N_5358,N_9116);
nand U13379 (N_13379,N_8822,N_5068);
nand U13380 (N_13380,N_8775,N_5910);
and U13381 (N_13381,N_7729,N_7297);
xnor U13382 (N_13382,N_8002,N_9402);
nor U13383 (N_13383,N_9027,N_6760);
xnor U13384 (N_13384,N_8738,N_5199);
or U13385 (N_13385,N_8375,N_5173);
and U13386 (N_13386,N_9581,N_9200);
or U13387 (N_13387,N_6634,N_6658);
nand U13388 (N_13388,N_5427,N_6659);
and U13389 (N_13389,N_8104,N_7166);
and U13390 (N_13390,N_5275,N_6007);
nor U13391 (N_13391,N_8542,N_7402);
and U13392 (N_13392,N_9027,N_7818);
and U13393 (N_13393,N_6192,N_8311);
nor U13394 (N_13394,N_6711,N_5225);
nor U13395 (N_13395,N_8747,N_7075);
nor U13396 (N_13396,N_6509,N_7798);
nand U13397 (N_13397,N_6059,N_5576);
or U13398 (N_13398,N_5924,N_9834);
and U13399 (N_13399,N_7868,N_9225);
xnor U13400 (N_13400,N_9287,N_8839);
or U13401 (N_13401,N_9408,N_6244);
or U13402 (N_13402,N_9729,N_6246);
xnor U13403 (N_13403,N_9130,N_7341);
xnor U13404 (N_13404,N_6555,N_6707);
nor U13405 (N_13405,N_8473,N_8675);
nand U13406 (N_13406,N_9576,N_9924);
nand U13407 (N_13407,N_5350,N_5906);
and U13408 (N_13408,N_7315,N_7673);
xor U13409 (N_13409,N_6169,N_8416);
nor U13410 (N_13410,N_9770,N_6698);
and U13411 (N_13411,N_8664,N_8930);
xor U13412 (N_13412,N_9832,N_7501);
xnor U13413 (N_13413,N_9121,N_7335);
nor U13414 (N_13414,N_5759,N_5610);
nor U13415 (N_13415,N_8507,N_9236);
nor U13416 (N_13416,N_6202,N_9404);
nand U13417 (N_13417,N_7165,N_6955);
and U13418 (N_13418,N_5929,N_9765);
nor U13419 (N_13419,N_5032,N_9157);
and U13420 (N_13420,N_5970,N_9324);
and U13421 (N_13421,N_8843,N_8098);
or U13422 (N_13422,N_6192,N_6760);
nor U13423 (N_13423,N_6966,N_7370);
nand U13424 (N_13424,N_9170,N_8401);
or U13425 (N_13425,N_5142,N_9969);
or U13426 (N_13426,N_7210,N_6186);
xnor U13427 (N_13427,N_8859,N_5103);
nor U13428 (N_13428,N_5353,N_7171);
or U13429 (N_13429,N_5317,N_8954);
and U13430 (N_13430,N_8042,N_8789);
or U13431 (N_13431,N_5643,N_8341);
or U13432 (N_13432,N_8796,N_9943);
nand U13433 (N_13433,N_8179,N_8999);
or U13434 (N_13434,N_5384,N_8152);
nor U13435 (N_13435,N_9728,N_9480);
or U13436 (N_13436,N_5806,N_6829);
nor U13437 (N_13437,N_8883,N_5889);
or U13438 (N_13438,N_6788,N_7124);
or U13439 (N_13439,N_7284,N_9159);
or U13440 (N_13440,N_8710,N_9063);
nand U13441 (N_13441,N_7246,N_5371);
and U13442 (N_13442,N_5484,N_5518);
xor U13443 (N_13443,N_7094,N_5143);
nand U13444 (N_13444,N_8676,N_7883);
nand U13445 (N_13445,N_9876,N_5487);
and U13446 (N_13446,N_6023,N_6469);
or U13447 (N_13447,N_7442,N_8686);
and U13448 (N_13448,N_8153,N_5933);
or U13449 (N_13449,N_9992,N_9126);
or U13450 (N_13450,N_8936,N_6082);
or U13451 (N_13451,N_9755,N_8926);
or U13452 (N_13452,N_7585,N_8009);
and U13453 (N_13453,N_9930,N_8532);
xor U13454 (N_13454,N_8677,N_6552);
nand U13455 (N_13455,N_9820,N_5581);
xnor U13456 (N_13456,N_6835,N_6246);
nor U13457 (N_13457,N_6105,N_7066);
nor U13458 (N_13458,N_9307,N_7883);
and U13459 (N_13459,N_7781,N_6290);
xor U13460 (N_13460,N_5181,N_9288);
nor U13461 (N_13461,N_6040,N_7294);
and U13462 (N_13462,N_5183,N_5450);
nor U13463 (N_13463,N_5424,N_5014);
and U13464 (N_13464,N_6214,N_6370);
nor U13465 (N_13465,N_8001,N_6753);
or U13466 (N_13466,N_5371,N_5098);
and U13467 (N_13467,N_8230,N_6212);
or U13468 (N_13468,N_6498,N_9034);
nand U13469 (N_13469,N_8330,N_6838);
and U13470 (N_13470,N_9466,N_8218);
nor U13471 (N_13471,N_7961,N_6042);
or U13472 (N_13472,N_9191,N_8928);
nor U13473 (N_13473,N_7215,N_6465);
and U13474 (N_13474,N_7944,N_5944);
nand U13475 (N_13475,N_8095,N_6800);
nor U13476 (N_13476,N_6199,N_5929);
xnor U13477 (N_13477,N_8113,N_5613);
nor U13478 (N_13478,N_8158,N_6465);
nand U13479 (N_13479,N_5899,N_8046);
nor U13480 (N_13480,N_8863,N_9792);
and U13481 (N_13481,N_5695,N_7614);
or U13482 (N_13482,N_8443,N_5975);
nand U13483 (N_13483,N_8297,N_8097);
nand U13484 (N_13484,N_7436,N_5118);
and U13485 (N_13485,N_9937,N_5323);
nor U13486 (N_13486,N_7387,N_9983);
and U13487 (N_13487,N_9525,N_5602);
or U13488 (N_13488,N_7997,N_9616);
and U13489 (N_13489,N_6781,N_6320);
nand U13490 (N_13490,N_7948,N_8614);
and U13491 (N_13491,N_8140,N_6635);
nand U13492 (N_13492,N_6515,N_6859);
nand U13493 (N_13493,N_7643,N_9242);
xor U13494 (N_13494,N_5613,N_9596);
nor U13495 (N_13495,N_8203,N_8060);
nand U13496 (N_13496,N_8312,N_8277);
and U13497 (N_13497,N_7895,N_8108);
nor U13498 (N_13498,N_5408,N_5244);
or U13499 (N_13499,N_9075,N_7044);
or U13500 (N_13500,N_8202,N_6291);
or U13501 (N_13501,N_5361,N_6641);
nand U13502 (N_13502,N_9813,N_8267);
or U13503 (N_13503,N_9770,N_6040);
nor U13504 (N_13504,N_6599,N_6602);
nor U13505 (N_13505,N_5579,N_8429);
or U13506 (N_13506,N_8822,N_9260);
nor U13507 (N_13507,N_8208,N_9853);
and U13508 (N_13508,N_5690,N_5146);
xnor U13509 (N_13509,N_7178,N_5228);
and U13510 (N_13510,N_5722,N_8126);
and U13511 (N_13511,N_8040,N_6415);
nand U13512 (N_13512,N_8744,N_9101);
nor U13513 (N_13513,N_5998,N_5568);
or U13514 (N_13514,N_6996,N_5703);
nand U13515 (N_13515,N_7839,N_8722);
nor U13516 (N_13516,N_8392,N_9268);
nor U13517 (N_13517,N_6347,N_8753);
nor U13518 (N_13518,N_9837,N_9363);
nor U13519 (N_13519,N_9077,N_8367);
and U13520 (N_13520,N_9103,N_9101);
nand U13521 (N_13521,N_8081,N_7235);
xnor U13522 (N_13522,N_6273,N_6931);
and U13523 (N_13523,N_5928,N_6920);
nor U13524 (N_13524,N_9567,N_9251);
or U13525 (N_13525,N_5918,N_9030);
nand U13526 (N_13526,N_5112,N_6904);
nand U13527 (N_13527,N_6483,N_8080);
xor U13528 (N_13528,N_9145,N_5894);
and U13529 (N_13529,N_5873,N_8486);
nor U13530 (N_13530,N_7879,N_9095);
and U13531 (N_13531,N_9706,N_7254);
nor U13532 (N_13532,N_8695,N_8872);
nor U13533 (N_13533,N_9329,N_9105);
nand U13534 (N_13534,N_8084,N_5997);
nand U13535 (N_13535,N_9866,N_6855);
nand U13536 (N_13536,N_9455,N_8488);
nand U13537 (N_13537,N_9236,N_9289);
nand U13538 (N_13538,N_6705,N_9277);
and U13539 (N_13539,N_9437,N_9827);
nor U13540 (N_13540,N_7042,N_6567);
xor U13541 (N_13541,N_7717,N_7721);
nand U13542 (N_13542,N_7474,N_5557);
or U13543 (N_13543,N_5479,N_7563);
nor U13544 (N_13544,N_8454,N_5631);
nor U13545 (N_13545,N_7283,N_7276);
nor U13546 (N_13546,N_6675,N_5853);
or U13547 (N_13547,N_9651,N_8949);
nor U13548 (N_13548,N_8082,N_6481);
and U13549 (N_13549,N_5634,N_5983);
nand U13550 (N_13550,N_6401,N_6486);
nand U13551 (N_13551,N_6006,N_8915);
and U13552 (N_13552,N_9579,N_8004);
and U13553 (N_13553,N_5264,N_7931);
xor U13554 (N_13554,N_9264,N_6637);
or U13555 (N_13555,N_5117,N_6121);
or U13556 (N_13556,N_6428,N_7079);
nor U13557 (N_13557,N_9418,N_6662);
nand U13558 (N_13558,N_5936,N_6547);
nor U13559 (N_13559,N_5320,N_6549);
xnor U13560 (N_13560,N_8647,N_9112);
and U13561 (N_13561,N_6522,N_6983);
or U13562 (N_13562,N_9713,N_7541);
nand U13563 (N_13563,N_7408,N_7832);
or U13564 (N_13564,N_8010,N_8144);
nand U13565 (N_13565,N_6951,N_5698);
and U13566 (N_13566,N_6264,N_5487);
or U13567 (N_13567,N_7894,N_9949);
or U13568 (N_13568,N_8588,N_9044);
nor U13569 (N_13569,N_7911,N_6246);
or U13570 (N_13570,N_7201,N_5265);
and U13571 (N_13571,N_5730,N_8368);
nor U13572 (N_13572,N_6760,N_6626);
nand U13573 (N_13573,N_5387,N_6579);
or U13574 (N_13574,N_9631,N_9445);
or U13575 (N_13575,N_9470,N_7937);
xnor U13576 (N_13576,N_7363,N_5751);
and U13577 (N_13577,N_6865,N_9378);
and U13578 (N_13578,N_8973,N_8784);
nor U13579 (N_13579,N_6625,N_8016);
or U13580 (N_13580,N_7944,N_9431);
nor U13581 (N_13581,N_9446,N_6819);
and U13582 (N_13582,N_8639,N_6711);
xor U13583 (N_13583,N_8266,N_7625);
nor U13584 (N_13584,N_5583,N_9280);
or U13585 (N_13585,N_6940,N_6936);
nand U13586 (N_13586,N_7074,N_7913);
nor U13587 (N_13587,N_5018,N_5484);
xor U13588 (N_13588,N_8808,N_8587);
and U13589 (N_13589,N_9800,N_9718);
nand U13590 (N_13590,N_5838,N_9329);
nand U13591 (N_13591,N_5213,N_6658);
xnor U13592 (N_13592,N_9315,N_9765);
nor U13593 (N_13593,N_5950,N_9345);
xnor U13594 (N_13594,N_5005,N_9952);
and U13595 (N_13595,N_9048,N_9077);
nand U13596 (N_13596,N_6405,N_6684);
and U13597 (N_13597,N_8910,N_9711);
nor U13598 (N_13598,N_6441,N_7243);
xor U13599 (N_13599,N_5650,N_6714);
xnor U13600 (N_13600,N_5374,N_9912);
and U13601 (N_13601,N_8775,N_9246);
nor U13602 (N_13602,N_7689,N_6618);
or U13603 (N_13603,N_5809,N_7808);
and U13604 (N_13604,N_8738,N_5044);
and U13605 (N_13605,N_5613,N_7144);
or U13606 (N_13606,N_5145,N_9675);
nand U13607 (N_13607,N_9460,N_7194);
nand U13608 (N_13608,N_9951,N_8446);
nor U13609 (N_13609,N_5301,N_6500);
nand U13610 (N_13610,N_5200,N_5674);
and U13611 (N_13611,N_6368,N_8164);
and U13612 (N_13612,N_9376,N_9732);
or U13613 (N_13613,N_6529,N_6690);
xor U13614 (N_13614,N_9359,N_7326);
nand U13615 (N_13615,N_7103,N_6530);
nand U13616 (N_13616,N_7474,N_5255);
xnor U13617 (N_13617,N_9500,N_9566);
or U13618 (N_13618,N_9324,N_7389);
nor U13619 (N_13619,N_9555,N_9499);
or U13620 (N_13620,N_6065,N_9128);
nand U13621 (N_13621,N_7892,N_7039);
or U13622 (N_13622,N_9205,N_5976);
and U13623 (N_13623,N_5914,N_8088);
or U13624 (N_13624,N_5484,N_6133);
or U13625 (N_13625,N_9847,N_8628);
nand U13626 (N_13626,N_8923,N_8100);
and U13627 (N_13627,N_7860,N_5633);
xnor U13628 (N_13628,N_5118,N_5832);
and U13629 (N_13629,N_8755,N_8411);
nand U13630 (N_13630,N_5256,N_5617);
and U13631 (N_13631,N_5620,N_8485);
nand U13632 (N_13632,N_5793,N_9754);
or U13633 (N_13633,N_6253,N_8924);
xor U13634 (N_13634,N_5038,N_5755);
nand U13635 (N_13635,N_6452,N_9882);
xor U13636 (N_13636,N_6373,N_8539);
nor U13637 (N_13637,N_8835,N_8456);
nand U13638 (N_13638,N_8964,N_6444);
nand U13639 (N_13639,N_9223,N_5797);
and U13640 (N_13640,N_5619,N_7763);
and U13641 (N_13641,N_7311,N_8191);
nand U13642 (N_13642,N_6237,N_6213);
or U13643 (N_13643,N_8273,N_8630);
or U13644 (N_13644,N_9411,N_5119);
nor U13645 (N_13645,N_5521,N_6030);
nor U13646 (N_13646,N_6778,N_9380);
nor U13647 (N_13647,N_8975,N_9337);
and U13648 (N_13648,N_9655,N_6488);
nor U13649 (N_13649,N_6535,N_6729);
nor U13650 (N_13650,N_9677,N_9269);
and U13651 (N_13651,N_8277,N_8380);
and U13652 (N_13652,N_6704,N_6786);
and U13653 (N_13653,N_9559,N_8433);
nor U13654 (N_13654,N_5889,N_7535);
nand U13655 (N_13655,N_7257,N_9289);
nor U13656 (N_13656,N_7743,N_9571);
nand U13657 (N_13657,N_6436,N_7757);
nor U13658 (N_13658,N_9238,N_5484);
nor U13659 (N_13659,N_8673,N_7676);
and U13660 (N_13660,N_9885,N_8963);
xnor U13661 (N_13661,N_5203,N_8496);
and U13662 (N_13662,N_5547,N_9907);
and U13663 (N_13663,N_5179,N_5797);
nor U13664 (N_13664,N_7292,N_9684);
xnor U13665 (N_13665,N_5124,N_6543);
or U13666 (N_13666,N_7946,N_7248);
nor U13667 (N_13667,N_5709,N_7525);
or U13668 (N_13668,N_9735,N_8748);
nand U13669 (N_13669,N_5879,N_5752);
or U13670 (N_13670,N_9105,N_8085);
nand U13671 (N_13671,N_8684,N_7773);
or U13672 (N_13672,N_5253,N_9009);
or U13673 (N_13673,N_6047,N_8958);
and U13674 (N_13674,N_5499,N_9991);
or U13675 (N_13675,N_6772,N_7359);
nor U13676 (N_13676,N_5540,N_6020);
nand U13677 (N_13677,N_7458,N_5039);
nor U13678 (N_13678,N_5336,N_9508);
nand U13679 (N_13679,N_8541,N_7212);
nor U13680 (N_13680,N_7196,N_8997);
nor U13681 (N_13681,N_5790,N_8057);
or U13682 (N_13682,N_8212,N_9237);
and U13683 (N_13683,N_9516,N_8551);
or U13684 (N_13684,N_6811,N_9670);
and U13685 (N_13685,N_5799,N_7630);
or U13686 (N_13686,N_9995,N_5391);
and U13687 (N_13687,N_6962,N_6883);
nor U13688 (N_13688,N_5497,N_6018);
nor U13689 (N_13689,N_9732,N_7744);
and U13690 (N_13690,N_6866,N_7521);
nor U13691 (N_13691,N_9309,N_8913);
nor U13692 (N_13692,N_6443,N_7210);
nand U13693 (N_13693,N_8980,N_9354);
or U13694 (N_13694,N_8018,N_8845);
nand U13695 (N_13695,N_6378,N_7880);
nand U13696 (N_13696,N_7695,N_9362);
or U13697 (N_13697,N_8028,N_5290);
and U13698 (N_13698,N_5259,N_5006);
nor U13699 (N_13699,N_9345,N_7394);
and U13700 (N_13700,N_5105,N_5111);
nor U13701 (N_13701,N_9103,N_9197);
and U13702 (N_13702,N_9061,N_7923);
and U13703 (N_13703,N_5452,N_9412);
and U13704 (N_13704,N_8926,N_5066);
or U13705 (N_13705,N_7422,N_5105);
nor U13706 (N_13706,N_8731,N_8618);
nand U13707 (N_13707,N_8807,N_5349);
xor U13708 (N_13708,N_9383,N_5022);
nand U13709 (N_13709,N_7030,N_7189);
and U13710 (N_13710,N_9945,N_7411);
or U13711 (N_13711,N_5939,N_7692);
and U13712 (N_13712,N_5721,N_9504);
nand U13713 (N_13713,N_8514,N_7408);
nor U13714 (N_13714,N_7110,N_6474);
or U13715 (N_13715,N_9262,N_6169);
nor U13716 (N_13716,N_8371,N_5251);
nand U13717 (N_13717,N_9957,N_9042);
and U13718 (N_13718,N_8692,N_8601);
nand U13719 (N_13719,N_8462,N_8572);
or U13720 (N_13720,N_6075,N_9432);
and U13721 (N_13721,N_9751,N_5290);
and U13722 (N_13722,N_9745,N_9256);
nand U13723 (N_13723,N_8820,N_9399);
nor U13724 (N_13724,N_9906,N_9592);
xnor U13725 (N_13725,N_5634,N_7195);
and U13726 (N_13726,N_5425,N_9669);
and U13727 (N_13727,N_8377,N_6007);
and U13728 (N_13728,N_7866,N_8161);
nand U13729 (N_13729,N_8384,N_7416);
nand U13730 (N_13730,N_5538,N_8784);
nand U13731 (N_13731,N_7992,N_5502);
and U13732 (N_13732,N_6456,N_9921);
or U13733 (N_13733,N_6407,N_9835);
and U13734 (N_13734,N_6696,N_5122);
or U13735 (N_13735,N_6619,N_9032);
nor U13736 (N_13736,N_9814,N_9212);
and U13737 (N_13737,N_9192,N_8382);
xnor U13738 (N_13738,N_6105,N_6137);
xnor U13739 (N_13739,N_7095,N_9370);
and U13740 (N_13740,N_8788,N_6425);
nor U13741 (N_13741,N_6921,N_9881);
and U13742 (N_13742,N_6654,N_8408);
xnor U13743 (N_13743,N_7283,N_7112);
nand U13744 (N_13744,N_5237,N_6848);
and U13745 (N_13745,N_6295,N_9554);
xor U13746 (N_13746,N_6133,N_8677);
nor U13747 (N_13747,N_5280,N_8041);
nor U13748 (N_13748,N_6597,N_6190);
xor U13749 (N_13749,N_6878,N_5582);
or U13750 (N_13750,N_6641,N_6442);
and U13751 (N_13751,N_7198,N_9641);
or U13752 (N_13752,N_5637,N_9418);
xor U13753 (N_13753,N_8930,N_7329);
nand U13754 (N_13754,N_9705,N_7188);
or U13755 (N_13755,N_8988,N_7749);
or U13756 (N_13756,N_6837,N_8247);
nand U13757 (N_13757,N_7796,N_7791);
and U13758 (N_13758,N_9692,N_7319);
or U13759 (N_13759,N_5714,N_9151);
or U13760 (N_13760,N_5133,N_8286);
nor U13761 (N_13761,N_5036,N_8056);
and U13762 (N_13762,N_6268,N_7973);
xnor U13763 (N_13763,N_7253,N_5214);
nor U13764 (N_13764,N_8662,N_5288);
nor U13765 (N_13765,N_5918,N_9708);
and U13766 (N_13766,N_8516,N_9867);
nand U13767 (N_13767,N_9609,N_7636);
nor U13768 (N_13768,N_5869,N_6179);
nand U13769 (N_13769,N_8529,N_8422);
and U13770 (N_13770,N_7236,N_9426);
nand U13771 (N_13771,N_8386,N_8231);
and U13772 (N_13772,N_6137,N_5382);
nor U13773 (N_13773,N_8654,N_8265);
and U13774 (N_13774,N_8561,N_8630);
or U13775 (N_13775,N_6529,N_6170);
or U13776 (N_13776,N_8032,N_6729);
nand U13777 (N_13777,N_6374,N_5978);
or U13778 (N_13778,N_6756,N_8192);
xnor U13779 (N_13779,N_9962,N_8657);
or U13780 (N_13780,N_7889,N_5238);
or U13781 (N_13781,N_8757,N_9414);
nor U13782 (N_13782,N_8650,N_9179);
xnor U13783 (N_13783,N_5865,N_5173);
and U13784 (N_13784,N_6164,N_9475);
and U13785 (N_13785,N_6386,N_5627);
or U13786 (N_13786,N_9189,N_5506);
and U13787 (N_13787,N_8531,N_7117);
xnor U13788 (N_13788,N_7884,N_5800);
nand U13789 (N_13789,N_9262,N_5886);
nor U13790 (N_13790,N_7081,N_7164);
xor U13791 (N_13791,N_9327,N_7170);
nor U13792 (N_13792,N_7769,N_8523);
and U13793 (N_13793,N_6560,N_6721);
or U13794 (N_13794,N_9152,N_7981);
nor U13795 (N_13795,N_5753,N_9697);
xor U13796 (N_13796,N_8762,N_6037);
or U13797 (N_13797,N_8650,N_9525);
nor U13798 (N_13798,N_9307,N_5664);
or U13799 (N_13799,N_7310,N_7518);
nor U13800 (N_13800,N_9903,N_7534);
or U13801 (N_13801,N_6247,N_7428);
nand U13802 (N_13802,N_9068,N_9104);
nand U13803 (N_13803,N_5298,N_9610);
or U13804 (N_13804,N_5355,N_7436);
or U13805 (N_13805,N_8233,N_7572);
and U13806 (N_13806,N_7143,N_7200);
nor U13807 (N_13807,N_6544,N_7598);
nand U13808 (N_13808,N_9307,N_7380);
nor U13809 (N_13809,N_8055,N_5271);
and U13810 (N_13810,N_9831,N_5179);
nor U13811 (N_13811,N_5012,N_8399);
and U13812 (N_13812,N_6731,N_8569);
xor U13813 (N_13813,N_9872,N_8859);
nor U13814 (N_13814,N_9148,N_7925);
nor U13815 (N_13815,N_8810,N_5366);
and U13816 (N_13816,N_7053,N_6474);
and U13817 (N_13817,N_5682,N_6898);
nor U13818 (N_13818,N_9238,N_5898);
and U13819 (N_13819,N_6322,N_5890);
or U13820 (N_13820,N_8825,N_9090);
or U13821 (N_13821,N_9610,N_7441);
and U13822 (N_13822,N_9985,N_9991);
and U13823 (N_13823,N_8938,N_5760);
and U13824 (N_13824,N_7387,N_9116);
and U13825 (N_13825,N_9653,N_7193);
nor U13826 (N_13826,N_5950,N_5653);
and U13827 (N_13827,N_6740,N_7624);
or U13828 (N_13828,N_6825,N_7696);
nor U13829 (N_13829,N_7542,N_9830);
and U13830 (N_13830,N_5409,N_8755);
and U13831 (N_13831,N_5463,N_7555);
nand U13832 (N_13832,N_6960,N_9015);
or U13833 (N_13833,N_5213,N_5982);
nand U13834 (N_13834,N_5677,N_5190);
or U13835 (N_13835,N_8534,N_5354);
nand U13836 (N_13836,N_9194,N_8408);
or U13837 (N_13837,N_9762,N_9222);
or U13838 (N_13838,N_9545,N_6955);
and U13839 (N_13839,N_6091,N_5657);
and U13840 (N_13840,N_6339,N_5199);
nand U13841 (N_13841,N_8452,N_5740);
or U13842 (N_13842,N_5146,N_6570);
or U13843 (N_13843,N_9675,N_7224);
nor U13844 (N_13844,N_7868,N_7333);
and U13845 (N_13845,N_8019,N_9937);
or U13846 (N_13846,N_8343,N_5968);
nand U13847 (N_13847,N_5491,N_7829);
nand U13848 (N_13848,N_7683,N_8352);
nand U13849 (N_13849,N_9155,N_7040);
or U13850 (N_13850,N_5795,N_5125);
and U13851 (N_13851,N_7781,N_5101);
and U13852 (N_13852,N_6476,N_7630);
xor U13853 (N_13853,N_8030,N_6793);
and U13854 (N_13854,N_6648,N_7669);
xor U13855 (N_13855,N_9341,N_5512);
nor U13856 (N_13856,N_9364,N_7988);
xnor U13857 (N_13857,N_8661,N_6642);
nand U13858 (N_13858,N_9203,N_7374);
nand U13859 (N_13859,N_5658,N_8764);
xor U13860 (N_13860,N_9823,N_5949);
nand U13861 (N_13861,N_7656,N_5127);
or U13862 (N_13862,N_5599,N_5495);
and U13863 (N_13863,N_8894,N_6298);
and U13864 (N_13864,N_9995,N_7060);
and U13865 (N_13865,N_7869,N_6074);
nor U13866 (N_13866,N_7985,N_9362);
nor U13867 (N_13867,N_7247,N_6257);
or U13868 (N_13868,N_5557,N_7176);
nor U13869 (N_13869,N_9808,N_7725);
nor U13870 (N_13870,N_9613,N_7514);
and U13871 (N_13871,N_8226,N_6906);
nor U13872 (N_13872,N_5484,N_9437);
xnor U13873 (N_13873,N_6824,N_9754);
nand U13874 (N_13874,N_5420,N_8513);
or U13875 (N_13875,N_8157,N_6642);
and U13876 (N_13876,N_7727,N_5278);
and U13877 (N_13877,N_5525,N_9697);
or U13878 (N_13878,N_7943,N_6147);
and U13879 (N_13879,N_9418,N_7822);
or U13880 (N_13880,N_8843,N_7719);
or U13881 (N_13881,N_7350,N_8728);
and U13882 (N_13882,N_5856,N_6911);
nor U13883 (N_13883,N_8893,N_6825);
and U13884 (N_13884,N_6710,N_9757);
and U13885 (N_13885,N_5857,N_8075);
xnor U13886 (N_13886,N_6278,N_6398);
nor U13887 (N_13887,N_6014,N_9195);
or U13888 (N_13888,N_9648,N_8286);
xor U13889 (N_13889,N_5484,N_6044);
and U13890 (N_13890,N_9201,N_8647);
and U13891 (N_13891,N_5801,N_8937);
and U13892 (N_13892,N_8125,N_8536);
or U13893 (N_13893,N_7000,N_8395);
and U13894 (N_13894,N_9480,N_6531);
and U13895 (N_13895,N_9461,N_6794);
nor U13896 (N_13896,N_7018,N_9024);
xnor U13897 (N_13897,N_7774,N_8829);
nor U13898 (N_13898,N_9051,N_7357);
nor U13899 (N_13899,N_7632,N_9906);
and U13900 (N_13900,N_8210,N_7037);
and U13901 (N_13901,N_5657,N_7866);
nand U13902 (N_13902,N_8784,N_5442);
nor U13903 (N_13903,N_8803,N_9483);
and U13904 (N_13904,N_9219,N_8337);
or U13905 (N_13905,N_9772,N_5158);
and U13906 (N_13906,N_5935,N_8682);
and U13907 (N_13907,N_8789,N_5937);
and U13908 (N_13908,N_5104,N_5390);
xnor U13909 (N_13909,N_9844,N_6610);
or U13910 (N_13910,N_7284,N_5129);
nand U13911 (N_13911,N_6656,N_6785);
and U13912 (N_13912,N_9784,N_6944);
nor U13913 (N_13913,N_9749,N_9607);
nand U13914 (N_13914,N_7867,N_7822);
xnor U13915 (N_13915,N_5635,N_5540);
and U13916 (N_13916,N_9852,N_7577);
xor U13917 (N_13917,N_8222,N_9135);
xnor U13918 (N_13918,N_8498,N_7259);
or U13919 (N_13919,N_9652,N_7538);
or U13920 (N_13920,N_8026,N_7002);
nand U13921 (N_13921,N_9625,N_5237);
nor U13922 (N_13922,N_7293,N_9036);
xnor U13923 (N_13923,N_6038,N_8602);
or U13924 (N_13924,N_9009,N_6115);
nand U13925 (N_13925,N_9603,N_9651);
nand U13926 (N_13926,N_6281,N_7508);
nor U13927 (N_13927,N_7960,N_9239);
or U13928 (N_13928,N_7665,N_5686);
nor U13929 (N_13929,N_5448,N_7601);
nand U13930 (N_13930,N_6851,N_9514);
nand U13931 (N_13931,N_6845,N_6522);
nor U13932 (N_13932,N_6132,N_8851);
xnor U13933 (N_13933,N_7708,N_7146);
nor U13934 (N_13934,N_6676,N_5505);
and U13935 (N_13935,N_5758,N_5271);
and U13936 (N_13936,N_6697,N_6224);
or U13937 (N_13937,N_9101,N_8488);
or U13938 (N_13938,N_6862,N_7190);
xor U13939 (N_13939,N_5554,N_8670);
nand U13940 (N_13940,N_6348,N_9274);
and U13941 (N_13941,N_7253,N_7256);
or U13942 (N_13942,N_9919,N_7027);
xnor U13943 (N_13943,N_8318,N_8562);
and U13944 (N_13944,N_5060,N_9339);
nand U13945 (N_13945,N_6511,N_9753);
and U13946 (N_13946,N_6406,N_5188);
and U13947 (N_13947,N_8228,N_7701);
nand U13948 (N_13948,N_9389,N_8364);
and U13949 (N_13949,N_5392,N_5705);
xnor U13950 (N_13950,N_7056,N_6435);
or U13951 (N_13951,N_6774,N_9571);
or U13952 (N_13952,N_9487,N_9023);
and U13953 (N_13953,N_8378,N_9407);
nand U13954 (N_13954,N_9849,N_8728);
or U13955 (N_13955,N_6797,N_8267);
and U13956 (N_13956,N_7999,N_7392);
and U13957 (N_13957,N_8735,N_5420);
nor U13958 (N_13958,N_6854,N_6733);
nor U13959 (N_13959,N_6236,N_5969);
xnor U13960 (N_13960,N_6746,N_8185);
nand U13961 (N_13961,N_6488,N_7845);
xnor U13962 (N_13962,N_7598,N_5611);
and U13963 (N_13963,N_7383,N_9467);
nand U13964 (N_13964,N_6099,N_7612);
nor U13965 (N_13965,N_9761,N_9411);
xor U13966 (N_13966,N_7882,N_5019);
nor U13967 (N_13967,N_7348,N_5611);
or U13968 (N_13968,N_9168,N_5593);
nor U13969 (N_13969,N_9330,N_6948);
or U13970 (N_13970,N_6376,N_5156);
or U13971 (N_13971,N_6787,N_7091);
or U13972 (N_13972,N_7736,N_9248);
nor U13973 (N_13973,N_5937,N_9359);
or U13974 (N_13974,N_7961,N_9708);
nand U13975 (N_13975,N_5756,N_8614);
or U13976 (N_13976,N_8693,N_9497);
and U13977 (N_13977,N_7183,N_6743);
xnor U13978 (N_13978,N_9817,N_9150);
or U13979 (N_13979,N_6505,N_6259);
nor U13980 (N_13980,N_9948,N_8600);
or U13981 (N_13981,N_7041,N_7712);
nor U13982 (N_13982,N_8623,N_6267);
nand U13983 (N_13983,N_9028,N_8631);
and U13984 (N_13984,N_6138,N_9151);
or U13985 (N_13985,N_5090,N_6411);
or U13986 (N_13986,N_5265,N_6729);
nand U13987 (N_13987,N_8268,N_8770);
nor U13988 (N_13988,N_8750,N_9942);
nand U13989 (N_13989,N_5987,N_5395);
nor U13990 (N_13990,N_7464,N_7699);
nor U13991 (N_13991,N_9843,N_7911);
and U13992 (N_13992,N_8049,N_8219);
nor U13993 (N_13993,N_6347,N_7122);
nand U13994 (N_13994,N_8099,N_8534);
nor U13995 (N_13995,N_6449,N_9657);
or U13996 (N_13996,N_5677,N_5349);
or U13997 (N_13997,N_8828,N_7765);
xor U13998 (N_13998,N_7931,N_8537);
and U13999 (N_13999,N_5317,N_5659);
or U14000 (N_14000,N_7603,N_8172);
or U14001 (N_14001,N_7558,N_5401);
nor U14002 (N_14002,N_6946,N_7054);
or U14003 (N_14003,N_8151,N_6952);
and U14004 (N_14004,N_5591,N_7056);
or U14005 (N_14005,N_7421,N_7738);
or U14006 (N_14006,N_7616,N_6439);
and U14007 (N_14007,N_8843,N_9220);
and U14008 (N_14008,N_8188,N_7534);
and U14009 (N_14009,N_6606,N_6552);
and U14010 (N_14010,N_6016,N_9512);
and U14011 (N_14011,N_8870,N_9515);
and U14012 (N_14012,N_8315,N_5225);
nand U14013 (N_14013,N_6673,N_9364);
nor U14014 (N_14014,N_9251,N_8802);
nor U14015 (N_14015,N_6915,N_6265);
and U14016 (N_14016,N_8540,N_9015);
nor U14017 (N_14017,N_9190,N_5428);
nor U14018 (N_14018,N_9659,N_5815);
or U14019 (N_14019,N_7510,N_7357);
or U14020 (N_14020,N_9657,N_6691);
nand U14021 (N_14021,N_9791,N_7377);
or U14022 (N_14022,N_8149,N_6197);
nand U14023 (N_14023,N_6457,N_7101);
and U14024 (N_14024,N_9885,N_7104);
or U14025 (N_14025,N_8791,N_5562);
and U14026 (N_14026,N_6180,N_8738);
nor U14027 (N_14027,N_6781,N_9385);
nor U14028 (N_14028,N_8952,N_8129);
or U14029 (N_14029,N_9106,N_8143);
nand U14030 (N_14030,N_7117,N_5382);
and U14031 (N_14031,N_6207,N_8521);
nor U14032 (N_14032,N_8014,N_7163);
nand U14033 (N_14033,N_6099,N_7394);
nor U14034 (N_14034,N_7248,N_7508);
nor U14035 (N_14035,N_8348,N_7611);
nor U14036 (N_14036,N_7212,N_8318);
and U14037 (N_14037,N_8894,N_6528);
nand U14038 (N_14038,N_7055,N_6817);
or U14039 (N_14039,N_6932,N_5443);
nor U14040 (N_14040,N_6634,N_9132);
nor U14041 (N_14041,N_8342,N_7923);
nor U14042 (N_14042,N_5541,N_6895);
and U14043 (N_14043,N_7388,N_5939);
or U14044 (N_14044,N_6615,N_9433);
nor U14045 (N_14045,N_8498,N_5991);
nand U14046 (N_14046,N_7328,N_5190);
or U14047 (N_14047,N_9268,N_9729);
nor U14048 (N_14048,N_8556,N_5704);
nor U14049 (N_14049,N_6510,N_9145);
nand U14050 (N_14050,N_8082,N_5458);
nand U14051 (N_14051,N_8853,N_5430);
nand U14052 (N_14052,N_8680,N_5388);
or U14053 (N_14053,N_7468,N_8404);
xor U14054 (N_14054,N_5780,N_9145);
or U14055 (N_14055,N_7771,N_6794);
nor U14056 (N_14056,N_9119,N_7962);
xor U14057 (N_14057,N_8261,N_9554);
nor U14058 (N_14058,N_8670,N_6710);
xor U14059 (N_14059,N_9966,N_5290);
and U14060 (N_14060,N_5989,N_6620);
nor U14061 (N_14061,N_8182,N_5311);
or U14062 (N_14062,N_6388,N_9714);
and U14063 (N_14063,N_7836,N_9424);
nand U14064 (N_14064,N_5570,N_5705);
nor U14065 (N_14065,N_6058,N_6401);
nand U14066 (N_14066,N_7667,N_8193);
nor U14067 (N_14067,N_8189,N_7419);
or U14068 (N_14068,N_5337,N_8657);
nor U14069 (N_14069,N_9326,N_9929);
nand U14070 (N_14070,N_8613,N_8572);
nand U14071 (N_14071,N_7317,N_5904);
or U14072 (N_14072,N_8837,N_7147);
or U14073 (N_14073,N_5438,N_8136);
nor U14074 (N_14074,N_5978,N_5400);
or U14075 (N_14075,N_7753,N_5954);
nand U14076 (N_14076,N_9523,N_8612);
nand U14077 (N_14077,N_7981,N_6077);
or U14078 (N_14078,N_6644,N_5384);
nor U14079 (N_14079,N_5259,N_5204);
nand U14080 (N_14080,N_5702,N_7853);
xnor U14081 (N_14081,N_5407,N_7569);
and U14082 (N_14082,N_8135,N_9253);
or U14083 (N_14083,N_8015,N_5031);
nand U14084 (N_14084,N_9166,N_6321);
nor U14085 (N_14085,N_7134,N_7112);
nand U14086 (N_14086,N_5644,N_5194);
nand U14087 (N_14087,N_6100,N_6825);
nor U14088 (N_14088,N_6214,N_8048);
nand U14089 (N_14089,N_7539,N_6638);
nor U14090 (N_14090,N_6162,N_7438);
nor U14091 (N_14091,N_7047,N_6737);
or U14092 (N_14092,N_8152,N_8658);
nor U14093 (N_14093,N_8265,N_6389);
xor U14094 (N_14094,N_9132,N_9184);
nor U14095 (N_14095,N_6085,N_8794);
and U14096 (N_14096,N_8059,N_9095);
or U14097 (N_14097,N_8100,N_8699);
nor U14098 (N_14098,N_6346,N_5451);
and U14099 (N_14099,N_5661,N_7021);
and U14100 (N_14100,N_5255,N_7119);
nor U14101 (N_14101,N_8807,N_5428);
and U14102 (N_14102,N_9372,N_5831);
or U14103 (N_14103,N_7667,N_7981);
and U14104 (N_14104,N_8020,N_7068);
nand U14105 (N_14105,N_6999,N_5784);
nand U14106 (N_14106,N_9396,N_7290);
and U14107 (N_14107,N_7198,N_7874);
nor U14108 (N_14108,N_7809,N_9226);
xnor U14109 (N_14109,N_5255,N_9503);
nand U14110 (N_14110,N_9842,N_5048);
nand U14111 (N_14111,N_6592,N_9638);
and U14112 (N_14112,N_5648,N_8952);
or U14113 (N_14113,N_9947,N_6013);
nand U14114 (N_14114,N_8310,N_7130);
nand U14115 (N_14115,N_6453,N_7153);
or U14116 (N_14116,N_9266,N_6062);
xor U14117 (N_14117,N_9339,N_8336);
or U14118 (N_14118,N_9378,N_7029);
xnor U14119 (N_14119,N_6968,N_6426);
and U14120 (N_14120,N_6020,N_6262);
or U14121 (N_14121,N_9529,N_7150);
or U14122 (N_14122,N_9655,N_6568);
and U14123 (N_14123,N_7002,N_9797);
nor U14124 (N_14124,N_8805,N_8197);
nor U14125 (N_14125,N_5779,N_9812);
nand U14126 (N_14126,N_7825,N_7997);
or U14127 (N_14127,N_5241,N_5283);
nand U14128 (N_14128,N_5160,N_8150);
nand U14129 (N_14129,N_5589,N_7254);
nand U14130 (N_14130,N_8492,N_7153);
nor U14131 (N_14131,N_5317,N_7849);
nand U14132 (N_14132,N_5759,N_6686);
or U14133 (N_14133,N_9208,N_8435);
nor U14134 (N_14134,N_8170,N_5438);
nor U14135 (N_14135,N_9307,N_8122);
nand U14136 (N_14136,N_7684,N_7926);
nand U14137 (N_14137,N_9526,N_9640);
nand U14138 (N_14138,N_8955,N_5219);
and U14139 (N_14139,N_7266,N_9235);
nor U14140 (N_14140,N_9710,N_8954);
and U14141 (N_14141,N_8901,N_8467);
and U14142 (N_14142,N_9205,N_8303);
and U14143 (N_14143,N_5210,N_9785);
nor U14144 (N_14144,N_8945,N_7374);
and U14145 (N_14145,N_7726,N_5043);
nor U14146 (N_14146,N_7453,N_8575);
or U14147 (N_14147,N_5416,N_7920);
xnor U14148 (N_14148,N_8408,N_5060);
nand U14149 (N_14149,N_9964,N_9439);
nor U14150 (N_14150,N_5422,N_6881);
nor U14151 (N_14151,N_7176,N_9492);
nor U14152 (N_14152,N_5486,N_5047);
nor U14153 (N_14153,N_7959,N_9606);
nor U14154 (N_14154,N_8009,N_7226);
nor U14155 (N_14155,N_5033,N_9330);
or U14156 (N_14156,N_6427,N_5067);
xor U14157 (N_14157,N_7500,N_8213);
nand U14158 (N_14158,N_9936,N_8083);
and U14159 (N_14159,N_9583,N_9427);
nand U14160 (N_14160,N_8167,N_5658);
nand U14161 (N_14161,N_7653,N_7220);
xnor U14162 (N_14162,N_9198,N_7246);
nor U14163 (N_14163,N_9947,N_6996);
and U14164 (N_14164,N_8606,N_8157);
xor U14165 (N_14165,N_9859,N_9356);
nor U14166 (N_14166,N_7767,N_9699);
or U14167 (N_14167,N_5250,N_5673);
nand U14168 (N_14168,N_5816,N_8022);
xor U14169 (N_14169,N_9791,N_6806);
nand U14170 (N_14170,N_9726,N_7832);
xor U14171 (N_14171,N_6021,N_5186);
and U14172 (N_14172,N_6875,N_7580);
nor U14173 (N_14173,N_8306,N_7780);
or U14174 (N_14174,N_5554,N_6760);
or U14175 (N_14175,N_6402,N_8848);
nor U14176 (N_14176,N_9961,N_5518);
nor U14177 (N_14177,N_7998,N_6523);
nand U14178 (N_14178,N_5074,N_7726);
nor U14179 (N_14179,N_8007,N_7706);
nand U14180 (N_14180,N_9374,N_7749);
and U14181 (N_14181,N_9013,N_7003);
and U14182 (N_14182,N_8266,N_9336);
or U14183 (N_14183,N_5071,N_9279);
nor U14184 (N_14184,N_5101,N_8609);
xor U14185 (N_14185,N_5701,N_7683);
nor U14186 (N_14186,N_9747,N_5693);
or U14187 (N_14187,N_8711,N_6186);
or U14188 (N_14188,N_5832,N_7630);
xnor U14189 (N_14189,N_7172,N_5246);
nor U14190 (N_14190,N_8478,N_9991);
or U14191 (N_14191,N_9848,N_5052);
and U14192 (N_14192,N_8465,N_6062);
or U14193 (N_14193,N_6814,N_9785);
nor U14194 (N_14194,N_8269,N_6292);
nand U14195 (N_14195,N_7194,N_9342);
and U14196 (N_14196,N_8073,N_7423);
and U14197 (N_14197,N_5977,N_5606);
nand U14198 (N_14198,N_5757,N_7111);
nand U14199 (N_14199,N_8251,N_5847);
or U14200 (N_14200,N_7463,N_7123);
and U14201 (N_14201,N_8778,N_8808);
or U14202 (N_14202,N_5897,N_5423);
nor U14203 (N_14203,N_8272,N_7564);
and U14204 (N_14204,N_8883,N_6302);
or U14205 (N_14205,N_6698,N_9326);
and U14206 (N_14206,N_6744,N_7409);
and U14207 (N_14207,N_7794,N_6698);
or U14208 (N_14208,N_5494,N_7480);
or U14209 (N_14209,N_7760,N_6334);
nor U14210 (N_14210,N_7515,N_8836);
nand U14211 (N_14211,N_7317,N_5007);
or U14212 (N_14212,N_5136,N_8982);
xnor U14213 (N_14213,N_9974,N_7089);
or U14214 (N_14214,N_7183,N_6257);
nand U14215 (N_14215,N_6158,N_8287);
nand U14216 (N_14216,N_5264,N_8766);
or U14217 (N_14217,N_9693,N_6277);
and U14218 (N_14218,N_7595,N_5386);
and U14219 (N_14219,N_5398,N_5680);
and U14220 (N_14220,N_8392,N_5883);
or U14221 (N_14221,N_9506,N_9811);
nor U14222 (N_14222,N_7343,N_7993);
or U14223 (N_14223,N_6684,N_9404);
nand U14224 (N_14224,N_5989,N_5866);
xnor U14225 (N_14225,N_8977,N_8855);
nor U14226 (N_14226,N_9429,N_9015);
nand U14227 (N_14227,N_7564,N_6787);
or U14228 (N_14228,N_5705,N_5691);
nor U14229 (N_14229,N_5826,N_7191);
and U14230 (N_14230,N_5461,N_5008);
nor U14231 (N_14231,N_6577,N_7850);
and U14232 (N_14232,N_7271,N_7680);
and U14233 (N_14233,N_5791,N_8948);
nand U14234 (N_14234,N_9626,N_7875);
nor U14235 (N_14235,N_6961,N_9405);
or U14236 (N_14236,N_5007,N_6600);
and U14237 (N_14237,N_7819,N_6048);
nand U14238 (N_14238,N_6763,N_6262);
nor U14239 (N_14239,N_8285,N_7920);
nor U14240 (N_14240,N_5356,N_8828);
nand U14241 (N_14241,N_8198,N_5554);
or U14242 (N_14242,N_6634,N_8318);
nor U14243 (N_14243,N_9588,N_6960);
nand U14244 (N_14244,N_7805,N_6256);
or U14245 (N_14245,N_8598,N_9757);
nand U14246 (N_14246,N_5053,N_5065);
and U14247 (N_14247,N_8311,N_8501);
and U14248 (N_14248,N_9889,N_8796);
nor U14249 (N_14249,N_9540,N_5454);
nor U14250 (N_14250,N_7352,N_5936);
and U14251 (N_14251,N_9356,N_6824);
nand U14252 (N_14252,N_5322,N_6199);
nand U14253 (N_14253,N_7363,N_8545);
xor U14254 (N_14254,N_6224,N_5369);
or U14255 (N_14255,N_7484,N_7030);
and U14256 (N_14256,N_9386,N_5384);
nand U14257 (N_14257,N_6772,N_7673);
and U14258 (N_14258,N_7975,N_6114);
nor U14259 (N_14259,N_7511,N_9354);
xor U14260 (N_14260,N_9875,N_9262);
nor U14261 (N_14261,N_9024,N_8836);
xor U14262 (N_14262,N_7737,N_8509);
nand U14263 (N_14263,N_9088,N_5825);
and U14264 (N_14264,N_6996,N_7531);
nor U14265 (N_14265,N_9818,N_8928);
or U14266 (N_14266,N_6627,N_5628);
nand U14267 (N_14267,N_8708,N_6365);
or U14268 (N_14268,N_9311,N_9544);
nand U14269 (N_14269,N_7195,N_6985);
nand U14270 (N_14270,N_7976,N_6083);
nand U14271 (N_14271,N_9517,N_7046);
and U14272 (N_14272,N_9561,N_6605);
nor U14273 (N_14273,N_5353,N_9986);
or U14274 (N_14274,N_7776,N_9698);
nand U14275 (N_14275,N_8182,N_5236);
nor U14276 (N_14276,N_8642,N_6091);
xnor U14277 (N_14277,N_7505,N_7398);
nor U14278 (N_14278,N_5992,N_5813);
and U14279 (N_14279,N_8018,N_6862);
and U14280 (N_14280,N_7354,N_9054);
or U14281 (N_14281,N_7733,N_6445);
nor U14282 (N_14282,N_8983,N_6874);
and U14283 (N_14283,N_9958,N_5792);
nand U14284 (N_14284,N_6968,N_6090);
and U14285 (N_14285,N_5818,N_8884);
and U14286 (N_14286,N_8216,N_6379);
nor U14287 (N_14287,N_8642,N_6006);
nand U14288 (N_14288,N_5995,N_7323);
and U14289 (N_14289,N_8354,N_6457);
nor U14290 (N_14290,N_6061,N_9265);
nor U14291 (N_14291,N_6350,N_7295);
or U14292 (N_14292,N_8992,N_5969);
and U14293 (N_14293,N_5624,N_5601);
or U14294 (N_14294,N_9568,N_6051);
or U14295 (N_14295,N_7002,N_9654);
xnor U14296 (N_14296,N_8441,N_6186);
and U14297 (N_14297,N_7484,N_9135);
nand U14298 (N_14298,N_7603,N_7483);
nand U14299 (N_14299,N_7972,N_9730);
nor U14300 (N_14300,N_8758,N_7802);
nor U14301 (N_14301,N_6094,N_7687);
or U14302 (N_14302,N_8260,N_9056);
xor U14303 (N_14303,N_7936,N_9021);
nor U14304 (N_14304,N_5006,N_8358);
nor U14305 (N_14305,N_7573,N_6698);
nor U14306 (N_14306,N_6116,N_6748);
nor U14307 (N_14307,N_7853,N_7856);
nand U14308 (N_14308,N_9450,N_5804);
or U14309 (N_14309,N_7760,N_7092);
xor U14310 (N_14310,N_8372,N_9812);
and U14311 (N_14311,N_8872,N_8140);
nor U14312 (N_14312,N_8129,N_7884);
and U14313 (N_14313,N_9045,N_6723);
nor U14314 (N_14314,N_6734,N_6682);
or U14315 (N_14315,N_8260,N_8421);
xnor U14316 (N_14316,N_8981,N_6938);
nor U14317 (N_14317,N_9716,N_6443);
nor U14318 (N_14318,N_8916,N_9076);
nor U14319 (N_14319,N_9920,N_5615);
xnor U14320 (N_14320,N_5182,N_5037);
and U14321 (N_14321,N_7338,N_8435);
nand U14322 (N_14322,N_7917,N_7760);
and U14323 (N_14323,N_8581,N_5676);
nor U14324 (N_14324,N_8918,N_6570);
xor U14325 (N_14325,N_7845,N_6294);
nor U14326 (N_14326,N_6463,N_7853);
or U14327 (N_14327,N_6895,N_7492);
and U14328 (N_14328,N_9605,N_9261);
and U14329 (N_14329,N_9326,N_7678);
or U14330 (N_14330,N_7414,N_7599);
nand U14331 (N_14331,N_6802,N_6273);
xnor U14332 (N_14332,N_5282,N_7191);
and U14333 (N_14333,N_7942,N_5225);
nor U14334 (N_14334,N_9382,N_7945);
or U14335 (N_14335,N_8777,N_9722);
or U14336 (N_14336,N_6107,N_5001);
nand U14337 (N_14337,N_9310,N_8911);
or U14338 (N_14338,N_5851,N_9206);
nor U14339 (N_14339,N_7968,N_9069);
nand U14340 (N_14340,N_8573,N_7239);
nand U14341 (N_14341,N_8385,N_5399);
and U14342 (N_14342,N_7451,N_7722);
xnor U14343 (N_14343,N_5002,N_9481);
nand U14344 (N_14344,N_5611,N_7149);
nor U14345 (N_14345,N_7688,N_5472);
xor U14346 (N_14346,N_8896,N_7627);
nor U14347 (N_14347,N_5338,N_8684);
or U14348 (N_14348,N_6098,N_6197);
or U14349 (N_14349,N_9645,N_9004);
and U14350 (N_14350,N_5151,N_5514);
xnor U14351 (N_14351,N_9290,N_6484);
nand U14352 (N_14352,N_9849,N_8129);
or U14353 (N_14353,N_8333,N_5188);
nand U14354 (N_14354,N_5550,N_5068);
and U14355 (N_14355,N_7326,N_9556);
or U14356 (N_14356,N_6834,N_5808);
nand U14357 (N_14357,N_5151,N_5220);
nand U14358 (N_14358,N_5811,N_6622);
and U14359 (N_14359,N_8550,N_5853);
and U14360 (N_14360,N_7173,N_5830);
or U14361 (N_14361,N_7254,N_9288);
and U14362 (N_14362,N_6206,N_8100);
xor U14363 (N_14363,N_7298,N_5486);
and U14364 (N_14364,N_5898,N_8152);
and U14365 (N_14365,N_6513,N_7867);
and U14366 (N_14366,N_8832,N_7381);
nand U14367 (N_14367,N_7125,N_6317);
xor U14368 (N_14368,N_6997,N_9097);
and U14369 (N_14369,N_9316,N_8971);
and U14370 (N_14370,N_6411,N_7270);
xor U14371 (N_14371,N_5765,N_6705);
or U14372 (N_14372,N_7580,N_5514);
or U14373 (N_14373,N_7733,N_9919);
nand U14374 (N_14374,N_6118,N_7998);
xor U14375 (N_14375,N_9113,N_5252);
nand U14376 (N_14376,N_8541,N_5705);
nor U14377 (N_14377,N_5431,N_9787);
nand U14378 (N_14378,N_8867,N_6748);
nor U14379 (N_14379,N_8575,N_6183);
or U14380 (N_14380,N_8296,N_9527);
nand U14381 (N_14381,N_8340,N_5407);
or U14382 (N_14382,N_7279,N_8866);
nor U14383 (N_14383,N_7663,N_8686);
nand U14384 (N_14384,N_5858,N_6061);
and U14385 (N_14385,N_9294,N_7028);
or U14386 (N_14386,N_9950,N_7791);
or U14387 (N_14387,N_7185,N_7372);
nand U14388 (N_14388,N_6824,N_9864);
or U14389 (N_14389,N_7464,N_8097);
nand U14390 (N_14390,N_9286,N_6330);
and U14391 (N_14391,N_5303,N_6036);
and U14392 (N_14392,N_9888,N_8988);
or U14393 (N_14393,N_5238,N_8637);
and U14394 (N_14394,N_7152,N_5315);
nor U14395 (N_14395,N_5739,N_5996);
xor U14396 (N_14396,N_9800,N_7459);
nand U14397 (N_14397,N_6517,N_7572);
and U14398 (N_14398,N_7656,N_9027);
and U14399 (N_14399,N_9812,N_6848);
and U14400 (N_14400,N_6842,N_8581);
nor U14401 (N_14401,N_9192,N_7164);
xor U14402 (N_14402,N_6532,N_7434);
or U14403 (N_14403,N_6404,N_9777);
and U14404 (N_14404,N_6173,N_9462);
and U14405 (N_14405,N_9572,N_5325);
nor U14406 (N_14406,N_9494,N_6111);
and U14407 (N_14407,N_6059,N_7574);
or U14408 (N_14408,N_6583,N_5944);
nor U14409 (N_14409,N_9622,N_9528);
and U14410 (N_14410,N_9193,N_9469);
or U14411 (N_14411,N_5440,N_8690);
nor U14412 (N_14412,N_6714,N_9484);
nand U14413 (N_14413,N_7555,N_8240);
or U14414 (N_14414,N_8396,N_8384);
or U14415 (N_14415,N_6931,N_5957);
or U14416 (N_14416,N_8559,N_5984);
nor U14417 (N_14417,N_9065,N_8484);
nor U14418 (N_14418,N_9177,N_6527);
nor U14419 (N_14419,N_8844,N_8126);
nor U14420 (N_14420,N_6657,N_9033);
nor U14421 (N_14421,N_7660,N_6303);
nand U14422 (N_14422,N_5910,N_6224);
xnor U14423 (N_14423,N_5515,N_9596);
and U14424 (N_14424,N_5209,N_8958);
nor U14425 (N_14425,N_5884,N_5689);
or U14426 (N_14426,N_9621,N_8000);
nand U14427 (N_14427,N_5685,N_7398);
nor U14428 (N_14428,N_5711,N_7632);
nor U14429 (N_14429,N_8851,N_8996);
nor U14430 (N_14430,N_6762,N_9430);
nor U14431 (N_14431,N_9941,N_9338);
nor U14432 (N_14432,N_7255,N_9397);
nor U14433 (N_14433,N_7184,N_6271);
and U14434 (N_14434,N_7086,N_9574);
nand U14435 (N_14435,N_7765,N_5393);
nand U14436 (N_14436,N_8087,N_5259);
nand U14437 (N_14437,N_7197,N_7402);
nor U14438 (N_14438,N_5686,N_6312);
and U14439 (N_14439,N_9867,N_9425);
nand U14440 (N_14440,N_8010,N_8509);
nor U14441 (N_14441,N_7066,N_7492);
nor U14442 (N_14442,N_9563,N_5967);
nor U14443 (N_14443,N_6420,N_9304);
nand U14444 (N_14444,N_9755,N_7444);
nand U14445 (N_14445,N_7999,N_7555);
or U14446 (N_14446,N_8042,N_7076);
and U14447 (N_14447,N_9198,N_9862);
nor U14448 (N_14448,N_8438,N_7998);
or U14449 (N_14449,N_6978,N_6864);
nor U14450 (N_14450,N_6393,N_6832);
nor U14451 (N_14451,N_9341,N_8282);
xnor U14452 (N_14452,N_5150,N_8979);
nor U14453 (N_14453,N_5245,N_8408);
nand U14454 (N_14454,N_9735,N_8784);
nand U14455 (N_14455,N_9999,N_9613);
nor U14456 (N_14456,N_9157,N_6961);
and U14457 (N_14457,N_9572,N_9982);
nor U14458 (N_14458,N_8717,N_6872);
and U14459 (N_14459,N_8548,N_7448);
or U14460 (N_14460,N_5977,N_8297);
nand U14461 (N_14461,N_7184,N_5339);
nor U14462 (N_14462,N_5283,N_9907);
or U14463 (N_14463,N_8187,N_6086);
nand U14464 (N_14464,N_5076,N_8885);
or U14465 (N_14465,N_5575,N_9445);
nand U14466 (N_14466,N_8797,N_9281);
and U14467 (N_14467,N_7163,N_9071);
nor U14468 (N_14468,N_5351,N_7626);
or U14469 (N_14469,N_9422,N_5453);
nand U14470 (N_14470,N_6194,N_6975);
nand U14471 (N_14471,N_5827,N_6496);
nand U14472 (N_14472,N_8760,N_7532);
or U14473 (N_14473,N_6524,N_6763);
nand U14474 (N_14474,N_5492,N_5891);
or U14475 (N_14475,N_9110,N_5032);
nand U14476 (N_14476,N_8066,N_5828);
and U14477 (N_14477,N_9878,N_8436);
nor U14478 (N_14478,N_7533,N_7915);
and U14479 (N_14479,N_9955,N_8114);
nand U14480 (N_14480,N_7090,N_6113);
or U14481 (N_14481,N_7102,N_6824);
nand U14482 (N_14482,N_5275,N_9931);
and U14483 (N_14483,N_5337,N_8130);
or U14484 (N_14484,N_5687,N_6749);
nand U14485 (N_14485,N_9016,N_5328);
xnor U14486 (N_14486,N_6430,N_9002);
nor U14487 (N_14487,N_5074,N_9702);
or U14488 (N_14488,N_8042,N_6492);
xor U14489 (N_14489,N_5098,N_5301);
xnor U14490 (N_14490,N_6686,N_9755);
and U14491 (N_14491,N_6913,N_7093);
nand U14492 (N_14492,N_6320,N_8593);
xor U14493 (N_14493,N_7158,N_9800);
and U14494 (N_14494,N_8251,N_9701);
or U14495 (N_14495,N_6955,N_9349);
or U14496 (N_14496,N_6091,N_8887);
and U14497 (N_14497,N_9304,N_9539);
and U14498 (N_14498,N_7283,N_7188);
xnor U14499 (N_14499,N_6413,N_9774);
or U14500 (N_14500,N_8605,N_8014);
and U14501 (N_14501,N_5720,N_8902);
or U14502 (N_14502,N_8297,N_6342);
or U14503 (N_14503,N_5585,N_8573);
nand U14504 (N_14504,N_5608,N_7235);
nor U14505 (N_14505,N_8917,N_7234);
nor U14506 (N_14506,N_6449,N_9231);
and U14507 (N_14507,N_9667,N_9286);
nand U14508 (N_14508,N_8980,N_6031);
nand U14509 (N_14509,N_6042,N_9846);
or U14510 (N_14510,N_9481,N_5514);
or U14511 (N_14511,N_7125,N_6725);
and U14512 (N_14512,N_6271,N_6166);
xor U14513 (N_14513,N_8101,N_8596);
nor U14514 (N_14514,N_6102,N_6546);
or U14515 (N_14515,N_6444,N_5180);
or U14516 (N_14516,N_8878,N_6222);
xnor U14517 (N_14517,N_6975,N_9829);
or U14518 (N_14518,N_9955,N_6050);
nor U14519 (N_14519,N_5085,N_6767);
and U14520 (N_14520,N_9441,N_8581);
or U14521 (N_14521,N_5489,N_7403);
or U14522 (N_14522,N_5652,N_8006);
nor U14523 (N_14523,N_6817,N_7007);
and U14524 (N_14524,N_6317,N_7286);
nand U14525 (N_14525,N_8008,N_9541);
or U14526 (N_14526,N_8283,N_7789);
nand U14527 (N_14527,N_5976,N_6354);
or U14528 (N_14528,N_7186,N_7488);
nand U14529 (N_14529,N_6005,N_6323);
nor U14530 (N_14530,N_9037,N_9791);
nand U14531 (N_14531,N_7513,N_5849);
xnor U14532 (N_14532,N_5887,N_8695);
and U14533 (N_14533,N_5563,N_5452);
or U14534 (N_14534,N_9115,N_6265);
and U14535 (N_14535,N_9825,N_6774);
xnor U14536 (N_14536,N_5577,N_9620);
and U14537 (N_14537,N_5912,N_7376);
nor U14538 (N_14538,N_8148,N_5535);
nand U14539 (N_14539,N_9709,N_9125);
or U14540 (N_14540,N_6704,N_8868);
or U14541 (N_14541,N_9833,N_5344);
or U14542 (N_14542,N_7482,N_6506);
xnor U14543 (N_14543,N_7850,N_9263);
nand U14544 (N_14544,N_9294,N_5635);
and U14545 (N_14545,N_5982,N_6345);
or U14546 (N_14546,N_8863,N_7497);
or U14547 (N_14547,N_5669,N_9837);
and U14548 (N_14548,N_7401,N_9788);
and U14549 (N_14549,N_7865,N_8295);
and U14550 (N_14550,N_9959,N_6861);
nor U14551 (N_14551,N_5786,N_8586);
and U14552 (N_14552,N_5775,N_9771);
nand U14553 (N_14553,N_6162,N_7278);
nor U14554 (N_14554,N_9881,N_8772);
xnor U14555 (N_14555,N_8928,N_8069);
and U14556 (N_14556,N_7159,N_7096);
or U14557 (N_14557,N_5054,N_5520);
or U14558 (N_14558,N_9629,N_9161);
or U14559 (N_14559,N_9747,N_8951);
nand U14560 (N_14560,N_6263,N_9311);
nor U14561 (N_14561,N_7670,N_8236);
or U14562 (N_14562,N_7002,N_9413);
or U14563 (N_14563,N_6139,N_7161);
nor U14564 (N_14564,N_7474,N_5647);
and U14565 (N_14565,N_7474,N_7164);
and U14566 (N_14566,N_5648,N_8370);
and U14567 (N_14567,N_5393,N_5475);
nand U14568 (N_14568,N_9619,N_7751);
or U14569 (N_14569,N_7799,N_8698);
and U14570 (N_14570,N_5331,N_9462);
or U14571 (N_14571,N_6098,N_5412);
and U14572 (N_14572,N_6136,N_5186);
nor U14573 (N_14573,N_6828,N_7571);
and U14574 (N_14574,N_9513,N_5704);
and U14575 (N_14575,N_7366,N_7309);
nor U14576 (N_14576,N_9201,N_6569);
and U14577 (N_14577,N_5286,N_5976);
nor U14578 (N_14578,N_5669,N_6456);
nand U14579 (N_14579,N_7477,N_9168);
nor U14580 (N_14580,N_5901,N_7096);
or U14581 (N_14581,N_5398,N_5572);
and U14582 (N_14582,N_6963,N_6116);
or U14583 (N_14583,N_5765,N_6769);
xor U14584 (N_14584,N_9817,N_7569);
nor U14585 (N_14585,N_9716,N_6415);
nor U14586 (N_14586,N_5887,N_9051);
or U14587 (N_14587,N_8881,N_5549);
or U14588 (N_14588,N_7657,N_6254);
or U14589 (N_14589,N_7651,N_5390);
or U14590 (N_14590,N_9393,N_5864);
nand U14591 (N_14591,N_7150,N_7259);
nor U14592 (N_14592,N_8506,N_7566);
xor U14593 (N_14593,N_5986,N_7267);
nand U14594 (N_14594,N_8909,N_8138);
nor U14595 (N_14595,N_9598,N_5053);
and U14596 (N_14596,N_7845,N_9730);
xor U14597 (N_14597,N_8322,N_6951);
or U14598 (N_14598,N_9131,N_7856);
and U14599 (N_14599,N_9220,N_6777);
and U14600 (N_14600,N_9084,N_6107);
nand U14601 (N_14601,N_7467,N_6075);
nand U14602 (N_14602,N_6983,N_6019);
or U14603 (N_14603,N_7161,N_6801);
and U14604 (N_14604,N_9392,N_9363);
or U14605 (N_14605,N_5493,N_5118);
or U14606 (N_14606,N_8018,N_8829);
nand U14607 (N_14607,N_5748,N_8480);
nand U14608 (N_14608,N_9834,N_8278);
and U14609 (N_14609,N_6703,N_6847);
xor U14610 (N_14610,N_6376,N_8281);
nand U14611 (N_14611,N_8686,N_5912);
nand U14612 (N_14612,N_9426,N_8464);
nor U14613 (N_14613,N_7361,N_7094);
nor U14614 (N_14614,N_7645,N_5762);
nand U14615 (N_14615,N_8438,N_5025);
and U14616 (N_14616,N_6145,N_5769);
or U14617 (N_14617,N_5806,N_7684);
or U14618 (N_14618,N_7244,N_7447);
and U14619 (N_14619,N_9040,N_8199);
xor U14620 (N_14620,N_9287,N_5977);
nand U14621 (N_14621,N_5109,N_8565);
or U14622 (N_14622,N_9149,N_5149);
nor U14623 (N_14623,N_8872,N_5173);
nor U14624 (N_14624,N_5699,N_9686);
or U14625 (N_14625,N_8288,N_9819);
and U14626 (N_14626,N_9325,N_9977);
xnor U14627 (N_14627,N_9777,N_8143);
xnor U14628 (N_14628,N_5025,N_7030);
and U14629 (N_14629,N_9802,N_9804);
and U14630 (N_14630,N_7922,N_8548);
or U14631 (N_14631,N_7003,N_5979);
xnor U14632 (N_14632,N_7396,N_6900);
or U14633 (N_14633,N_6404,N_5027);
or U14634 (N_14634,N_9831,N_8040);
or U14635 (N_14635,N_8591,N_8769);
nand U14636 (N_14636,N_6059,N_9840);
and U14637 (N_14637,N_5288,N_7326);
and U14638 (N_14638,N_5429,N_5039);
nor U14639 (N_14639,N_7939,N_6631);
or U14640 (N_14640,N_7755,N_5314);
nand U14641 (N_14641,N_5151,N_5435);
and U14642 (N_14642,N_6745,N_7131);
nand U14643 (N_14643,N_7430,N_6815);
nor U14644 (N_14644,N_5011,N_7511);
xnor U14645 (N_14645,N_9160,N_6430);
and U14646 (N_14646,N_6818,N_5487);
xor U14647 (N_14647,N_6886,N_5079);
nor U14648 (N_14648,N_5678,N_9489);
nor U14649 (N_14649,N_8688,N_9287);
nor U14650 (N_14650,N_7199,N_5386);
xnor U14651 (N_14651,N_6654,N_6097);
nor U14652 (N_14652,N_8503,N_7065);
xor U14653 (N_14653,N_8599,N_8903);
or U14654 (N_14654,N_8777,N_9839);
xnor U14655 (N_14655,N_6737,N_8190);
nor U14656 (N_14656,N_8213,N_8166);
and U14657 (N_14657,N_8143,N_7247);
or U14658 (N_14658,N_7723,N_6193);
xnor U14659 (N_14659,N_8132,N_6463);
nand U14660 (N_14660,N_8749,N_5935);
nand U14661 (N_14661,N_5846,N_8135);
nor U14662 (N_14662,N_6585,N_6672);
or U14663 (N_14663,N_9580,N_5942);
xor U14664 (N_14664,N_5504,N_9675);
nand U14665 (N_14665,N_7685,N_6215);
nor U14666 (N_14666,N_8393,N_6014);
and U14667 (N_14667,N_9040,N_7555);
nand U14668 (N_14668,N_7853,N_6972);
nand U14669 (N_14669,N_9406,N_5746);
and U14670 (N_14670,N_6255,N_9469);
nand U14671 (N_14671,N_6597,N_9244);
or U14672 (N_14672,N_7165,N_6681);
or U14673 (N_14673,N_7765,N_9828);
nand U14674 (N_14674,N_8395,N_7111);
nand U14675 (N_14675,N_8421,N_7292);
or U14676 (N_14676,N_7578,N_8154);
and U14677 (N_14677,N_7319,N_8637);
or U14678 (N_14678,N_9019,N_9531);
nor U14679 (N_14679,N_8597,N_6515);
nand U14680 (N_14680,N_9379,N_8265);
or U14681 (N_14681,N_5153,N_9530);
nand U14682 (N_14682,N_5185,N_9245);
nor U14683 (N_14683,N_5018,N_5272);
and U14684 (N_14684,N_7859,N_6055);
and U14685 (N_14685,N_6170,N_9717);
and U14686 (N_14686,N_6272,N_5521);
or U14687 (N_14687,N_7240,N_6679);
nor U14688 (N_14688,N_8686,N_8534);
and U14689 (N_14689,N_5014,N_8811);
and U14690 (N_14690,N_8426,N_6748);
and U14691 (N_14691,N_6961,N_7058);
nand U14692 (N_14692,N_5378,N_6687);
and U14693 (N_14693,N_7787,N_8023);
nand U14694 (N_14694,N_8109,N_6739);
or U14695 (N_14695,N_8402,N_8166);
nand U14696 (N_14696,N_6325,N_5628);
nand U14697 (N_14697,N_7566,N_8693);
nand U14698 (N_14698,N_9682,N_6167);
or U14699 (N_14699,N_5449,N_9156);
and U14700 (N_14700,N_6713,N_9845);
and U14701 (N_14701,N_6020,N_6836);
and U14702 (N_14702,N_6891,N_8483);
or U14703 (N_14703,N_8224,N_6737);
nand U14704 (N_14704,N_8299,N_5143);
and U14705 (N_14705,N_6529,N_8067);
nand U14706 (N_14706,N_7479,N_8744);
and U14707 (N_14707,N_9523,N_6924);
nand U14708 (N_14708,N_9658,N_8600);
and U14709 (N_14709,N_9007,N_9161);
and U14710 (N_14710,N_9131,N_6071);
or U14711 (N_14711,N_9145,N_7750);
nand U14712 (N_14712,N_9220,N_7793);
or U14713 (N_14713,N_8456,N_6399);
and U14714 (N_14714,N_5412,N_6835);
nand U14715 (N_14715,N_7644,N_5927);
nor U14716 (N_14716,N_7458,N_5741);
nand U14717 (N_14717,N_8156,N_6787);
nand U14718 (N_14718,N_8186,N_5859);
nand U14719 (N_14719,N_6320,N_7809);
and U14720 (N_14720,N_6637,N_8720);
and U14721 (N_14721,N_6695,N_6770);
nor U14722 (N_14722,N_7877,N_8761);
or U14723 (N_14723,N_8949,N_7940);
or U14724 (N_14724,N_6398,N_9322);
or U14725 (N_14725,N_8869,N_8279);
nor U14726 (N_14726,N_5026,N_8888);
and U14727 (N_14727,N_5279,N_7445);
nand U14728 (N_14728,N_5397,N_8223);
or U14729 (N_14729,N_9020,N_9583);
nand U14730 (N_14730,N_7822,N_8481);
and U14731 (N_14731,N_6926,N_8046);
and U14732 (N_14732,N_9979,N_6334);
nand U14733 (N_14733,N_7206,N_8052);
and U14734 (N_14734,N_7310,N_5363);
or U14735 (N_14735,N_8373,N_8902);
and U14736 (N_14736,N_8565,N_6428);
or U14737 (N_14737,N_7999,N_6104);
and U14738 (N_14738,N_8162,N_9489);
nand U14739 (N_14739,N_8112,N_6964);
and U14740 (N_14740,N_7650,N_5467);
and U14741 (N_14741,N_8402,N_6368);
nand U14742 (N_14742,N_5200,N_8972);
xnor U14743 (N_14743,N_6156,N_7778);
or U14744 (N_14744,N_7773,N_7892);
and U14745 (N_14745,N_6558,N_5718);
nor U14746 (N_14746,N_8867,N_9073);
and U14747 (N_14747,N_6751,N_8684);
nand U14748 (N_14748,N_7878,N_5951);
nor U14749 (N_14749,N_9014,N_5578);
and U14750 (N_14750,N_5003,N_7696);
nor U14751 (N_14751,N_9861,N_5050);
nand U14752 (N_14752,N_5591,N_8047);
or U14753 (N_14753,N_9092,N_7904);
or U14754 (N_14754,N_5958,N_6670);
nor U14755 (N_14755,N_5361,N_7209);
nor U14756 (N_14756,N_6851,N_6051);
nor U14757 (N_14757,N_7999,N_5127);
nand U14758 (N_14758,N_6117,N_9222);
and U14759 (N_14759,N_7812,N_6716);
xnor U14760 (N_14760,N_5710,N_7334);
and U14761 (N_14761,N_8561,N_5812);
nor U14762 (N_14762,N_7407,N_8710);
and U14763 (N_14763,N_5134,N_6965);
nand U14764 (N_14764,N_8416,N_7806);
and U14765 (N_14765,N_5267,N_8152);
and U14766 (N_14766,N_5824,N_8204);
nor U14767 (N_14767,N_5351,N_9856);
nand U14768 (N_14768,N_5944,N_6618);
nor U14769 (N_14769,N_6039,N_8021);
or U14770 (N_14770,N_5306,N_9498);
nand U14771 (N_14771,N_9472,N_9383);
xor U14772 (N_14772,N_8573,N_5876);
or U14773 (N_14773,N_7549,N_8975);
and U14774 (N_14774,N_7056,N_6643);
nand U14775 (N_14775,N_7668,N_5474);
xnor U14776 (N_14776,N_8854,N_6551);
and U14777 (N_14777,N_5822,N_6259);
nand U14778 (N_14778,N_5518,N_9856);
nor U14779 (N_14779,N_7581,N_6144);
nor U14780 (N_14780,N_7616,N_5236);
and U14781 (N_14781,N_8717,N_8053);
nand U14782 (N_14782,N_7328,N_7172);
or U14783 (N_14783,N_8793,N_8169);
nand U14784 (N_14784,N_9638,N_7055);
nor U14785 (N_14785,N_5885,N_9365);
and U14786 (N_14786,N_8784,N_6495);
xor U14787 (N_14787,N_7566,N_9332);
nor U14788 (N_14788,N_8597,N_7530);
or U14789 (N_14789,N_9747,N_6934);
xor U14790 (N_14790,N_9714,N_5332);
or U14791 (N_14791,N_7365,N_7292);
nor U14792 (N_14792,N_7353,N_7680);
and U14793 (N_14793,N_9521,N_5821);
xnor U14794 (N_14794,N_6955,N_7110);
or U14795 (N_14795,N_5155,N_6762);
or U14796 (N_14796,N_5418,N_6041);
nor U14797 (N_14797,N_7419,N_8858);
xnor U14798 (N_14798,N_7971,N_6901);
or U14799 (N_14799,N_5010,N_9547);
nand U14800 (N_14800,N_9507,N_6053);
nand U14801 (N_14801,N_8127,N_6340);
nor U14802 (N_14802,N_8055,N_7223);
nor U14803 (N_14803,N_5697,N_9223);
or U14804 (N_14804,N_7177,N_7085);
or U14805 (N_14805,N_8491,N_7296);
and U14806 (N_14806,N_7726,N_9206);
and U14807 (N_14807,N_5970,N_8061);
and U14808 (N_14808,N_6862,N_8209);
nor U14809 (N_14809,N_8355,N_8046);
xor U14810 (N_14810,N_5069,N_9892);
and U14811 (N_14811,N_8717,N_8589);
xor U14812 (N_14812,N_8594,N_6951);
or U14813 (N_14813,N_6290,N_9370);
or U14814 (N_14814,N_7836,N_7230);
xor U14815 (N_14815,N_6175,N_9954);
or U14816 (N_14816,N_7753,N_7349);
xnor U14817 (N_14817,N_7972,N_9352);
nand U14818 (N_14818,N_8692,N_8746);
or U14819 (N_14819,N_9975,N_7717);
and U14820 (N_14820,N_6007,N_7847);
nand U14821 (N_14821,N_8632,N_7182);
and U14822 (N_14822,N_8831,N_7132);
or U14823 (N_14823,N_9497,N_8910);
and U14824 (N_14824,N_6000,N_8184);
nand U14825 (N_14825,N_6321,N_7954);
and U14826 (N_14826,N_9127,N_7572);
xor U14827 (N_14827,N_8219,N_8097);
nand U14828 (N_14828,N_7331,N_6470);
and U14829 (N_14829,N_8120,N_5426);
nand U14830 (N_14830,N_8416,N_6051);
nand U14831 (N_14831,N_6720,N_5247);
nor U14832 (N_14832,N_5893,N_9094);
nor U14833 (N_14833,N_6071,N_8454);
or U14834 (N_14834,N_5963,N_7335);
and U14835 (N_14835,N_9480,N_7834);
or U14836 (N_14836,N_9456,N_9363);
nand U14837 (N_14837,N_7755,N_6313);
nor U14838 (N_14838,N_7692,N_9281);
nor U14839 (N_14839,N_6203,N_9402);
and U14840 (N_14840,N_9847,N_8765);
nand U14841 (N_14841,N_9173,N_9575);
and U14842 (N_14842,N_8453,N_8192);
nor U14843 (N_14843,N_9276,N_6509);
and U14844 (N_14844,N_6057,N_5459);
or U14845 (N_14845,N_6562,N_6149);
xor U14846 (N_14846,N_7351,N_8216);
nand U14847 (N_14847,N_9633,N_7605);
and U14848 (N_14848,N_5243,N_6900);
nand U14849 (N_14849,N_9038,N_6835);
nor U14850 (N_14850,N_8667,N_8331);
and U14851 (N_14851,N_6366,N_7417);
nand U14852 (N_14852,N_5539,N_9541);
nand U14853 (N_14853,N_9471,N_5688);
nand U14854 (N_14854,N_9732,N_6929);
nand U14855 (N_14855,N_8090,N_5897);
and U14856 (N_14856,N_7185,N_6200);
and U14857 (N_14857,N_6255,N_6302);
or U14858 (N_14858,N_9936,N_9791);
nor U14859 (N_14859,N_9406,N_9153);
or U14860 (N_14860,N_7665,N_6971);
xnor U14861 (N_14861,N_9181,N_7118);
or U14862 (N_14862,N_7546,N_6747);
nand U14863 (N_14863,N_5299,N_8818);
nand U14864 (N_14864,N_6988,N_9052);
nor U14865 (N_14865,N_7941,N_9511);
nor U14866 (N_14866,N_6840,N_7552);
xnor U14867 (N_14867,N_6980,N_8479);
xnor U14868 (N_14868,N_7967,N_7452);
or U14869 (N_14869,N_9526,N_8040);
and U14870 (N_14870,N_9164,N_5267);
and U14871 (N_14871,N_8320,N_5435);
and U14872 (N_14872,N_5125,N_8294);
nor U14873 (N_14873,N_9670,N_6530);
nand U14874 (N_14874,N_6838,N_6385);
nand U14875 (N_14875,N_9969,N_8388);
xnor U14876 (N_14876,N_6415,N_8702);
nor U14877 (N_14877,N_9896,N_8871);
and U14878 (N_14878,N_6368,N_9274);
or U14879 (N_14879,N_7716,N_5852);
or U14880 (N_14880,N_8783,N_6615);
nor U14881 (N_14881,N_5838,N_7386);
and U14882 (N_14882,N_9946,N_5703);
nand U14883 (N_14883,N_6948,N_6788);
nand U14884 (N_14884,N_6986,N_8390);
nand U14885 (N_14885,N_6469,N_7668);
or U14886 (N_14886,N_8371,N_5769);
xnor U14887 (N_14887,N_5963,N_7183);
nand U14888 (N_14888,N_9285,N_7261);
nor U14889 (N_14889,N_5171,N_8063);
or U14890 (N_14890,N_6139,N_5335);
or U14891 (N_14891,N_9991,N_8718);
nand U14892 (N_14892,N_9455,N_5223);
nand U14893 (N_14893,N_6364,N_7726);
nand U14894 (N_14894,N_5981,N_9465);
or U14895 (N_14895,N_7148,N_7142);
nor U14896 (N_14896,N_8223,N_5420);
nand U14897 (N_14897,N_8575,N_9303);
and U14898 (N_14898,N_6192,N_7229);
nor U14899 (N_14899,N_7419,N_8357);
nor U14900 (N_14900,N_5236,N_5142);
or U14901 (N_14901,N_9792,N_8552);
and U14902 (N_14902,N_7403,N_8270);
and U14903 (N_14903,N_9475,N_7168);
or U14904 (N_14904,N_7705,N_5182);
or U14905 (N_14905,N_5886,N_6152);
and U14906 (N_14906,N_5696,N_9310);
or U14907 (N_14907,N_8642,N_8695);
nand U14908 (N_14908,N_9449,N_7767);
and U14909 (N_14909,N_7251,N_7456);
xor U14910 (N_14910,N_9164,N_8262);
nor U14911 (N_14911,N_7417,N_6983);
nor U14912 (N_14912,N_6591,N_6930);
nand U14913 (N_14913,N_6602,N_7191);
nor U14914 (N_14914,N_5615,N_8711);
and U14915 (N_14915,N_6438,N_8572);
nand U14916 (N_14916,N_9163,N_5119);
nor U14917 (N_14917,N_8902,N_8234);
xnor U14918 (N_14918,N_8370,N_6133);
or U14919 (N_14919,N_5067,N_6478);
or U14920 (N_14920,N_9373,N_9715);
nand U14921 (N_14921,N_5174,N_5636);
xor U14922 (N_14922,N_7329,N_8002);
or U14923 (N_14923,N_7329,N_7201);
or U14924 (N_14924,N_5851,N_5788);
or U14925 (N_14925,N_6337,N_6907);
or U14926 (N_14926,N_5097,N_8190);
nor U14927 (N_14927,N_6966,N_9458);
nor U14928 (N_14928,N_7851,N_6508);
nor U14929 (N_14929,N_6953,N_5095);
nand U14930 (N_14930,N_5865,N_8761);
nor U14931 (N_14931,N_5505,N_9050);
xor U14932 (N_14932,N_7220,N_5359);
and U14933 (N_14933,N_5428,N_5052);
nor U14934 (N_14934,N_5974,N_7158);
or U14935 (N_14935,N_6748,N_7008);
nor U14936 (N_14936,N_5890,N_6020);
and U14937 (N_14937,N_9694,N_5529);
nor U14938 (N_14938,N_8802,N_6394);
nor U14939 (N_14939,N_7890,N_6624);
nor U14940 (N_14940,N_6122,N_5458);
nor U14941 (N_14941,N_8403,N_5765);
and U14942 (N_14942,N_9660,N_6156);
or U14943 (N_14943,N_5892,N_6848);
nand U14944 (N_14944,N_8699,N_6519);
and U14945 (N_14945,N_5185,N_9550);
or U14946 (N_14946,N_7760,N_7058);
or U14947 (N_14947,N_9569,N_5891);
nor U14948 (N_14948,N_6717,N_6207);
or U14949 (N_14949,N_7481,N_8107);
nand U14950 (N_14950,N_7783,N_6678);
nor U14951 (N_14951,N_9369,N_7893);
and U14952 (N_14952,N_6837,N_9142);
and U14953 (N_14953,N_6751,N_5622);
and U14954 (N_14954,N_5179,N_8415);
nor U14955 (N_14955,N_5106,N_6755);
and U14956 (N_14956,N_9108,N_9504);
nor U14957 (N_14957,N_6081,N_8448);
nor U14958 (N_14958,N_9664,N_6744);
and U14959 (N_14959,N_7604,N_8624);
or U14960 (N_14960,N_7095,N_9396);
and U14961 (N_14961,N_8227,N_5149);
or U14962 (N_14962,N_8021,N_8457);
nor U14963 (N_14963,N_5823,N_5733);
nor U14964 (N_14964,N_9957,N_5138);
or U14965 (N_14965,N_6778,N_5699);
nor U14966 (N_14966,N_9839,N_8657);
or U14967 (N_14967,N_6873,N_7900);
and U14968 (N_14968,N_9508,N_8649);
or U14969 (N_14969,N_8214,N_7265);
nor U14970 (N_14970,N_7891,N_6891);
nand U14971 (N_14971,N_5317,N_5242);
nor U14972 (N_14972,N_6133,N_7981);
and U14973 (N_14973,N_6043,N_5404);
xor U14974 (N_14974,N_8688,N_7144);
xor U14975 (N_14975,N_8708,N_8024);
xnor U14976 (N_14976,N_6698,N_8037);
and U14977 (N_14977,N_9542,N_9906);
nor U14978 (N_14978,N_5095,N_9983);
nor U14979 (N_14979,N_7152,N_9440);
and U14980 (N_14980,N_8055,N_8065);
nand U14981 (N_14981,N_8411,N_7508);
nand U14982 (N_14982,N_7677,N_8641);
or U14983 (N_14983,N_7669,N_7432);
nand U14984 (N_14984,N_6094,N_6870);
nor U14985 (N_14985,N_7247,N_7219);
nor U14986 (N_14986,N_7804,N_6643);
nor U14987 (N_14987,N_7505,N_6946);
xnor U14988 (N_14988,N_8566,N_8000);
or U14989 (N_14989,N_9462,N_7163);
nor U14990 (N_14990,N_5427,N_9554);
or U14991 (N_14991,N_7650,N_5362);
nor U14992 (N_14992,N_6201,N_5367);
nor U14993 (N_14993,N_9251,N_8856);
nand U14994 (N_14994,N_9404,N_7632);
or U14995 (N_14995,N_9698,N_9678);
and U14996 (N_14996,N_5326,N_8738);
nor U14997 (N_14997,N_6606,N_9236);
and U14998 (N_14998,N_6260,N_8245);
nand U14999 (N_14999,N_7286,N_9230);
and U15000 (N_15000,N_14426,N_14004);
nor U15001 (N_15001,N_10118,N_11019);
and U15002 (N_15002,N_12203,N_14574);
or U15003 (N_15003,N_10780,N_14363);
and U15004 (N_15004,N_11062,N_10439);
or U15005 (N_15005,N_13197,N_12641);
nand U15006 (N_15006,N_12884,N_12951);
xnor U15007 (N_15007,N_13145,N_10239);
nor U15008 (N_15008,N_10444,N_11191);
or U15009 (N_15009,N_12300,N_14793);
nand U15010 (N_15010,N_12405,N_13712);
nand U15011 (N_15011,N_11307,N_12936);
or U15012 (N_15012,N_14951,N_14115);
xnor U15013 (N_15013,N_14029,N_10116);
xnor U15014 (N_15014,N_14428,N_14932);
nand U15015 (N_15015,N_14403,N_10272);
nand U15016 (N_15016,N_13074,N_12858);
nand U15017 (N_15017,N_10809,N_11247);
or U15018 (N_15018,N_10174,N_14388);
nor U15019 (N_15019,N_13891,N_10996);
nor U15020 (N_15020,N_13165,N_13771);
or U15021 (N_15021,N_14696,N_10514);
nor U15022 (N_15022,N_12989,N_13623);
and U15023 (N_15023,N_14617,N_12607);
nand U15024 (N_15024,N_13783,N_10521);
or U15025 (N_15025,N_13268,N_13386);
and U15026 (N_15026,N_13099,N_10518);
or U15027 (N_15027,N_11477,N_14781);
or U15028 (N_15028,N_10900,N_11718);
and U15029 (N_15029,N_12412,N_11230);
and U15030 (N_15030,N_14745,N_13740);
nor U15031 (N_15031,N_12679,N_13034);
or U15032 (N_15032,N_12584,N_14087);
nor U15033 (N_15033,N_13897,N_10488);
nand U15034 (N_15034,N_13104,N_12207);
and U15035 (N_15035,N_14083,N_13028);
nor U15036 (N_15036,N_11172,N_14066);
nor U15037 (N_15037,N_13179,N_10123);
nor U15038 (N_15038,N_14643,N_10148);
or U15039 (N_15039,N_13300,N_10534);
or U15040 (N_15040,N_14054,N_12236);
and U15041 (N_15041,N_12482,N_13661);
xnor U15042 (N_15042,N_11156,N_10293);
nor U15043 (N_15043,N_10924,N_14436);
or U15044 (N_15044,N_10867,N_10283);
xor U15045 (N_15045,N_10258,N_11335);
nor U15046 (N_15046,N_11023,N_11933);
nand U15047 (N_15047,N_12291,N_13142);
nor U15048 (N_15048,N_14693,N_11236);
xor U15049 (N_15049,N_10397,N_14190);
nand U15050 (N_15050,N_11492,N_13143);
and U15051 (N_15051,N_11640,N_12760);
nand U15052 (N_15052,N_13285,N_14979);
nand U15053 (N_15053,N_10964,N_11356);
nor U15054 (N_15054,N_14369,N_10940);
nor U15055 (N_15055,N_11420,N_10250);
nor U15056 (N_15056,N_11138,N_10413);
nand U15057 (N_15057,N_13475,N_14763);
or U15058 (N_15058,N_10385,N_14233);
nand U15059 (N_15059,N_10192,N_13789);
or U15060 (N_15060,N_10510,N_12504);
and U15061 (N_15061,N_12838,N_11700);
xnor U15062 (N_15062,N_10628,N_11692);
nor U15063 (N_15063,N_10841,N_13177);
nor U15064 (N_15064,N_10898,N_10217);
nand U15065 (N_15065,N_11174,N_10794);
nor U15066 (N_15066,N_10237,N_13080);
and U15067 (N_15067,N_10117,N_10374);
xor U15068 (N_15068,N_10332,N_11865);
xor U15069 (N_15069,N_12536,N_12588);
nand U15070 (N_15070,N_11800,N_13590);
nor U15071 (N_15071,N_11665,N_11158);
nand U15072 (N_15072,N_14479,N_12010);
and U15073 (N_15073,N_14117,N_14450);
xnor U15074 (N_15074,N_10008,N_11602);
nor U15075 (N_15075,N_11581,N_10960);
nand U15076 (N_15076,N_10540,N_13108);
or U15077 (N_15077,N_14618,N_11040);
nor U15078 (N_15078,N_13322,N_13186);
and U15079 (N_15079,N_10543,N_13530);
or U15080 (N_15080,N_11292,N_14179);
xor U15081 (N_15081,N_14641,N_14442);
and U15082 (N_15082,N_11661,N_10705);
xor U15083 (N_15083,N_10456,N_14760);
nand U15084 (N_15084,N_12923,N_10464);
nor U15085 (N_15085,N_12514,N_14331);
or U15086 (N_15086,N_10222,N_11945);
and U15087 (N_15087,N_14678,N_12628);
nor U15088 (N_15088,N_12888,N_13121);
or U15089 (N_15089,N_13470,N_10766);
xor U15090 (N_15090,N_10104,N_12998);
nor U15091 (N_15091,N_13782,N_14989);
or U15092 (N_15092,N_13601,N_12167);
xor U15093 (N_15093,N_11784,N_14882);
nand U15094 (N_15094,N_11900,N_11251);
nand U15095 (N_15095,N_11862,N_12810);
nor U15096 (N_15096,N_12900,N_11810);
and U15097 (N_15097,N_10015,N_13125);
nor U15098 (N_15098,N_11179,N_11636);
or U15099 (N_15099,N_10102,N_12154);
nand U15100 (N_15100,N_14326,N_10695);
nand U15101 (N_15101,N_13954,N_10531);
nor U15102 (N_15102,N_12052,N_12713);
and U15103 (N_15103,N_10496,N_14782);
or U15104 (N_15104,N_14024,N_14431);
nor U15105 (N_15105,N_12809,N_11280);
and U15106 (N_15106,N_10775,N_13428);
xor U15107 (N_15107,N_12460,N_11978);
nand U15108 (N_15108,N_14320,N_11165);
nand U15109 (N_15109,N_13249,N_14134);
nand U15110 (N_15110,N_12078,N_13633);
nor U15111 (N_15111,N_11697,N_13335);
nor U15112 (N_15112,N_11837,N_13963);
nand U15113 (N_15113,N_12781,N_12136);
xnor U15114 (N_15114,N_11791,N_11631);
nor U15115 (N_15115,N_10181,N_13657);
or U15116 (N_15116,N_10714,N_14988);
nor U15117 (N_15117,N_12107,N_10090);
or U15118 (N_15118,N_11128,N_10952);
nand U15119 (N_15119,N_14525,N_10536);
and U15120 (N_15120,N_12689,N_11396);
nand U15121 (N_15121,N_12761,N_10732);
nand U15122 (N_15122,N_12876,N_10834);
or U15123 (N_15123,N_11495,N_10939);
and U15124 (N_15124,N_12083,N_13224);
and U15125 (N_15125,N_13372,N_11599);
nand U15126 (N_15126,N_11888,N_13157);
xnor U15127 (N_15127,N_13962,N_10388);
nor U15128 (N_15128,N_12750,N_10870);
or U15129 (N_15129,N_11662,N_13917);
or U15130 (N_15130,N_11695,N_12836);
nand U15131 (N_15131,N_10314,N_14173);
or U15132 (N_15132,N_11184,N_14018);
nand U15133 (N_15133,N_10596,N_12963);
or U15134 (N_15134,N_11159,N_10369);
nor U15135 (N_15135,N_14516,N_10143);
nand U15136 (N_15136,N_13815,N_12293);
or U15137 (N_15137,N_14182,N_10055);
and U15138 (N_15138,N_10083,N_10031);
xnor U15139 (N_15139,N_14774,N_14455);
nand U15140 (N_15140,N_12341,N_13799);
nand U15141 (N_15141,N_12674,N_14315);
and U15142 (N_15142,N_12583,N_14299);
nor U15143 (N_15143,N_13884,N_12671);
nor U15144 (N_15144,N_12979,N_14538);
nand U15145 (N_15145,N_12687,N_11099);
or U15146 (N_15146,N_11368,N_13619);
nand U15147 (N_15147,N_10884,N_12110);
and U15148 (N_15148,N_11459,N_10773);
and U15149 (N_15149,N_12946,N_12443);
or U15150 (N_15150,N_11821,N_10264);
or U15151 (N_15151,N_12498,N_10709);
nand U15152 (N_15152,N_11219,N_10934);
or U15153 (N_15153,N_12099,N_11234);
or U15154 (N_15154,N_11067,N_11827);
and U15155 (N_15155,N_10538,N_12673);
and U15156 (N_15156,N_13925,N_12367);
or U15157 (N_15157,N_12731,N_11095);
nand U15158 (N_15158,N_13187,N_10893);
and U15159 (N_15159,N_13902,N_11507);
nor U15160 (N_15160,N_13461,N_11363);
nand U15161 (N_15161,N_11135,N_14500);
nor U15162 (N_15162,N_10615,N_14990);
nor U15163 (N_15163,N_13120,N_12200);
nor U15164 (N_15164,N_12224,N_14832);
or U15165 (N_15165,N_11373,N_12666);
and U15166 (N_15166,N_13752,N_11263);
or U15167 (N_15167,N_14602,N_14293);
nor U15168 (N_15168,N_11160,N_14692);
nand U15169 (N_15169,N_14681,N_12239);
nor U15170 (N_15170,N_12407,N_13246);
nor U15171 (N_15171,N_13026,N_11444);
and U15172 (N_15172,N_14942,N_11087);
nor U15173 (N_15173,N_14999,N_14568);
xor U15174 (N_15174,N_12592,N_10390);
nand U15175 (N_15175,N_14978,N_13149);
or U15176 (N_15176,N_13214,N_12327);
nor U15177 (N_15177,N_11613,N_11090);
and U15178 (N_15178,N_10600,N_11327);
or U15179 (N_15179,N_11248,N_11468);
nand U15180 (N_15180,N_14532,N_13404);
nand U15181 (N_15181,N_12304,N_13959);
and U15182 (N_15182,N_12613,N_11555);
nand U15183 (N_15183,N_13083,N_14583);
nand U15184 (N_15184,N_12863,N_13573);
nor U15185 (N_15185,N_14223,N_13044);
nand U15186 (N_15186,N_10172,N_13556);
xnor U15187 (N_15187,N_12318,N_13443);
or U15188 (N_15188,N_13260,N_10001);
nand U15189 (N_15189,N_11673,N_10259);
or U15190 (N_15190,N_12508,N_11473);
and U15191 (N_15191,N_14160,N_12262);
and U15192 (N_15192,N_11809,N_12567);
or U15193 (N_15193,N_12399,N_13881);
nor U15194 (N_15194,N_13585,N_11134);
xor U15195 (N_15195,N_10957,N_12901);
nand U15196 (N_15196,N_11104,N_14171);
and U15197 (N_15197,N_12438,N_13354);
and U15198 (N_15198,N_10970,N_11276);
and U15199 (N_15199,N_10204,N_10299);
and U15200 (N_15200,N_12701,N_12112);
or U15201 (N_15201,N_13856,N_14199);
and U15202 (N_15202,N_11007,N_12181);
and U15203 (N_15203,N_10356,N_10120);
nand U15204 (N_15204,N_11180,N_12094);
nand U15205 (N_15205,N_10618,N_14755);
nor U15206 (N_15206,N_13073,N_13251);
or U15207 (N_15207,N_11188,N_10214);
nor U15208 (N_15208,N_12379,N_12226);
or U15209 (N_15209,N_13489,N_10096);
xor U15210 (N_15210,N_10985,N_14127);
nand U15211 (N_15211,N_11683,N_10159);
nand U15212 (N_15212,N_10820,N_10489);
nor U15213 (N_15213,N_13367,N_11585);
nor U15214 (N_15214,N_13781,N_11163);
nand U15215 (N_15215,N_13818,N_10984);
nor U15216 (N_15216,N_14048,N_14256);
or U15217 (N_15217,N_11565,N_14178);
nor U15218 (N_15218,N_12287,N_12615);
nand U15219 (N_15219,N_11947,N_13445);
nor U15220 (N_15220,N_11445,N_10682);
nor U15221 (N_15221,N_12550,N_10410);
or U15222 (N_15222,N_11244,N_10650);
nand U15223 (N_15223,N_13040,N_13765);
nor U15224 (N_15224,N_14174,N_13022);
and U15225 (N_15225,N_10469,N_14187);
and U15226 (N_15226,N_10125,N_13773);
or U15227 (N_15227,N_11824,N_12736);
nand U15228 (N_15228,N_10247,N_11469);
xnor U15229 (N_15229,N_14152,N_13613);
nand U15230 (N_15230,N_11657,N_12012);
and U15231 (N_15231,N_12416,N_14820);
nand U15232 (N_15232,N_14950,N_11975);
nand U15233 (N_15233,N_11534,N_11932);
or U15234 (N_15234,N_10895,N_13020);
nand U15235 (N_15235,N_12845,N_10516);
nand U15236 (N_15236,N_10022,N_10178);
nand U15237 (N_15237,N_13532,N_12653);
nor U15238 (N_15238,N_13518,N_14579);
nand U15239 (N_15239,N_11702,N_12138);
xor U15240 (N_15240,N_10923,N_11788);
nor U15241 (N_15241,N_11488,N_13041);
or U15242 (N_15242,N_12530,N_11301);
nand U15243 (N_15243,N_12120,N_13628);
or U15244 (N_15244,N_12437,N_14778);
nand U15245 (N_15245,N_11310,N_14414);
nor U15246 (N_15246,N_14281,N_12101);
nand U15247 (N_15247,N_10045,N_14305);
and U15248 (N_15248,N_12413,N_14239);
xor U15249 (N_15249,N_12074,N_12216);
nand U15250 (N_15250,N_14056,N_12204);
nor U15251 (N_15251,N_11034,N_12883);
nor U15252 (N_15252,N_14548,N_14580);
and U15253 (N_15253,N_13229,N_10325);
or U15254 (N_15254,N_11238,N_11653);
nand U15255 (N_15255,N_12077,N_14886);
and U15256 (N_15256,N_10784,N_11740);
nand U15257 (N_15257,N_14298,N_12543);
and U15258 (N_15258,N_14786,N_12643);
or U15259 (N_15259,N_12507,N_11408);
and U15260 (N_15260,N_12213,N_11890);
and U15261 (N_15261,N_12091,N_12685);
nor U15262 (N_15262,N_13349,N_13792);
nand U15263 (N_15263,N_12335,N_14013);
or U15264 (N_15264,N_10868,N_13727);
xor U15265 (N_15265,N_14228,N_13172);
nor U15266 (N_15266,N_11765,N_11329);
nand U15267 (N_15267,N_14207,N_12124);
nand U15268 (N_15268,N_10508,N_12307);
and U15269 (N_15269,N_11604,N_10943);
and U15270 (N_15270,N_14433,N_13930);
and U15271 (N_15271,N_12055,N_11915);
nand U15272 (N_15272,N_13469,N_14615);
nand U15273 (N_15273,N_14992,N_10737);
and U15274 (N_15274,N_12886,N_12002);
nor U15275 (N_15275,N_10630,N_12965);
or U15276 (N_15276,N_13648,N_12813);
nor U15277 (N_15277,N_10589,N_14088);
xor U15278 (N_15278,N_14789,N_12904);
nor U15279 (N_15279,N_10739,N_12126);
nor U15280 (N_15280,N_10762,N_10954);
nor U15281 (N_15281,N_13943,N_11762);
xor U15282 (N_15282,N_11232,N_13638);
nand U15283 (N_15283,N_11588,N_10398);
xor U15284 (N_15284,N_11654,N_13766);
or U15285 (N_15285,N_11037,N_10209);
or U15286 (N_15286,N_12991,N_12678);
xnor U15287 (N_15287,N_10046,N_14954);
or U15288 (N_15288,N_14032,N_10885);
xnor U15289 (N_15289,N_11305,N_12113);
nor U15290 (N_15290,N_12920,N_10224);
or U15291 (N_15291,N_11928,N_14716);
xor U15292 (N_15292,N_13205,N_13013);
nand U15293 (N_15293,N_10016,N_10462);
and U15294 (N_15294,N_14652,N_10335);
nand U15295 (N_15295,N_10161,N_10294);
or U15296 (N_15296,N_11253,N_10476);
nand U15297 (N_15297,N_10065,N_13018);
and U15298 (N_15298,N_13745,N_10207);
and U15299 (N_15299,N_10763,N_11167);
nand U15300 (N_15300,N_13284,N_13681);
nor U15301 (N_15301,N_10504,N_14116);
and U15302 (N_15302,N_12425,N_14855);
nand U15303 (N_15303,N_13868,N_11887);
xnor U15304 (N_15304,N_14427,N_13112);
nor U15305 (N_15305,N_14588,N_12048);
and U15306 (N_15306,N_14219,N_14539);
nor U15307 (N_15307,N_12245,N_10837);
nor U15308 (N_15308,N_13595,N_14661);
and U15309 (N_15309,N_12746,N_11993);
and U15310 (N_15310,N_12131,N_14959);
nor U15311 (N_15311,N_10134,N_14265);
or U15312 (N_15312,N_12569,N_10640);
and U15313 (N_15313,N_11794,N_11027);
nor U15314 (N_15314,N_14139,N_14873);
nand U15315 (N_15315,N_12468,N_13786);
nor U15316 (N_15316,N_12410,N_14845);
nand U15317 (N_15317,N_11761,N_12987);
nand U15318 (N_15318,N_13291,N_13705);
nor U15319 (N_15319,N_13975,N_11483);
nor U15320 (N_15320,N_14600,N_12559);
nor U15321 (N_15321,N_12452,N_11691);
or U15322 (N_15322,N_10481,N_10583);
nand U15323 (N_15323,N_12414,N_11807);
and U15324 (N_15324,N_13473,N_13694);
xor U15325 (N_15325,N_13821,N_10030);
nor U15326 (N_15326,N_11851,N_12068);
nor U15327 (N_15327,N_14266,N_13506);
and U15328 (N_15328,N_13813,N_13846);
and U15329 (N_15329,N_11484,N_13418);
and U15330 (N_15330,N_12800,N_13690);
nand U15331 (N_15331,N_10693,N_12576);
nand U15332 (N_15332,N_13774,N_12037);
nand U15333 (N_15333,N_11460,N_14475);
nand U15334 (N_15334,N_13071,N_11053);
xor U15335 (N_15335,N_14451,N_14561);
or U15336 (N_15336,N_13547,N_12486);
or U15337 (N_15337,N_10344,N_12422);
and U15338 (N_15338,N_14853,N_13275);
nand U15339 (N_15339,N_12669,N_12652);
nor U15340 (N_15340,N_10563,N_11441);
nor U15341 (N_15341,N_10855,N_11709);
or U15342 (N_15342,N_13222,N_10231);
or U15343 (N_15343,N_13934,N_12342);
nand U15344 (N_15344,N_13411,N_13751);
nor U15345 (N_15345,N_13841,N_13524);
nand U15346 (N_15346,N_11437,N_12523);
nand U15347 (N_15347,N_12476,N_10770);
nand U15348 (N_15348,N_11514,N_13481);
or U15349 (N_15349,N_12839,N_14981);
nor U15350 (N_15350,N_10429,N_10494);
or U15351 (N_15351,N_11557,N_11463);
and U15352 (N_15352,N_13696,N_14260);
and U15353 (N_15353,N_11024,N_10017);
or U15354 (N_15354,N_13167,N_11838);
and U15355 (N_15355,N_11717,N_12457);
and U15356 (N_15356,N_11619,N_10499);
or U15357 (N_15357,N_14161,N_13414);
or U15358 (N_15358,N_12996,N_12006);
xnor U15359 (N_15359,N_12034,N_10570);
nor U15360 (N_15360,N_13769,N_12295);
xor U15361 (N_15361,N_13181,N_11752);
or U15362 (N_15362,N_13651,N_14371);
nor U15363 (N_15363,N_11202,N_10533);
or U15364 (N_15364,N_11705,N_12784);
and U15365 (N_15365,N_12719,N_14841);
nor U15366 (N_15366,N_13989,N_12390);
nand U15367 (N_15367,N_11586,N_14528);
nor U15368 (N_15368,N_11913,N_12690);
or U15369 (N_15369,N_13265,N_11927);
nor U15370 (N_15370,N_13049,N_12696);
and U15371 (N_15371,N_11750,N_14237);
nor U15372 (N_15372,N_11907,N_13931);
or U15373 (N_15373,N_10180,N_14708);
or U15374 (N_15374,N_11112,N_11073);
and U15375 (N_15375,N_10613,N_12029);
or U15376 (N_15376,N_12645,N_11001);
nor U15377 (N_15377,N_13327,N_12532);
nand U15378 (N_15378,N_13816,N_14075);
nand U15379 (N_15379,N_10111,N_13425);
nand U15380 (N_15380,N_13134,N_10882);
or U15381 (N_15381,N_10480,N_11342);
nor U15382 (N_15382,N_12235,N_13641);
or U15383 (N_15383,N_11031,N_14498);
or U15384 (N_15384,N_13620,N_10070);
nand U15385 (N_15385,N_12521,N_10292);
nor U15386 (N_15386,N_13070,N_10158);
nor U15387 (N_15387,N_12528,N_13048);
nand U15388 (N_15388,N_13699,N_14278);
nand U15389 (N_15389,N_14731,N_11245);
xnor U15390 (N_15390,N_14404,N_10750);
or U15391 (N_15391,N_12714,N_13598);
nor U15392 (N_15392,N_10389,N_12419);
nor U15393 (N_15393,N_11523,N_13755);
nand U15394 (N_15394,N_14819,N_14076);
and U15395 (N_15395,N_12925,N_13296);
nor U15396 (N_15396,N_12475,N_12357);
and U15397 (N_15397,N_11898,N_12531);
nor U15398 (N_15398,N_11412,N_10297);
and U15399 (N_15399,N_12111,N_14750);
nor U15400 (N_15400,N_13981,N_10745);
nor U15401 (N_15401,N_14595,N_10561);
or U15402 (N_15402,N_12539,N_14499);
or U15403 (N_15403,N_10170,N_10564);
nand U15404 (N_15404,N_11689,N_14826);
and U15405 (N_15405,N_11286,N_10490);
nand U15406 (N_15406,N_14672,N_12095);
or U15407 (N_15407,N_10680,N_11340);
nor U15408 (N_15408,N_11883,N_11341);
nand U15409 (N_15409,N_11686,N_13715);
or U15410 (N_15410,N_10616,N_10273);
or U15411 (N_15411,N_12620,N_14858);
or U15412 (N_15412,N_13767,N_13419);
and U15413 (N_15413,N_12082,N_14700);
or U15414 (N_15414,N_14145,N_10189);
or U15415 (N_15415,N_11731,N_11541);
nor U15416 (N_15416,N_10528,N_14245);
nor U15417 (N_15417,N_11980,N_10131);
and U15418 (N_15418,N_10727,N_13310);
and U15419 (N_15419,N_10326,N_10696);
and U15420 (N_15420,N_14898,N_14202);
nor U15421 (N_15421,N_12887,N_11852);
nor U15422 (N_15422,N_10691,N_11061);
and U15423 (N_15423,N_11083,N_11597);
nand U15424 (N_15424,N_12032,N_12171);
nand U15425 (N_15425,N_13045,N_14146);
nand U15426 (N_15426,N_12593,N_12747);
nand U15427 (N_15427,N_12259,N_10077);
nor U15428 (N_15428,N_14509,N_11096);
nor U15429 (N_15429,N_12162,N_11777);
xnor U15430 (N_15430,N_12088,N_11759);
and U15431 (N_15431,N_12520,N_12743);
and U15432 (N_15432,N_13169,N_13163);
nand U15433 (N_15433,N_14552,N_11211);
and U15434 (N_15434,N_10886,N_11311);
and U15435 (N_15435,N_13117,N_14495);
nand U15436 (N_15436,N_14365,N_12054);
and U15437 (N_15437,N_14586,N_14476);
nor U15438 (N_15438,N_13288,N_11707);
or U15439 (N_15439,N_12166,N_11331);
and U15440 (N_15440,N_13242,N_10132);
nand U15441 (N_15441,N_11434,N_12090);
nor U15442 (N_15442,N_11751,N_12591);
or U15443 (N_15443,N_10874,N_14733);
nand U15444 (N_15444,N_14271,N_14645);
or U15445 (N_15445,N_13379,N_13314);
nand U15446 (N_15446,N_10274,N_11598);
nor U15447 (N_15447,N_11231,N_14412);
or U15448 (N_15448,N_12336,N_12121);
and U15449 (N_15449,N_13225,N_14947);
nand U15450 (N_15450,N_11387,N_12815);
or U15451 (N_15451,N_14550,N_10427);
or U15452 (N_15452,N_12629,N_13286);
nand U15453 (N_15453,N_13665,N_12829);
nand U15454 (N_15454,N_14135,N_10721);
and U15455 (N_15455,N_12169,N_14071);
and U15456 (N_15456,N_12982,N_13678);
nor U15457 (N_15457,N_12477,N_10251);
xnor U15458 (N_15458,N_10415,N_12223);
or U15459 (N_15459,N_12267,N_14776);
and U15460 (N_15460,N_14554,N_11461);
or U15461 (N_15461,N_13682,N_14148);
or U15462 (N_15462,N_13780,N_10730);
or U15463 (N_15463,N_13292,N_11351);
nor U15464 (N_15464,N_11935,N_12377);
or U15465 (N_15465,N_12408,N_10084);
or U15466 (N_15466,N_13199,N_14168);
and U15467 (N_15467,N_13184,N_13339);
nand U15468 (N_15468,N_13869,N_14899);
or U15469 (N_15469,N_13733,N_13521);
nand U15470 (N_15470,N_10553,N_12970);
nand U15471 (N_15471,N_10002,N_14710);
nand U15472 (N_15472,N_11267,N_12465);
or U15473 (N_15473,N_11166,N_13534);
nand U15474 (N_15474,N_14732,N_10162);
and U15475 (N_15475,N_13876,N_12495);
nor U15476 (N_15476,N_14280,N_14683);
nor U15477 (N_15477,N_13173,N_10992);
or U15478 (N_15478,N_13839,N_12041);
and U15479 (N_15479,N_11770,N_10312);
and U15480 (N_15480,N_11446,N_11485);
and U15481 (N_15481,N_13840,N_11415);
or U15482 (N_15482,N_12197,N_12400);
or U15483 (N_15483,N_10422,N_11257);
or U15484 (N_15484,N_13323,N_10287);
and U15485 (N_15485,N_10086,N_14839);
or U15486 (N_15486,N_12777,N_13564);
nor U15487 (N_15487,N_11498,N_10590);
nor U15488 (N_15488,N_12463,N_11476);
or U15489 (N_15489,N_10642,N_12503);
and U15490 (N_15490,N_10505,N_10064);
nor U15491 (N_15491,N_10127,N_14566);
nand U15492 (N_15492,N_13560,N_14409);
xnor U15493 (N_15493,N_10289,N_11906);
nand U15494 (N_15494,N_14395,N_12106);
and U15495 (N_15495,N_10334,N_12004);
and U15496 (N_15496,N_11222,N_11317);
nor U15497 (N_15497,N_11634,N_11394);
nand U15498 (N_15498,N_11902,N_10021);
nand U15499 (N_15499,N_11013,N_14236);
or U15500 (N_15500,N_13448,N_11401);
or U15501 (N_15501,N_11330,N_10654);
and U15502 (N_15502,N_12681,N_11922);
nor U15503 (N_15503,N_11760,N_12619);
and U15504 (N_15504,N_10075,N_10927);
nand U15505 (N_15505,N_10253,N_10449);
nand U15506 (N_15506,N_14768,N_13449);
and U15507 (N_15507,N_14279,N_11643);
or U15508 (N_15508,N_12605,N_12305);
nor U15509 (N_15509,N_14741,N_13746);
nor U15510 (N_15510,N_14540,N_10999);
nand U15511 (N_15511,N_11479,N_13984);
and U15512 (N_15512,N_11551,N_13264);
or U15513 (N_15513,N_13955,N_12955);
and U15514 (N_15514,N_12961,N_10813);
nor U15515 (N_15515,N_10926,N_11482);
or U15516 (N_15516,N_11382,N_10382);
nand U15517 (N_15517,N_13543,N_14098);
nor U15518 (N_15518,N_14481,N_14756);
and U15519 (N_15519,N_14578,N_12439);
and U15520 (N_15520,N_12225,N_12788);
nand U15521 (N_15521,N_11439,N_13575);
nor U15522 (N_15522,N_14356,N_12911);
and U15523 (N_15523,N_13146,N_13887);
xor U15524 (N_15524,N_10445,N_12692);
and U15525 (N_15525,N_11798,N_11934);
nor U15526 (N_15526,N_11600,N_12145);
and U15527 (N_15527,N_10216,N_14757);
xnor U15528 (N_15528,N_11524,N_11984);
and U15529 (N_15529,N_10498,N_10135);
or U15530 (N_15530,N_10541,N_10798);
nor U15531 (N_15531,N_13873,N_12244);
nor U15532 (N_15532,N_12252,N_10483);
nand U15533 (N_15533,N_11834,N_12114);
xor U15534 (N_15534,N_12423,N_14053);
nor U15535 (N_15535,N_11549,N_12233);
xnor U15536 (N_15536,N_10585,N_14192);
nand U15537 (N_15537,N_12365,N_11375);
or U15538 (N_15538,N_12192,N_10663);
nor U15539 (N_15539,N_12016,N_11754);
or U15540 (N_15540,N_11775,N_11436);
xor U15541 (N_15541,N_10629,N_14506);
and U15542 (N_15542,N_12933,N_11361);
xnor U15543 (N_15543,N_14226,N_12027);
xnor U15544 (N_15544,N_13653,N_12526);
and U15545 (N_15545,N_14631,N_11719);
nand U15546 (N_15546,N_13939,N_13190);
nor U15547 (N_15547,N_13153,N_14047);
nor U15548 (N_15548,N_10225,N_10205);
nor U15549 (N_15549,N_10119,N_10255);
or U15550 (N_15550,N_12975,N_11982);
nor U15551 (N_15551,N_13646,N_13063);
nand U15552 (N_15552,N_10238,N_10281);
nand U15553 (N_15553,N_14930,N_12022);
or U15554 (N_15554,N_14944,N_14015);
nor U15555 (N_15555,N_12066,N_13457);
nor U15556 (N_15556,N_10994,N_11012);
or U15557 (N_15557,N_12686,N_14702);
nor U15558 (N_15558,N_13308,N_13491);
and U15559 (N_15559,N_14940,N_11835);
and U15560 (N_15560,N_14915,N_11215);
or U15561 (N_15561,N_10171,N_12237);
nor U15562 (N_15562,N_12721,N_11388);
xnor U15563 (N_15563,N_13731,N_11201);
xor U15564 (N_15564,N_13208,N_14463);
or U15565 (N_15565,N_10789,N_14423);
nand U15566 (N_15566,N_12733,N_10669);
and U15567 (N_15567,N_14064,N_12974);
nor U15568 (N_15568,N_13706,N_11414);
nand U15569 (N_15569,N_12424,N_10342);
nand U15570 (N_15570,N_12568,N_13378);
nand U15571 (N_15571,N_13858,N_12971);
nand U15572 (N_15572,N_14938,N_14939);
or U15573 (N_15573,N_13062,N_10903);
and U15574 (N_15574,N_14195,N_14364);
nand U15575 (N_15575,N_14799,N_13822);
nand U15576 (N_15576,N_11758,N_13067);
nand U15577 (N_15577,N_13937,N_13719);
or U15578 (N_15578,N_13166,N_12394);
or U15579 (N_15579,N_10019,N_13807);
or U15580 (N_15580,N_13433,N_14767);
and U15581 (N_15581,N_11052,N_13313);
nor U15582 (N_15582,N_12734,N_10690);
nand U15583 (N_15583,N_13245,N_13940);
xnor U15584 (N_15584,N_14042,N_14828);
xor U15585 (N_15585,N_11676,N_14158);
nor U15586 (N_15586,N_12856,N_10656);
nand U15587 (N_15587,N_12711,N_12290);
or U15588 (N_15588,N_10552,N_14458);
nor U15589 (N_15589,N_12383,N_10066);
or U15590 (N_15590,N_14314,N_14770);
or U15591 (N_15591,N_14128,N_13750);
nand U15592 (N_15592,N_10011,N_12749);
xnor U15593 (N_15593,N_13985,N_12140);
and U15594 (N_15594,N_13015,N_14402);
xnor U15595 (N_15595,N_10500,N_13790);
nand U15596 (N_15596,N_13948,N_12381);
nor U15597 (N_15597,N_10333,N_13837);
and U15598 (N_15598,N_10425,N_10810);
nor U15599 (N_15599,N_12045,N_13319);
and U15600 (N_15600,N_10777,N_14036);
and U15601 (N_15601,N_11080,N_13307);
nor U15602 (N_15602,N_13437,N_11092);
nand U15603 (N_15603,N_11874,N_11994);
xor U15604 (N_15604,N_10877,N_12623);
and U15605 (N_15605,N_11046,N_14856);
nand U15606 (N_15606,N_12966,N_13155);
nor U15607 (N_15607,N_12442,N_13753);
or U15608 (N_15608,N_13565,N_14872);
and U15609 (N_15609,N_11371,N_14212);
or U15610 (N_15610,N_13226,N_14283);
nand U15611 (N_15611,N_12757,N_13156);
nor U15612 (N_15612,N_13133,N_13211);
and U15613 (N_15613,N_10408,N_14925);
nand U15614 (N_15614,N_10542,N_14316);
nand U15615 (N_15615,N_12984,N_13874);
nor U15616 (N_15616,N_11010,N_10896);
nor U15617 (N_15617,N_14103,N_11442);
nand U15618 (N_15618,N_12626,N_10948);
or U15619 (N_15619,N_13631,N_11147);
or U15620 (N_15620,N_13794,N_13115);
and U15621 (N_15621,N_11277,N_11859);
or U15622 (N_15622,N_10593,N_14061);
nor U15623 (N_15623,N_11730,N_11208);
or U15624 (N_15624,N_12729,N_14227);
nor U15625 (N_15625,N_10967,N_10966);
nor U15626 (N_15626,N_14665,N_13928);
and U15627 (N_15627,N_13047,N_10215);
xnor U15628 (N_15628,N_13509,N_11533);
nor U15629 (N_15629,N_12994,N_10373);
and U15630 (N_15630,N_11826,N_11106);
and U15631 (N_15631,N_13207,N_12878);
nand U15632 (N_15632,N_13845,N_10814);
and U15633 (N_15633,N_13949,N_11304);
and U15634 (N_15634,N_14060,N_11785);
and U15635 (N_15635,N_14963,N_10438);
nand U15636 (N_15636,N_10704,N_10836);
or U15637 (N_15637,N_11288,N_10917);
nand U15638 (N_15638,N_10580,N_11196);
or U15639 (N_15639,N_10675,N_12050);
nand U15640 (N_15640,N_11711,N_14842);
nor U15641 (N_15641,N_13369,N_10962);
xnor U15642 (N_15642,N_14558,N_11512);
nand U15643 (N_15643,N_11753,N_13513);
or U15644 (N_15644,N_12962,N_13064);
nor U15645 (N_15645,N_14180,N_12610);
nand U15646 (N_15646,N_14557,N_14201);
nor U15647 (N_15647,N_14691,N_13150);
nor U15648 (N_15648,N_13720,N_12675);
or U15649 (N_15649,N_13387,N_14802);
nand U15650 (N_15650,N_13990,N_14382);
xor U15651 (N_15651,N_10482,N_14438);
nor U15652 (N_15652,N_14067,N_11885);
nand U15653 (N_15653,N_14688,N_12771);
nor U15654 (N_15654,N_11646,N_10646);
nand U15655 (N_15655,N_10687,N_10853);
or U15656 (N_15656,N_11823,N_11098);
nand U15657 (N_15657,N_10269,N_13272);
and U15658 (N_15658,N_11564,N_14387);
or U15659 (N_15659,N_14564,N_13973);
or U15660 (N_15660,N_14795,N_13465);
and U15661 (N_15661,N_14050,N_12130);
and U15662 (N_15662,N_14012,N_10701);
nand U15663 (N_15663,N_12648,N_14934);
nor U15664 (N_15664,N_12378,N_11068);
or U15665 (N_15665,N_14474,N_12954);
nand U15666 (N_15666,N_11323,N_10565);
nand U15667 (N_15667,N_10574,N_12448);
nor U15668 (N_15668,N_14883,N_12801);
nand U15669 (N_15669,N_12180,N_14425);
xnor U15670 (N_15670,N_13704,N_12773);
nand U15671 (N_15671,N_14157,N_13735);
xnor U15672 (N_15672,N_14467,N_10720);
or U15673 (N_15673,N_10949,N_10594);
or U15674 (N_15674,N_13434,N_11879);
nand U15675 (N_15675,N_10511,N_12511);
or U15676 (N_15676,N_13757,N_11528);
xor U15677 (N_15677,N_12176,N_10486);
and U15678 (N_15678,N_11189,N_11918);
and U15679 (N_15679,N_14897,N_11326);
nor U15680 (N_15680,N_13879,N_12667);
xor U15681 (N_15681,N_11298,N_12895);
nand U15682 (N_15682,N_11958,N_11542);
and U15683 (N_15683,N_13918,N_13916);
and U15684 (N_15684,N_10435,N_13276);
and U15685 (N_15685,N_12491,N_13212);
or U15686 (N_15686,N_11675,N_12358);
xnor U15687 (N_15687,N_14244,N_14810);
xor U15688 (N_15688,N_14055,N_14200);
and U15689 (N_15689,N_13867,N_12277);
or U15690 (N_15690,N_12638,N_11558);
nor U15691 (N_15691,N_14788,N_12123);
nor U15692 (N_15692,N_14531,N_10559);
nand U15693 (N_15693,N_14653,N_13860);
and U15694 (N_15694,N_12924,N_11968);
nand U15695 (N_15695,N_13538,N_13679);
nand U15696 (N_15696,N_14165,N_13775);
and U15697 (N_15697,N_10442,N_12949);
nor U15698 (N_15698,N_13003,N_13677);
nand U15699 (N_15699,N_11976,N_13315);
nand U15700 (N_15700,N_14037,N_13127);
and U15701 (N_15701,N_13784,N_13559);
nand U15702 (N_15702,N_12704,N_10267);
nand U15703 (N_15703,N_14787,N_10761);
xor U15704 (N_15704,N_13611,N_14508);
xnor U15705 (N_15705,N_12627,N_13863);
and U15706 (N_15706,N_14304,N_10492);
nand U15707 (N_15707,N_14141,N_12501);
nor U15708 (N_15708,N_14248,N_12945);
or U15709 (N_15709,N_14461,N_13911);
and U15710 (N_15710,N_11732,N_11405);
or U15711 (N_15711,N_10157,N_14888);
nand U15712 (N_15712,N_11570,N_12700);
or U15713 (N_15713,N_12340,N_14286);
xnor U15714 (N_15714,N_10980,N_13200);
nand U15715 (N_15715,N_12190,N_14512);
or U15716 (N_15716,N_11367,N_11171);
nand U15717 (N_15717,N_13920,N_11416);
nand U15718 (N_15718,N_14867,N_11071);
nand U15719 (N_15719,N_11109,N_11582);
and U15720 (N_15720,N_13287,N_10200);
nor U15721 (N_15721,N_12401,N_11877);
and U15722 (N_15722,N_10503,N_12049);
and U15723 (N_15723,N_14333,N_10602);
and U15724 (N_15724,N_11440,N_12472);
or U15725 (N_15725,N_14862,N_14385);
nand U15726 (N_15726,N_12505,N_13553);
and U15727 (N_15727,N_12693,N_10800);
and U15728 (N_15728,N_11720,N_14625);
nand U15729 (N_15729,N_14273,N_14095);
nand U15730 (N_15730,N_14660,N_14874);
nor U15731 (N_15731,N_10527,N_10130);
xnor U15732 (N_15732,N_13561,N_14573);
and U15733 (N_15733,N_12374,N_14045);
nand U15734 (N_15734,N_14659,N_13896);
and U15735 (N_15735,N_13684,N_13689);
or U15736 (N_15736,N_10988,N_11650);
nand U15737 (N_15737,N_14703,N_14808);
nor U15738 (N_15738,N_12270,N_14958);
nor U15739 (N_15739,N_14923,N_14381);
or U15740 (N_15740,N_10728,N_11457);
or U15741 (N_15741,N_13912,N_14622);
or U15742 (N_15742,N_11795,N_10579);
nor U15743 (N_15743,N_10155,N_10218);
nor U15744 (N_15744,N_14251,N_14572);
or U15745 (N_15745,N_14232,N_11568);
and U15746 (N_15746,N_12433,N_12563);
nor U15747 (N_15747,N_12228,N_14639);
nor U15748 (N_15748,N_13957,N_14276);
nor U15749 (N_15749,N_10756,N_13152);
nor U15750 (N_15750,N_14974,N_13890);
and U15751 (N_15751,N_11573,N_14341);
nor U15752 (N_15752,N_11051,N_13600);
or U15753 (N_15753,N_11871,N_14234);
nand U15754 (N_15754,N_14956,N_13188);
nor U15755 (N_15755,N_11682,N_14309);
and U15756 (N_15756,N_12792,N_13033);
nor U15757 (N_15757,N_12102,N_10169);
or U15758 (N_15758,N_10341,N_12684);
or U15759 (N_15759,N_10153,N_14765);
nor U15760 (N_15760,N_13416,N_11124);
nor U15761 (N_15761,N_11380,N_11618);
and U15762 (N_15762,N_10797,N_10653);
and U15763 (N_15763,N_11470,N_10857);
or U15764 (N_15764,N_10271,N_12072);
nor U15765 (N_15765,N_12269,N_10290);
and U15766 (N_15766,N_10951,N_13621);
nor U15767 (N_15767,N_13341,N_11016);
nor U15768 (N_15768,N_10113,N_10981);
nor U15769 (N_15769,N_11332,N_14758);
nand U15770 (N_15770,N_11070,N_13154);
and U15771 (N_15771,N_14651,N_10915);
nor U15772 (N_15772,N_10478,N_13072);
or U15773 (N_15773,N_11525,N_14991);
and U15774 (N_15774,N_12624,N_14021);
nand U15775 (N_15775,N_12431,N_13938);
and U15776 (N_15776,N_10437,N_11005);
nand U15777 (N_15777,N_10941,N_13643);
nand U15778 (N_15778,N_14697,N_13399);
and U15779 (N_15779,N_11239,N_11028);
nor U15780 (N_15780,N_11407,N_14971);
nand U15781 (N_15781,N_10513,N_14282);
nand U15782 (N_15782,N_12343,N_14358);
or U15783 (N_15783,N_11129,N_12938);
and U15784 (N_15784,N_13992,N_12242);
and U15785 (N_15785,N_14454,N_12752);
nor U15786 (N_15786,N_10710,N_14255);
nor U15787 (N_15787,N_14590,N_11609);
and U15788 (N_15788,N_13987,N_10950);
or U15789 (N_15789,N_13511,N_14511);
or U15790 (N_15790,N_11082,N_12393);
nand U15791 (N_15791,N_10230,N_12980);
or U15792 (N_15792,N_11246,N_14337);
nor U15793 (N_15793,N_13979,N_13843);
or U15794 (N_15794,N_13371,N_12011);
and U15795 (N_15795,N_10454,N_14677);
xor U15796 (N_15796,N_13698,N_13346);
or U15797 (N_15797,N_12934,N_11045);
nand U15798 (N_15798,N_11450,N_10961);
and U15799 (N_15799,N_10010,N_13348);
nand U15800 (N_15800,N_13834,N_11860);
and U15801 (N_15801,N_14114,N_12208);
or U15802 (N_15802,N_14945,N_14614);
nand U15803 (N_15803,N_10904,N_10423);
or U15804 (N_15804,N_13329,N_13068);
and U15805 (N_15805,N_11033,N_11268);
or U15806 (N_15806,N_11428,N_13861);
xnor U15807 (N_15807,N_13135,N_13754);
nor U15808 (N_15808,N_10331,N_11337);
and U15809 (N_15809,N_11376,N_11079);
nor U15810 (N_15810,N_13946,N_14868);
nor U15811 (N_15811,N_12058,N_10004);
nand U15812 (N_15812,N_14737,N_14466);
and U15813 (N_15813,N_12581,N_10160);
xor U15814 (N_15814,N_13965,N_14321);
nand U15815 (N_15815,N_11644,N_10817);
nor U15816 (N_15816,N_12128,N_14943);
nand U15817 (N_15817,N_12406,N_13079);
nand U15818 (N_15818,N_12206,N_13557);
or U15819 (N_15819,N_11660,N_10301);
or U15820 (N_15820,N_14023,N_14931);
and U15821 (N_15821,N_11393,N_10888);
xnor U15822 (N_15822,N_11379,N_14699);
or U15823 (N_15823,N_13505,N_11677);
nor U15824 (N_15824,N_14869,N_11701);
and U15825 (N_15825,N_11513,N_14549);
or U15826 (N_15826,N_13439,N_13360);
nand U15827 (N_15827,N_12724,N_11977);
nor U15828 (N_15828,N_10826,N_12261);
nor U15829 (N_15829,N_14049,N_10212);
nor U15830 (N_15830,N_11929,N_10530);
nor U15831 (N_15831,N_10473,N_12769);
and U15832 (N_15832,N_11041,N_14773);
nor U15833 (N_15833,N_13562,N_11017);
nor U15834 (N_15834,N_10348,N_10459);
or U15835 (N_15835,N_11493,N_13978);
nor U15836 (N_15836,N_14739,N_13695);
nor U15837 (N_15837,N_11951,N_10517);
nand U15838 (N_15838,N_10968,N_12564);
nand U15839 (N_15839,N_14338,N_13081);
nor U15840 (N_15840,N_12632,N_12250);
or U15841 (N_15841,N_11716,N_13710);
or U15842 (N_15842,N_13088,N_13801);
nand U15843 (N_15843,N_14243,N_13692);
xor U15844 (N_15844,N_11793,N_12868);
nand U15845 (N_15845,N_14759,N_11433);
nor U15846 (N_15846,N_10706,N_13358);
xnor U15847 (N_15847,N_13809,N_13759);
or U15848 (N_15848,N_11050,N_12404);
and U15849 (N_15849,N_12601,N_11392);
and U15850 (N_15850,N_12008,N_10786);
or U15851 (N_15851,N_10576,N_13194);
and U15852 (N_15852,N_10520,N_14144);
or U15853 (N_15853,N_13877,N_10227);
nand U15854 (N_15854,N_13527,N_13274);
nor U15855 (N_15855,N_14524,N_13103);
and U15856 (N_15856,N_12513,N_13488);
or U15857 (N_15857,N_11227,N_14430);
xor U15858 (N_15858,N_10485,N_10975);
or U15859 (N_15859,N_10095,N_11259);
xor U15860 (N_15860,N_13256,N_12778);
or U15861 (N_15861,N_13097,N_14547);
nand U15862 (N_15862,N_13914,N_11633);
and U15863 (N_15863,N_11515,N_10370);
nand U15864 (N_15864,N_10911,N_14636);
or U15865 (N_15865,N_14721,N_14949);
or U15866 (N_15866,N_11339,N_10288);
and U15867 (N_15867,N_10087,N_12695);
nand U15868 (N_15868,N_11967,N_11856);
nor U15869 (N_15869,N_10614,N_13403);
and U15870 (N_15870,N_13722,N_11764);
nor U15871 (N_15871,N_12395,N_14796);
xnor U15872 (N_15872,N_13798,N_13415);
and U15873 (N_15873,N_13828,N_13545);
and U15874 (N_15874,N_12231,N_13636);
and U15875 (N_15875,N_10295,N_13405);
nor U15876 (N_15876,N_14247,N_13397);
nor U15877 (N_15877,N_11505,N_11628);
xnor U15878 (N_15878,N_13578,N_12043);
and U15879 (N_15879,N_14746,N_14077);
or U15880 (N_15880,N_10698,N_12085);
or U15881 (N_15881,N_13717,N_12392);
or U15882 (N_15882,N_13654,N_11348);
nand U15883 (N_15883,N_10024,N_14390);
nand U15884 (N_15884,N_12791,N_12430);
xnor U15885 (N_15885,N_10243,N_12636);
or U15886 (N_15886,N_14964,N_13401);
nor U15887 (N_15887,N_12859,N_13913);
nor U15888 (N_15888,N_12510,N_11830);
xnor U15889 (N_15889,N_10586,N_12910);
or U15890 (N_15890,N_14560,N_14121);
nand U15891 (N_15891,N_10069,N_11642);
and U15892 (N_15892,N_14035,N_13458);
nor U15893 (N_15893,N_14735,N_14400);
and U15894 (N_15894,N_13007,N_13922);
and U15895 (N_15895,N_13412,N_12273);
nand U15896 (N_15896,N_14424,N_12549);
nand U15897 (N_15897,N_14058,N_11909);
xor U15898 (N_15898,N_14608,N_12188);
nor U15899 (N_15899,N_12944,N_12209);
nor U15900 (N_15900,N_13193,N_12164);
nor U15901 (N_15901,N_12765,N_10448);
or U15902 (N_15902,N_12346,N_13228);
and U15903 (N_15903,N_10188,N_13131);
and U15904 (N_15904,N_13898,N_13435);
or U15905 (N_15905,N_10897,N_10673);
nand U15906 (N_15906,N_10688,N_13295);
nor U15907 (N_15907,N_11094,N_13396);
or U15908 (N_15908,N_12783,N_13355);
nand U15909 (N_15909,N_11058,N_10712);
nor U15910 (N_15910,N_14118,N_10956);
or U15911 (N_15911,N_10925,N_11608);
or U15912 (N_15912,N_14307,N_14575);
or U15913 (N_15913,N_11250,N_12260);
xor U15914 (N_15914,N_12079,N_13580);
or U15915 (N_15915,N_11990,N_13340);
or U15916 (N_15916,N_11456,N_13541);
and U15917 (N_15917,N_10044,N_10025);
and U15918 (N_15918,N_10402,N_13459);
and U15919 (N_15919,N_14948,N_10375);
nand U15920 (N_15920,N_11491,N_10315);
nand U15921 (N_15921,N_14740,N_10942);
xnor U15922 (N_15922,N_13566,N_10946);
xnor U15923 (N_15923,N_13098,N_14186);
nand U15924 (N_15924,N_10151,N_11844);
nor U15925 (N_15925,N_11991,N_10043);
nand U15926 (N_15926,N_11435,N_11819);
and U15927 (N_15927,N_12007,N_10573);
nor U15928 (N_15928,N_13238,N_13306);
nor U15929 (N_15929,N_12864,N_12705);
and U15930 (N_15930,N_13391,N_11841);
and U15931 (N_15931,N_10343,N_11546);
nand U15932 (N_15932,N_13763,N_12364);
nand U15933 (N_15933,N_12642,N_10092);
and U15934 (N_15934,N_10568,N_14567);
nor U15935 (N_15935,N_14840,N_13886);
or U15936 (N_15936,N_13114,N_10037);
nand U15937 (N_15937,N_14728,N_13961);
nand U15938 (N_15938,N_10751,N_13370);
or U15939 (N_15939,N_14846,N_14714);
or U15940 (N_15940,N_14362,N_10515);
nand U15941 (N_15941,N_14091,N_11948);
and U15942 (N_15942,N_10246,N_11153);
or U15943 (N_15943,N_10684,N_10578);
and U15944 (N_15944,N_11734,N_12506);
nand U15945 (N_15945,N_10566,N_10937);
or U15946 (N_15946,N_11175,N_14616);
and U15947 (N_15947,N_13056,N_14911);
or U15948 (N_15948,N_11241,N_14611);
or U15949 (N_15949,N_14877,N_11395);
and U15950 (N_15950,N_13424,N_12751);
nand U15951 (N_15951,N_10812,N_13838);
xnor U15952 (N_15952,N_11538,N_14530);
nor U15953 (N_15953,N_14571,N_11278);
and U15954 (N_15954,N_10768,N_12265);
nand U15955 (N_15955,N_14252,N_12061);
nor U15956 (N_15956,N_10257,N_10424);
nor U15957 (N_15957,N_14312,N_13927);
or U15958 (N_15958,N_14729,N_13471);
or U15959 (N_15959,N_14837,N_13995);
or U15960 (N_15960,N_12174,N_10349);
or U15961 (N_15961,N_12851,N_11580);
xor U15962 (N_15962,N_10686,N_14073);
and U15963 (N_15963,N_10453,N_13092);
nor U15964 (N_15964,N_13362,N_14446);
nand U15965 (N_15965,N_14010,N_11199);
or U15966 (N_15966,N_11336,N_13005);
or U15967 (N_15967,N_13785,N_10219);
or U15968 (N_15968,N_13586,N_12115);
or U15969 (N_15969,N_14379,N_12230);
or U15970 (N_15970,N_11403,N_11377);
or U15971 (N_15971,N_14821,N_10213);
nand U15972 (N_15972,N_13880,N_13942);
nor U15973 (N_15973,N_11181,N_13674);
nand U15974 (N_15974,N_11853,N_12649);
or U15975 (N_15975,N_10873,N_12199);
nor U15976 (N_15976,N_12840,N_10097);
and U15977 (N_15977,N_12952,N_13021);
or U15978 (N_15978,N_14638,N_14607);
and U15979 (N_15979,N_10452,N_14679);
nor U15980 (N_15980,N_10003,N_14440);
nor U15981 (N_15981,N_13749,N_10177);
or U15982 (N_15982,N_12639,N_11713);
xnor U15983 (N_15983,N_13787,N_10150);
nor U15984 (N_15984,N_11510,N_10063);
and U15985 (N_15985,N_14429,N_10982);
and U15986 (N_15986,N_10569,N_13683);
and U15987 (N_15987,N_13085,N_12227);
or U15988 (N_15988,N_12268,N_12575);
nand U15989 (N_15989,N_12363,N_10138);
nor U15990 (N_15990,N_10495,N_12152);
or U15991 (N_15991,N_14453,N_13968);
nand U15992 (N_15992,N_14908,N_14441);
and U15993 (N_15993,N_10361,N_12009);
nor U15994 (N_15994,N_13823,N_12308);
and U15995 (N_15995,N_13383,N_13271);
or U15996 (N_15996,N_10697,N_10384);
nor U15997 (N_15997,N_13337,N_12718);
or U15998 (N_15998,N_12618,N_11869);
or U15999 (N_15999,N_13554,N_12362);
nand U16000 (N_16000,N_13262,N_11805);
nand U16001 (N_16001,N_10816,N_10270);
nand U16002 (N_16002,N_12284,N_14663);
and U16003 (N_16003,N_11678,N_12953);
and U16004 (N_16004,N_13010,N_10577);
nand U16005 (N_16005,N_11995,N_10321);
nor U16006 (N_16006,N_11786,N_12735);
nand U16007 (N_16007,N_12183,N_12816);
and U16008 (N_16008,N_11889,N_12978);
or U16009 (N_16009,N_11334,N_14203);
xor U16010 (N_16010,N_11745,N_11354);
nand U16011 (N_16011,N_14912,N_12464);
nor U16012 (N_16012,N_10689,N_13084);
and U16013 (N_16013,N_13001,N_14452);
nand U16014 (N_16014,N_13384,N_11009);
or U16015 (N_16015,N_10048,N_13854);
or U16016 (N_16016,N_13137,N_14065);
and U16017 (N_16017,N_14183,N_14983);
nand U16018 (N_16018,N_12471,N_13451);
nor U16019 (N_16019,N_13298,N_11789);
and U16020 (N_16020,N_12659,N_13158);
and U16021 (N_16021,N_14241,N_12818);
or U16022 (N_16022,N_13027,N_10428);
and U16023 (N_16023,N_11773,N_12656);
nor U16024 (N_16024,N_12017,N_13304);
nor U16025 (N_16025,N_12834,N_12772);
nand U16026 (N_16026,N_12780,N_14416);
nor U16027 (N_16027,N_13862,N_11517);
xnor U16028 (N_16028,N_13066,N_14749);
or U16029 (N_16029,N_13851,N_12658);
or U16030 (N_16030,N_14890,N_11797);
nor U16031 (N_16031,N_13533,N_13711);
xnor U16032 (N_16032,N_10754,N_11345);
and U16033 (N_16033,N_12373,N_11866);
or U16034 (N_16034,N_10649,N_10279);
or U16035 (N_16035,N_12019,N_13988);
or U16036 (N_16036,N_12148,N_14843);
nor U16037 (N_16037,N_11384,N_12033);
or U16038 (N_16038,N_14086,N_11490);
and U16039 (N_16039,N_13512,N_10599);
or U16040 (N_16040,N_11155,N_11941);
and U16041 (N_16041,N_11926,N_10865);
nor U16042 (N_16042,N_14527,N_10729);
nor U16043 (N_16043,N_13870,N_11223);
or U16044 (N_16044,N_12873,N_11669);
and U16045 (N_16045,N_12603,N_12820);
or U16046 (N_16046,N_14551,N_11029);
or U16047 (N_16047,N_10626,N_14875);
or U16048 (N_16048,N_12282,N_10317);
and U16049 (N_16049,N_14535,N_10047);
and U16050 (N_16050,N_11638,N_13582);
and U16051 (N_16051,N_11260,N_10067);
nor U16052 (N_16052,N_14613,N_13100);
nand U16053 (N_16053,N_14005,N_11535);
nand U16054 (N_16054,N_14039,N_13647);
nand U16055 (N_16055,N_12368,N_11481);
or U16056 (N_16056,N_13095,N_11314);
or U16057 (N_16057,N_13237,N_10799);
or U16058 (N_16058,N_12995,N_13128);
nand U16059 (N_16059,N_14712,N_14125);
nor U16060 (N_16060,N_12861,N_13919);
nand U16061 (N_16061,N_13182,N_13279);
xnor U16062 (N_16062,N_12803,N_11313);
nand U16063 (N_16063,N_14378,N_11997);
or U16064 (N_16064,N_14465,N_14330);
nor U16065 (N_16065,N_14797,N_14725);
or U16066 (N_16066,N_13305,N_11177);
nor U16067 (N_16067,N_14394,N_14680);
or U16068 (N_16068,N_14921,N_10197);
or U16069 (N_16069,N_14584,N_13817);
and U16070 (N_16070,N_13106,N_14123);
nor U16071 (N_16071,N_12210,N_14917);
and U16072 (N_16072,N_12104,N_12348);
nand U16073 (N_16073,N_13758,N_12828);
nand U16074 (N_16074,N_12220,N_12258);
and U16075 (N_16075,N_10512,N_13053);
nor U16076 (N_16076,N_14094,N_10525);
nand U16077 (N_16077,N_10376,N_14189);
nor U16078 (N_16078,N_10223,N_11254);
nor U16079 (N_16079,N_13676,N_13039);
or U16080 (N_16080,N_14968,N_10736);
or U16081 (N_16081,N_13607,N_11612);
nand U16082 (N_16082,N_13576,N_11622);
or U16083 (N_16083,N_13591,N_12597);
nand U16084 (N_16084,N_13991,N_10265);
nand U16085 (N_16085,N_10781,N_14772);
xnor U16086 (N_16086,N_14386,N_13257);
nor U16087 (N_16087,N_12311,N_13096);
nor U16088 (N_16088,N_12411,N_12170);
and U16089 (N_16089,N_12421,N_14687);
and U16090 (N_16090,N_14825,N_14300);
nand U16091 (N_16091,N_11242,N_12677);
xnor U16092 (N_16092,N_12533,N_10194);
or U16093 (N_16093,N_12434,N_11075);
nor U16094 (N_16094,N_10367,N_11592);
nor U16095 (N_16095,N_10560,N_11833);
nand U16096 (N_16096,N_14852,N_12986);
nor U16097 (N_16097,N_11855,N_13241);
nand U16098 (N_16098,N_12345,N_10360);
or U16099 (N_16099,N_10471,N_13004);
and U16100 (N_16100,N_13101,N_13882);
nand U16101 (N_16101,N_12015,N_14107);
nor U16102 (N_16102,N_10202,N_14270);
xor U16103 (N_16103,N_13593,N_12827);
or U16104 (N_16104,N_14439,N_10394);
and U16105 (N_16105,N_11820,N_12297);
or U16106 (N_16106,N_11983,N_11207);
nor U16107 (N_16107,N_14327,N_14656);
and U16108 (N_16108,N_11036,N_14262);
nor U16109 (N_16109,N_12872,N_11192);
xor U16110 (N_16110,N_14849,N_13388);
or U16111 (N_16111,N_13480,N_10601);
xnor U16112 (N_16112,N_11743,N_10105);
nand U16113 (N_16113,N_10802,N_11708);
nor U16114 (N_16114,N_12302,N_11458);
nand U16115 (N_16115,N_11076,N_14838);
xnor U16116 (N_16116,N_12908,N_13855);
or U16117 (N_16117,N_11043,N_10082);
nor U16118 (N_16118,N_13539,N_13630);
nor U16119 (N_16119,N_11766,N_14864);
nand U16120 (N_16120,N_11021,N_10535);
or U16121 (N_16121,N_13476,N_12717);
nand U16122 (N_16122,N_11370,N_12350);
nand U16123 (N_16123,N_14933,N_11409);
nand U16124 (N_16124,N_13744,N_12779);
xor U16125 (N_16125,N_14965,N_13398);
nand U16126 (N_16126,N_12432,N_10724);
xnor U16127 (N_16127,N_13417,N_11566);
nand U16128 (N_16128,N_11813,N_13872);
and U16129 (N_16129,N_12894,N_13293);
nand U16130 (N_16130,N_12000,N_11611);
xor U16131 (N_16131,N_14513,N_12420);
and U16132 (N_16132,N_13544,N_13635);
and U16133 (N_16133,N_12560,N_13483);
nand U16134 (N_16134,N_14224,N_13025);
or U16135 (N_16135,N_10871,N_12196);
and U16136 (N_16136,N_11543,N_12545);
and U16137 (N_16137,N_10863,N_10185);
nor U16138 (N_16138,N_10353,N_10278);
nand U16139 (N_16139,N_14747,N_10849);
nor U16140 (N_16140,N_12352,N_14827);
nor U16141 (N_16141,N_14977,N_13209);
and U16142 (N_16142,N_11266,N_11648);
nand U16143 (N_16143,N_10261,N_14896);
nand U16144 (N_16144,N_14294,N_11108);
nor U16145 (N_16145,N_12582,N_11229);
nand U16146 (N_16146,N_12384,N_10029);
nor U16147 (N_16147,N_13364,N_11639);
nor U16148 (N_16148,N_10906,N_12712);
nor U16149 (N_16149,N_10339,N_13178);
or U16150 (N_16150,N_11074,N_10027);
or U16151 (N_16151,N_14928,N_10537);
nand U16152 (N_16152,N_14994,N_12356);
xor U16153 (N_16153,N_10322,N_12723);
nor U16154 (N_16154,N_10232,N_14918);
or U16155 (N_16155,N_12798,N_10089);
nor U16156 (N_16156,N_14082,N_12942);
nor U16157 (N_16157,N_10383,N_10989);
nor U16158 (N_16158,N_12880,N_13756);
nor U16159 (N_16159,N_13043,N_12775);
and U16160 (N_16160,N_11696,N_14706);
nor U16161 (N_16161,N_14470,N_11672);
nand U16162 (N_16162,N_10539,N_14469);
nor U16163 (N_16163,N_10685,N_14001);
or U16164 (N_16164,N_12612,N_13472);
nand U16165 (N_16165,N_10847,N_11679);
nor U16166 (N_16166,N_14122,N_12254);
nand U16167 (N_16167,N_12320,N_13820);
nand U16168 (N_16168,N_11496,N_12787);
nor U16169 (N_16169,N_10972,N_10203);
nand U16170 (N_16170,N_10053,N_13494);
and U16171 (N_16171,N_12403,N_12552);
xnor U16172 (N_16172,N_10244,N_12137);
or U16173 (N_16173,N_13707,N_12370);
nor U16174 (N_16174,N_13734,N_13998);
or U16175 (N_16175,N_10592,N_11756);
or U16176 (N_16176,N_13610,N_13587);
or U16177 (N_16177,N_14302,N_10935);
nor U16178 (N_16178,N_12499,N_14556);
nand U16179 (N_16179,N_11953,N_11419);
xnor U16180 (N_16180,N_14328,N_10801);
and U16181 (N_16181,N_14880,N_13057);
or U16182 (N_16182,N_10328,N_12014);
or U16183 (N_16183,N_10359,N_13666);
or U16184 (N_16184,N_14997,N_11107);
nor U16185 (N_16185,N_14132,N_10606);
xnor U16186 (N_16186,N_12515,N_12795);
nand U16187 (N_16187,N_10676,N_10549);
nor U16188 (N_16188,N_11903,N_12186);
or U16189 (N_16189,N_10458,N_11423);
or U16190 (N_16190,N_11449,N_11121);
and U16191 (N_16191,N_10758,N_11858);
xnor U16192 (N_16192,N_11563,N_13189);
nor U16193 (N_16193,N_10436,N_10655);
nor U16194 (N_16194,N_12312,N_13368);
nand U16195 (N_16195,N_14443,N_14408);
nand U16196 (N_16196,N_12080,N_10759);
or U16197 (N_16197,N_11540,N_12726);
nor U16198 (N_16198,N_12489,N_12144);
and U16199 (N_16199,N_13283,N_12271);
and U16200 (N_16200,N_11897,N_13685);
nor U16201 (N_16201,N_10000,N_13709);
and U16202 (N_16202,N_12806,N_10327);
and U16203 (N_16203,N_14503,N_10955);
nand U16204 (N_16204,N_13667,N_14000);
or U16205 (N_16205,N_12967,N_11938);
and U16206 (N_16206,N_14941,N_13907);
or U16207 (N_16207,N_13255,N_11426);
nand U16208 (N_16208,N_13395,N_11002);
nand U16209 (N_16209,N_14209,N_11272);
or U16210 (N_16210,N_11338,N_12651);
nor U16211 (N_16211,N_11472,N_13701);
and U16212 (N_16212,N_13889,N_12122);
or U16213 (N_16213,N_12306,N_12739);
nand U16214 (N_16214,N_13440,N_10142);
nand U16215 (N_16215,N_11025,N_11355);
or U16216 (N_16216,N_10771,N_11658);
or U16217 (N_16217,N_13468,N_14292);
xnor U16218 (N_16218,N_10823,N_10324);
and U16219 (N_16219,N_10631,N_11427);
nor U16220 (N_16220,N_12948,N_13357);
or U16221 (N_16221,N_12309,N_11868);
and U16222 (N_16222,N_14779,N_13496);
or U16223 (N_16223,N_14596,N_11681);
nor U16224 (N_16224,N_14285,N_12767);
nor U16225 (N_16225,N_10969,N_14887);
and U16226 (N_16226,N_11959,N_10041);
nor U16227 (N_16227,N_10093,N_10582);
nor U16228 (N_16228,N_14126,N_10298);
nand U16229 (N_16229,N_10466,N_14919);
nor U16230 (N_16230,N_14818,N_12135);
nand U16231 (N_16231,N_13467,N_12038);
or U16232 (N_16232,N_11185,N_13737);
nand U16233 (N_16233,N_11233,N_13900);
nor U16234 (N_16234,N_10403,N_13011);
nand U16235 (N_16235,N_12635,N_13558);
and U16236 (N_16236,N_10049,N_10101);
or U16237 (N_16237,N_10098,N_13947);
nor U16238 (N_16238,N_11733,N_12542);
nand U16239 (N_16239,N_14359,N_14340);
nand U16240 (N_16240,N_12647,N_13408);
or U16241 (N_16241,N_10146,N_13390);
or U16242 (N_16242,N_14924,N_11085);
and U16243 (N_16243,N_12480,N_11605);
and U16244 (N_16244,N_12947,N_10487);
or U16245 (N_16245,N_11811,N_13952);
nand U16246 (N_16246,N_11312,N_11173);
and U16247 (N_16247,N_12571,N_14635);
or U16248 (N_16248,N_11896,N_11962);
xor U16249 (N_16249,N_10938,N_11240);
nor U16250 (N_16250,N_12380,N_13906);
and U16251 (N_16251,N_12338,N_11891);
and U16252 (N_16252,N_12426,N_13141);
nand U16253 (N_16253,N_11137,N_14847);
and U16254 (N_16254,N_11279,N_12875);
and U16255 (N_16255,N_10112,N_11399);
nor U16256 (N_16256,N_14213,N_13960);
and U16257 (N_16257,N_13721,N_12276);
nor U16258 (N_16258,N_14332,N_12445);
nand U16259 (N_16259,N_14184,N_12915);
or U16260 (N_16260,N_13546,N_12676);
nand U16261 (N_16261,N_12825,N_13664);
and U16262 (N_16262,N_12981,N_14240);
nand U16263 (N_16263,N_12741,N_10009);
nand U16264 (N_16264,N_13687,N_13510);
nand U16265 (N_16265,N_11161,N_13206);
nor U16266 (N_16266,N_14881,N_10811);
nor U16267 (N_16267,N_10805,N_14214);
or U16268 (N_16268,N_10665,N_12329);
and U16269 (N_16269,N_14096,N_12232);
or U16270 (N_16270,N_14405,N_10742);
and U16271 (N_16271,N_10944,N_10523);
nand U16272 (N_16272,N_10263,N_13060);
nor U16273 (N_16273,N_10973,N_12579);
nor U16274 (N_16274,N_14457,N_10551);
and U16275 (N_16275,N_12814,N_13980);
or U16276 (N_16276,N_10300,N_11778);
and U16277 (N_16277,N_11999,N_10038);
nor U16278 (N_16278,N_10139,N_14008);
nor U16279 (N_16279,N_13159,N_11455);
nand U16280 (N_16280,N_10554,N_14301);
nor U16281 (N_16281,N_10891,N_14526);
nand U16282 (N_16282,N_11601,N_14803);
nor U16283 (N_16283,N_10262,N_11552);
nand U16284 (N_16284,N_13738,N_12753);
nor U16285 (N_16285,N_13055,N_13250);
nand U16286 (N_16286,N_12353,N_14486);
and U16287 (N_16287,N_10109,N_12903);
or U16288 (N_16288,N_12766,N_10351);
nand U16289 (N_16289,N_14471,N_11011);
nor U16290 (N_16290,N_13462,N_14599);
nand U16291 (N_16291,N_14084,N_12315);
nor U16292 (N_16292,N_12324,N_14383);
or U16293 (N_16293,N_11294,N_10959);
nor U16294 (N_16294,N_13726,N_13464);
nor U16295 (N_16295,N_14478,N_14753);
nor U16296 (N_16296,N_12770,N_10735);
nand U16297 (N_16297,N_13191,N_12473);
nor U16298 (N_16298,N_13215,N_14140);
and U16299 (N_16299,N_14242,N_12294);
and U16300 (N_16300,N_12595,N_12565);
or U16301 (N_16301,N_12682,N_13389);
and U16302 (N_16302,N_12490,N_10091);
or U16303 (N_16303,N_12097,N_10501);
nor U16304 (N_16304,N_12621,N_14120);
or U16305 (N_16305,N_14955,N_11790);
nand U16306 (N_16306,N_13993,N_10921);
nand U16307 (N_16307,N_13549,N_14419);
nor U16308 (N_16308,N_10400,N_10406);
nor U16309 (N_16309,N_12127,N_11362);
nand U16310 (N_16310,N_12548,N_11989);
nand U16311 (N_16311,N_13680,N_14962);
or U16312 (N_16312,N_10866,N_11316);
xnor U16313 (N_16313,N_10556,N_14907);
nor U16314 (N_16314,N_11321,N_13857);
xnor U16315 (N_16315,N_10722,N_13668);
or U16316 (N_16316,N_11308,N_13094);
nor U16317 (N_16317,N_10661,N_13139);
and U16318 (N_16318,N_10235,N_13500);
nand U16319 (N_16319,N_13148,N_14514);
nand U16320 (N_16320,N_13791,N_10971);
or U16321 (N_16321,N_12182,N_14637);
nor U16322 (N_16322,N_11398,N_13844);
nand U16323 (N_16323,N_13352,N_12558);
or U16324 (N_16324,N_10252,N_10910);
nand U16325 (N_16325,N_10305,N_10472);
or U16326 (N_16326,N_14592,N_11996);
nor U16327 (N_16327,N_14895,N_11218);
and U16328 (N_16328,N_14421,N_12785);
nand U16329 (N_16329,N_11151,N_10455);
and U16330 (N_16330,N_12762,N_11782);
and U16331 (N_16331,N_12912,N_13303);
or U16332 (N_16332,N_14343,N_11500);
and U16333 (N_16333,N_13832,N_14866);
nand U16334 (N_16334,N_12737,N_12322);
nor U16335 (N_16335,N_12698,N_12248);
nor U16336 (N_16336,N_12241,N_11228);
or U16337 (N_16337,N_11193,N_13945);
nor U16338 (N_16338,N_13800,N_13866);
nor U16339 (N_16339,N_10991,N_11026);
nor U16340 (N_16340,N_14360,N_10286);
nand U16341 (N_16341,N_10723,N_13233);
or U16342 (N_16342,N_14167,N_14484);
nand U16343 (N_16343,N_12039,N_13454);
or U16344 (N_16344,N_12706,N_11774);
nor U16345 (N_16345,N_13261,N_13431);
or U16346 (N_16346,N_14410,N_14070);
and U16347 (N_16347,N_11901,N_10099);
or U16348 (N_16348,N_11737,N_13589);
and U16349 (N_16349,N_10018,N_10782);
nor U16350 (N_16350,N_14581,N_14675);
xnor U16351 (N_16351,N_13507,N_13627);
nor U16352 (N_16352,N_10078,N_11006);
nor U16353 (N_16353,N_14310,N_10164);
nand U16354 (N_16354,N_10154,N_14510);
and U16355 (N_16355,N_11116,N_13484);
nand U16356 (N_16356,N_10827,N_11567);
nor U16357 (N_16357,N_14254,N_13713);
or U16358 (N_16358,N_12326,N_14730);
nand U16359 (N_16359,N_12319,N_13023);
and U16360 (N_16360,N_14102,N_13550);
or U16361 (N_16361,N_13944,N_14563);
nand U16362 (N_16362,N_14375,N_14253);
or U16363 (N_16363,N_14792,N_14973);
nand U16364 (N_16364,N_11746,N_13220);
or U16365 (N_16365,N_11299,N_13050);
or U16366 (N_16366,N_10993,N_14844);
and U16367 (N_16367,N_12728,N_14417);
and U16368 (N_16368,N_12841,N_10639);
or U16369 (N_16369,N_13036,N_10313);
nor U16370 (N_16370,N_13616,N_13086);
and U16371 (N_16371,N_13299,N_10358);
or U16372 (N_16372,N_12585,N_10133);
or U16373 (N_16373,N_10892,N_12288);
and U16374 (N_16374,N_11867,N_12042);
nand U16375 (N_16375,N_10103,N_11814);
xnor U16376 (N_16376,N_10899,N_14231);
nor U16377 (N_16377,N_13376,N_10059);
or U16378 (N_16378,N_14092,N_13602);
and U16379 (N_16379,N_13243,N_14468);
nor U16380 (N_16380,N_10526,N_14718);
or U16381 (N_16381,N_14634,N_14970);
or U16382 (N_16382,N_10479,N_14261);
nand U16383 (N_16383,N_10330,N_14334);
xor U16384 (N_16384,N_14522,N_12053);
and U16385 (N_16385,N_12035,N_11815);
and U16386 (N_16386,N_10772,N_11195);
xnor U16387 (N_16387,N_10054,N_11710);
nand U16388 (N_16388,N_11270,N_14295);
xnor U16389 (N_16389,N_14860,N_14670);
nor U16390 (N_16390,N_13827,N_11143);
and U16391 (N_16391,N_10719,N_11487);
nand U16392 (N_16392,N_12020,N_14515);
or U16393 (N_16393,N_11956,N_12517);
or U16394 (N_16394,N_14154,N_12249);
nor U16395 (N_16395,N_11261,N_11562);
nand U16396 (N_16396,N_10718,N_12916);
xnor U16397 (N_16397,N_12793,N_10608);
xor U16398 (N_16398,N_14961,N_14878);
nor U16399 (N_16399,N_11589,N_13116);
nor U16400 (N_16400,N_10226,N_14533);
and U16401 (N_16401,N_12382,N_12046);
nor U16402 (N_16402,N_13278,N_11603);
nand U16403 (N_16403,N_11204,N_13542);
or U16404 (N_16404,N_10137,N_14319);
and U16405 (N_16405,N_12898,N_14349);
nand U16406 (N_16406,N_11103,N_12617);
and U16407 (N_16407,N_11522,N_13009);
or U16408 (N_16408,N_11848,N_11300);
nor U16409 (N_16409,N_12960,N_14553);
and U16410 (N_16410,N_13185,N_12194);
nand U16411 (N_16411,N_13363,N_10660);
nor U16412 (N_16412,N_12417,N_14545);
nor U16413 (N_16413,N_10529,N_10302);
nand U16414 (N_16414,N_10562,N_14543);
nand U16415 (N_16415,N_11358,N_14376);
and U16416 (N_16416,N_10240,N_11290);
or U16417 (N_16417,N_13198,N_14689);
nand U16418 (N_16418,N_11462,N_14268);
nand U16419 (N_16419,N_13811,N_14626);
or U16420 (N_16420,N_12609,N_11674);
and U16421 (N_16421,N_11937,N_10431);
nor U16422 (N_16422,N_14984,N_11666);
and U16423 (N_16423,N_11319,N_14711);
or U16424 (N_16424,N_13716,N_12913);
or U16425 (N_16425,N_10774,N_12157);
nor U16426 (N_16426,N_12129,N_12502);
nor U16427 (N_16427,N_10296,N_14722);
nand U16428 (N_16428,N_14633,N_13997);
nand U16429 (N_16429,N_14097,N_14682);
nor U16430 (N_16430,N_14163,N_11346);
and U16431 (N_16431,N_14766,N_12187);
or U16432 (N_16432,N_12105,N_12103);
or U16433 (N_16433,N_12021,N_11119);
and U16434 (N_16434,N_12822,N_14258);
or U16435 (N_16435,N_13660,N_14257);
or U16436 (N_16436,N_11876,N_14900);
nand U16437 (N_16437,N_13923,N_13492);
or U16438 (N_16438,N_13520,N_11347);
nor U16439 (N_16439,N_11133,N_12023);
nand U16440 (N_16440,N_10340,N_12644);
nor U16441 (N_16441,N_13447,N_10440);
nand U16442 (N_16442,N_11783,N_10726);
nor U16443 (N_16443,N_10806,N_14627);
nor U16444 (N_16444,N_13892,N_14658);
nor U16445 (N_16445,N_14007,N_10567);
nand U16446 (N_16446,N_12654,N_12069);
xnor U16447 (N_16447,N_13482,N_12314);
nor U16448 (N_16448,N_13102,N_14863);
and U16449 (N_16449,N_14488,N_11374);
xor U16450 (N_16450,N_10460,N_11152);
nor U16451 (N_16451,N_14009,N_11863);
and U16452 (N_16452,N_12347,N_13069);
nor U16453 (N_16453,N_14017,N_11486);
nand U16454 (N_16454,N_12458,N_11727);
nor U16455 (N_16455,N_12133,N_10210);
nand U16456 (N_16456,N_10753,N_11685);
and U16457 (N_16457,N_10713,N_10434);
nand U16458 (N_16458,N_13373,N_13350);
and U16459 (N_16459,N_11688,N_11728);
or U16460 (N_16460,N_11400,N_10913);
nor U16461 (N_16461,N_10667,N_14559);
and U16462 (N_16462,N_10670,N_11369);
xor U16463 (N_16463,N_12087,N_12683);
nor U16464 (N_16464,N_10785,N_12059);
nand U16465 (N_16465,N_11504,N_11120);
nor U16466 (N_16466,N_12281,N_13375);
xnor U16467 (N_16467,N_10420,N_13254);
or U16468 (N_16468,N_14291,N_10591);
and U16469 (N_16469,N_10700,N_13201);
nor U16470 (N_16470,N_12973,N_12359);
nand U16471 (N_16471,N_11693,N_11126);
nor U16472 (N_16472,N_10411,N_13330);
xnor U16473 (N_16473,N_11944,N_10622);
nand U16474 (N_16474,N_10778,N_11893);
nor U16475 (N_16475,N_10229,N_14249);
or U16476 (N_16476,N_11501,N_12195);
nor U16477 (N_16477,N_14110,N_12756);
nand U16478 (N_16478,N_13762,N_10363);
xnor U16479 (N_16479,N_10198,N_12835);
and U16480 (N_16480,N_14870,N_13893);
xor U16481 (N_16481,N_10042,N_10767);
and U16482 (N_16482,N_13640,N_10752);
and U16483 (N_16483,N_13614,N_12529);
nor U16484 (N_16484,N_14325,N_11873);
xnor U16485 (N_16485,N_13087,N_11649);
nand U16486 (N_16486,N_10818,N_13406);
or U16487 (N_16487,N_14288,N_13742);
or U16488 (N_16488,N_12483,N_12790);
and U16489 (N_16489,N_14717,N_10931);
or U16490 (N_16490,N_11287,N_11545);
or U16491 (N_16491,N_12397,N_12375);
nor U16492 (N_16492,N_13240,N_11110);
and U16493 (N_16493,N_11623,N_12939);
nor U16494 (N_16494,N_13217,N_12100);
nand U16495 (N_16495,N_12385,N_13523);
and U16496 (N_16496,N_10715,N_12497);
or U16497 (N_16497,N_13269,N_10319);
and U16498 (N_16498,N_12738,N_11771);
and U16499 (N_16499,N_14493,N_13612);
nor U16500 (N_16500,N_14743,N_12450);
nand U16501 (N_16501,N_14569,N_12292);
or U16502 (N_16502,N_14068,N_10879);
or U16503 (N_16503,N_12257,N_10079);
nor U16504 (N_16504,N_12882,N_13356);
or U16505 (N_16505,N_12163,N_11894);
or U16506 (N_16506,N_14507,N_14910);
nor U16507 (N_16507,N_13430,N_13670);
nor U16508 (N_16508,N_11150,N_10076);
and U16509 (N_16509,N_10858,N_12189);
nand U16510 (N_16510,N_11624,N_11917);
nor U16511 (N_16511,N_10354,N_14805);
nand U16512 (N_16512,N_12301,N_14662);
nor U16513 (N_16513,N_12680,N_11849);
or U16514 (N_16514,N_10405,N_11187);
and U16515 (N_16515,N_13526,N_10557);
and U16516 (N_16516,N_12622,N_11102);
or U16517 (N_16517,N_12360,N_10497);
xor U16518 (N_16518,N_10945,N_11285);
and U16519 (N_16519,N_10234,N_12655);
nor U16520 (N_16520,N_13014,N_12333);
nor U16521 (N_16521,N_11583,N_11418);
nand U16522 (N_16522,N_14518,N_13637);
xor U16523 (N_16523,N_12222,N_12234);
nand U16524 (N_16524,N_12817,N_14336);
nand U16525 (N_16525,N_11647,N_12849);
nor U16526 (N_16526,N_11610,N_14397);
and U16527 (N_16527,N_10026,N_11365);
and U16528 (N_16528,N_14605,N_14657);
and U16529 (N_16529,N_12453,N_12860);
nand U16530 (N_16530,N_10666,N_14529);
nand U16531 (N_16531,N_13393,N_11870);
or U16532 (N_16532,N_14879,N_13270);
and U16533 (N_16533,N_13230,N_13446);
nand U16534 (N_16534,N_12018,N_12871);
or U16535 (N_16535,N_14829,N_11554);
xor U16536 (N_16536,N_13597,N_13147);
nor U16537 (N_16537,N_10658,N_14396);
or U16538 (N_16538,N_11063,N_14445);
nor U16539 (N_16539,N_13479,N_10441);
or U16540 (N_16540,N_12843,N_12073);
and U16541 (N_16541,N_10193,N_10167);
nand U16542 (N_16542,N_10641,N_12160);
nand U16543 (N_16543,N_12096,N_11091);
nor U16544 (N_16544,N_12071,N_14373);
xor U16545 (N_16545,N_11142,N_13231);
nand U16546 (N_16546,N_13632,N_13126);
or U16547 (N_16547,N_11748,N_10468);
nor U16548 (N_16548,N_10145,N_12031);
or U16549 (N_16549,N_12494,N_10386);
xnor U16550 (N_16550,N_10977,N_14851);
or U16551 (N_16551,N_13536,N_11914);
or U16552 (N_16552,N_11579,N_10692);
and U16553 (N_16553,N_10638,N_12455);
nand U16554 (N_16554,N_10371,N_11144);
nand U16555 (N_16555,N_14811,N_13054);
nand U16556 (N_16556,N_13498,N_12070);
nand U16557 (N_16557,N_14217,N_14489);
or U16558 (N_16558,N_13777,N_14034);
nand U16559 (N_16559,N_13956,N_14311);
or U16560 (N_16560,N_13052,N_11209);
and U16561 (N_16561,N_13109,N_11413);
nor U16562 (N_16562,N_14079,N_13111);
and U16563 (N_16563,N_11243,N_11302);
or U16564 (N_16564,N_11164,N_13353);
xor U16565 (N_16565,N_12263,N_11169);
nand U16566 (N_16566,N_10433,N_14905);
nand U16567 (N_16567,N_13502,N_13596);
or U16568 (N_16568,N_12555,N_13328);
and U16569 (N_16569,N_14576,N_11987);
nand U16570 (N_16570,N_11769,N_10979);
xnor U16571 (N_16571,N_11385,N_14594);
nor U16572 (N_16572,N_10179,N_14377);
nand U16573 (N_16573,N_10717,N_14669);
nor U16574 (N_16574,N_13921,N_14411);
xnor U16575 (N_16575,N_12977,N_14090);
xor U16576 (N_16576,N_14074,N_13441);
nor U16577 (N_16577,N_13569,N_12201);
nor U16578 (N_16578,N_10350,N_14885);
or U16579 (N_16579,N_14742,N_14780);
or U16580 (N_16580,N_13966,N_12064);
and U16581 (N_16581,N_14355,N_13210);
nor U16582 (N_16582,N_14674,N_14987);
or U16583 (N_16583,N_12193,N_13497);
or U16584 (N_16584,N_12546,N_13802);
or U16585 (N_16585,N_11295,N_14922);
or U16586 (N_16586,N_14204,N_13515);
nor U16587 (N_16587,N_10852,N_11911);
nand U16588 (N_16588,N_13267,N_13618);
xnor U16589 (N_16589,N_14577,N_11544);
nor U16590 (N_16590,N_10558,N_11157);
or U16591 (N_16591,N_14449,N_12819);
nor U16592 (N_16592,N_14206,N_13365);
and U16593 (N_16593,N_11768,N_13124);
or U16594 (N_16594,N_11100,N_12334);
nor U16595 (N_16595,N_11742,N_12598);
and U16596 (N_16596,N_13579,N_12918);
nor U16597 (N_16597,N_13528,N_14374);
and U16598 (N_16598,N_11880,N_13776);
xnor U16599 (N_16599,N_11306,N_11799);
and U16600 (N_16600,N_11123,N_13282);
and U16601 (N_16601,N_10588,N_11620);
and U16602 (N_16602,N_14339,N_13407);
xor U16603 (N_16603,N_13796,N_10474);
nand U16604 (N_16604,N_14909,N_13788);
nor U16605 (N_16605,N_12478,N_13221);
and U16606 (N_16606,N_11130,N_14175);
xor U16607 (N_16607,N_11183,N_14052);
nand U16608 (N_16608,N_13019,N_14598);
nand U16609 (N_16609,N_14993,N_11787);
and U16610 (N_16610,N_10249,N_10532);
nor U16611 (N_16611,N_11093,N_11060);
nand U16612 (N_16612,N_13932,N_11584);
xor U16613 (N_16613,N_14771,N_11736);
and U16614 (N_16614,N_11747,N_10100);
or U16615 (N_16615,N_12371,N_10187);
nand U16616 (N_16616,N_13144,N_13908);
or U16617 (N_16617,N_13588,N_11274);
xor U16618 (N_16618,N_11792,N_12484);
and U16619 (N_16619,N_12158,N_13604);
xnor U16620 (N_16620,N_14348,N_14494);
xnor U16621 (N_16621,N_14904,N_12928);
xnor U16622 (N_16622,N_12240,N_10610);
nor U16623 (N_16623,N_11553,N_11296);
nand U16624 (N_16624,N_10907,N_10581);
and U16625 (N_16625,N_14646,N_12467);
nand U16626 (N_16626,N_13718,N_12694);
and U16627 (N_16627,N_13302,N_10141);
nor U16628 (N_16628,N_12740,N_14597);
or U16629 (N_16629,N_10168,N_10401);
nand U16630 (N_16630,N_10266,N_11998);
or U16631 (N_16631,N_13848,N_11226);
nand U16632 (N_16632,N_14025,N_11220);
nand U16633 (N_16633,N_10206,N_12275);
and U16634 (N_16634,N_10822,N_14222);
or U16635 (N_16635,N_10679,N_10308);
nand U16636 (N_16636,N_14798,N_10149);
or U16637 (N_16637,N_11635,N_12143);
nor U16638 (N_16638,N_13736,N_11381);
xor U16639 (N_16639,N_14814,N_11954);
xor U16640 (N_16640,N_12663,N_11453);
nand U16641 (N_16641,N_11593,N_14969);
or U16642 (N_16642,N_11957,N_13519);
nor U16643 (N_16643,N_10364,N_13351);
nor U16644 (N_16644,N_11904,N_13252);
xor U16645 (N_16645,N_13904,N_12537);
xor U16646 (N_16646,N_14246,N_10509);
nor U16647 (N_16647,N_10571,N_10467);
or U16648 (N_16648,N_10417,N_14694);
and U16649 (N_16649,N_12289,N_12600);
nand U16650 (N_16650,N_14031,N_14920);
nor U16651 (N_16651,N_12519,N_14420);
nor U16652 (N_16652,N_12914,N_12754);
nor U16653 (N_16653,N_10052,N_14698);
xnor U16654 (N_16654,N_12742,N_11596);
xor U16655 (N_16655,N_12561,N_14391);
nor U16656 (N_16656,N_13474,N_11537);
nand U16657 (N_16657,N_10862,N_10484);
and U16658 (N_16658,N_13385,N_11960);
nor U16659 (N_16659,N_12415,N_13162);
and U16660 (N_16660,N_13118,N_12125);
nor U16661 (N_16661,N_13176,N_10627);
or U16662 (N_16662,N_13244,N_11659);
or U16663 (N_16663,N_10734,N_12566);
nor U16664 (N_16664,N_10260,N_10890);
nand U16665 (N_16665,N_11065,N_11656);
nand U16666 (N_16666,N_13122,N_11706);
or U16667 (N_16667,N_11923,N_13432);
and U16668 (N_16668,N_13626,N_13140);
nand U16669 (N_16669,N_14623,N_14106);
and U16670 (N_16670,N_12748,N_13584);
or U16671 (N_16671,N_13743,N_14303);
and U16672 (N_16672,N_14603,N_12084);
nor U16673 (N_16673,N_11168,N_13452);
or U16674 (N_16674,N_13059,N_12608);
and U16675 (N_16675,N_12997,N_13301);
and U16676 (N_16676,N_12337,N_14713);
nand U16677 (N_16677,N_11576,N_10872);
nor U16678 (N_16678,N_12509,N_14080);
nor U16679 (N_16679,N_14630,N_11466);
and U16680 (N_16680,N_14250,N_12119);
nor U16681 (N_16681,N_11406,N_14975);
nand U16682 (N_16682,N_10544,N_13728);
nand U16683 (N_16683,N_11284,N_14744);
nor U16684 (N_16684,N_11464,N_13204);
nor U16685 (N_16685,N_10106,N_10080);
nor U16686 (N_16686,N_13202,N_12596);
and U16687 (N_16687,N_11499,N_13552);
nand U16688 (N_16688,N_14715,N_11200);
or U16689 (N_16689,N_13078,N_14072);
and U16690 (N_16690,N_14848,N_11511);
nand U16691 (N_16691,N_12722,N_10081);
nand U16692 (N_16692,N_12866,N_13175);
xor U16693 (N_16693,N_14859,N_13924);
or U16694 (N_16694,N_12065,N_10275);
or U16695 (N_16695,N_12844,N_11008);
or U16696 (N_16696,N_11042,N_12745);
or U16697 (N_16697,N_14738,N_14736);
xor U16698 (N_16698,N_12013,N_14644);
and U16699 (N_16699,N_14322,N_14619);
nand U16700 (N_16700,N_11808,N_11632);
or U16701 (N_16701,N_10624,N_11115);
nand U16702 (N_16702,N_13429,N_11812);
and U16703 (N_16703,N_10824,N_14815);
and U16704 (N_16704,N_13986,N_13247);
nand U16705 (N_16705,N_11145,N_14536);
nand U16706 (N_16706,N_10677,N_13971);
nor U16707 (N_16707,N_14727,N_14437);
or U16708 (N_16708,N_13729,N_13779);
or U16709 (N_16709,N_14783,N_11735);
or U16710 (N_16710,N_14119,N_12727);
xor U16711 (N_16711,N_13567,N_11273);
and U16712 (N_16712,N_12274,N_12574);
nor U16713 (N_16713,N_14491,N_11404);
nor U16714 (N_16714,N_11621,N_14057);
nand U16715 (N_16715,N_11714,N_11652);
and U16716 (N_16716,N_12853,N_10379);
xnor U16717 (N_16717,N_11655,N_12310);
nand U16718 (N_16718,N_10320,N_13693);
nor U16719 (N_16719,N_10636,N_10788);
nor U16720 (N_16720,N_13675,N_13836);
and U16721 (N_16721,N_10623,N_14761);
nor U16722 (N_16722,N_14668,N_13649);
nor U16723 (N_16723,N_10854,N_11574);
nand U16724 (N_16724,N_14435,N_10963);
nand U16725 (N_16725,N_14014,N_11578);
or U16726 (N_16726,N_12932,N_12156);
or U16727 (N_16727,N_11489,N_14794);
or U16728 (N_16728,N_11828,N_13024);
nor U16729 (N_16729,N_10595,N_10201);
nand U16730 (N_16730,N_14830,N_10276);
nor U16731 (N_16731,N_13967,N_10110);
nand U16732 (N_16732,N_12075,N_11105);
nand U16733 (N_16733,N_12116,N_12551);
nor U16734 (N_16734,N_14306,N_10648);
nand U16735 (N_16735,N_11744,N_12108);
nand U16736 (N_16736,N_12720,N_14368);
nand U16737 (N_16737,N_13658,N_14267);
and U16738 (N_16738,N_12117,N_10835);
nand U16739 (N_16739,N_11970,N_11283);
xnor U16740 (N_16740,N_11429,N_12826);
nand U16741 (N_16741,N_11818,N_11822);
and U16742 (N_16742,N_12253,N_13289);
or U16743 (N_16743,N_10634,N_14407);
and U16744 (N_16744,N_10741,N_11536);
and U16745 (N_16745,N_10743,N_13577);
or U16746 (N_16746,N_11749,N_11467);
and U16747 (N_16747,N_13730,N_14308);
and U16748 (N_16748,N_11776,N_14648);
and U16749 (N_16749,N_10277,N_10073);
and U16750 (N_16750,N_14523,N_10880);
or U16751 (N_16751,N_10914,N_11081);
and U16752 (N_16752,N_11088,N_11343);
nand U16753 (N_16753,N_11629,N_13732);
nor U16754 (N_16754,N_14610,N_14129);
nand U16755 (N_16755,N_13002,N_11899);
nor U16756 (N_16756,N_10842,N_11816);
xor U16757 (N_16757,N_14459,N_14980);
nor U16758 (N_16758,N_14884,N_11663);
and U16759 (N_16759,N_14834,N_12449);
xor U16760 (N_16760,N_14655,N_14482);
nand U16761 (N_16761,N_13051,N_12823);
nand U16762 (N_16762,N_14041,N_13263);
and U16763 (N_16763,N_12330,N_14752);
or U16764 (N_16764,N_14415,N_14166);
and U16765 (N_16765,N_14342,N_14354);
nand U16766 (N_16766,N_13570,N_11494);
nand U16767 (N_16767,N_12402,N_12768);
xnor U16768 (N_16768,N_12436,N_12699);
nand U16769 (N_16769,N_14967,N_14323);
or U16770 (N_16770,N_12833,N_14502);
nor U16771 (N_16771,N_12602,N_12535);
or U16772 (N_16772,N_14520,N_13969);
nor U16773 (N_16773,N_12299,N_14191);
and U16774 (N_16774,N_10191,N_12668);
xnor U16775 (N_16775,N_13977,N_12481);
nand U16776 (N_16776,N_12958,N_10905);
xnor U16777 (N_16777,N_13572,N_14748);
nor U16778 (N_16778,N_13089,N_13688);
xor U16779 (N_16779,N_13290,N_13336);
nor U16780 (N_16780,N_12794,N_10451);
and U16781 (N_16781,N_12935,N_14002);
and U16782 (N_16782,N_14807,N_10165);
nor U16783 (N_16783,N_11919,N_10387);
or U16784 (N_16784,N_14914,N_11594);
or U16785 (N_16785,N_12852,N_14504);
nand U16786 (N_16786,N_13650,N_11048);
nor U16787 (N_16787,N_12657,N_13864);
nand U16788 (N_16788,N_11670,N_13174);
xnor U16789 (N_16789,N_10184,N_14208);
and U16790 (N_16790,N_14422,N_14352);
or U16791 (N_16791,N_10242,N_10058);
nor U16792 (N_16792,N_11328,N_10107);
nor U16793 (N_16793,N_12298,N_14906);
xnor U16794 (N_16794,N_11389,N_13061);
xor U16795 (N_16795,N_10825,N_13615);
or U16796 (N_16796,N_14649,N_11687);
or U16797 (N_16797,N_11454,N_11432);
or U16798 (N_16798,N_14263,N_12030);
xor U16799 (N_16799,N_13501,N_10740);
nor U16800 (N_16800,N_13516,N_11503);
nor U16801 (N_16801,N_14221,N_14444);
nand U16802 (N_16802,N_10755,N_12172);
nor U16803 (N_16803,N_14801,N_13345);
nor U16804 (N_16804,N_14654,N_12847);
nand U16805 (N_16805,N_12804,N_13926);
or U16806 (N_16806,N_14705,N_11961);
or U16807 (N_16807,N_11324,N_11194);
or U16808 (N_16808,N_10461,N_13366);
nor U16809 (N_16809,N_12488,N_10747);
xor U16810 (N_16810,N_13853,N_10545);
xnor U16811 (N_16811,N_10491,N_12178);
or U16812 (N_16812,N_14078,N_14473);
and U16813 (N_16813,N_12212,N_12703);
or U16814 (N_16814,N_14216,N_12927);
nor U16815 (N_16815,N_10395,N_10647);
nor U16816 (N_16816,N_12524,N_13951);
xor U16817 (N_16817,N_11293,N_12028);
and U16818 (N_16818,N_10245,N_12139);
or U16819 (N_16819,N_11303,N_10068);
nand U16820 (N_16820,N_13982,N_12132);
and U16821 (N_16821,N_12527,N_13903);
xnor U16822 (N_16822,N_13426,N_12906);
and U16823 (N_16823,N_10336,N_10832);
nor U16824 (N_16824,N_12003,N_11715);
nand U16825 (N_16825,N_10071,N_13535);
xor U16826 (N_16826,N_14684,N_12303);
and U16827 (N_16827,N_12198,N_14582);
or U16828 (N_16828,N_13000,N_13970);
or U16829 (N_16829,N_11806,N_11206);
or U16830 (N_16830,N_11015,N_10674);
and U16831 (N_16831,N_13634,N_13107);
nand U16832 (N_16832,N_10668,N_11974);
nor U16833 (N_16833,N_11443,N_12889);
or U16834 (N_16834,N_13672,N_10050);
and U16835 (N_16835,N_11575,N_10399);
and U16836 (N_16836,N_14960,N_10519);
nand U16837 (N_16837,N_12177,N_11722);
nand U16838 (N_16838,N_13042,N_10920);
or U16839 (N_16839,N_12776,N_13076);
nor U16840 (N_16840,N_10869,N_14624);
nor U16841 (N_16841,N_13321,N_12214);
nand U16842 (N_16842,N_12921,N_14044);
nand U16843 (N_16843,N_12391,N_14181);
nand U16844 (N_16844,N_14350,N_10597);
and U16845 (N_16845,N_11344,N_12715);
nand U16846 (N_16846,N_14769,N_11118);
xnor U16847 (N_16847,N_13006,N_10790);
nor U16848 (N_16848,N_14413,N_11291);
and U16849 (N_16849,N_11526,N_11146);
or U16850 (N_16850,N_13514,N_13421);
and U16851 (N_16851,N_11190,N_13132);
and U16852 (N_16852,N_12544,N_14113);
and U16853 (N_16853,N_12247,N_10208);
or U16854 (N_16854,N_11803,N_11281);
nand U16855 (N_16855,N_13700,N_10020);
or U16856 (N_16856,N_13895,N_13333);
nor U16857 (N_16857,N_14640,N_11097);
nor U16858 (N_16858,N_14667,N_11667);
nand U16859 (N_16859,N_10929,N_14274);
or U16860 (N_16860,N_13380,N_11022);
nor U16861 (N_16861,N_13442,N_14089);
nor U16862 (N_16862,N_14344,N_12165);
nor U16863 (N_16863,N_11258,N_12444);
nand U16864 (N_16864,N_10645,N_13486);
nand U16865 (N_16865,N_11516,N_10804);
nand U16866 (N_16866,N_12147,N_12789);
or U16867 (N_16867,N_14671,N_12151);
nand U16868 (N_16868,N_13392,N_14367);
and U16869 (N_16869,N_13994,N_10446);
or U16870 (N_16870,N_12349,N_13770);
and U16871 (N_16871,N_13130,N_11839);
nor U16872 (N_16872,N_10953,N_14483);
and U16873 (N_16873,N_10432,N_11847);
nand U16874 (N_16874,N_11383,N_14153);
and U16875 (N_16875,N_14995,N_12427);
or U16876 (N_16876,N_14133,N_11895);
or U16877 (N_16877,N_14235,N_10702);
and U16878 (N_16878,N_13878,N_12755);
nand U16879 (N_16879,N_11739,N_13499);
and U16880 (N_16880,N_11366,N_14935);
or U16881 (N_16881,N_13460,N_10450);
and U16882 (N_16882,N_11478,N_10256);
nand U16883 (N_16883,N_11965,N_11430);
nand U16884 (N_16884,N_12205,N_10783);
or U16885 (N_16885,N_11950,N_13427);
nand U16886 (N_16886,N_12398,N_10285);
xor U16887 (N_16887,N_12474,N_11804);
nor U16888 (N_16888,N_10166,N_13996);
nor U16889 (N_16889,N_11402,N_11162);
and U16890 (N_16890,N_14764,N_14366);
nand U16891 (N_16891,N_11550,N_12990);
and U16892 (N_16892,N_12328,N_14606);
xor U16893 (N_16893,N_13008,N_11333);
nor U16894 (N_16894,N_14946,N_10430);
and U16895 (N_16895,N_11509,N_11249);
nor U16896 (N_16896,N_12926,N_11262);
nand U16897 (N_16897,N_14177,N_13825);
nand U16898 (N_16898,N_14861,N_11069);
and U16899 (N_16899,N_13058,N_13075);
and U16900 (N_16900,N_13983,N_13581);
and U16901 (N_16901,N_14555,N_11547);
or U16902 (N_16902,N_12580,N_11936);
or U16903 (N_16903,N_13608,N_10958);
nor U16904 (N_16904,N_14521,N_13662);
nor U16905 (N_16905,N_14972,N_10607);
and U16906 (N_16906,N_10635,N_10346);
nor U16907 (N_16907,N_12943,N_13317);
or U16908 (N_16908,N_14131,N_10304);
or U16909 (N_16909,N_12459,N_14156);
or U16910 (N_16910,N_10129,N_14824);
nor U16911 (N_16911,N_14143,N_14393);
nor U16912 (N_16912,N_10760,N_11559);
nor U16913 (N_16913,N_13065,N_10036);
or U16914 (N_16914,N_10671,N_11560);
or U16915 (N_16915,N_13865,N_13795);
xor U16916 (N_16916,N_14353,N_14800);
and U16917 (N_16917,N_11875,N_12877);
nor U16918 (N_16918,N_13603,N_11122);
nor U16919 (N_16919,N_12672,N_12893);
and U16920 (N_16920,N_11969,N_11615);
and U16921 (N_16921,N_11475,N_11723);
nor U16922 (N_16922,N_10828,N_11518);
nor U16923 (N_16923,N_12937,N_10156);
nor U16924 (N_16924,N_12376,N_14916);
nand U16925 (N_16925,N_11939,N_13859);
nand U16926 (N_16926,N_13964,N_14809);
or U16927 (N_16927,N_14976,N_10057);
nand U16928 (N_16928,N_11572,N_10546);
or U16929 (N_16929,N_13377,N_13950);
nor U16930 (N_16930,N_11850,N_10792);
and U16931 (N_16931,N_11049,N_13113);
nor U16932 (N_16932,N_11448,N_11910);
nand U16933 (N_16933,N_13659,N_13899);
nor U16934 (N_16934,N_12992,N_10657);
nor U16935 (N_16935,N_12959,N_12388);
or U16936 (N_16936,N_11607,N_13091);
and U16937 (N_16937,N_14194,N_13030);
and U16938 (N_16938,N_13410,N_12161);
and U16939 (N_16939,N_10074,N_11113);
xor U16940 (N_16940,N_10859,N_12246);
nor U16941 (N_16941,N_12086,N_10173);
and U16942 (N_16942,N_14230,N_11057);
and U16943 (N_16943,N_11921,N_13504);
or U16944 (N_16944,N_10329,N_12093);
nand U16945 (N_16945,N_11447,N_13138);
nand U16946 (N_16946,N_10477,N_10023);
or U16947 (N_16947,N_14085,N_12317);
or U16948 (N_16948,N_11521,N_12646);
or U16949 (N_16949,N_11704,N_14003);
and U16950 (N_16950,N_10121,N_13450);
nor U16951 (N_16951,N_10922,N_13046);
xnor U16952 (N_16952,N_14497,N_11637);
nand U16953 (N_16953,N_10878,N_11884);
and U16954 (N_16954,N_12586,N_12846);
or U16955 (N_16955,N_12985,N_14775);
nand U16956 (N_16956,N_13093,N_13161);
and U16957 (N_16957,N_13490,N_10447);
nand U16958 (N_16958,N_10085,N_12285);
nand U16959 (N_16959,N_13171,N_10062);
and U16960 (N_16960,N_14998,N_13324);
nor U16961 (N_16961,N_12854,N_10381);
or U16962 (N_16962,N_14865,N_12633);
and U16963 (N_16963,N_11309,N_10765);
nand U16964 (N_16964,N_12730,N_12286);
and U16965 (N_16965,N_12057,N_11699);
nor U16966 (N_16966,N_13311,N_10377);
nand U16967 (N_16967,N_14612,N_14632);
nand U16968 (N_16968,N_11101,N_10933);
nand U16969 (N_16969,N_13797,N_12661);
nand U16970 (N_16970,N_11421,N_10284);
or U16971 (N_16971,N_14628,N_10769);
nor U16972 (N_16972,N_13332,N_10902);
or U16973 (N_16973,N_13236,N_13702);
and U16974 (N_16974,N_11988,N_10307);
nor U16975 (N_16975,N_11451,N_13974);
nor U16976 (N_16976,N_13606,N_13170);
and U16977 (N_16977,N_11726,N_13760);
nand U16978 (N_16978,N_11872,N_14176);
xor U16979 (N_16979,N_14791,N_14104);
nor U16980 (N_16980,N_13123,N_12540);
and U16981 (N_16981,N_14069,N_12272);
nand U16982 (N_16982,N_11422,N_10547);
and U16983 (N_16983,N_12485,N_11971);
nor U16984 (N_16984,N_12660,N_13574);
and U16985 (N_16985,N_12573,N_10072);
nor U16986 (N_16986,N_10147,N_14046);
nand U16987 (N_16987,N_13629,N_10986);
or U16988 (N_16988,N_13487,N_10418);
and U16989 (N_16989,N_13625,N_14275);
xnor U16990 (N_16990,N_10060,N_10612);
or U16991 (N_16991,N_11411,N_11038);
nor U16992 (N_16992,N_12702,N_12387);
and U16993 (N_16993,N_10831,N_10012);
and U16994 (N_16994,N_13381,N_12278);
and U16995 (N_16995,N_12892,N_12179);
nor U16996 (N_16996,N_10637,N_11973);
nand U16997 (N_16997,N_14019,N_11985);
xor U16998 (N_16998,N_12134,N_10703);
and U16999 (N_16999,N_13344,N_12331);
and U17000 (N_17000,N_12081,N_10347);
or U17001 (N_17001,N_14953,N_10040);
nand U17002 (N_17002,N_13819,N_14093);
or U17003 (N_17003,N_12707,N_14384);
xnor U17004 (N_17004,N_13929,N_11892);
nand U17005 (N_17005,N_12725,N_13850);
and U17006 (N_17006,N_10997,N_11952);
or U17007 (N_17007,N_14647,N_13232);
nand U17008 (N_17008,N_10803,N_12848);
xor U17009 (N_17009,N_14929,N_13203);
or U17010 (N_17010,N_12256,N_14149);
and U17011 (N_17011,N_14434,N_14269);
nor U17012 (N_17012,N_10039,N_13652);
and U17013 (N_17013,N_11322,N_13227);
and U17014 (N_17014,N_10124,N_12922);
and U17015 (N_17015,N_13105,N_13599);
nand U17016 (N_17016,N_12710,N_14813);
or U17017 (N_17017,N_12184,N_13077);
or U17018 (N_17018,N_14197,N_14130);
or U17019 (N_17019,N_13438,N_10572);
nor U17020 (N_17020,N_13110,N_14892);
nor U17021 (N_17021,N_13266,N_11625);
nor U17022 (N_17022,N_10426,N_13219);
and U17023 (N_17023,N_12089,N_11916);
xnor U17024 (N_17024,N_10550,N_14734);
or U17025 (N_17025,N_13548,N_11569);
or U17026 (N_17026,N_14033,N_14464);
nor U17027 (N_17027,N_13617,N_10749);
and U17028 (N_17028,N_12808,N_11577);
or U17029 (N_17029,N_13422,N_10392);
or U17030 (N_17030,N_12051,N_13031);
nand U17031 (N_17031,N_11721,N_11548);
nand U17032 (N_17032,N_12897,N_13622);
nor U17033 (N_17033,N_10932,N_11054);
and U17034 (N_17034,N_10470,N_10672);
nand U17035 (N_17035,N_10746,N_12056);
nor U17036 (N_17036,N_11424,N_11908);
nor U17037 (N_17037,N_13082,N_11350);
nand U17038 (N_17038,N_11520,N_14264);
and U17039 (N_17039,N_10846,N_13508);
nand U17040 (N_17040,N_14587,N_10796);
xor U17041 (N_17041,N_11943,N_10808);
nor U17042 (N_17042,N_12957,N_12440);
nand U17043 (N_17043,N_11930,N_12429);
and U17044 (N_17044,N_12355,N_13958);
or U17045 (N_17045,N_12589,N_10795);
and U17046 (N_17046,N_14620,N_13571);
nor U17047 (N_17047,N_13478,N_14609);
nor U17048 (N_17048,N_10241,N_11626);
nand U17049 (N_17049,N_13537,N_10620);
nand U17050 (N_17050,N_13778,N_11949);
nor U17051 (N_17051,N_10175,N_13936);
xor U17052 (N_17052,N_13805,N_14517);
xor U17053 (N_17053,N_14188,N_11271);
xor U17054 (N_17054,N_12869,N_13455);
nor U17055 (N_17055,N_14664,N_11132);
or U17056 (N_17056,N_10861,N_12824);
and U17057 (N_17057,N_12060,N_12832);
and U17058 (N_17058,N_14022,N_13768);
nand U17059 (N_17059,N_13669,N_10708);
xnor U17060 (N_17060,N_14361,N_10006);
nand U17061 (N_17061,N_14902,N_12538);
and U17062 (N_17062,N_14501,N_14936);
and U17063 (N_17063,N_12850,N_14806);
or U17064 (N_17064,N_11182,N_10748);
xor U17065 (N_17065,N_10936,N_10643);
nand U17066 (N_17066,N_10901,N_10032);
or U17067 (N_17067,N_14296,N_14026);
nand U17068 (N_17068,N_12525,N_13708);
xor U17069 (N_17069,N_11221,N_14351);
and U17070 (N_17070,N_11741,N_10733);
xor U17071 (N_17071,N_14913,N_14290);
nor U17072 (N_17072,N_10114,N_10056);
and U17073 (N_17073,N_13656,N_12456);
nor U17074 (N_17074,N_12428,N_10136);
or U17075 (N_17075,N_12036,N_14996);
nor U17076 (N_17076,N_12146,N_10311);
and U17077 (N_17077,N_14777,N_12150);
or U17078 (N_17078,N_10916,N_11056);
and U17079 (N_17079,N_10609,N_12470);
nand U17080 (N_17080,N_10919,N_14406);
nand U17081 (N_17081,N_10407,N_12764);
nand U17082 (N_17082,N_11352,N_14544);
or U17083 (N_17083,N_14028,N_12625);
or U17084 (N_17084,N_13359,N_12964);
xnor U17085 (N_17085,N_13239,N_13976);
and U17086 (N_17086,N_10604,N_14519);
and U17087 (N_17087,N_13842,N_10974);
or U17088 (N_17088,N_14287,N_13999);
nor U17089 (N_17089,N_10186,N_14480);
or U17090 (N_17090,N_12479,N_10372);
nor U17091 (N_17091,N_11886,N_11829);
or U17092 (N_17092,N_13213,N_11539);
and U17093 (N_17093,N_10662,N_13456);
nor U17094 (N_17094,N_10221,N_12518);
nor U17095 (N_17095,N_14164,N_10416);
nand U17096 (N_17096,N_10368,N_13029);
xor U17097 (N_17097,N_11364,N_14399);
nor U17098 (N_17098,N_12732,N_13223);
nand U17099 (N_17099,N_11802,N_12611);
and U17100 (N_17100,N_10965,N_10338);
nor U17101 (N_17101,N_14723,N_11780);
and U17102 (N_17102,N_12369,N_10421);
nor U17103 (N_17103,N_13522,N_10791);
nor U17104 (N_17104,N_12361,N_10419);
nand U17105 (N_17105,N_14259,N_14903);
and U17106 (N_17106,N_13739,N_12688);
nand U17107 (N_17107,N_11320,N_11571);
and U17108 (N_17108,N_13216,N_12118);
nand U17109 (N_17109,N_13334,N_12896);
and U17110 (N_17110,N_12142,N_14081);
or U17111 (N_17111,N_12983,N_11840);
nand U17112 (N_17112,N_12155,N_13320);
nand U17113 (N_17113,N_11963,N_10310);
nand U17114 (N_17114,N_11252,N_13747);
nand U17115 (N_17115,N_12447,N_14099);
nand U17116 (N_17116,N_12396,N_13180);
nor U17117 (N_17117,N_10391,N_14172);
or U17118 (N_17118,N_11878,N_12763);
and U17119 (N_17119,N_11255,N_13806);
or U17120 (N_17120,N_10821,N_12665);
nor U17121 (N_17121,N_12865,N_13933);
or U17122 (N_17122,N_12441,N_14317);
or U17123 (N_17123,N_12554,N_10493);
and U17124 (N_17124,N_12899,N_12469);
nand U17125 (N_17125,N_11529,N_13517);
nand U17126 (N_17126,N_12697,N_11882);
and U17127 (N_17127,N_13849,N_12025);
and U17128 (N_17128,N_14205,N_10228);
or U17129 (N_17129,N_10522,N_10983);
and U17130 (N_17130,N_13772,N_13812);
or U17131 (N_17131,N_13347,N_10845);
and U17132 (N_17132,N_11039,N_12857);
and U17133 (N_17133,N_13294,N_12905);
and U17134 (N_17134,N_11857,N_10843);
nand U17135 (N_17135,N_12451,N_12976);
and U17136 (N_17136,N_11864,N_13297);
nand U17137 (N_17137,N_13309,N_14804);
xor U17138 (N_17138,N_13485,N_14051);
and U17139 (N_17139,N_13847,N_14835);
or U17140 (N_17140,N_12862,N_12500);
or U17141 (N_17141,N_14812,N_10507);
nor U17142 (N_17142,N_12606,N_14831);
nor U17143 (N_17143,N_11217,N_14816);
nand U17144 (N_17144,N_12062,N_11530);
nand U17145 (N_17145,N_12466,N_13248);
nand U17146 (N_17146,N_11055,N_10829);
nor U17147 (N_17147,N_14220,N_12758);
and U17148 (N_17148,N_10196,N_12175);
nand U17149 (N_17149,N_14485,N_12604);
nand U17150 (N_17150,N_11269,N_14142);
or U17151 (N_17151,N_11531,N_10199);
nor U17152 (N_17152,N_13888,N_12807);
or U17153 (N_17153,N_13644,N_13218);
and U17154 (N_17154,N_11078,N_14448);
nand U17155 (N_17155,N_14447,N_10506);
xor U17156 (N_17156,N_14666,N_11452);
or U17157 (N_17157,N_11289,N_11020);
and U17158 (N_17158,N_10617,N_14218);
nor U17159 (N_17159,N_12812,N_14695);
and U17160 (N_17160,N_11077,N_12493);
or U17161 (N_17161,N_12999,N_10211);
nand U17162 (N_17162,N_14398,N_13824);
and U17163 (N_17163,N_10659,N_10851);
or U17164 (N_17164,N_14894,N_13592);
xor U17165 (N_17165,N_10282,N_14372);
nand U17166 (N_17166,N_11846,N_13691);
xnor U17167 (N_17167,N_11925,N_11237);
nand U17168 (N_17168,N_11972,N_11315);
or U17169 (N_17169,N_11213,N_10182);
or U17170 (N_17170,N_13568,N_11139);
nand U17171 (N_17171,N_14389,N_11059);
nor U17172 (N_17172,N_14059,N_14650);
nor U17173 (N_17173,N_14370,N_13724);
or U17174 (N_17174,N_12874,N_14101);
nor U17175 (N_17175,N_12811,N_10807);
nand U17176 (N_17176,N_11527,N_13803);
or U17177 (N_17177,N_12616,N_14927);
nor U17178 (N_17178,N_12149,N_11712);
nand U17179 (N_17179,N_10393,N_11617);
nand U17180 (N_17180,N_11390,N_12344);
nor U17181 (N_17181,N_12435,N_13915);
nor U17182 (N_17182,N_13420,N_14462);
nor U17183 (N_17183,N_11519,N_12516);
nor U17184 (N_17184,N_11779,N_12238);
nor U17185 (N_17185,N_12670,N_12389);
and U17186 (N_17186,N_12076,N_11471);
and U17187 (N_17187,N_13714,N_13645);
nor U17188 (N_17188,N_10463,N_12219);
nand U17189 (N_17189,N_12323,N_14062);
nand U17190 (N_17190,N_13529,N_10291);
nand U17191 (N_17191,N_14196,N_11587);
nand U17192 (N_17192,N_12885,N_10947);
nor U17193 (N_17193,N_11595,N_12879);
or U17194 (N_17194,N_11203,N_10061);
nand U17195 (N_17195,N_11627,N_12522);
and U17196 (N_17196,N_12759,N_12221);
nand U17197 (N_17197,N_11801,N_12890);
nand U17198 (N_17198,N_12578,N_10793);
nand U17199 (N_17199,N_12553,N_14472);
nor U17200 (N_17200,N_12650,N_11684);
nor U17201 (N_17201,N_12446,N_13160);
nor U17202 (N_17202,N_11018,N_11131);
nor U17203 (N_17203,N_11966,N_12215);
nor U17204 (N_17204,N_12044,N_13871);
nor U17205 (N_17205,N_10883,N_11668);
or U17206 (N_17206,N_13463,N_10318);
xor U17207 (N_17207,N_14836,N_10830);
nand U17208 (N_17208,N_12919,N_11282);
or U17209 (N_17209,N_11127,N_12557);
or U17210 (N_17210,N_10183,N_14063);
or U17211 (N_17211,N_11724,N_12098);
nor U17212 (N_17212,N_10443,N_11825);
nand U17213 (N_17213,N_14225,N_11140);
and U17214 (N_17214,N_14020,N_11353);
nor U17215 (N_17215,N_13793,N_14926);
nor U17216 (N_17216,N_10716,N_13835);
xnor U17217 (N_17217,N_10887,N_12870);
nand U17218 (N_17218,N_13382,N_10611);
or U17219 (N_17219,N_11003,N_13409);
or U17220 (N_17220,N_10652,N_11035);
nor U17221 (N_17221,N_11178,N_14229);
or U17222 (N_17222,N_12372,N_10007);
and U17223 (N_17223,N_13830,N_14982);
nor U17224 (N_17224,N_14707,N_12040);
nor U17225 (N_17225,N_10409,N_11297);
or U17226 (N_17226,N_10309,N_11912);
nand U17227 (N_17227,N_14754,N_11004);
nor U17228 (N_17228,N_14857,N_13493);
and U17229 (N_17229,N_14185,N_13090);
and U17230 (N_17230,N_11000,N_12168);
or U17231 (N_17231,N_10248,N_12796);
nor U17232 (N_17232,N_10190,N_10412);
nand U17233 (N_17233,N_11141,N_10819);
nand U17234 (N_17234,N_10707,N_13273);
nand U17235 (N_17235,N_13583,N_13935);
nor U17236 (N_17236,N_14346,N_11645);
and U17237 (N_17237,N_10345,N_11832);
and U17238 (N_17238,N_11842,N_12941);
and U17239 (N_17239,N_12541,N_14477);
and U17240 (N_17240,N_10176,N_14198);
xnor U17241 (N_17241,N_13741,N_13875);
nor U17242 (N_17242,N_10894,N_10362);
nand U17243 (N_17243,N_13804,N_14676);
xnor U17244 (N_17244,N_11508,N_14686);
and U17245 (N_17245,N_14790,N_10833);
nor U17246 (N_17246,N_14460,N_12316);
and U17247 (N_17247,N_12218,N_14690);
xor U17248 (N_17248,N_13642,N_12577);
and U17249 (N_17249,N_10414,N_12562);
nand U17250 (N_17250,N_14876,N_14345);
and U17251 (N_17251,N_10694,N_12492);
and U17252 (N_17252,N_14297,N_14784);
and U17253 (N_17253,N_12831,N_11265);
nor U17254 (N_17254,N_11089,N_10115);
and U17255 (N_17255,N_12454,N_11372);
and U17256 (N_17256,N_12830,N_10930);
nor U17257 (N_17257,N_10280,N_12950);
or U17258 (N_17258,N_11942,N_13235);
or U17259 (N_17259,N_14537,N_11210);
nand U17260 (N_17260,N_12972,N_13312);
or U17261 (N_17261,N_14100,N_13129);
or U17262 (N_17262,N_11386,N_11235);
and U17263 (N_17263,N_14357,N_14817);
or U17264 (N_17264,N_12587,N_12556);
and U17265 (N_17265,N_11032,N_11186);
nand U17266 (N_17266,N_10254,N_14238);
nand U17267 (N_17267,N_11198,N_12662);
nor U17268 (N_17268,N_14891,N_11438);
and U17269 (N_17269,N_14108,N_14589);
or U17270 (N_17270,N_13883,N_12063);
or U17271 (N_17271,N_10126,N_13814);
xnor U17272 (N_17272,N_11506,N_10625);
and U17273 (N_17273,N_10035,N_11931);
nand U17274 (N_17274,N_14038,N_14193);
and U17275 (N_17275,N_10352,N_10838);
and U17276 (N_17276,N_10651,N_11397);
nand U17277 (N_17277,N_13503,N_12159);
nand U17278 (N_17278,N_14724,N_13761);
xor U17279 (N_17279,N_11030,N_11170);
or U17280 (N_17280,N_12024,N_14043);
or U17281 (N_17281,N_11651,N_14889);
nor U17282 (N_17282,N_12321,N_11212);
xnor U17283 (N_17283,N_11556,N_13136);
xor U17284 (N_17284,N_13326,N_10365);
and U17285 (N_17285,N_11176,N_13525);
nand U17286 (N_17286,N_14534,N_14546);
xor U17287 (N_17287,N_10316,N_13183);
or U17288 (N_17288,N_11044,N_10366);
or U17289 (N_17289,N_12264,N_14601);
nand U17290 (N_17290,N_10457,N_10990);
nor U17291 (N_17291,N_10094,N_12631);
nand U17292 (N_17292,N_10908,N_10108);
and U17293 (N_17293,N_13563,N_10632);
nor U17294 (N_17294,N_13413,N_13012);
and U17295 (N_17295,N_14505,N_14593);
and U17296 (N_17296,N_12774,N_11905);
and U17297 (N_17297,N_10357,N_10764);
xor U17298 (N_17298,N_10404,N_10605);
and U17299 (N_17299,N_14318,N_10051);
or U17300 (N_17300,N_13477,N_11831);
and U17301 (N_17301,N_11725,N_14111);
nor U17302 (N_17302,N_13325,N_13905);
or U17303 (N_17303,N_12782,N_13168);
and U17304 (N_17304,N_10725,N_14150);
nand U17305 (N_17305,N_12821,N_11275);
nand U17306 (N_17306,N_14719,N_14542);
nor U17307 (N_17307,N_10122,N_14854);
or U17308 (N_17308,N_13831,N_13038);
and U17309 (N_17309,N_10909,N_13234);
nor U17310 (N_17310,N_14496,N_11772);
nand U17311 (N_17311,N_11796,N_10757);
nor U17312 (N_17312,N_11154,N_13901);
nand U17313 (N_17313,N_10815,N_14169);
nor U17314 (N_17314,N_13119,N_10584);
xor U17315 (N_17315,N_13686,N_11843);
or U17316 (N_17316,N_14986,N_13605);
and U17317 (N_17317,N_12634,N_12092);
nor U17318 (N_17318,N_13624,N_13037);
nand U17319 (N_17319,N_12005,N_12909);
nor U17320 (N_17320,N_14642,N_13594);
nand U17321 (N_17321,N_10744,N_12211);
or U17322 (N_17322,N_11845,N_10711);
or U17323 (N_17323,N_13808,N_13531);
nand U17324 (N_17324,N_12279,N_11881);
and U17325 (N_17325,N_12026,N_12255);
nor U17326 (N_17326,N_12599,N_10396);
xnor U17327 (N_17327,N_11264,N_11359);
and U17328 (N_17328,N_13609,N_10323);
nor U17329 (N_17329,N_10731,N_11606);
xor U17330 (N_17330,N_10787,N_13703);
nand U17331 (N_17331,N_10912,N_14155);
and U17332 (N_17332,N_10603,N_11940);
xor U17333 (N_17333,N_11836,N_11964);
or U17334 (N_17334,N_11955,N_13258);
nand U17335 (N_17335,N_14347,N_14329);
or U17336 (N_17336,N_13673,N_12354);
nor U17337 (N_17337,N_12842,N_12630);
nor U17338 (N_17338,N_11360,N_13277);
or U17339 (N_17339,N_13639,N_12487);
and U17340 (N_17340,N_10876,N_11698);
nor U17341 (N_17341,N_10465,N_10850);
xor U17342 (N_17342,N_11425,N_12339);
or U17343 (N_17343,N_12664,N_10195);
nand U17344 (N_17344,N_11703,N_13342);
nand U17345 (N_17345,N_13394,N_13833);
and U17346 (N_17346,N_13910,N_11136);
xor U17347 (N_17347,N_14685,N_14893);
nand U17348 (N_17348,N_13697,N_13764);
xor U17349 (N_17349,N_14726,N_12691);
and U17350 (N_17350,N_12993,N_11755);
nor U17351 (N_17351,N_13723,N_10987);
nand U17352 (N_17352,N_13725,N_12325);
nor U17353 (N_17353,N_12512,N_12931);
xnor U17354 (N_17354,N_14272,N_11680);
and U17355 (N_17355,N_13035,N_11641);
or U17356 (N_17356,N_13972,N_11047);
nor U17357 (N_17357,N_14277,N_10303);
or U17358 (N_17358,N_12930,N_13495);
nor U17359 (N_17359,N_14380,N_11216);
or U17360 (N_17360,N_14709,N_12251);
or U17361 (N_17361,N_13894,N_11084);
or U17362 (N_17362,N_12940,N_10840);
nor U17363 (N_17363,N_13555,N_11763);
and U17364 (N_17364,N_12185,N_12001);
nand U17365 (N_17365,N_12547,N_11117);
and U17366 (N_17366,N_14621,N_10337);
nor U17367 (N_17367,N_12243,N_12496);
or U17368 (N_17368,N_14016,N_14487);
and U17369 (N_17369,N_14006,N_13466);
nor U17370 (N_17370,N_14937,N_11205);
or U17371 (N_17371,N_11986,N_13281);
xnor U17372 (N_17372,N_14138,N_14604);
and U17373 (N_17373,N_12141,N_10889);
nand U17374 (N_17374,N_13400,N_13343);
nor U17375 (N_17375,N_12280,N_11920);
and U17376 (N_17376,N_12805,N_14562);
nor U17377 (N_17377,N_13331,N_10848);
nor U17378 (N_17378,N_14823,N_10268);
or U17379 (N_17379,N_14901,N_10918);
nor U17380 (N_17380,N_13810,N_10598);
nand U17381 (N_17381,N_11214,N_14833);
nor U17382 (N_17382,N_13164,N_10683);
nand U17383 (N_17383,N_10587,N_10644);
nor U17384 (N_17384,N_12837,N_13909);
nand U17385 (N_17385,N_13017,N_13402);
or U17386 (N_17386,N_12572,N_11197);
and U17387 (N_17387,N_10881,N_10998);
or U17388 (N_17388,N_11664,N_12614);
nor U17389 (N_17389,N_11861,N_10633);
nor U17390 (N_17390,N_14490,N_12969);
nor U17391 (N_17391,N_12802,N_11410);
or U17392 (N_17392,N_12461,N_10664);
nand U17393 (N_17393,N_14215,N_14211);
or U17394 (N_17394,N_10502,N_12191);
or U17395 (N_17395,N_10013,N_12902);
nor U17396 (N_17396,N_14957,N_12570);
nor U17397 (N_17397,N_13671,N_11224);
xnor U17398 (N_17398,N_11502,N_11497);
nand U17399 (N_17399,N_14952,N_12173);
and U17400 (N_17400,N_13192,N_11757);
xnor U17401 (N_17401,N_11431,N_11616);
nand U17402 (N_17402,N_13540,N_12855);
nor U17403 (N_17403,N_14871,N_12153);
nand U17404 (N_17404,N_10014,N_11729);
nand U17405 (N_17405,N_12594,N_13032);
and U17406 (N_17406,N_14289,N_10621);
nor U17407 (N_17407,N_11325,N_14170);
nand U17408 (N_17408,N_13280,N_13444);
or U17409 (N_17409,N_11256,N_12266);
nand U17410 (N_17410,N_11480,N_10005);
and U17411 (N_17411,N_10128,N_10034);
or U17412 (N_17412,N_10860,N_10779);
and U17413 (N_17413,N_14704,N_11125);
xor U17414 (N_17414,N_12799,N_11064);
nor U17415 (N_17415,N_13318,N_14966);
and U17416 (N_17416,N_10555,N_12351);
nor U17417 (N_17417,N_14701,N_12296);
and U17418 (N_17418,N_14151,N_10976);
nand U17419 (N_17419,N_10875,N_14850);
nor U17420 (N_17420,N_10699,N_11817);
nand U17421 (N_17421,N_12786,N_10355);
nor U17422 (N_17422,N_14492,N_11690);
or U17423 (N_17423,N_12418,N_12047);
nor U17424 (N_17424,N_10864,N_10033);
and U17425 (N_17425,N_10575,N_11694);
and U17426 (N_17426,N_11318,N_12744);
xnor U17427 (N_17427,N_11378,N_13453);
and U17428 (N_17428,N_12313,N_11591);
or U17429 (N_17429,N_12929,N_11349);
nand U17430 (N_17430,N_11561,N_13826);
or U17431 (N_17431,N_14040,N_14324);
or U17432 (N_17432,N_11767,N_10776);
nor U17433 (N_17433,N_10839,N_12109);
nand U17434 (N_17434,N_12988,N_12217);
xor U17435 (N_17435,N_11532,N_13151);
nor U17436 (N_17436,N_11781,N_11630);
and U17437 (N_17437,N_12709,N_11225);
and U17438 (N_17438,N_14105,N_11391);
nand U17439 (N_17439,N_12956,N_14027);
or U17440 (N_17440,N_11671,N_14284);
or U17441 (N_17441,N_13196,N_11014);
nand U17442 (N_17442,N_14822,N_11149);
nand U17443 (N_17443,N_13941,N_12386);
and U17444 (N_17444,N_14109,N_12462);
and U17445 (N_17445,N_13423,N_10475);
xor U17446 (N_17446,N_14541,N_14112);
or U17447 (N_17447,N_14030,N_14432);
and U17448 (N_17448,N_10928,N_12917);
or U17449 (N_17449,N_10220,N_13829);
nand U17450 (N_17450,N_12590,N_10995);
and U17451 (N_17451,N_12968,N_11474);
or U17452 (N_17452,N_14570,N_11992);
nor U17453 (N_17453,N_14456,N_14335);
or U17454 (N_17454,N_12366,N_14137);
or U17455 (N_17455,N_12283,N_11148);
nand U17456 (N_17456,N_14762,N_12067);
nor U17457 (N_17457,N_13655,N_13253);
or U17458 (N_17458,N_10378,N_13953);
and U17459 (N_17459,N_13374,N_10681);
nand U17460 (N_17460,N_13436,N_13852);
nor U17461 (N_17461,N_10619,N_11114);
and U17462 (N_17462,N_14392,N_10844);
or U17463 (N_17463,N_12797,N_12409);
and U17464 (N_17464,N_14147,N_11111);
nor U17465 (N_17465,N_10978,N_14585);
or U17466 (N_17466,N_14673,N_10678);
and U17467 (N_17467,N_12708,N_11465);
and U17468 (N_17468,N_11072,N_11066);
nor U17469 (N_17469,N_11614,N_12716);
nand U17470 (N_17470,N_14985,N_11357);
or U17471 (N_17471,N_12534,N_13551);
and U17472 (N_17472,N_14785,N_13748);
or U17473 (N_17473,N_13338,N_13885);
nor U17474 (N_17474,N_11738,N_10548);
nand U17475 (N_17475,N_12891,N_12867);
nor U17476 (N_17476,N_13361,N_10380);
nor U17477 (N_17477,N_12881,N_10028);
nand U17478 (N_17478,N_11981,N_14136);
or U17479 (N_17479,N_11979,N_13016);
or U17480 (N_17480,N_11854,N_14162);
nor U17481 (N_17481,N_11946,N_10236);
or U17482 (N_17482,N_10140,N_14565);
xnor U17483 (N_17483,N_14011,N_14629);
or U17484 (N_17484,N_10163,N_14159);
nor U17485 (N_17485,N_12907,N_14313);
or U17486 (N_17486,N_13195,N_13663);
nor U17487 (N_17487,N_13316,N_10524);
nor U17488 (N_17488,N_10088,N_12202);
or U17489 (N_17489,N_10144,N_12637);
and U17490 (N_17490,N_12332,N_13259);
nor U17491 (N_17491,N_12640,N_14591);
or U17492 (N_17492,N_10306,N_10738);
nand U17493 (N_17493,N_11924,N_11417);
nor U17494 (N_17494,N_14124,N_10233);
or U17495 (N_17495,N_14210,N_12229);
xor U17496 (N_17496,N_14401,N_14418);
or U17497 (N_17497,N_14751,N_10152);
or U17498 (N_17498,N_11086,N_14720);
nor U17499 (N_17499,N_11590,N_10856);
and U17500 (N_17500,N_14561,N_12817);
xnor U17501 (N_17501,N_11830,N_11194);
nor U17502 (N_17502,N_11104,N_14268);
or U17503 (N_17503,N_12101,N_13153);
and U17504 (N_17504,N_11818,N_10532);
nor U17505 (N_17505,N_14768,N_10544);
xnor U17506 (N_17506,N_12956,N_13896);
nor U17507 (N_17507,N_11760,N_11575);
xor U17508 (N_17508,N_12015,N_12522);
and U17509 (N_17509,N_14158,N_13334);
or U17510 (N_17510,N_14761,N_13658);
xor U17511 (N_17511,N_13036,N_10311);
nor U17512 (N_17512,N_13387,N_10748);
and U17513 (N_17513,N_10471,N_13985);
nand U17514 (N_17514,N_12901,N_11026);
nand U17515 (N_17515,N_13359,N_13687);
or U17516 (N_17516,N_12545,N_11276);
nand U17517 (N_17517,N_14455,N_13719);
xor U17518 (N_17518,N_10279,N_11440);
nor U17519 (N_17519,N_11733,N_10581);
or U17520 (N_17520,N_10391,N_12490);
or U17521 (N_17521,N_14218,N_10192);
nand U17522 (N_17522,N_11454,N_14087);
or U17523 (N_17523,N_11964,N_11761);
nand U17524 (N_17524,N_13087,N_10477);
or U17525 (N_17525,N_14076,N_14531);
or U17526 (N_17526,N_12711,N_10349);
or U17527 (N_17527,N_13705,N_13156);
or U17528 (N_17528,N_11997,N_10466);
nand U17529 (N_17529,N_13555,N_12686);
or U17530 (N_17530,N_10108,N_14834);
nand U17531 (N_17531,N_14861,N_11359);
and U17532 (N_17532,N_11969,N_13726);
and U17533 (N_17533,N_11435,N_11125);
xor U17534 (N_17534,N_10106,N_13932);
and U17535 (N_17535,N_12295,N_10215);
nand U17536 (N_17536,N_13291,N_11895);
nand U17537 (N_17537,N_12874,N_10865);
nor U17538 (N_17538,N_11498,N_14693);
nor U17539 (N_17539,N_14594,N_13510);
nor U17540 (N_17540,N_14137,N_14988);
or U17541 (N_17541,N_14884,N_14469);
or U17542 (N_17542,N_12449,N_13439);
or U17543 (N_17543,N_13866,N_12145);
or U17544 (N_17544,N_12295,N_11914);
nand U17545 (N_17545,N_11480,N_14376);
nor U17546 (N_17546,N_11682,N_12999);
xor U17547 (N_17547,N_12951,N_10364);
xor U17548 (N_17548,N_14869,N_14374);
and U17549 (N_17549,N_13148,N_13890);
nand U17550 (N_17550,N_11071,N_14089);
and U17551 (N_17551,N_13705,N_12493);
nor U17552 (N_17552,N_10509,N_12054);
nor U17553 (N_17553,N_14130,N_10426);
nand U17554 (N_17554,N_11365,N_11018);
nor U17555 (N_17555,N_13034,N_12768);
nand U17556 (N_17556,N_11512,N_10256);
nand U17557 (N_17557,N_10911,N_10789);
and U17558 (N_17558,N_13981,N_14147);
or U17559 (N_17559,N_11573,N_12111);
and U17560 (N_17560,N_11688,N_12274);
or U17561 (N_17561,N_10673,N_14155);
nor U17562 (N_17562,N_12742,N_13831);
and U17563 (N_17563,N_11149,N_13404);
and U17564 (N_17564,N_12160,N_12910);
xnor U17565 (N_17565,N_12279,N_10570);
and U17566 (N_17566,N_11048,N_14704);
and U17567 (N_17567,N_10231,N_10301);
and U17568 (N_17568,N_10313,N_12164);
nand U17569 (N_17569,N_14554,N_10270);
nor U17570 (N_17570,N_11298,N_14619);
nand U17571 (N_17571,N_13029,N_13957);
or U17572 (N_17572,N_10508,N_12836);
nor U17573 (N_17573,N_11834,N_11815);
xor U17574 (N_17574,N_10223,N_14973);
or U17575 (N_17575,N_12717,N_10647);
and U17576 (N_17576,N_10715,N_12537);
nor U17577 (N_17577,N_11344,N_14712);
nor U17578 (N_17578,N_14425,N_10506);
and U17579 (N_17579,N_11209,N_11098);
nor U17580 (N_17580,N_13546,N_13002);
nand U17581 (N_17581,N_12801,N_10752);
nand U17582 (N_17582,N_13324,N_13464);
and U17583 (N_17583,N_14351,N_13008);
xor U17584 (N_17584,N_13948,N_12145);
nand U17585 (N_17585,N_10144,N_10782);
or U17586 (N_17586,N_13911,N_14682);
nand U17587 (N_17587,N_11605,N_14264);
xnor U17588 (N_17588,N_14735,N_10335);
nand U17589 (N_17589,N_14708,N_11997);
and U17590 (N_17590,N_12709,N_10819);
or U17591 (N_17591,N_11594,N_10522);
nand U17592 (N_17592,N_13778,N_14274);
nand U17593 (N_17593,N_13651,N_11854);
nand U17594 (N_17594,N_14204,N_10668);
or U17595 (N_17595,N_12733,N_14311);
and U17596 (N_17596,N_14451,N_14369);
and U17597 (N_17597,N_14147,N_10829);
or U17598 (N_17598,N_11388,N_13146);
and U17599 (N_17599,N_12498,N_12094);
or U17600 (N_17600,N_10674,N_10794);
and U17601 (N_17601,N_13370,N_13102);
or U17602 (N_17602,N_12454,N_11652);
nor U17603 (N_17603,N_12262,N_14912);
nor U17604 (N_17604,N_12331,N_12240);
xor U17605 (N_17605,N_12520,N_14330);
or U17606 (N_17606,N_13074,N_12521);
and U17607 (N_17607,N_14325,N_14375);
and U17608 (N_17608,N_12636,N_12566);
nand U17609 (N_17609,N_13835,N_12466);
or U17610 (N_17610,N_13102,N_14341);
or U17611 (N_17611,N_13770,N_14803);
and U17612 (N_17612,N_12124,N_11210);
nor U17613 (N_17613,N_13057,N_12611);
or U17614 (N_17614,N_13730,N_12686);
and U17615 (N_17615,N_12466,N_13574);
and U17616 (N_17616,N_11417,N_11867);
and U17617 (N_17617,N_12744,N_10204);
and U17618 (N_17618,N_14366,N_13664);
nand U17619 (N_17619,N_13027,N_14825);
xnor U17620 (N_17620,N_14000,N_10400);
and U17621 (N_17621,N_14957,N_12579);
xor U17622 (N_17622,N_12713,N_12246);
nand U17623 (N_17623,N_12771,N_13362);
nor U17624 (N_17624,N_10646,N_12250);
nor U17625 (N_17625,N_14559,N_13721);
and U17626 (N_17626,N_12547,N_13971);
nor U17627 (N_17627,N_11125,N_11463);
or U17628 (N_17628,N_12378,N_13681);
nor U17629 (N_17629,N_11694,N_13701);
or U17630 (N_17630,N_14388,N_13309);
nand U17631 (N_17631,N_13408,N_10246);
xnor U17632 (N_17632,N_14601,N_14899);
or U17633 (N_17633,N_13617,N_11810);
or U17634 (N_17634,N_11483,N_10823);
nor U17635 (N_17635,N_11335,N_13120);
xnor U17636 (N_17636,N_13440,N_13527);
nor U17637 (N_17637,N_12988,N_10859);
or U17638 (N_17638,N_12101,N_10721);
or U17639 (N_17639,N_10670,N_11466);
or U17640 (N_17640,N_14321,N_12234);
nand U17641 (N_17641,N_10936,N_11904);
nor U17642 (N_17642,N_14132,N_11819);
nor U17643 (N_17643,N_12482,N_13354);
nand U17644 (N_17644,N_11803,N_13585);
or U17645 (N_17645,N_10098,N_13641);
xor U17646 (N_17646,N_10579,N_14818);
and U17647 (N_17647,N_14319,N_11299);
nor U17648 (N_17648,N_12772,N_10328);
or U17649 (N_17649,N_14768,N_11438);
nand U17650 (N_17650,N_12450,N_10115);
or U17651 (N_17651,N_12572,N_11142);
and U17652 (N_17652,N_13779,N_11936);
and U17653 (N_17653,N_10158,N_11941);
and U17654 (N_17654,N_13449,N_12186);
nor U17655 (N_17655,N_14538,N_13838);
nor U17656 (N_17656,N_13352,N_13332);
or U17657 (N_17657,N_13498,N_14795);
or U17658 (N_17658,N_11258,N_14846);
or U17659 (N_17659,N_14640,N_10168);
or U17660 (N_17660,N_14014,N_10023);
nor U17661 (N_17661,N_10386,N_12407);
nand U17662 (N_17662,N_13626,N_11843);
and U17663 (N_17663,N_10229,N_14990);
and U17664 (N_17664,N_11393,N_10090);
or U17665 (N_17665,N_12473,N_14553);
nand U17666 (N_17666,N_11518,N_12521);
and U17667 (N_17667,N_14871,N_13516);
nand U17668 (N_17668,N_10308,N_10312);
or U17669 (N_17669,N_13468,N_12947);
and U17670 (N_17670,N_11912,N_14929);
and U17671 (N_17671,N_11639,N_13434);
nor U17672 (N_17672,N_13493,N_11647);
or U17673 (N_17673,N_13362,N_13137);
nand U17674 (N_17674,N_12519,N_12913);
xnor U17675 (N_17675,N_12412,N_13792);
nor U17676 (N_17676,N_12065,N_10312);
or U17677 (N_17677,N_11279,N_12582);
or U17678 (N_17678,N_13679,N_13605);
nor U17679 (N_17679,N_10658,N_14028);
nor U17680 (N_17680,N_12701,N_10694);
and U17681 (N_17681,N_11589,N_13827);
or U17682 (N_17682,N_10126,N_13119);
nand U17683 (N_17683,N_11797,N_13329);
nor U17684 (N_17684,N_13369,N_14941);
nand U17685 (N_17685,N_12831,N_14891);
nor U17686 (N_17686,N_13567,N_12310);
or U17687 (N_17687,N_10519,N_14387);
nand U17688 (N_17688,N_13396,N_10869);
or U17689 (N_17689,N_11016,N_11002);
nand U17690 (N_17690,N_12798,N_12713);
or U17691 (N_17691,N_11260,N_11988);
or U17692 (N_17692,N_13421,N_14542);
nand U17693 (N_17693,N_10888,N_10275);
or U17694 (N_17694,N_10310,N_12012);
and U17695 (N_17695,N_12851,N_14534);
nand U17696 (N_17696,N_11952,N_12388);
xor U17697 (N_17697,N_14192,N_11446);
nor U17698 (N_17698,N_10191,N_12478);
nand U17699 (N_17699,N_13399,N_12434);
nand U17700 (N_17700,N_12684,N_11381);
or U17701 (N_17701,N_11805,N_10433);
nand U17702 (N_17702,N_12178,N_14632);
or U17703 (N_17703,N_12096,N_14211);
nand U17704 (N_17704,N_14835,N_11415);
nand U17705 (N_17705,N_10693,N_14957);
and U17706 (N_17706,N_11210,N_12966);
nor U17707 (N_17707,N_13567,N_12047);
nor U17708 (N_17708,N_13988,N_13072);
or U17709 (N_17709,N_13742,N_13163);
and U17710 (N_17710,N_13662,N_13804);
nor U17711 (N_17711,N_10014,N_12245);
or U17712 (N_17712,N_11002,N_14261);
nor U17713 (N_17713,N_13977,N_11508);
xor U17714 (N_17714,N_12860,N_12664);
or U17715 (N_17715,N_13777,N_12622);
and U17716 (N_17716,N_12210,N_10085);
nor U17717 (N_17717,N_12483,N_13406);
nor U17718 (N_17718,N_13305,N_10568);
and U17719 (N_17719,N_12138,N_10537);
xor U17720 (N_17720,N_13510,N_11569);
and U17721 (N_17721,N_10495,N_11493);
and U17722 (N_17722,N_10363,N_14100);
nand U17723 (N_17723,N_11422,N_10203);
or U17724 (N_17724,N_10890,N_11334);
or U17725 (N_17725,N_14054,N_10350);
and U17726 (N_17726,N_12224,N_14993);
nor U17727 (N_17727,N_10027,N_11902);
nor U17728 (N_17728,N_12673,N_10493);
xnor U17729 (N_17729,N_11704,N_11579);
nand U17730 (N_17730,N_11700,N_14026);
nand U17731 (N_17731,N_12471,N_12848);
xor U17732 (N_17732,N_12602,N_11857);
or U17733 (N_17733,N_14049,N_14459);
xnor U17734 (N_17734,N_12441,N_12925);
nand U17735 (N_17735,N_14256,N_13340);
nand U17736 (N_17736,N_14131,N_11480);
nor U17737 (N_17737,N_12418,N_12862);
nand U17738 (N_17738,N_14321,N_14522);
and U17739 (N_17739,N_14938,N_10289);
nand U17740 (N_17740,N_10617,N_14754);
nor U17741 (N_17741,N_14776,N_13261);
nor U17742 (N_17742,N_13223,N_12692);
nand U17743 (N_17743,N_14894,N_14818);
nor U17744 (N_17744,N_13084,N_11891);
nor U17745 (N_17745,N_10793,N_12338);
nor U17746 (N_17746,N_14125,N_12533);
or U17747 (N_17747,N_12055,N_12308);
or U17748 (N_17748,N_13474,N_12445);
nor U17749 (N_17749,N_13348,N_13857);
or U17750 (N_17750,N_14256,N_14424);
xor U17751 (N_17751,N_12855,N_12589);
and U17752 (N_17752,N_14899,N_11634);
nand U17753 (N_17753,N_13043,N_11275);
nand U17754 (N_17754,N_11725,N_11477);
nand U17755 (N_17755,N_10713,N_11346);
nor U17756 (N_17756,N_13752,N_14962);
or U17757 (N_17757,N_14669,N_10193);
or U17758 (N_17758,N_10539,N_10134);
nand U17759 (N_17759,N_13109,N_13303);
and U17760 (N_17760,N_12604,N_13043);
nand U17761 (N_17761,N_14896,N_12114);
nand U17762 (N_17762,N_12523,N_14554);
nor U17763 (N_17763,N_12639,N_13048);
nand U17764 (N_17764,N_14311,N_10921);
nor U17765 (N_17765,N_12655,N_13366);
nor U17766 (N_17766,N_14584,N_10657);
nand U17767 (N_17767,N_11969,N_14562);
nor U17768 (N_17768,N_14618,N_10622);
or U17769 (N_17769,N_13560,N_14040);
and U17770 (N_17770,N_11265,N_10183);
and U17771 (N_17771,N_14182,N_11359);
nand U17772 (N_17772,N_14655,N_14582);
nand U17773 (N_17773,N_11464,N_12907);
nand U17774 (N_17774,N_11691,N_12930);
or U17775 (N_17775,N_12817,N_12406);
nor U17776 (N_17776,N_11434,N_13278);
or U17777 (N_17777,N_12989,N_13879);
and U17778 (N_17778,N_11743,N_14323);
nor U17779 (N_17779,N_13496,N_10392);
or U17780 (N_17780,N_11221,N_11551);
xnor U17781 (N_17781,N_10201,N_13985);
or U17782 (N_17782,N_11040,N_12377);
or U17783 (N_17783,N_10921,N_13400);
or U17784 (N_17784,N_11808,N_11138);
or U17785 (N_17785,N_10121,N_13358);
nor U17786 (N_17786,N_12217,N_14007);
nor U17787 (N_17787,N_13105,N_10650);
or U17788 (N_17788,N_13060,N_10187);
or U17789 (N_17789,N_14344,N_13375);
nor U17790 (N_17790,N_10724,N_13951);
nor U17791 (N_17791,N_12586,N_14097);
nand U17792 (N_17792,N_10868,N_12065);
nor U17793 (N_17793,N_11496,N_11515);
xnor U17794 (N_17794,N_12946,N_12493);
and U17795 (N_17795,N_12173,N_14236);
and U17796 (N_17796,N_12131,N_10206);
and U17797 (N_17797,N_13102,N_12075);
nand U17798 (N_17798,N_10227,N_12143);
xnor U17799 (N_17799,N_14645,N_14582);
or U17800 (N_17800,N_12049,N_13046);
nor U17801 (N_17801,N_10086,N_14438);
and U17802 (N_17802,N_14619,N_12973);
or U17803 (N_17803,N_12320,N_12139);
or U17804 (N_17804,N_12579,N_10219);
nor U17805 (N_17805,N_14997,N_13922);
nand U17806 (N_17806,N_14182,N_10329);
or U17807 (N_17807,N_13486,N_14226);
and U17808 (N_17808,N_10135,N_10356);
nand U17809 (N_17809,N_12397,N_13556);
and U17810 (N_17810,N_12915,N_13058);
nor U17811 (N_17811,N_13001,N_12309);
and U17812 (N_17812,N_12573,N_11467);
or U17813 (N_17813,N_11412,N_11123);
nand U17814 (N_17814,N_11879,N_14934);
nor U17815 (N_17815,N_11629,N_12065);
and U17816 (N_17816,N_11019,N_11917);
nand U17817 (N_17817,N_11279,N_14377);
nand U17818 (N_17818,N_14042,N_12661);
nand U17819 (N_17819,N_14108,N_13859);
and U17820 (N_17820,N_11979,N_13496);
or U17821 (N_17821,N_11398,N_11584);
xnor U17822 (N_17822,N_11397,N_10533);
or U17823 (N_17823,N_14018,N_13119);
or U17824 (N_17824,N_11421,N_11682);
nand U17825 (N_17825,N_11423,N_10421);
nor U17826 (N_17826,N_12265,N_14834);
xnor U17827 (N_17827,N_12614,N_10594);
nand U17828 (N_17828,N_14329,N_13575);
and U17829 (N_17829,N_12033,N_12522);
and U17830 (N_17830,N_12118,N_13260);
nor U17831 (N_17831,N_10673,N_12420);
or U17832 (N_17832,N_11007,N_12017);
nor U17833 (N_17833,N_11154,N_11788);
and U17834 (N_17834,N_12853,N_13446);
and U17835 (N_17835,N_10600,N_13932);
xor U17836 (N_17836,N_11160,N_10720);
or U17837 (N_17837,N_13835,N_13041);
nor U17838 (N_17838,N_11954,N_14108);
nand U17839 (N_17839,N_10961,N_11969);
or U17840 (N_17840,N_14181,N_14898);
or U17841 (N_17841,N_13084,N_14309);
and U17842 (N_17842,N_10019,N_11989);
nand U17843 (N_17843,N_13202,N_11553);
nand U17844 (N_17844,N_10783,N_11455);
xor U17845 (N_17845,N_10040,N_11151);
nor U17846 (N_17846,N_12254,N_10765);
or U17847 (N_17847,N_10618,N_12289);
nand U17848 (N_17848,N_13507,N_13679);
nor U17849 (N_17849,N_11549,N_10272);
and U17850 (N_17850,N_13431,N_14683);
or U17851 (N_17851,N_12956,N_10421);
nor U17852 (N_17852,N_11617,N_11715);
or U17853 (N_17853,N_12213,N_11575);
and U17854 (N_17854,N_10520,N_12846);
or U17855 (N_17855,N_14577,N_13731);
nand U17856 (N_17856,N_10394,N_11174);
nand U17857 (N_17857,N_13823,N_14555);
nand U17858 (N_17858,N_10183,N_11327);
nand U17859 (N_17859,N_10939,N_12404);
or U17860 (N_17860,N_14016,N_13937);
xnor U17861 (N_17861,N_11680,N_12728);
or U17862 (N_17862,N_12094,N_14042);
and U17863 (N_17863,N_10589,N_13453);
nor U17864 (N_17864,N_10084,N_12126);
nand U17865 (N_17865,N_12934,N_12416);
and U17866 (N_17866,N_11609,N_11674);
or U17867 (N_17867,N_12065,N_13934);
or U17868 (N_17868,N_13638,N_12575);
xor U17869 (N_17869,N_12766,N_13465);
and U17870 (N_17870,N_13215,N_12708);
or U17871 (N_17871,N_13881,N_12681);
nor U17872 (N_17872,N_12721,N_11819);
nand U17873 (N_17873,N_12263,N_14300);
nand U17874 (N_17874,N_10552,N_14828);
nand U17875 (N_17875,N_10829,N_14089);
nand U17876 (N_17876,N_13856,N_13957);
nand U17877 (N_17877,N_11343,N_12992);
or U17878 (N_17878,N_10759,N_10392);
nor U17879 (N_17879,N_13569,N_14834);
and U17880 (N_17880,N_14725,N_13223);
nor U17881 (N_17881,N_13489,N_11185);
or U17882 (N_17882,N_11407,N_11604);
and U17883 (N_17883,N_13453,N_12298);
nor U17884 (N_17884,N_12412,N_14417);
or U17885 (N_17885,N_13955,N_13119);
and U17886 (N_17886,N_14519,N_10398);
or U17887 (N_17887,N_10838,N_13024);
or U17888 (N_17888,N_11175,N_14830);
and U17889 (N_17889,N_11281,N_12474);
and U17890 (N_17890,N_11144,N_10216);
and U17891 (N_17891,N_14139,N_11365);
xor U17892 (N_17892,N_11776,N_10014);
or U17893 (N_17893,N_13845,N_14270);
nand U17894 (N_17894,N_11366,N_12658);
nand U17895 (N_17895,N_11894,N_10211);
or U17896 (N_17896,N_14043,N_13293);
nor U17897 (N_17897,N_14941,N_13801);
and U17898 (N_17898,N_11649,N_11206);
or U17899 (N_17899,N_11271,N_12001);
or U17900 (N_17900,N_13084,N_12321);
and U17901 (N_17901,N_13216,N_12081);
nor U17902 (N_17902,N_10510,N_10250);
and U17903 (N_17903,N_14840,N_11290);
and U17904 (N_17904,N_13874,N_14590);
nor U17905 (N_17905,N_10990,N_10600);
nand U17906 (N_17906,N_14750,N_11165);
nand U17907 (N_17907,N_10610,N_12099);
nor U17908 (N_17908,N_10869,N_14551);
and U17909 (N_17909,N_10236,N_10634);
and U17910 (N_17910,N_14547,N_12320);
xnor U17911 (N_17911,N_13986,N_14717);
or U17912 (N_17912,N_10887,N_14890);
and U17913 (N_17913,N_12378,N_13722);
or U17914 (N_17914,N_12466,N_10839);
xor U17915 (N_17915,N_13435,N_12704);
and U17916 (N_17916,N_14028,N_13867);
nor U17917 (N_17917,N_11019,N_11344);
or U17918 (N_17918,N_14257,N_13251);
or U17919 (N_17919,N_10862,N_12290);
nor U17920 (N_17920,N_11447,N_13639);
nand U17921 (N_17921,N_11329,N_10070);
nand U17922 (N_17922,N_11369,N_13149);
and U17923 (N_17923,N_12597,N_11981);
nand U17924 (N_17924,N_14001,N_11908);
nor U17925 (N_17925,N_13244,N_14742);
or U17926 (N_17926,N_11123,N_12037);
nand U17927 (N_17927,N_10321,N_12115);
and U17928 (N_17928,N_10881,N_14686);
nor U17929 (N_17929,N_11441,N_10569);
xor U17930 (N_17930,N_12074,N_14392);
and U17931 (N_17931,N_11336,N_11229);
and U17932 (N_17932,N_14353,N_12241);
and U17933 (N_17933,N_13411,N_11005);
and U17934 (N_17934,N_12116,N_10036);
nor U17935 (N_17935,N_10137,N_11512);
nor U17936 (N_17936,N_10038,N_10328);
nand U17937 (N_17937,N_10321,N_10503);
and U17938 (N_17938,N_13481,N_11117);
nor U17939 (N_17939,N_14930,N_14873);
or U17940 (N_17940,N_10663,N_14942);
nand U17941 (N_17941,N_14515,N_12307);
or U17942 (N_17942,N_13853,N_12669);
nor U17943 (N_17943,N_14417,N_13399);
or U17944 (N_17944,N_12828,N_12898);
nor U17945 (N_17945,N_14700,N_11273);
xor U17946 (N_17946,N_12545,N_13779);
nand U17947 (N_17947,N_10818,N_14884);
or U17948 (N_17948,N_10189,N_11777);
nor U17949 (N_17949,N_13210,N_11153);
nand U17950 (N_17950,N_14767,N_13395);
nand U17951 (N_17951,N_12409,N_10574);
and U17952 (N_17952,N_12716,N_11067);
nor U17953 (N_17953,N_11702,N_10775);
nor U17954 (N_17954,N_10161,N_12191);
and U17955 (N_17955,N_10528,N_11973);
nand U17956 (N_17956,N_12144,N_13052);
and U17957 (N_17957,N_14722,N_11307);
nor U17958 (N_17958,N_10025,N_10742);
nor U17959 (N_17959,N_11035,N_11122);
xnor U17960 (N_17960,N_13658,N_14143);
or U17961 (N_17961,N_13813,N_12319);
nor U17962 (N_17962,N_14698,N_10984);
nand U17963 (N_17963,N_10456,N_12999);
nor U17964 (N_17964,N_14155,N_13594);
nor U17965 (N_17965,N_10836,N_13622);
nor U17966 (N_17966,N_14025,N_11400);
nand U17967 (N_17967,N_14651,N_10560);
and U17968 (N_17968,N_10820,N_10104);
nor U17969 (N_17969,N_14007,N_11701);
nand U17970 (N_17970,N_12739,N_13953);
or U17971 (N_17971,N_10965,N_12196);
and U17972 (N_17972,N_14454,N_10375);
and U17973 (N_17973,N_14995,N_10207);
nor U17974 (N_17974,N_14526,N_10383);
nand U17975 (N_17975,N_13092,N_10807);
or U17976 (N_17976,N_11161,N_13875);
nand U17977 (N_17977,N_12224,N_14208);
nand U17978 (N_17978,N_12681,N_13860);
xor U17979 (N_17979,N_10746,N_10795);
nor U17980 (N_17980,N_11876,N_14640);
nand U17981 (N_17981,N_10074,N_10052);
or U17982 (N_17982,N_11306,N_12567);
xnor U17983 (N_17983,N_13113,N_13450);
or U17984 (N_17984,N_14713,N_12739);
or U17985 (N_17985,N_11774,N_12145);
nand U17986 (N_17986,N_13583,N_10879);
xor U17987 (N_17987,N_11705,N_12770);
nand U17988 (N_17988,N_10991,N_13528);
nor U17989 (N_17989,N_10609,N_11978);
or U17990 (N_17990,N_13417,N_14196);
nand U17991 (N_17991,N_14537,N_11198);
or U17992 (N_17992,N_10351,N_11084);
and U17993 (N_17993,N_13326,N_10682);
or U17994 (N_17994,N_14187,N_13777);
nand U17995 (N_17995,N_12034,N_12902);
nor U17996 (N_17996,N_11402,N_13332);
nor U17997 (N_17997,N_14592,N_10363);
xor U17998 (N_17998,N_12240,N_10486);
nor U17999 (N_17999,N_13733,N_14617);
xnor U18000 (N_18000,N_14699,N_12061);
and U18001 (N_18001,N_13347,N_13036);
nor U18002 (N_18002,N_11842,N_12516);
nor U18003 (N_18003,N_12514,N_11640);
and U18004 (N_18004,N_12906,N_13957);
nor U18005 (N_18005,N_14648,N_12607);
nor U18006 (N_18006,N_12780,N_13225);
nand U18007 (N_18007,N_10857,N_10037);
nor U18008 (N_18008,N_14529,N_10556);
nand U18009 (N_18009,N_13591,N_11560);
or U18010 (N_18010,N_12946,N_13398);
and U18011 (N_18011,N_11927,N_13590);
and U18012 (N_18012,N_12201,N_14145);
nor U18013 (N_18013,N_13242,N_13265);
nand U18014 (N_18014,N_14455,N_14242);
nor U18015 (N_18015,N_14291,N_10312);
and U18016 (N_18016,N_10686,N_13283);
nor U18017 (N_18017,N_14089,N_14123);
nand U18018 (N_18018,N_12321,N_12903);
and U18019 (N_18019,N_10542,N_11098);
xor U18020 (N_18020,N_11773,N_14152);
nor U18021 (N_18021,N_14704,N_12355);
nand U18022 (N_18022,N_13574,N_11340);
and U18023 (N_18023,N_11559,N_14929);
nor U18024 (N_18024,N_12343,N_13796);
or U18025 (N_18025,N_12702,N_14574);
or U18026 (N_18026,N_13293,N_13337);
nor U18027 (N_18027,N_12086,N_13944);
nor U18028 (N_18028,N_13797,N_12840);
and U18029 (N_18029,N_10171,N_13612);
nand U18030 (N_18030,N_13563,N_13208);
and U18031 (N_18031,N_12063,N_11713);
xor U18032 (N_18032,N_13129,N_12462);
or U18033 (N_18033,N_12797,N_11219);
nor U18034 (N_18034,N_11161,N_14780);
xnor U18035 (N_18035,N_13232,N_14008);
nand U18036 (N_18036,N_11362,N_11796);
and U18037 (N_18037,N_13764,N_12805);
and U18038 (N_18038,N_13373,N_12681);
nor U18039 (N_18039,N_10488,N_12555);
nor U18040 (N_18040,N_12081,N_10242);
or U18041 (N_18041,N_14001,N_14941);
xor U18042 (N_18042,N_12295,N_12350);
nor U18043 (N_18043,N_11285,N_10270);
nand U18044 (N_18044,N_11149,N_10819);
nor U18045 (N_18045,N_11431,N_14114);
nor U18046 (N_18046,N_10120,N_12781);
and U18047 (N_18047,N_14090,N_11468);
nand U18048 (N_18048,N_10680,N_11932);
and U18049 (N_18049,N_13048,N_10908);
and U18050 (N_18050,N_10886,N_10206);
nor U18051 (N_18051,N_13382,N_11207);
nor U18052 (N_18052,N_10055,N_12460);
or U18053 (N_18053,N_13843,N_12069);
and U18054 (N_18054,N_13883,N_11843);
nor U18055 (N_18055,N_10982,N_14153);
nand U18056 (N_18056,N_14485,N_11240);
or U18057 (N_18057,N_13454,N_11134);
nand U18058 (N_18058,N_14092,N_11691);
or U18059 (N_18059,N_14409,N_13305);
nor U18060 (N_18060,N_11142,N_11995);
nand U18061 (N_18061,N_10151,N_11907);
and U18062 (N_18062,N_11605,N_13874);
and U18063 (N_18063,N_11038,N_11372);
or U18064 (N_18064,N_10526,N_11274);
or U18065 (N_18065,N_10801,N_13925);
nor U18066 (N_18066,N_13339,N_13420);
and U18067 (N_18067,N_13876,N_11584);
and U18068 (N_18068,N_12697,N_14941);
xor U18069 (N_18069,N_11380,N_12003);
or U18070 (N_18070,N_14164,N_13504);
and U18071 (N_18071,N_13449,N_13531);
nor U18072 (N_18072,N_12886,N_11671);
and U18073 (N_18073,N_11531,N_12555);
xnor U18074 (N_18074,N_11935,N_12434);
nor U18075 (N_18075,N_10649,N_11066);
or U18076 (N_18076,N_13731,N_10156);
nand U18077 (N_18077,N_10125,N_11118);
xor U18078 (N_18078,N_12379,N_11753);
or U18079 (N_18079,N_11322,N_13947);
or U18080 (N_18080,N_11573,N_14075);
and U18081 (N_18081,N_10216,N_11160);
nor U18082 (N_18082,N_13689,N_10868);
nor U18083 (N_18083,N_14863,N_12901);
xor U18084 (N_18084,N_14947,N_10061);
and U18085 (N_18085,N_14525,N_14071);
nor U18086 (N_18086,N_12005,N_10001);
nand U18087 (N_18087,N_10079,N_13789);
nand U18088 (N_18088,N_10591,N_14460);
nor U18089 (N_18089,N_14574,N_14368);
and U18090 (N_18090,N_10391,N_12211);
and U18091 (N_18091,N_11325,N_11600);
nand U18092 (N_18092,N_11512,N_13299);
nand U18093 (N_18093,N_13656,N_12859);
nor U18094 (N_18094,N_14440,N_13689);
and U18095 (N_18095,N_10522,N_12251);
nor U18096 (N_18096,N_13882,N_12488);
or U18097 (N_18097,N_13666,N_12101);
or U18098 (N_18098,N_11380,N_12854);
nand U18099 (N_18099,N_11960,N_13468);
nor U18100 (N_18100,N_11366,N_12736);
or U18101 (N_18101,N_12618,N_11796);
or U18102 (N_18102,N_10388,N_12874);
xor U18103 (N_18103,N_11695,N_10571);
nand U18104 (N_18104,N_10027,N_11208);
xnor U18105 (N_18105,N_13479,N_12792);
nand U18106 (N_18106,N_12488,N_11238);
nand U18107 (N_18107,N_14546,N_11785);
and U18108 (N_18108,N_14756,N_13790);
or U18109 (N_18109,N_14682,N_14811);
nor U18110 (N_18110,N_12434,N_12476);
and U18111 (N_18111,N_10801,N_12777);
nor U18112 (N_18112,N_11686,N_14980);
nand U18113 (N_18113,N_11699,N_10541);
or U18114 (N_18114,N_11920,N_12111);
nor U18115 (N_18115,N_10436,N_11720);
and U18116 (N_18116,N_12265,N_10066);
or U18117 (N_18117,N_11909,N_10234);
nor U18118 (N_18118,N_10735,N_10143);
and U18119 (N_18119,N_11619,N_13630);
nor U18120 (N_18120,N_14720,N_12837);
and U18121 (N_18121,N_12333,N_13077);
or U18122 (N_18122,N_14403,N_14112);
nand U18123 (N_18123,N_11757,N_13583);
nor U18124 (N_18124,N_10666,N_12826);
or U18125 (N_18125,N_13271,N_10489);
xnor U18126 (N_18126,N_10077,N_13939);
and U18127 (N_18127,N_12366,N_12293);
nand U18128 (N_18128,N_12266,N_11091);
and U18129 (N_18129,N_14147,N_11959);
or U18130 (N_18130,N_10988,N_12150);
and U18131 (N_18131,N_13565,N_11889);
and U18132 (N_18132,N_14038,N_14880);
or U18133 (N_18133,N_14356,N_10281);
or U18134 (N_18134,N_13120,N_10245);
and U18135 (N_18135,N_10587,N_12771);
or U18136 (N_18136,N_14480,N_10069);
nor U18137 (N_18137,N_12671,N_13673);
nand U18138 (N_18138,N_13341,N_10386);
and U18139 (N_18139,N_14295,N_11571);
and U18140 (N_18140,N_12339,N_12863);
nor U18141 (N_18141,N_11222,N_13456);
and U18142 (N_18142,N_14342,N_13395);
nand U18143 (N_18143,N_13547,N_14681);
xor U18144 (N_18144,N_14307,N_13314);
or U18145 (N_18145,N_11797,N_14205);
xor U18146 (N_18146,N_12654,N_12418);
or U18147 (N_18147,N_14310,N_11555);
nor U18148 (N_18148,N_11492,N_14955);
xnor U18149 (N_18149,N_10959,N_14240);
or U18150 (N_18150,N_10945,N_11469);
and U18151 (N_18151,N_13406,N_11364);
or U18152 (N_18152,N_11559,N_14992);
or U18153 (N_18153,N_10600,N_11440);
nor U18154 (N_18154,N_13838,N_10883);
or U18155 (N_18155,N_12363,N_14312);
nor U18156 (N_18156,N_13210,N_13198);
nand U18157 (N_18157,N_13530,N_14031);
and U18158 (N_18158,N_12911,N_13081);
nand U18159 (N_18159,N_10233,N_13335);
and U18160 (N_18160,N_13427,N_12802);
nand U18161 (N_18161,N_13355,N_10415);
nor U18162 (N_18162,N_13877,N_12294);
nor U18163 (N_18163,N_14500,N_10736);
or U18164 (N_18164,N_12760,N_12589);
nand U18165 (N_18165,N_13917,N_13306);
nor U18166 (N_18166,N_14268,N_13086);
or U18167 (N_18167,N_12215,N_13539);
xor U18168 (N_18168,N_14880,N_10660);
and U18169 (N_18169,N_11359,N_12687);
nand U18170 (N_18170,N_14295,N_10629);
nor U18171 (N_18171,N_11487,N_10979);
nor U18172 (N_18172,N_11866,N_13545);
nor U18173 (N_18173,N_10889,N_11600);
and U18174 (N_18174,N_13356,N_11663);
and U18175 (N_18175,N_13745,N_13139);
or U18176 (N_18176,N_14871,N_14151);
xnor U18177 (N_18177,N_14649,N_11779);
or U18178 (N_18178,N_13819,N_14463);
nand U18179 (N_18179,N_11214,N_13677);
nand U18180 (N_18180,N_11661,N_12006);
or U18181 (N_18181,N_13531,N_13111);
nor U18182 (N_18182,N_14231,N_14153);
xnor U18183 (N_18183,N_13071,N_12853);
nor U18184 (N_18184,N_13848,N_11925);
nor U18185 (N_18185,N_14141,N_12607);
or U18186 (N_18186,N_14829,N_12217);
nand U18187 (N_18187,N_14668,N_13829);
or U18188 (N_18188,N_13926,N_12967);
or U18189 (N_18189,N_11855,N_11422);
and U18190 (N_18190,N_10456,N_11943);
nand U18191 (N_18191,N_11653,N_14925);
nor U18192 (N_18192,N_13477,N_12220);
nand U18193 (N_18193,N_13402,N_13094);
nor U18194 (N_18194,N_10560,N_10281);
nor U18195 (N_18195,N_14620,N_12486);
or U18196 (N_18196,N_10721,N_12189);
and U18197 (N_18197,N_12905,N_10208);
nand U18198 (N_18198,N_11244,N_13411);
nor U18199 (N_18199,N_10264,N_10696);
nand U18200 (N_18200,N_14699,N_10857);
nor U18201 (N_18201,N_14842,N_10342);
nand U18202 (N_18202,N_12534,N_12019);
nand U18203 (N_18203,N_11771,N_12334);
nor U18204 (N_18204,N_10126,N_14573);
or U18205 (N_18205,N_10969,N_14330);
and U18206 (N_18206,N_12604,N_11218);
xor U18207 (N_18207,N_10937,N_12819);
or U18208 (N_18208,N_12067,N_13835);
nand U18209 (N_18209,N_11717,N_10826);
xnor U18210 (N_18210,N_14598,N_12940);
nand U18211 (N_18211,N_13011,N_14401);
nand U18212 (N_18212,N_12402,N_13850);
or U18213 (N_18213,N_13710,N_12218);
and U18214 (N_18214,N_10532,N_12079);
or U18215 (N_18215,N_10849,N_11907);
nand U18216 (N_18216,N_12441,N_13421);
nand U18217 (N_18217,N_14632,N_14534);
and U18218 (N_18218,N_14031,N_12575);
nand U18219 (N_18219,N_11891,N_10059);
nor U18220 (N_18220,N_10442,N_13456);
nor U18221 (N_18221,N_11697,N_11203);
and U18222 (N_18222,N_12261,N_10526);
and U18223 (N_18223,N_12418,N_14970);
nand U18224 (N_18224,N_13088,N_11173);
or U18225 (N_18225,N_11246,N_11008);
nor U18226 (N_18226,N_12898,N_10973);
or U18227 (N_18227,N_11333,N_12688);
and U18228 (N_18228,N_12546,N_13135);
or U18229 (N_18229,N_14476,N_10699);
and U18230 (N_18230,N_11332,N_12862);
or U18231 (N_18231,N_14574,N_13437);
nand U18232 (N_18232,N_11716,N_14388);
nor U18233 (N_18233,N_14186,N_10897);
nand U18234 (N_18234,N_14775,N_14905);
or U18235 (N_18235,N_14752,N_11696);
or U18236 (N_18236,N_13422,N_10591);
xor U18237 (N_18237,N_14710,N_11996);
nor U18238 (N_18238,N_10544,N_10504);
xnor U18239 (N_18239,N_10983,N_13145);
and U18240 (N_18240,N_11832,N_12728);
nor U18241 (N_18241,N_13353,N_10810);
nor U18242 (N_18242,N_11238,N_14627);
nand U18243 (N_18243,N_12044,N_13407);
xor U18244 (N_18244,N_11226,N_14005);
nand U18245 (N_18245,N_12050,N_12829);
and U18246 (N_18246,N_11918,N_12432);
nand U18247 (N_18247,N_10685,N_11108);
and U18248 (N_18248,N_10021,N_14721);
nand U18249 (N_18249,N_14774,N_11724);
and U18250 (N_18250,N_11080,N_11874);
or U18251 (N_18251,N_10006,N_12213);
nor U18252 (N_18252,N_14724,N_11379);
or U18253 (N_18253,N_14207,N_14705);
nand U18254 (N_18254,N_11678,N_12587);
and U18255 (N_18255,N_11530,N_10636);
or U18256 (N_18256,N_14601,N_11486);
nor U18257 (N_18257,N_10944,N_12678);
xnor U18258 (N_18258,N_13937,N_11358);
nand U18259 (N_18259,N_11001,N_14608);
or U18260 (N_18260,N_11323,N_13291);
and U18261 (N_18261,N_12823,N_12336);
nand U18262 (N_18262,N_10958,N_12481);
and U18263 (N_18263,N_10101,N_12350);
nand U18264 (N_18264,N_13062,N_12928);
nor U18265 (N_18265,N_11969,N_11784);
nand U18266 (N_18266,N_12135,N_14615);
nand U18267 (N_18267,N_14293,N_10419);
and U18268 (N_18268,N_14635,N_12477);
nand U18269 (N_18269,N_11652,N_12487);
nor U18270 (N_18270,N_14524,N_11358);
nand U18271 (N_18271,N_11456,N_10117);
and U18272 (N_18272,N_12991,N_12756);
or U18273 (N_18273,N_14185,N_13890);
or U18274 (N_18274,N_10717,N_10705);
nand U18275 (N_18275,N_14170,N_12455);
and U18276 (N_18276,N_14473,N_11479);
nand U18277 (N_18277,N_14337,N_13749);
xnor U18278 (N_18278,N_12842,N_12103);
and U18279 (N_18279,N_12388,N_13541);
or U18280 (N_18280,N_11856,N_12425);
nor U18281 (N_18281,N_14244,N_12352);
xnor U18282 (N_18282,N_12648,N_12193);
and U18283 (N_18283,N_12973,N_10256);
or U18284 (N_18284,N_11787,N_12854);
or U18285 (N_18285,N_13710,N_11011);
nor U18286 (N_18286,N_10684,N_10788);
nand U18287 (N_18287,N_14183,N_14735);
and U18288 (N_18288,N_10757,N_11508);
nand U18289 (N_18289,N_10751,N_10103);
nor U18290 (N_18290,N_13338,N_13186);
xor U18291 (N_18291,N_13497,N_14745);
nand U18292 (N_18292,N_11396,N_10213);
nand U18293 (N_18293,N_13651,N_14471);
nor U18294 (N_18294,N_10564,N_14994);
nand U18295 (N_18295,N_12568,N_13927);
nor U18296 (N_18296,N_12438,N_13746);
nor U18297 (N_18297,N_12842,N_13935);
or U18298 (N_18298,N_14784,N_10315);
and U18299 (N_18299,N_13718,N_11203);
nor U18300 (N_18300,N_11349,N_14001);
or U18301 (N_18301,N_12141,N_13664);
xor U18302 (N_18302,N_12634,N_14138);
nor U18303 (N_18303,N_13652,N_11593);
nand U18304 (N_18304,N_10330,N_14437);
nor U18305 (N_18305,N_12920,N_10180);
nand U18306 (N_18306,N_13130,N_13820);
nor U18307 (N_18307,N_12164,N_11377);
or U18308 (N_18308,N_13358,N_10806);
nand U18309 (N_18309,N_10876,N_10989);
nand U18310 (N_18310,N_13551,N_14488);
and U18311 (N_18311,N_10587,N_12238);
nor U18312 (N_18312,N_13689,N_12766);
nor U18313 (N_18313,N_11142,N_13557);
nand U18314 (N_18314,N_13881,N_10456);
nand U18315 (N_18315,N_12767,N_12234);
and U18316 (N_18316,N_14676,N_10717);
nor U18317 (N_18317,N_14037,N_13746);
nor U18318 (N_18318,N_10526,N_11121);
or U18319 (N_18319,N_11467,N_10015);
nor U18320 (N_18320,N_11293,N_11361);
nand U18321 (N_18321,N_11548,N_13208);
nor U18322 (N_18322,N_13340,N_13134);
nand U18323 (N_18323,N_12136,N_11741);
and U18324 (N_18324,N_12367,N_12401);
or U18325 (N_18325,N_11185,N_11900);
nand U18326 (N_18326,N_14078,N_12204);
nand U18327 (N_18327,N_14699,N_14290);
or U18328 (N_18328,N_10314,N_12057);
nor U18329 (N_18329,N_13693,N_12339);
xnor U18330 (N_18330,N_13342,N_10208);
nand U18331 (N_18331,N_13276,N_12907);
nand U18332 (N_18332,N_12996,N_11262);
or U18333 (N_18333,N_10212,N_10766);
or U18334 (N_18334,N_14174,N_11252);
xnor U18335 (N_18335,N_13282,N_14127);
nor U18336 (N_18336,N_12159,N_10260);
nor U18337 (N_18337,N_11049,N_11626);
nand U18338 (N_18338,N_13304,N_12317);
nand U18339 (N_18339,N_12881,N_11663);
nand U18340 (N_18340,N_14398,N_11165);
nor U18341 (N_18341,N_14269,N_10090);
nand U18342 (N_18342,N_11504,N_10639);
xnor U18343 (N_18343,N_11286,N_12220);
or U18344 (N_18344,N_12589,N_13002);
or U18345 (N_18345,N_10870,N_13016);
or U18346 (N_18346,N_13168,N_12406);
or U18347 (N_18347,N_14674,N_12240);
xnor U18348 (N_18348,N_10426,N_14966);
or U18349 (N_18349,N_13654,N_10413);
and U18350 (N_18350,N_14901,N_12660);
nand U18351 (N_18351,N_10421,N_13034);
xor U18352 (N_18352,N_12455,N_13035);
and U18353 (N_18353,N_11223,N_10328);
xor U18354 (N_18354,N_13085,N_10817);
nand U18355 (N_18355,N_10480,N_13853);
nor U18356 (N_18356,N_12869,N_11683);
and U18357 (N_18357,N_12234,N_12814);
nor U18358 (N_18358,N_10546,N_11398);
or U18359 (N_18359,N_14034,N_11112);
nand U18360 (N_18360,N_10759,N_14745);
nand U18361 (N_18361,N_11326,N_14974);
nand U18362 (N_18362,N_11115,N_10494);
and U18363 (N_18363,N_12341,N_10743);
nand U18364 (N_18364,N_14453,N_12085);
or U18365 (N_18365,N_12927,N_11978);
nor U18366 (N_18366,N_13905,N_13801);
or U18367 (N_18367,N_14687,N_11607);
and U18368 (N_18368,N_13746,N_12316);
nand U18369 (N_18369,N_10069,N_14682);
or U18370 (N_18370,N_12827,N_12668);
or U18371 (N_18371,N_14412,N_11909);
nand U18372 (N_18372,N_12631,N_13782);
and U18373 (N_18373,N_10275,N_11728);
or U18374 (N_18374,N_12701,N_13694);
nor U18375 (N_18375,N_10824,N_13386);
and U18376 (N_18376,N_10685,N_14817);
and U18377 (N_18377,N_11088,N_14519);
or U18378 (N_18378,N_14197,N_10780);
and U18379 (N_18379,N_12552,N_14101);
xnor U18380 (N_18380,N_13327,N_10623);
nand U18381 (N_18381,N_12050,N_10672);
and U18382 (N_18382,N_13842,N_11694);
and U18383 (N_18383,N_13253,N_11513);
xnor U18384 (N_18384,N_12369,N_11038);
or U18385 (N_18385,N_11653,N_12215);
or U18386 (N_18386,N_13307,N_12196);
and U18387 (N_18387,N_14383,N_14082);
xnor U18388 (N_18388,N_11867,N_13417);
or U18389 (N_18389,N_14372,N_10222);
or U18390 (N_18390,N_12867,N_14899);
xnor U18391 (N_18391,N_13722,N_12896);
and U18392 (N_18392,N_14656,N_14171);
and U18393 (N_18393,N_14953,N_10640);
and U18394 (N_18394,N_14175,N_10905);
nor U18395 (N_18395,N_10144,N_13326);
or U18396 (N_18396,N_13387,N_14807);
and U18397 (N_18397,N_10774,N_14882);
nor U18398 (N_18398,N_10597,N_11289);
nor U18399 (N_18399,N_11839,N_10770);
nand U18400 (N_18400,N_14144,N_14684);
nor U18401 (N_18401,N_14334,N_14214);
nand U18402 (N_18402,N_10860,N_13367);
nor U18403 (N_18403,N_12539,N_14993);
nand U18404 (N_18404,N_12686,N_10424);
or U18405 (N_18405,N_14496,N_11685);
and U18406 (N_18406,N_11214,N_13846);
and U18407 (N_18407,N_12048,N_14530);
nor U18408 (N_18408,N_10254,N_10370);
or U18409 (N_18409,N_13361,N_12177);
nor U18410 (N_18410,N_12465,N_13874);
and U18411 (N_18411,N_13939,N_10242);
nand U18412 (N_18412,N_10779,N_10809);
nor U18413 (N_18413,N_14848,N_14048);
nand U18414 (N_18414,N_12114,N_13010);
nor U18415 (N_18415,N_10974,N_13466);
nor U18416 (N_18416,N_13551,N_13133);
and U18417 (N_18417,N_14287,N_14965);
nand U18418 (N_18418,N_12086,N_13298);
and U18419 (N_18419,N_12695,N_14284);
and U18420 (N_18420,N_11765,N_14924);
nor U18421 (N_18421,N_11213,N_12078);
or U18422 (N_18422,N_11454,N_11873);
or U18423 (N_18423,N_12118,N_13972);
nand U18424 (N_18424,N_11699,N_10058);
and U18425 (N_18425,N_11765,N_12840);
or U18426 (N_18426,N_14871,N_12198);
nor U18427 (N_18427,N_14202,N_11774);
or U18428 (N_18428,N_10266,N_12546);
nand U18429 (N_18429,N_10672,N_12830);
or U18430 (N_18430,N_12641,N_12622);
nand U18431 (N_18431,N_14641,N_11323);
or U18432 (N_18432,N_14859,N_12991);
or U18433 (N_18433,N_13813,N_11375);
nand U18434 (N_18434,N_11894,N_10171);
and U18435 (N_18435,N_13183,N_11877);
or U18436 (N_18436,N_11189,N_13078);
xnor U18437 (N_18437,N_12005,N_11060);
or U18438 (N_18438,N_12878,N_10896);
and U18439 (N_18439,N_12371,N_14830);
or U18440 (N_18440,N_12696,N_14813);
and U18441 (N_18441,N_11421,N_14165);
and U18442 (N_18442,N_12006,N_11245);
or U18443 (N_18443,N_10310,N_11959);
and U18444 (N_18444,N_14987,N_12868);
nand U18445 (N_18445,N_10784,N_13627);
nand U18446 (N_18446,N_14343,N_10358);
nor U18447 (N_18447,N_10906,N_12982);
nor U18448 (N_18448,N_12519,N_14150);
nor U18449 (N_18449,N_11445,N_11068);
nor U18450 (N_18450,N_14692,N_13323);
or U18451 (N_18451,N_13124,N_12137);
and U18452 (N_18452,N_12339,N_14566);
or U18453 (N_18453,N_14172,N_11708);
or U18454 (N_18454,N_12938,N_11519);
and U18455 (N_18455,N_14977,N_13010);
or U18456 (N_18456,N_12391,N_14585);
and U18457 (N_18457,N_13884,N_11081);
nor U18458 (N_18458,N_12873,N_13856);
nor U18459 (N_18459,N_10850,N_12308);
nor U18460 (N_18460,N_13072,N_12020);
or U18461 (N_18461,N_13861,N_10312);
or U18462 (N_18462,N_13098,N_12578);
nor U18463 (N_18463,N_12876,N_11536);
or U18464 (N_18464,N_14055,N_14600);
and U18465 (N_18465,N_10556,N_11057);
or U18466 (N_18466,N_14610,N_14540);
nor U18467 (N_18467,N_10710,N_14173);
or U18468 (N_18468,N_11654,N_13648);
or U18469 (N_18469,N_13399,N_12952);
or U18470 (N_18470,N_11102,N_11451);
nor U18471 (N_18471,N_11995,N_12919);
xor U18472 (N_18472,N_10362,N_12383);
nor U18473 (N_18473,N_13584,N_11255);
nor U18474 (N_18474,N_10428,N_11843);
and U18475 (N_18475,N_11379,N_13687);
nand U18476 (N_18476,N_13353,N_14247);
nor U18477 (N_18477,N_14664,N_12446);
nor U18478 (N_18478,N_14300,N_12053);
nor U18479 (N_18479,N_10861,N_10565);
or U18480 (N_18480,N_12327,N_14498);
nand U18481 (N_18481,N_13744,N_10805);
nand U18482 (N_18482,N_13501,N_13491);
nand U18483 (N_18483,N_10884,N_14669);
nor U18484 (N_18484,N_12476,N_11435);
or U18485 (N_18485,N_13084,N_13177);
and U18486 (N_18486,N_13685,N_12275);
or U18487 (N_18487,N_12388,N_13564);
and U18488 (N_18488,N_11896,N_12264);
nand U18489 (N_18489,N_14568,N_11991);
nand U18490 (N_18490,N_12429,N_14745);
nor U18491 (N_18491,N_10918,N_12252);
nand U18492 (N_18492,N_12197,N_11591);
nand U18493 (N_18493,N_11475,N_10562);
nand U18494 (N_18494,N_11122,N_12227);
and U18495 (N_18495,N_11280,N_10422);
nor U18496 (N_18496,N_14430,N_11957);
xnor U18497 (N_18497,N_14291,N_11770);
or U18498 (N_18498,N_10872,N_14253);
nor U18499 (N_18499,N_13685,N_14502);
nor U18500 (N_18500,N_12546,N_12782);
nand U18501 (N_18501,N_14480,N_10515);
or U18502 (N_18502,N_14833,N_14257);
and U18503 (N_18503,N_11140,N_14838);
nand U18504 (N_18504,N_12102,N_14125);
or U18505 (N_18505,N_13407,N_11080);
xnor U18506 (N_18506,N_14422,N_11366);
and U18507 (N_18507,N_13576,N_14440);
and U18508 (N_18508,N_12463,N_14165);
nand U18509 (N_18509,N_10698,N_14503);
nand U18510 (N_18510,N_13924,N_11112);
and U18511 (N_18511,N_13393,N_10178);
nor U18512 (N_18512,N_12473,N_14583);
or U18513 (N_18513,N_10607,N_13896);
nor U18514 (N_18514,N_13374,N_14462);
or U18515 (N_18515,N_12653,N_11671);
or U18516 (N_18516,N_11583,N_14373);
nor U18517 (N_18517,N_11953,N_11361);
or U18518 (N_18518,N_13301,N_13720);
and U18519 (N_18519,N_14225,N_13586);
nand U18520 (N_18520,N_11300,N_12457);
and U18521 (N_18521,N_13385,N_13429);
nor U18522 (N_18522,N_13170,N_12476);
nor U18523 (N_18523,N_11101,N_10798);
and U18524 (N_18524,N_11755,N_12590);
nand U18525 (N_18525,N_10412,N_14018);
and U18526 (N_18526,N_12781,N_10328);
nor U18527 (N_18527,N_12780,N_14780);
xnor U18528 (N_18528,N_14931,N_12085);
nand U18529 (N_18529,N_10618,N_14398);
or U18530 (N_18530,N_12721,N_13830);
and U18531 (N_18531,N_11675,N_11021);
xnor U18532 (N_18532,N_13838,N_10585);
or U18533 (N_18533,N_13403,N_10799);
or U18534 (N_18534,N_14304,N_11079);
and U18535 (N_18535,N_13961,N_10069);
nor U18536 (N_18536,N_10197,N_10574);
and U18537 (N_18537,N_10439,N_14242);
and U18538 (N_18538,N_10150,N_14198);
nand U18539 (N_18539,N_12620,N_13488);
nor U18540 (N_18540,N_11686,N_11027);
and U18541 (N_18541,N_14898,N_14334);
nand U18542 (N_18542,N_11208,N_11155);
nand U18543 (N_18543,N_10191,N_11300);
nor U18544 (N_18544,N_13684,N_14017);
or U18545 (N_18545,N_13922,N_13319);
nor U18546 (N_18546,N_11319,N_11015);
and U18547 (N_18547,N_12530,N_14348);
nor U18548 (N_18548,N_12364,N_11675);
and U18549 (N_18549,N_11600,N_10700);
nand U18550 (N_18550,N_14301,N_11212);
and U18551 (N_18551,N_14568,N_14747);
or U18552 (N_18552,N_10845,N_14090);
nand U18553 (N_18553,N_10594,N_11816);
nor U18554 (N_18554,N_14535,N_11936);
and U18555 (N_18555,N_12124,N_10478);
nand U18556 (N_18556,N_10350,N_11408);
nor U18557 (N_18557,N_13611,N_10450);
or U18558 (N_18558,N_10436,N_10902);
nand U18559 (N_18559,N_12526,N_11865);
nor U18560 (N_18560,N_14390,N_12672);
and U18561 (N_18561,N_12131,N_12009);
nand U18562 (N_18562,N_14427,N_12099);
and U18563 (N_18563,N_14584,N_13866);
nand U18564 (N_18564,N_12899,N_12489);
and U18565 (N_18565,N_11317,N_10740);
and U18566 (N_18566,N_12440,N_13289);
and U18567 (N_18567,N_14484,N_12980);
or U18568 (N_18568,N_14260,N_10295);
xor U18569 (N_18569,N_14880,N_14795);
and U18570 (N_18570,N_10096,N_14043);
or U18571 (N_18571,N_10693,N_12168);
and U18572 (N_18572,N_13532,N_14058);
nor U18573 (N_18573,N_11274,N_12162);
or U18574 (N_18574,N_12176,N_14039);
nand U18575 (N_18575,N_10462,N_14614);
nor U18576 (N_18576,N_13767,N_10574);
and U18577 (N_18577,N_14233,N_14587);
or U18578 (N_18578,N_11308,N_10756);
xnor U18579 (N_18579,N_10904,N_14854);
nand U18580 (N_18580,N_11462,N_11991);
nand U18581 (N_18581,N_11610,N_10090);
and U18582 (N_18582,N_13000,N_12052);
and U18583 (N_18583,N_10496,N_10285);
nor U18584 (N_18584,N_11803,N_13287);
nor U18585 (N_18585,N_13038,N_12227);
and U18586 (N_18586,N_14805,N_11450);
nor U18587 (N_18587,N_10155,N_14496);
or U18588 (N_18588,N_14920,N_14150);
or U18589 (N_18589,N_11799,N_11331);
and U18590 (N_18590,N_13059,N_11218);
nand U18591 (N_18591,N_10681,N_11593);
nand U18592 (N_18592,N_14867,N_13107);
and U18593 (N_18593,N_10745,N_13993);
nand U18594 (N_18594,N_14007,N_11670);
xor U18595 (N_18595,N_13789,N_14564);
or U18596 (N_18596,N_14969,N_12305);
nor U18597 (N_18597,N_14317,N_11190);
xnor U18598 (N_18598,N_11716,N_12503);
nor U18599 (N_18599,N_13403,N_13569);
xor U18600 (N_18600,N_13204,N_12019);
nor U18601 (N_18601,N_14510,N_11248);
nor U18602 (N_18602,N_11656,N_14303);
nand U18603 (N_18603,N_14136,N_14656);
nand U18604 (N_18604,N_13246,N_10054);
nor U18605 (N_18605,N_12025,N_13402);
nor U18606 (N_18606,N_10612,N_14102);
or U18607 (N_18607,N_12099,N_14483);
and U18608 (N_18608,N_12065,N_14759);
nand U18609 (N_18609,N_14043,N_13853);
nor U18610 (N_18610,N_12066,N_13532);
nand U18611 (N_18611,N_12830,N_11158);
or U18612 (N_18612,N_10314,N_11809);
or U18613 (N_18613,N_13037,N_11060);
nand U18614 (N_18614,N_10287,N_11942);
and U18615 (N_18615,N_14771,N_13387);
nand U18616 (N_18616,N_10531,N_10512);
or U18617 (N_18617,N_13824,N_13254);
nand U18618 (N_18618,N_12250,N_11517);
and U18619 (N_18619,N_13561,N_12374);
or U18620 (N_18620,N_10824,N_14591);
nor U18621 (N_18621,N_10604,N_11127);
nor U18622 (N_18622,N_12488,N_11674);
nor U18623 (N_18623,N_14850,N_14001);
xor U18624 (N_18624,N_12637,N_13477);
or U18625 (N_18625,N_10964,N_11782);
nor U18626 (N_18626,N_10537,N_10650);
and U18627 (N_18627,N_12382,N_13482);
and U18628 (N_18628,N_11699,N_10116);
or U18629 (N_18629,N_12207,N_14538);
or U18630 (N_18630,N_10204,N_11907);
nand U18631 (N_18631,N_11632,N_12125);
or U18632 (N_18632,N_14918,N_11435);
and U18633 (N_18633,N_11945,N_14977);
nor U18634 (N_18634,N_12599,N_14076);
and U18635 (N_18635,N_11187,N_13695);
nor U18636 (N_18636,N_13846,N_12760);
nor U18637 (N_18637,N_11658,N_10966);
xor U18638 (N_18638,N_10140,N_14998);
nand U18639 (N_18639,N_12152,N_11470);
nor U18640 (N_18640,N_12713,N_13948);
nand U18641 (N_18641,N_14879,N_11100);
and U18642 (N_18642,N_14256,N_14114);
nor U18643 (N_18643,N_10029,N_14635);
and U18644 (N_18644,N_13525,N_12315);
or U18645 (N_18645,N_12789,N_10684);
xnor U18646 (N_18646,N_10340,N_11798);
or U18647 (N_18647,N_13089,N_14443);
nor U18648 (N_18648,N_14327,N_10367);
nand U18649 (N_18649,N_12259,N_12673);
or U18650 (N_18650,N_13913,N_14955);
nor U18651 (N_18651,N_14493,N_10940);
nor U18652 (N_18652,N_11380,N_12886);
nor U18653 (N_18653,N_10910,N_13556);
nor U18654 (N_18654,N_14184,N_12831);
and U18655 (N_18655,N_14162,N_12538);
or U18656 (N_18656,N_14122,N_14363);
nand U18657 (N_18657,N_12202,N_11252);
xnor U18658 (N_18658,N_12941,N_11386);
xor U18659 (N_18659,N_11164,N_14214);
nand U18660 (N_18660,N_14726,N_10562);
nor U18661 (N_18661,N_12364,N_12556);
or U18662 (N_18662,N_12322,N_10446);
nand U18663 (N_18663,N_13781,N_11442);
nand U18664 (N_18664,N_12210,N_13666);
nand U18665 (N_18665,N_13133,N_10858);
nor U18666 (N_18666,N_13353,N_12811);
or U18667 (N_18667,N_13571,N_11304);
and U18668 (N_18668,N_13920,N_14252);
or U18669 (N_18669,N_14037,N_12267);
or U18670 (N_18670,N_12411,N_12912);
nand U18671 (N_18671,N_13912,N_11835);
xnor U18672 (N_18672,N_13379,N_10286);
and U18673 (N_18673,N_12272,N_10077);
nor U18674 (N_18674,N_12753,N_14737);
and U18675 (N_18675,N_11425,N_10887);
or U18676 (N_18676,N_12163,N_13055);
nand U18677 (N_18677,N_10810,N_11509);
nand U18678 (N_18678,N_10825,N_12585);
nand U18679 (N_18679,N_14734,N_11222);
nand U18680 (N_18680,N_12857,N_13626);
nand U18681 (N_18681,N_13918,N_12060);
and U18682 (N_18682,N_12274,N_12365);
or U18683 (N_18683,N_14706,N_14531);
nand U18684 (N_18684,N_14472,N_10492);
nor U18685 (N_18685,N_12897,N_10073);
xor U18686 (N_18686,N_13917,N_11398);
xnor U18687 (N_18687,N_11860,N_14048);
or U18688 (N_18688,N_13803,N_14826);
or U18689 (N_18689,N_12852,N_10614);
nor U18690 (N_18690,N_10366,N_10327);
xor U18691 (N_18691,N_11126,N_14396);
xnor U18692 (N_18692,N_10232,N_13640);
xor U18693 (N_18693,N_12431,N_11548);
or U18694 (N_18694,N_10222,N_10314);
nand U18695 (N_18695,N_10410,N_14047);
nor U18696 (N_18696,N_11863,N_13449);
and U18697 (N_18697,N_11193,N_11790);
and U18698 (N_18698,N_13638,N_10958);
or U18699 (N_18699,N_10580,N_10667);
or U18700 (N_18700,N_13822,N_13195);
nor U18701 (N_18701,N_14666,N_13887);
and U18702 (N_18702,N_13582,N_10196);
nand U18703 (N_18703,N_13612,N_10025);
nor U18704 (N_18704,N_12695,N_11189);
nor U18705 (N_18705,N_10822,N_13725);
nor U18706 (N_18706,N_13797,N_12431);
and U18707 (N_18707,N_14185,N_13395);
xnor U18708 (N_18708,N_11555,N_14111);
and U18709 (N_18709,N_13020,N_14938);
and U18710 (N_18710,N_12962,N_12545);
nand U18711 (N_18711,N_11106,N_11206);
nand U18712 (N_18712,N_14880,N_11220);
nor U18713 (N_18713,N_11891,N_14336);
or U18714 (N_18714,N_10935,N_14473);
xnor U18715 (N_18715,N_11962,N_14424);
or U18716 (N_18716,N_13516,N_12661);
nand U18717 (N_18717,N_13849,N_13651);
and U18718 (N_18718,N_10005,N_12045);
and U18719 (N_18719,N_13047,N_12499);
and U18720 (N_18720,N_11032,N_10596);
and U18721 (N_18721,N_12867,N_12849);
or U18722 (N_18722,N_13668,N_11354);
nor U18723 (N_18723,N_10071,N_14739);
nand U18724 (N_18724,N_13753,N_14887);
xor U18725 (N_18725,N_12254,N_10213);
nor U18726 (N_18726,N_13418,N_12045);
nor U18727 (N_18727,N_14535,N_12717);
nor U18728 (N_18728,N_14677,N_10582);
nor U18729 (N_18729,N_13572,N_11686);
or U18730 (N_18730,N_13151,N_13903);
nand U18731 (N_18731,N_12640,N_12495);
nor U18732 (N_18732,N_12544,N_10174);
nand U18733 (N_18733,N_12688,N_13518);
xor U18734 (N_18734,N_10074,N_13664);
or U18735 (N_18735,N_11798,N_14887);
or U18736 (N_18736,N_14793,N_14615);
or U18737 (N_18737,N_13741,N_10176);
nor U18738 (N_18738,N_14660,N_13663);
nor U18739 (N_18739,N_11068,N_11630);
nor U18740 (N_18740,N_10960,N_12209);
or U18741 (N_18741,N_11634,N_13781);
and U18742 (N_18742,N_14098,N_11103);
nand U18743 (N_18743,N_12489,N_11703);
nor U18744 (N_18744,N_13895,N_14925);
and U18745 (N_18745,N_10862,N_12752);
nand U18746 (N_18746,N_11178,N_13582);
xnor U18747 (N_18747,N_10556,N_10996);
nor U18748 (N_18748,N_13011,N_10239);
xor U18749 (N_18749,N_14517,N_14775);
or U18750 (N_18750,N_12247,N_12988);
and U18751 (N_18751,N_10096,N_12416);
nor U18752 (N_18752,N_12207,N_11870);
nand U18753 (N_18753,N_14978,N_14567);
nor U18754 (N_18754,N_12525,N_13508);
or U18755 (N_18755,N_13171,N_11035);
nor U18756 (N_18756,N_13109,N_12778);
nor U18757 (N_18757,N_13929,N_11396);
xor U18758 (N_18758,N_14903,N_12338);
nor U18759 (N_18759,N_12225,N_14429);
xnor U18760 (N_18760,N_13342,N_12387);
nand U18761 (N_18761,N_12075,N_13921);
and U18762 (N_18762,N_13221,N_12329);
xor U18763 (N_18763,N_14465,N_14309);
xor U18764 (N_18764,N_11760,N_10494);
or U18765 (N_18765,N_10146,N_12118);
and U18766 (N_18766,N_12860,N_11852);
nor U18767 (N_18767,N_10685,N_11111);
nand U18768 (N_18768,N_10117,N_11562);
and U18769 (N_18769,N_13356,N_11474);
or U18770 (N_18770,N_11359,N_10691);
or U18771 (N_18771,N_12310,N_11354);
and U18772 (N_18772,N_13390,N_13863);
nor U18773 (N_18773,N_11685,N_10354);
or U18774 (N_18774,N_14632,N_12106);
xnor U18775 (N_18775,N_14077,N_13164);
nand U18776 (N_18776,N_11907,N_11324);
and U18777 (N_18777,N_14810,N_11443);
and U18778 (N_18778,N_14002,N_14878);
nor U18779 (N_18779,N_14835,N_11568);
nor U18780 (N_18780,N_12122,N_13394);
nor U18781 (N_18781,N_14342,N_10119);
nand U18782 (N_18782,N_11200,N_10775);
and U18783 (N_18783,N_11056,N_13004);
nand U18784 (N_18784,N_13484,N_10406);
or U18785 (N_18785,N_11454,N_11305);
nor U18786 (N_18786,N_13588,N_13643);
and U18787 (N_18787,N_10882,N_14626);
nor U18788 (N_18788,N_12110,N_13408);
nor U18789 (N_18789,N_10592,N_12196);
or U18790 (N_18790,N_10111,N_13428);
or U18791 (N_18791,N_10973,N_12516);
nor U18792 (N_18792,N_10203,N_11335);
nand U18793 (N_18793,N_10013,N_12873);
nor U18794 (N_18794,N_13524,N_10777);
nor U18795 (N_18795,N_12692,N_14340);
and U18796 (N_18796,N_13527,N_12252);
nand U18797 (N_18797,N_14756,N_12140);
nor U18798 (N_18798,N_13265,N_13114);
nor U18799 (N_18799,N_10506,N_14740);
and U18800 (N_18800,N_11735,N_14665);
nor U18801 (N_18801,N_14320,N_13955);
or U18802 (N_18802,N_12151,N_11535);
nand U18803 (N_18803,N_14118,N_12434);
nand U18804 (N_18804,N_10471,N_11864);
or U18805 (N_18805,N_12681,N_11239);
nand U18806 (N_18806,N_10105,N_11164);
or U18807 (N_18807,N_12779,N_11717);
nand U18808 (N_18808,N_14369,N_10031);
nor U18809 (N_18809,N_14497,N_13169);
nand U18810 (N_18810,N_14606,N_14196);
or U18811 (N_18811,N_10779,N_13268);
and U18812 (N_18812,N_11756,N_11731);
xnor U18813 (N_18813,N_11047,N_12825);
nor U18814 (N_18814,N_14686,N_12014);
xor U18815 (N_18815,N_12246,N_14052);
xor U18816 (N_18816,N_12999,N_12621);
nand U18817 (N_18817,N_11364,N_12322);
nand U18818 (N_18818,N_10628,N_14226);
nand U18819 (N_18819,N_11172,N_11425);
nand U18820 (N_18820,N_14348,N_11707);
and U18821 (N_18821,N_11543,N_13832);
xor U18822 (N_18822,N_12680,N_13226);
xor U18823 (N_18823,N_10711,N_14423);
xnor U18824 (N_18824,N_13700,N_10648);
nor U18825 (N_18825,N_12220,N_13699);
nand U18826 (N_18826,N_13078,N_11782);
or U18827 (N_18827,N_11662,N_11327);
nand U18828 (N_18828,N_10950,N_10295);
or U18829 (N_18829,N_11459,N_14823);
and U18830 (N_18830,N_14153,N_12647);
nand U18831 (N_18831,N_10288,N_12219);
xor U18832 (N_18832,N_11938,N_13387);
or U18833 (N_18833,N_14767,N_12398);
nor U18834 (N_18834,N_11953,N_10002);
and U18835 (N_18835,N_10382,N_14148);
or U18836 (N_18836,N_11115,N_14044);
nand U18837 (N_18837,N_14845,N_11208);
xor U18838 (N_18838,N_11516,N_12962);
or U18839 (N_18839,N_10232,N_14211);
or U18840 (N_18840,N_10333,N_10211);
nor U18841 (N_18841,N_11402,N_11990);
or U18842 (N_18842,N_11358,N_11518);
nor U18843 (N_18843,N_13383,N_10107);
nor U18844 (N_18844,N_11777,N_11431);
nor U18845 (N_18845,N_11793,N_12844);
nor U18846 (N_18846,N_12432,N_10798);
nor U18847 (N_18847,N_10841,N_11781);
nand U18848 (N_18848,N_10288,N_13750);
nor U18849 (N_18849,N_11982,N_12019);
or U18850 (N_18850,N_11013,N_13282);
or U18851 (N_18851,N_12641,N_13465);
and U18852 (N_18852,N_10564,N_14355);
nand U18853 (N_18853,N_13655,N_12028);
nand U18854 (N_18854,N_10902,N_10614);
and U18855 (N_18855,N_11527,N_14822);
and U18856 (N_18856,N_11400,N_14839);
or U18857 (N_18857,N_12782,N_10605);
nor U18858 (N_18858,N_14062,N_11393);
or U18859 (N_18859,N_14978,N_13328);
nor U18860 (N_18860,N_13553,N_14358);
xnor U18861 (N_18861,N_11286,N_14861);
nand U18862 (N_18862,N_14781,N_13237);
xnor U18863 (N_18863,N_11558,N_10130);
and U18864 (N_18864,N_14206,N_10374);
nor U18865 (N_18865,N_10913,N_10343);
or U18866 (N_18866,N_14578,N_11567);
and U18867 (N_18867,N_10107,N_11380);
nor U18868 (N_18868,N_12213,N_11060);
nand U18869 (N_18869,N_12158,N_14876);
nand U18870 (N_18870,N_13237,N_10231);
or U18871 (N_18871,N_12330,N_14248);
nand U18872 (N_18872,N_11796,N_13388);
and U18873 (N_18873,N_13916,N_11392);
nand U18874 (N_18874,N_12156,N_11412);
and U18875 (N_18875,N_13266,N_11052);
and U18876 (N_18876,N_12793,N_11677);
and U18877 (N_18877,N_12573,N_11750);
nand U18878 (N_18878,N_14568,N_11556);
nor U18879 (N_18879,N_12581,N_14414);
or U18880 (N_18880,N_11687,N_14705);
and U18881 (N_18881,N_12040,N_14941);
or U18882 (N_18882,N_10863,N_10298);
or U18883 (N_18883,N_14063,N_11692);
or U18884 (N_18884,N_11402,N_11603);
and U18885 (N_18885,N_10430,N_13738);
and U18886 (N_18886,N_13086,N_13807);
nor U18887 (N_18887,N_14627,N_12666);
xnor U18888 (N_18888,N_13855,N_10413);
nor U18889 (N_18889,N_12950,N_10769);
nand U18890 (N_18890,N_11910,N_10035);
and U18891 (N_18891,N_10558,N_10148);
nand U18892 (N_18892,N_11213,N_11056);
xor U18893 (N_18893,N_10173,N_11630);
or U18894 (N_18894,N_12578,N_11629);
and U18895 (N_18895,N_11474,N_14225);
nand U18896 (N_18896,N_12850,N_11106);
nand U18897 (N_18897,N_14292,N_12739);
nand U18898 (N_18898,N_11900,N_13949);
or U18899 (N_18899,N_12062,N_13947);
and U18900 (N_18900,N_10053,N_13029);
and U18901 (N_18901,N_14251,N_13507);
nor U18902 (N_18902,N_12222,N_10928);
and U18903 (N_18903,N_12117,N_12426);
nand U18904 (N_18904,N_10965,N_14453);
or U18905 (N_18905,N_12793,N_10016);
nand U18906 (N_18906,N_14796,N_13004);
nand U18907 (N_18907,N_11519,N_14148);
nor U18908 (N_18908,N_14501,N_12484);
nand U18909 (N_18909,N_14268,N_13912);
and U18910 (N_18910,N_10176,N_10631);
and U18911 (N_18911,N_11254,N_14550);
and U18912 (N_18912,N_13083,N_10595);
and U18913 (N_18913,N_12520,N_13477);
or U18914 (N_18914,N_12455,N_12557);
nor U18915 (N_18915,N_11950,N_10295);
or U18916 (N_18916,N_12124,N_12684);
or U18917 (N_18917,N_10418,N_12451);
nand U18918 (N_18918,N_14499,N_12278);
or U18919 (N_18919,N_13918,N_11094);
nor U18920 (N_18920,N_10645,N_10604);
or U18921 (N_18921,N_13904,N_13076);
or U18922 (N_18922,N_10693,N_11253);
nand U18923 (N_18923,N_11768,N_10844);
nand U18924 (N_18924,N_12340,N_11461);
or U18925 (N_18925,N_11119,N_11262);
nand U18926 (N_18926,N_11582,N_10178);
nor U18927 (N_18927,N_14450,N_14503);
xor U18928 (N_18928,N_14731,N_10843);
nor U18929 (N_18929,N_13572,N_13413);
xnor U18930 (N_18930,N_14541,N_10982);
nand U18931 (N_18931,N_12383,N_10897);
nand U18932 (N_18932,N_14773,N_14416);
nand U18933 (N_18933,N_10848,N_12585);
nand U18934 (N_18934,N_11052,N_10484);
xnor U18935 (N_18935,N_11416,N_12127);
or U18936 (N_18936,N_10305,N_10906);
and U18937 (N_18937,N_13703,N_11478);
or U18938 (N_18938,N_13678,N_10528);
nor U18939 (N_18939,N_10322,N_14633);
xnor U18940 (N_18940,N_11605,N_10437);
or U18941 (N_18941,N_10505,N_13984);
or U18942 (N_18942,N_10348,N_11781);
nand U18943 (N_18943,N_11936,N_11619);
or U18944 (N_18944,N_12115,N_13558);
or U18945 (N_18945,N_12173,N_14699);
nand U18946 (N_18946,N_14049,N_12593);
nor U18947 (N_18947,N_14517,N_12244);
or U18948 (N_18948,N_14803,N_14612);
nand U18949 (N_18949,N_14718,N_12013);
or U18950 (N_18950,N_14642,N_12479);
and U18951 (N_18951,N_14601,N_11617);
nor U18952 (N_18952,N_14460,N_13904);
nand U18953 (N_18953,N_11214,N_10406);
nor U18954 (N_18954,N_12408,N_11152);
nor U18955 (N_18955,N_11612,N_10528);
and U18956 (N_18956,N_14530,N_14195);
and U18957 (N_18957,N_14686,N_14516);
and U18958 (N_18958,N_10777,N_13768);
nand U18959 (N_18959,N_12630,N_10080);
nand U18960 (N_18960,N_12070,N_10379);
nor U18961 (N_18961,N_13353,N_10872);
or U18962 (N_18962,N_13968,N_14478);
or U18963 (N_18963,N_14571,N_11387);
or U18964 (N_18964,N_13078,N_11804);
nor U18965 (N_18965,N_12470,N_14610);
nand U18966 (N_18966,N_14012,N_10537);
xnor U18967 (N_18967,N_11383,N_10398);
or U18968 (N_18968,N_14800,N_13178);
or U18969 (N_18969,N_11307,N_11659);
and U18970 (N_18970,N_13412,N_14396);
nand U18971 (N_18971,N_11532,N_11778);
and U18972 (N_18972,N_12971,N_11437);
xor U18973 (N_18973,N_12802,N_11627);
and U18974 (N_18974,N_12700,N_13981);
nand U18975 (N_18975,N_11123,N_14184);
nor U18976 (N_18976,N_13580,N_14239);
nor U18977 (N_18977,N_14391,N_13371);
or U18978 (N_18978,N_10013,N_14125);
or U18979 (N_18979,N_11861,N_11548);
or U18980 (N_18980,N_10580,N_10905);
or U18981 (N_18981,N_14465,N_10432);
or U18982 (N_18982,N_10490,N_10567);
xnor U18983 (N_18983,N_10716,N_11547);
nand U18984 (N_18984,N_12536,N_13005);
or U18985 (N_18985,N_11876,N_14697);
xnor U18986 (N_18986,N_11479,N_14388);
nand U18987 (N_18987,N_14917,N_13577);
or U18988 (N_18988,N_14817,N_14902);
and U18989 (N_18989,N_13479,N_12960);
nand U18990 (N_18990,N_14630,N_13406);
nor U18991 (N_18991,N_12879,N_12628);
xor U18992 (N_18992,N_13011,N_14642);
and U18993 (N_18993,N_11563,N_10329);
nand U18994 (N_18994,N_13914,N_10863);
or U18995 (N_18995,N_12685,N_10544);
nand U18996 (N_18996,N_10086,N_10635);
nor U18997 (N_18997,N_13530,N_14868);
nor U18998 (N_18998,N_12744,N_11518);
nand U18999 (N_18999,N_10390,N_11470);
nor U19000 (N_19000,N_12725,N_12680);
or U19001 (N_19001,N_12577,N_10771);
nand U19002 (N_19002,N_11692,N_12476);
and U19003 (N_19003,N_14983,N_14288);
nor U19004 (N_19004,N_10351,N_10345);
or U19005 (N_19005,N_14899,N_12495);
xnor U19006 (N_19006,N_12883,N_11584);
and U19007 (N_19007,N_12870,N_14736);
nand U19008 (N_19008,N_12269,N_11559);
and U19009 (N_19009,N_14507,N_12093);
and U19010 (N_19010,N_14825,N_13291);
nor U19011 (N_19011,N_10871,N_11236);
and U19012 (N_19012,N_12590,N_14031);
and U19013 (N_19013,N_10160,N_10492);
or U19014 (N_19014,N_11667,N_11967);
or U19015 (N_19015,N_14425,N_12898);
nand U19016 (N_19016,N_12746,N_14596);
nand U19017 (N_19017,N_11923,N_12129);
xnor U19018 (N_19018,N_11204,N_11666);
nor U19019 (N_19019,N_14680,N_11536);
or U19020 (N_19020,N_10648,N_10179);
xor U19021 (N_19021,N_11792,N_12659);
nor U19022 (N_19022,N_11217,N_14045);
and U19023 (N_19023,N_12005,N_10484);
nand U19024 (N_19024,N_13691,N_10449);
nand U19025 (N_19025,N_14385,N_12987);
nand U19026 (N_19026,N_10859,N_13713);
or U19027 (N_19027,N_14142,N_10954);
nand U19028 (N_19028,N_12927,N_11110);
and U19029 (N_19029,N_11502,N_10562);
nand U19030 (N_19030,N_12097,N_14751);
and U19031 (N_19031,N_11161,N_10072);
or U19032 (N_19032,N_10081,N_10588);
nand U19033 (N_19033,N_11805,N_11813);
or U19034 (N_19034,N_11106,N_10815);
nor U19035 (N_19035,N_10391,N_12909);
or U19036 (N_19036,N_13433,N_10556);
nor U19037 (N_19037,N_11449,N_12412);
and U19038 (N_19038,N_11917,N_10634);
and U19039 (N_19039,N_11994,N_10513);
nand U19040 (N_19040,N_11049,N_13806);
nor U19041 (N_19041,N_12616,N_11550);
or U19042 (N_19042,N_10054,N_14921);
nor U19043 (N_19043,N_13293,N_10894);
or U19044 (N_19044,N_14256,N_14023);
or U19045 (N_19045,N_14373,N_12797);
and U19046 (N_19046,N_12069,N_12924);
nand U19047 (N_19047,N_10515,N_12087);
nand U19048 (N_19048,N_10671,N_14620);
nor U19049 (N_19049,N_10851,N_13000);
and U19050 (N_19050,N_10435,N_11834);
or U19051 (N_19051,N_10201,N_10466);
xnor U19052 (N_19052,N_12760,N_11324);
or U19053 (N_19053,N_12381,N_12176);
nor U19054 (N_19054,N_11174,N_13299);
or U19055 (N_19055,N_12932,N_10277);
and U19056 (N_19056,N_13256,N_14105);
nand U19057 (N_19057,N_14600,N_14160);
and U19058 (N_19058,N_14685,N_14711);
and U19059 (N_19059,N_14652,N_12925);
and U19060 (N_19060,N_11992,N_10830);
nor U19061 (N_19061,N_10954,N_10113);
or U19062 (N_19062,N_14152,N_14048);
nand U19063 (N_19063,N_13550,N_12514);
nand U19064 (N_19064,N_13643,N_12205);
nand U19065 (N_19065,N_14089,N_11910);
nor U19066 (N_19066,N_11773,N_11060);
and U19067 (N_19067,N_11030,N_13646);
xnor U19068 (N_19068,N_14342,N_14899);
or U19069 (N_19069,N_14256,N_11176);
and U19070 (N_19070,N_13263,N_12880);
or U19071 (N_19071,N_13409,N_14251);
and U19072 (N_19072,N_12977,N_13157);
and U19073 (N_19073,N_13628,N_11340);
nand U19074 (N_19074,N_12955,N_10768);
nor U19075 (N_19075,N_13943,N_14420);
nor U19076 (N_19076,N_12830,N_14496);
nand U19077 (N_19077,N_10506,N_10855);
and U19078 (N_19078,N_11605,N_14733);
nand U19079 (N_19079,N_10829,N_12336);
or U19080 (N_19080,N_14498,N_14056);
nand U19081 (N_19081,N_10515,N_13619);
nor U19082 (N_19082,N_10257,N_12013);
nor U19083 (N_19083,N_10456,N_13295);
nor U19084 (N_19084,N_12168,N_14467);
nor U19085 (N_19085,N_12710,N_12153);
or U19086 (N_19086,N_11824,N_11566);
nor U19087 (N_19087,N_12949,N_11016);
or U19088 (N_19088,N_13996,N_13789);
nand U19089 (N_19089,N_13331,N_13374);
or U19090 (N_19090,N_13217,N_10405);
and U19091 (N_19091,N_14566,N_11162);
xnor U19092 (N_19092,N_10814,N_12048);
xnor U19093 (N_19093,N_13591,N_14487);
xor U19094 (N_19094,N_13430,N_12058);
or U19095 (N_19095,N_10720,N_14425);
nand U19096 (N_19096,N_11582,N_11352);
and U19097 (N_19097,N_14601,N_10839);
or U19098 (N_19098,N_11478,N_10415);
and U19099 (N_19099,N_11611,N_11524);
nand U19100 (N_19100,N_11242,N_12385);
nor U19101 (N_19101,N_11349,N_14911);
nand U19102 (N_19102,N_14130,N_12851);
and U19103 (N_19103,N_10330,N_12741);
xor U19104 (N_19104,N_12380,N_13064);
and U19105 (N_19105,N_10124,N_10502);
xor U19106 (N_19106,N_14907,N_13576);
or U19107 (N_19107,N_11891,N_11469);
nor U19108 (N_19108,N_11413,N_13959);
or U19109 (N_19109,N_12350,N_10200);
and U19110 (N_19110,N_14260,N_11402);
and U19111 (N_19111,N_13078,N_13609);
xnor U19112 (N_19112,N_10253,N_13861);
or U19113 (N_19113,N_14055,N_14101);
and U19114 (N_19114,N_14139,N_11278);
xnor U19115 (N_19115,N_11206,N_13891);
or U19116 (N_19116,N_14557,N_10296);
and U19117 (N_19117,N_14090,N_12955);
or U19118 (N_19118,N_12227,N_11935);
nor U19119 (N_19119,N_13787,N_10680);
and U19120 (N_19120,N_10791,N_10676);
nand U19121 (N_19121,N_12279,N_10797);
xor U19122 (N_19122,N_12937,N_10380);
and U19123 (N_19123,N_13063,N_10309);
nand U19124 (N_19124,N_12441,N_13146);
nor U19125 (N_19125,N_14924,N_10607);
nor U19126 (N_19126,N_10979,N_12199);
nand U19127 (N_19127,N_11496,N_12074);
nand U19128 (N_19128,N_13053,N_11595);
nor U19129 (N_19129,N_13261,N_14782);
nand U19130 (N_19130,N_11384,N_13404);
nand U19131 (N_19131,N_11433,N_14336);
nor U19132 (N_19132,N_11710,N_14220);
nor U19133 (N_19133,N_14518,N_11552);
or U19134 (N_19134,N_11891,N_11585);
nor U19135 (N_19135,N_13765,N_11863);
xnor U19136 (N_19136,N_14341,N_12106);
nand U19137 (N_19137,N_11393,N_12718);
xor U19138 (N_19138,N_11702,N_12733);
nor U19139 (N_19139,N_14404,N_10359);
or U19140 (N_19140,N_11833,N_13790);
nor U19141 (N_19141,N_14502,N_14438);
or U19142 (N_19142,N_12704,N_11374);
nor U19143 (N_19143,N_11215,N_13870);
nand U19144 (N_19144,N_10694,N_12725);
nor U19145 (N_19145,N_11255,N_13051);
or U19146 (N_19146,N_13646,N_11828);
nand U19147 (N_19147,N_11737,N_10144);
nor U19148 (N_19148,N_12508,N_14753);
nor U19149 (N_19149,N_11826,N_12373);
and U19150 (N_19150,N_11904,N_11614);
and U19151 (N_19151,N_13562,N_10448);
and U19152 (N_19152,N_13936,N_12261);
or U19153 (N_19153,N_13299,N_14809);
or U19154 (N_19154,N_10787,N_14582);
nor U19155 (N_19155,N_10973,N_10630);
or U19156 (N_19156,N_12022,N_10039);
and U19157 (N_19157,N_11940,N_11034);
nor U19158 (N_19158,N_10614,N_10865);
nand U19159 (N_19159,N_11050,N_14397);
nor U19160 (N_19160,N_12269,N_12458);
or U19161 (N_19161,N_12133,N_10524);
nand U19162 (N_19162,N_14198,N_12608);
nor U19163 (N_19163,N_12536,N_12357);
and U19164 (N_19164,N_11174,N_12369);
and U19165 (N_19165,N_13462,N_10906);
and U19166 (N_19166,N_14148,N_14453);
nor U19167 (N_19167,N_14357,N_12592);
nor U19168 (N_19168,N_10162,N_13434);
nor U19169 (N_19169,N_10823,N_13859);
or U19170 (N_19170,N_10954,N_10114);
and U19171 (N_19171,N_10130,N_12091);
or U19172 (N_19172,N_11964,N_13285);
or U19173 (N_19173,N_12023,N_10557);
and U19174 (N_19174,N_13062,N_12897);
or U19175 (N_19175,N_11374,N_10458);
nand U19176 (N_19176,N_11903,N_11615);
nand U19177 (N_19177,N_14744,N_13472);
nor U19178 (N_19178,N_11624,N_12835);
and U19179 (N_19179,N_14496,N_12362);
xnor U19180 (N_19180,N_13308,N_13766);
xnor U19181 (N_19181,N_14615,N_14163);
and U19182 (N_19182,N_14108,N_10993);
nor U19183 (N_19183,N_11742,N_14813);
and U19184 (N_19184,N_13347,N_14473);
and U19185 (N_19185,N_13058,N_14212);
or U19186 (N_19186,N_12852,N_14240);
or U19187 (N_19187,N_13377,N_14940);
nor U19188 (N_19188,N_13900,N_10545);
or U19189 (N_19189,N_11271,N_10293);
nor U19190 (N_19190,N_11557,N_12650);
or U19191 (N_19191,N_13878,N_12673);
or U19192 (N_19192,N_11030,N_11991);
nor U19193 (N_19193,N_12307,N_11077);
and U19194 (N_19194,N_14540,N_12632);
and U19195 (N_19195,N_12908,N_11146);
nand U19196 (N_19196,N_10766,N_14340);
or U19197 (N_19197,N_10258,N_11504);
nand U19198 (N_19198,N_10117,N_13445);
xor U19199 (N_19199,N_14507,N_12098);
nand U19200 (N_19200,N_12328,N_12539);
nand U19201 (N_19201,N_10566,N_12667);
or U19202 (N_19202,N_12317,N_14011);
or U19203 (N_19203,N_14004,N_14790);
nor U19204 (N_19204,N_13623,N_10062);
and U19205 (N_19205,N_12655,N_12133);
and U19206 (N_19206,N_10871,N_11942);
and U19207 (N_19207,N_11834,N_13122);
xor U19208 (N_19208,N_14328,N_10996);
and U19209 (N_19209,N_12531,N_11167);
nand U19210 (N_19210,N_11675,N_11606);
or U19211 (N_19211,N_11190,N_12089);
nor U19212 (N_19212,N_14205,N_14533);
nor U19213 (N_19213,N_13848,N_13284);
or U19214 (N_19214,N_13648,N_14537);
and U19215 (N_19215,N_14501,N_12237);
and U19216 (N_19216,N_14714,N_13777);
or U19217 (N_19217,N_12767,N_12369);
xnor U19218 (N_19218,N_14260,N_14086);
or U19219 (N_19219,N_13052,N_14173);
or U19220 (N_19220,N_12770,N_13470);
and U19221 (N_19221,N_12806,N_13244);
nor U19222 (N_19222,N_10555,N_14481);
xor U19223 (N_19223,N_10525,N_13311);
nor U19224 (N_19224,N_12869,N_12572);
nand U19225 (N_19225,N_11601,N_11794);
or U19226 (N_19226,N_12778,N_14217);
or U19227 (N_19227,N_13048,N_10504);
xor U19228 (N_19228,N_13008,N_14937);
or U19229 (N_19229,N_10535,N_13771);
nor U19230 (N_19230,N_14072,N_11622);
and U19231 (N_19231,N_12122,N_10436);
xor U19232 (N_19232,N_12953,N_12376);
and U19233 (N_19233,N_12015,N_11279);
and U19234 (N_19234,N_13031,N_11335);
nand U19235 (N_19235,N_12456,N_13566);
or U19236 (N_19236,N_11085,N_14408);
and U19237 (N_19237,N_12862,N_10263);
nor U19238 (N_19238,N_14803,N_10898);
or U19239 (N_19239,N_14556,N_13246);
nor U19240 (N_19240,N_12916,N_11761);
nor U19241 (N_19241,N_12442,N_12497);
nand U19242 (N_19242,N_14888,N_13637);
nor U19243 (N_19243,N_12310,N_13337);
and U19244 (N_19244,N_13076,N_10817);
or U19245 (N_19245,N_10557,N_12066);
nand U19246 (N_19246,N_12438,N_10513);
nor U19247 (N_19247,N_11355,N_12034);
or U19248 (N_19248,N_13435,N_13703);
xor U19249 (N_19249,N_10677,N_12546);
nand U19250 (N_19250,N_14364,N_11181);
nand U19251 (N_19251,N_12207,N_10030);
xor U19252 (N_19252,N_12983,N_13531);
and U19253 (N_19253,N_13737,N_14831);
or U19254 (N_19254,N_13698,N_13273);
xnor U19255 (N_19255,N_14797,N_10200);
and U19256 (N_19256,N_11427,N_12655);
nor U19257 (N_19257,N_12015,N_13006);
nand U19258 (N_19258,N_11012,N_11785);
nor U19259 (N_19259,N_12729,N_11874);
nand U19260 (N_19260,N_13174,N_14377);
nand U19261 (N_19261,N_12070,N_10245);
nand U19262 (N_19262,N_14732,N_12243);
xor U19263 (N_19263,N_14358,N_11838);
nand U19264 (N_19264,N_14068,N_12371);
nand U19265 (N_19265,N_13831,N_14451);
nor U19266 (N_19266,N_12032,N_10247);
xnor U19267 (N_19267,N_12996,N_13852);
and U19268 (N_19268,N_12532,N_14977);
nor U19269 (N_19269,N_14910,N_12506);
or U19270 (N_19270,N_13998,N_12796);
or U19271 (N_19271,N_10958,N_13054);
or U19272 (N_19272,N_12027,N_10003);
and U19273 (N_19273,N_14678,N_10574);
or U19274 (N_19274,N_12325,N_11873);
nor U19275 (N_19275,N_14429,N_14103);
or U19276 (N_19276,N_14414,N_14045);
nor U19277 (N_19277,N_13953,N_10575);
nor U19278 (N_19278,N_14838,N_14153);
nand U19279 (N_19279,N_13448,N_11649);
nand U19280 (N_19280,N_12737,N_10495);
nand U19281 (N_19281,N_13229,N_11716);
xnor U19282 (N_19282,N_11959,N_11339);
xnor U19283 (N_19283,N_13822,N_14692);
and U19284 (N_19284,N_12455,N_13455);
or U19285 (N_19285,N_14136,N_10298);
and U19286 (N_19286,N_12510,N_11313);
nand U19287 (N_19287,N_12747,N_12631);
nor U19288 (N_19288,N_11499,N_14874);
or U19289 (N_19289,N_13339,N_12623);
xnor U19290 (N_19290,N_11426,N_14914);
nor U19291 (N_19291,N_12197,N_11976);
or U19292 (N_19292,N_10291,N_10167);
and U19293 (N_19293,N_14862,N_10109);
nor U19294 (N_19294,N_12520,N_13664);
and U19295 (N_19295,N_12575,N_14243);
or U19296 (N_19296,N_14561,N_11659);
and U19297 (N_19297,N_13109,N_11793);
nand U19298 (N_19298,N_12456,N_12611);
and U19299 (N_19299,N_12517,N_12100);
nor U19300 (N_19300,N_10240,N_12709);
xor U19301 (N_19301,N_13368,N_10248);
or U19302 (N_19302,N_10325,N_10961);
or U19303 (N_19303,N_12841,N_12574);
nand U19304 (N_19304,N_12954,N_13866);
nand U19305 (N_19305,N_11194,N_13646);
nand U19306 (N_19306,N_14116,N_10832);
and U19307 (N_19307,N_12864,N_14521);
nand U19308 (N_19308,N_12781,N_11652);
nor U19309 (N_19309,N_12388,N_14144);
or U19310 (N_19310,N_10535,N_12568);
xor U19311 (N_19311,N_11078,N_13157);
and U19312 (N_19312,N_11839,N_12854);
xnor U19313 (N_19313,N_13622,N_14719);
or U19314 (N_19314,N_12206,N_10420);
nand U19315 (N_19315,N_14987,N_13026);
xor U19316 (N_19316,N_12231,N_13249);
xor U19317 (N_19317,N_13396,N_12311);
nor U19318 (N_19318,N_10008,N_13721);
and U19319 (N_19319,N_14953,N_13494);
nor U19320 (N_19320,N_14326,N_13872);
nor U19321 (N_19321,N_11730,N_14389);
or U19322 (N_19322,N_13938,N_11180);
nand U19323 (N_19323,N_10895,N_14641);
nor U19324 (N_19324,N_14195,N_13392);
nand U19325 (N_19325,N_12855,N_13925);
and U19326 (N_19326,N_12045,N_12783);
nand U19327 (N_19327,N_10073,N_10984);
xnor U19328 (N_19328,N_14990,N_12150);
and U19329 (N_19329,N_14117,N_12228);
nor U19330 (N_19330,N_11522,N_12779);
nor U19331 (N_19331,N_11825,N_10027);
nor U19332 (N_19332,N_12100,N_11346);
or U19333 (N_19333,N_13715,N_10133);
nand U19334 (N_19334,N_14353,N_12606);
xor U19335 (N_19335,N_10764,N_14509);
and U19336 (N_19336,N_12989,N_13727);
and U19337 (N_19337,N_12135,N_12253);
or U19338 (N_19338,N_12452,N_11632);
xnor U19339 (N_19339,N_14944,N_12143);
and U19340 (N_19340,N_13038,N_10196);
and U19341 (N_19341,N_11355,N_14775);
xor U19342 (N_19342,N_11297,N_10081);
nand U19343 (N_19343,N_13074,N_11449);
nor U19344 (N_19344,N_10215,N_13728);
and U19345 (N_19345,N_14934,N_14247);
and U19346 (N_19346,N_11150,N_13256);
or U19347 (N_19347,N_12373,N_13979);
nand U19348 (N_19348,N_14666,N_12242);
and U19349 (N_19349,N_13867,N_11239);
xor U19350 (N_19350,N_13434,N_12826);
and U19351 (N_19351,N_12198,N_13257);
or U19352 (N_19352,N_11793,N_13588);
and U19353 (N_19353,N_10513,N_12928);
nor U19354 (N_19354,N_14350,N_11508);
xor U19355 (N_19355,N_10737,N_14029);
nor U19356 (N_19356,N_11228,N_10362);
xor U19357 (N_19357,N_10806,N_11323);
or U19358 (N_19358,N_14372,N_12648);
nor U19359 (N_19359,N_13000,N_11964);
xnor U19360 (N_19360,N_14601,N_13573);
or U19361 (N_19361,N_11421,N_11531);
nand U19362 (N_19362,N_13138,N_13912);
and U19363 (N_19363,N_14746,N_12736);
nand U19364 (N_19364,N_11297,N_11895);
nand U19365 (N_19365,N_13573,N_11259);
or U19366 (N_19366,N_12685,N_12462);
nand U19367 (N_19367,N_14769,N_10679);
nor U19368 (N_19368,N_13659,N_11441);
nor U19369 (N_19369,N_13864,N_12097);
and U19370 (N_19370,N_12387,N_11260);
and U19371 (N_19371,N_12181,N_14872);
and U19372 (N_19372,N_12819,N_11829);
or U19373 (N_19373,N_12694,N_13290);
nor U19374 (N_19374,N_13997,N_11095);
and U19375 (N_19375,N_10155,N_12739);
and U19376 (N_19376,N_10745,N_10656);
nor U19377 (N_19377,N_10167,N_10844);
nor U19378 (N_19378,N_11677,N_13618);
and U19379 (N_19379,N_13504,N_12708);
nor U19380 (N_19380,N_10544,N_13788);
nor U19381 (N_19381,N_10354,N_13706);
and U19382 (N_19382,N_10095,N_14246);
xnor U19383 (N_19383,N_14437,N_13031);
nand U19384 (N_19384,N_12421,N_10907);
nor U19385 (N_19385,N_11640,N_14979);
nor U19386 (N_19386,N_13727,N_13331);
nand U19387 (N_19387,N_13656,N_13827);
or U19388 (N_19388,N_12647,N_14082);
or U19389 (N_19389,N_10533,N_14333);
or U19390 (N_19390,N_13895,N_11292);
nor U19391 (N_19391,N_13563,N_10349);
and U19392 (N_19392,N_14483,N_14929);
and U19393 (N_19393,N_10154,N_11807);
and U19394 (N_19394,N_11767,N_14811);
or U19395 (N_19395,N_12174,N_12818);
and U19396 (N_19396,N_14436,N_12194);
and U19397 (N_19397,N_14575,N_14361);
nor U19398 (N_19398,N_10128,N_14594);
and U19399 (N_19399,N_13952,N_14805);
nor U19400 (N_19400,N_13351,N_13755);
nand U19401 (N_19401,N_10583,N_12780);
and U19402 (N_19402,N_14513,N_12304);
nand U19403 (N_19403,N_14705,N_11217);
and U19404 (N_19404,N_10273,N_13716);
or U19405 (N_19405,N_10280,N_14486);
or U19406 (N_19406,N_12833,N_13239);
nand U19407 (N_19407,N_12089,N_13640);
nor U19408 (N_19408,N_14478,N_12355);
or U19409 (N_19409,N_14705,N_11371);
nand U19410 (N_19410,N_14334,N_10909);
nor U19411 (N_19411,N_12977,N_14923);
nor U19412 (N_19412,N_11009,N_11499);
nand U19413 (N_19413,N_13424,N_13485);
xnor U19414 (N_19414,N_12815,N_12644);
nand U19415 (N_19415,N_14788,N_12287);
nor U19416 (N_19416,N_12826,N_13010);
nor U19417 (N_19417,N_14605,N_13851);
and U19418 (N_19418,N_13913,N_10238);
or U19419 (N_19419,N_10003,N_11476);
or U19420 (N_19420,N_14080,N_10145);
xor U19421 (N_19421,N_12541,N_14718);
nand U19422 (N_19422,N_10501,N_12090);
xor U19423 (N_19423,N_12588,N_14211);
or U19424 (N_19424,N_14188,N_14238);
xnor U19425 (N_19425,N_13678,N_14632);
or U19426 (N_19426,N_13079,N_11972);
nand U19427 (N_19427,N_12933,N_12544);
xnor U19428 (N_19428,N_14751,N_13885);
and U19429 (N_19429,N_11258,N_13080);
nor U19430 (N_19430,N_12616,N_12847);
or U19431 (N_19431,N_12625,N_11940);
nor U19432 (N_19432,N_12300,N_10000);
nand U19433 (N_19433,N_13470,N_10649);
nand U19434 (N_19434,N_13605,N_11218);
or U19435 (N_19435,N_10081,N_12099);
nor U19436 (N_19436,N_10406,N_10560);
and U19437 (N_19437,N_10553,N_14953);
nor U19438 (N_19438,N_14571,N_10472);
or U19439 (N_19439,N_12407,N_11449);
and U19440 (N_19440,N_14600,N_13100);
and U19441 (N_19441,N_14194,N_14266);
and U19442 (N_19442,N_14371,N_13040);
or U19443 (N_19443,N_14781,N_10058);
or U19444 (N_19444,N_14009,N_14212);
nand U19445 (N_19445,N_12784,N_14613);
nand U19446 (N_19446,N_11101,N_11961);
nor U19447 (N_19447,N_12144,N_13138);
and U19448 (N_19448,N_12062,N_10494);
and U19449 (N_19449,N_12029,N_12963);
xor U19450 (N_19450,N_12496,N_13343);
nor U19451 (N_19451,N_10374,N_14192);
nor U19452 (N_19452,N_14294,N_12859);
and U19453 (N_19453,N_14269,N_12648);
nor U19454 (N_19454,N_12593,N_11102);
nand U19455 (N_19455,N_12701,N_10196);
nor U19456 (N_19456,N_14951,N_10201);
nand U19457 (N_19457,N_11131,N_12683);
or U19458 (N_19458,N_14981,N_10840);
nand U19459 (N_19459,N_12832,N_12408);
or U19460 (N_19460,N_11534,N_13135);
nand U19461 (N_19461,N_14015,N_12959);
nand U19462 (N_19462,N_14043,N_10605);
and U19463 (N_19463,N_12549,N_12426);
nand U19464 (N_19464,N_14217,N_10106);
and U19465 (N_19465,N_10874,N_10656);
and U19466 (N_19466,N_13617,N_11714);
nand U19467 (N_19467,N_13222,N_14521);
or U19468 (N_19468,N_10810,N_12878);
nor U19469 (N_19469,N_12056,N_10226);
nor U19470 (N_19470,N_14583,N_10098);
nand U19471 (N_19471,N_13059,N_12463);
and U19472 (N_19472,N_13607,N_12130);
or U19473 (N_19473,N_10399,N_12663);
or U19474 (N_19474,N_12720,N_11421);
and U19475 (N_19475,N_12728,N_11809);
nand U19476 (N_19476,N_11958,N_14117);
or U19477 (N_19477,N_10392,N_14433);
and U19478 (N_19478,N_13271,N_10433);
or U19479 (N_19479,N_11031,N_14425);
or U19480 (N_19480,N_13928,N_10903);
or U19481 (N_19481,N_11907,N_13762);
nor U19482 (N_19482,N_14398,N_13413);
nor U19483 (N_19483,N_11296,N_13709);
nand U19484 (N_19484,N_13920,N_12738);
or U19485 (N_19485,N_10023,N_12285);
or U19486 (N_19486,N_12986,N_10622);
and U19487 (N_19487,N_11347,N_14264);
and U19488 (N_19488,N_10284,N_10804);
and U19489 (N_19489,N_11149,N_13233);
nor U19490 (N_19490,N_10743,N_11564);
nand U19491 (N_19491,N_14093,N_14055);
nand U19492 (N_19492,N_10150,N_14899);
nor U19493 (N_19493,N_12488,N_14956);
nand U19494 (N_19494,N_10750,N_12705);
nor U19495 (N_19495,N_13602,N_10030);
or U19496 (N_19496,N_10801,N_10586);
nand U19497 (N_19497,N_14202,N_12738);
nor U19498 (N_19498,N_11830,N_14884);
or U19499 (N_19499,N_13774,N_10221);
nor U19500 (N_19500,N_11782,N_11483);
and U19501 (N_19501,N_13340,N_12462);
or U19502 (N_19502,N_12450,N_12052);
and U19503 (N_19503,N_11626,N_10539);
nand U19504 (N_19504,N_13350,N_10664);
and U19505 (N_19505,N_14772,N_13468);
or U19506 (N_19506,N_11989,N_12863);
xnor U19507 (N_19507,N_14953,N_10360);
and U19508 (N_19508,N_14880,N_10546);
and U19509 (N_19509,N_13750,N_11215);
xor U19510 (N_19510,N_10836,N_10621);
and U19511 (N_19511,N_14607,N_11397);
xnor U19512 (N_19512,N_14078,N_12987);
nand U19513 (N_19513,N_11259,N_11820);
and U19514 (N_19514,N_13085,N_14637);
nor U19515 (N_19515,N_10065,N_10940);
xor U19516 (N_19516,N_13780,N_13078);
or U19517 (N_19517,N_11844,N_14490);
nand U19518 (N_19518,N_13216,N_11614);
nor U19519 (N_19519,N_13124,N_11696);
nand U19520 (N_19520,N_14473,N_12842);
or U19521 (N_19521,N_13297,N_13307);
nor U19522 (N_19522,N_12320,N_11940);
nor U19523 (N_19523,N_11002,N_13909);
nand U19524 (N_19524,N_10828,N_13870);
or U19525 (N_19525,N_14420,N_13030);
or U19526 (N_19526,N_10851,N_13660);
xnor U19527 (N_19527,N_10964,N_13793);
nor U19528 (N_19528,N_12927,N_12370);
nand U19529 (N_19529,N_11749,N_11492);
xnor U19530 (N_19530,N_14215,N_13898);
and U19531 (N_19531,N_10780,N_12922);
and U19532 (N_19532,N_10445,N_11529);
and U19533 (N_19533,N_10184,N_12509);
nand U19534 (N_19534,N_10733,N_11427);
nand U19535 (N_19535,N_14807,N_11758);
and U19536 (N_19536,N_11226,N_14342);
and U19537 (N_19537,N_11576,N_13373);
nor U19538 (N_19538,N_14646,N_14815);
and U19539 (N_19539,N_11188,N_12259);
nand U19540 (N_19540,N_14059,N_12110);
and U19541 (N_19541,N_10393,N_10698);
nand U19542 (N_19542,N_11599,N_12220);
and U19543 (N_19543,N_10187,N_10140);
nor U19544 (N_19544,N_14584,N_11240);
nor U19545 (N_19545,N_14821,N_11290);
or U19546 (N_19546,N_14974,N_14243);
xnor U19547 (N_19547,N_14657,N_12104);
nor U19548 (N_19548,N_11811,N_13649);
and U19549 (N_19549,N_11434,N_12430);
and U19550 (N_19550,N_14332,N_12909);
and U19551 (N_19551,N_10246,N_13592);
nor U19552 (N_19552,N_14089,N_10497);
and U19553 (N_19553,N_13933,N_14758);
nor U19554 (N_19554,N_11945,N_11303);
xnor U19555 (N_19555,N_10529,N_14333);
and U19556 (N_19556,N_10774,N_14508);
xnor U19557 (N_19557,N_11674,N_11587);
nand U19558 (N_19558,N_10215,N_14854);
and U19559 (N_19559,N_14559,N_10442);
nor U19560 (N_19560,N_14161,N_14106);
nor U19561 (N_19561,N_14954,N_11137);
nor U19562 (N_19562,N_13980,N_10857);
or U19563 (N_19563,N_12806,N_13457);
or U19564 (N_19564,N_12077,N_12563);
nand U19565 (N_19565,N_10427,N_10523);
nand U19566 (N_19566,N_13131,N_10080);
or U19567 (N_19567,N_12263,N_12768);
and U19568 (N_19568,N_11962,N_11506);
nand U19569 (N_19569,N_13358,N_11569);
nor U19570 (N_19570,N_14971,N_12873);
nand U19571 (N_19571,N_12952,N_14025);
nor U19572 (N_19572,N_10655,N_14680);
nor U19573 (N_19573,N_12594,N_11719);
or U19574 (N_19574,N_12281,N_12269);
and U19575 (N_19575,N_10509,N_11506);
xor U19576 (N_19576,N_14296,N_13377);
or U19577 (N_19577,N_10521,N_14096);
nor U19578 (N_19578,N_13806,N_12107);
nor U19579 (N_19579,N_10065,N_12908);
nand U19580 (N_19580,N_14543,N_11121);
or U19581 (N_19581,N_11986,N_12760);
or U19582 (N_19582,N_11342,N_10029);
and U19583 (N_19583,N_10209,N_14437);
nand U19584 (N_19584,N_11833,N_13438);
and U19585 (N_19585,N_13841,N_14270);
nand U19586 (N_19586,N_13514,N_10635);
and U19587 (N_19587,N_11732,N_14582);
or U19588 (N_19588,N_10416,N_10214);
or U19589 (N_19589,N_11075,N_12533);
nand U19590 (N_19590,N_11157,N_10929);
or U19591 (N_19591,N_12425,N_10591);
and U19592 (N_19592,N_14443,N_13821);
or U19593 (N_19593,N_10857,N_10756);
nand U19594 (N_19594,N_11614,N_12162);
and U19595 (N_19595,N_10761,N_12610);
and U19596 (N_19596,N_10196,N_14967);
nor U19597 (N_19597,N_10416,N_14190);
and U19598 (N_19598,N_11091,N_10905);
nor U19599 (N_19599,N_14986,N_11644);
xor U19600 (N_19600,N_14435,N_13413);
nor U19601 (N_19601,N_11323,N_10174);
nor U19602 (N_19602,N_13025,N_10038);
or U19603 (N_19603,N_10313,N_11426);
nand U19604 (N_19604,N_14345,N_14225);
nor U19605 (N_19605,N_10183,N_10640);
and U19606 (N_19606,N_14066,N_10882);
nand U19607 (N_19607,N_13941,N_14678);
and U19608 (N_19608,N_12406,N_13405);
nand U19609 (N_19609,N_14428,N_13925);
and U19610 (N_19610,N_12926,N_13744);
and U19611 (N_19611,N_10072,N_13681);
and U19612 (N_19612,N_13289,N_10548);
nand U19613 (N_19613,N_13348,N_12148);
and U19614 (N_19614,N_12843,N_14831);
or U19615 (N_19615,N_14953,N_10007);
or U19616 (N_19616,N_12779,N_10266);
nand U19617 (N_19617,N_11610,N_14401);
nor U19618 (N_19618,N_10188,N_13553);
and U19619 (N_19619,N_10207,N_14143);
nor U19620 (N_19620,N_10633,N_12248);
or U19621 (N_19621,N_12852,N_14349);
nor U19622 (N_19622,N_11486,N_12711);
nand U19623 (N_19623,N_14289,N_11873);
and U19624 (N_19624,N_11063,N_11872);
nand U19625 (N_19625,N_14379,N_14671);
nor U19626 (N_19626,N_10317,N_12589);
and U19627 (N_19627,N_13239,N_14595);
nor U19628 (N_19628,N_13306,N_12619);
nand U19629 (N_19629,N_13827,N_11581);
xor U19630 (N_19630,N_13345,N_11050);
nand U19631 (N_19631,N_13911,N_13138);
nand U19632 (N_19632,N_13100,N_13577);
nand U19633 (N_19633,N_14869,N_11892);
xnor U19634 (N_19634,N_12841,N_11581);
or U19635 (N_19635,N_10077,N_14028);
and U19636 (N_19636,N_10940,N_12937);
and U19637 (N_19637,N_13200,N_14364);
or U19638 (N_19638,N_13395,N_11049);
and U19639 (N_19639,N_10723,N_10021);
nor U19640 (N_19640,N_13147,N_12639);
xor U19641 (N_19641,N_13320,N_14131);
xnor U19642 (N_19642,N_11808,N_11616);
nor U19643 (N_19643,N_12201,N_10715);
xnor U19644 (N_19644,N_11816,N_11867);
nand U19645 (N_19645,N_12762,N_14035);
nand U19646 (N_19646,N_12782,N_14603);
nor U19647 (N_19647,N_11370,N_13595);
and U19648 (N_19648,N_12104,N_12548);
nand U19649 (N_19649,N_12118,N_10450);
or U19650 (N_19650,N_14891,N_11953);
or U19651 (N_19651,N_11104,N_12272);
xor U19652 (N_19652,N_13339,N_13034);
nor U19653 (N_19653,N_14553,N_11520);
nand U19654 (N_19654,N_10508,N_14419);
nand U19655 (N_19655,N_10674,N_13962);
and U19656 (N_19656,N_10359,N_10823);
and U19657 (N_19657,N_12724,N_11291);
nand U19658 (N_19658,N_14117,N_11232);
xnor U19659 (N_19659,N_10571,N_12385);
nand U19660 (N_19660,N_14995,N_10966);
or U19661 (N_19661,N_10519,N_14901);
nor U19662 (N_19662,N_11978,N_14988);
and U19663 (N_19663,N_11792,N_12292);
nand U19664 (N_19664,N_10870,N_14696);
or U19665 (N_19665,N_14078,N_14955);
and U19666 (N_19666,N_10010,N_10837);
or U19667 (N_19667,N_12613,N_12994);
nor U19668 (N_19668,N_12654,N_10478);
nor U19669 (N_19669,N_11989,N_14429);
or U19670 (N_19670,N_14647,N_12383);
nor U19671 (N_19671,N_11283,N_14862);
and U19672 (N_19672,N_11499,N_10109);
and U19673 (N_19673,N_11062,N_10925);
xnor U19674 (N_19674,N_12022,N_11985);
and U19675 (N_19675,N_11793,N_10178);
nand U19676 (N_19676,N_11345,N_14104);
or U19677 (N_19677,N_14904,N_11527);
and U19678 (N_19678,N_10905,N_10635);
nand U19679 (N_19679,N_10881,N_10054);
or U19680 (N_19680,N_11928,N_12744);
and U19681 (N_19681,N_11080,N_10272);
nand U19682 (N_19682,N_14804,N_13612);
or U19683 (N_19683,N_11975,N_14912);
and U19684 (N_19684,N_12520,N_10301);
or U19685 (N_19685,N_10206,N_10357);
or U19686 (N_19686,N_11048,N_11881);
or U19687 (N_19687,N_11806,N_11220);
or U19688 (N_19688,N_12011,N_12813);
or U19689 (N_19689,N_12471,N_14463);
or U19690 (N_19690,N_13689,N_10064);
nor U19691 (N_19691,N_11094,N_10273);
nor U19692 (N_19692,N_10274,N_13217);
nand U19693 (N_19693,N_14086,N_12265);
and U19694 (N_19694,N_11572,N_14365);
or U19695 (N_19695,N_12567,N_11181);
nor U19696 (N_19696,N_14130,N_13959);
and U19697 (N_19697,N_11974,N_11698);
nand U19698 (N_19698,N_10116,N_13813);
xor U19699 (N_19699,N_12358,N_14392);
or U19700 (N_19700,N_12186,N_14067);
or U19701 (N_19701,N_10828,N_10688);
or U19702 (N_19702,N_14879,N_10726);
nand U19703 (N_19703,N_14239,N_13464);
or U19704 (N_19704,N_14737,N_12122);
and U19705 (N_19705,N_13923,N_13258);
or U19706 (N_19706,N_13141,N_13680);
or U19707 (N_19707,N_11007,N_12969);
xnor U19708 (N_19708,N_12577,N_10573);
nand U19709 (N_19709,N_11721,N_10664);
and U19710 (N_19710,N_10500,N_11553);
nand U19711 (N_19711,N_13605,N_14849);
nand U19712 (N_19712,N_13567,N_10788);
or U19713 (N_19713,N_10499,N_14461);
and U19714 (N_19714,N_10386,N_12531);
or U19715 (N_19715,N_12821,N_10082);
and U19716 (N_19716,N_11650,N_12044);
and U19717 (N_19717,N_14672,N_14518);
nor U19718 (N_19718,N_10479,N_11190);
and U19719 (N_19719,N_14922,N_10785);
and U19720 (N_19720,N_10555,N_10376);
and U19721 (N_19721,N_12686,N_11474);
nand U19722 (N_19722,N_11989,N_13333);
or U19723 (N_19723,N_10031,N_14955);
nand U19724 (N_19724,N_13203,N_12002);
or U19725 (N_19725,N_10441,N_14022);
and U19726 (N_19726,N_10490,N_11927);
and U19727 (N_19727,N_13279,N_11868);
nor U19728 (N_19728,N_14578,N_13970);
nand U19729 (N_19729,N_11072,N_10167);
nand U19730 (N_19730,N_13197,N_12318);
nor U19731 (N_19731,N_11236,N_13665);
or U19732 (N_19732,N_10756,N_11347);
nand U19733 (N_19733,N_10612,N_11503);
or U19734 (N_19734,N_13925,N_12162);
and U19735 (N_19735,N_12326,N_12135);
nor U19736 (N_19736,N_14181,N_12544);
nor U19737 (N_19737,N_13468,N_11344);
nor U19738 (N_19738,N_12289,N_12126);
nand U19739 (N_19739,N_13820,N_11845);
nand U19740 (N_19740,N_11078,N_13609);
nor U19741 (N_19741,N_10404,N_12048);
nand U19742 (N_19742,N_10790,N_10488);
and U19743 (N_19743,N_12919,N_14367);
nor U19744 (N_19744,N_14395,N_11125);
nand U19745 (N_19745,N_12422,N_10013);
and U19746 (N_19746,N_12811,N_14601);
and U19747 (N_19747,N_13394,N_10197);
nand U19748 (N_19748,N_13132,N_13585);
nand U19749 (N_19749,N_14757,N_13580);
and U19750 (N_19750,N_10655,N_10815);
nor U19751 (N_19751,N_14805,N_14477);
or U19752 (N_19752,N_10660,N_14342);
nand U19753 (N_19753,N_14333,N_10915);
nor U19754 (N_19754,N_14781,N_13733);
or U19755 (N_19755,N_12251,N_11213);
and U19756 (N_19756,N_14000,N_11573);
or U19757 (N_19757,N_11839,N_13506);
nand U19758 (N_19758,N_11209,N_13606);
nand U19759 (N_19759,N_14449,N_13672);
and U19760 (N_19760,N_12871,N_12378);
nor U19761 (N_19761,N_13397,N_12067);
nand U19762 (N_19762,N_11333,N_13201);
nand U19763 (N_19763,N_11269,N_10708);
and U19764 (N_19764,N_11665,N_11155);
nand U19765 (N_19765,N_11037,N_13889);
or U19766 (N_19766,N_10746,N_13298);
nand U19767 (N_19767,N_14889,N_12952);
and U19768 (N_19768,N_14834,N_13919);
nor U19769 (N_19769,N_10723,N_13446);
or U19770 (N_19770,N_14593,N_11203);
nor U19771 (N_19771,N_11520,N_11454);
nand U19772 (N_19772,N_14442,N_12443);
nor U19773 (N_19773,N_11259,N_10946);
xor U19774 (N_19774,N_13545,N_12035);
or U19775 (N_19775,N_10397,N_14548);
nor U19776 (N_19776,N_12828,N_13341);
xor U19777 (N_19777,N_14041,N_10796);
nand U19778 (N_19778,N_13122,N_11527);
or U19779 (N_19779,N_13199,N_10179);
or U19780 (N_19780,N_11265,N_14115);
xnor U19781 (N_19781,N_10194,N_14895);
and U19782 (N_19782,N_12141,N_11763);
nand U19783 (N_19783,N_14654,N_14366);
nor U19784 (N_19784,N_12813,N_11290);
or U19785 (N_19785,N_14697,N_10714);
nand U19786 (N_19786,N_12686,N_12507);
or U19787 (N_19787,N_11234,N_12338);
nand U19788 (N_19788,N_13678,N_11459);
and U19789 (N_19789,N_14189,N_12659);
nor U19790 (N_19790,N_11802,N_11179);
xnor U19791 (N_19791,N_10709,N_11876);
nor U19792 (N_19792,N_14890,N_14523);
nand U19793 (N_19793,N_10467,N_12794);
or U19794 (N_19794,N_14170,N_12779);
xor U19795 (N_19795,N_13255,N_14888);
or U19796 (N_19796,N_13511,N_11102);
xnor U19797 (N_19797,N_11148,N_10172);
nor U19798 (N_19798,N_12578,N_12172);
nand U19799 (N_19799,N_13138,N_10089);
and U19800 (N_19800,N_14623,N_12243);
xnor U19801 (N_19801,N_12456,N_14582);
and U19802 (N_19802,N_10678,N_11471);
and U19803 (N_19803,N_12460,N_11972);
or U19804 (N_19804,N_14766,N_10957);
nor U19805 (N_19805,N_12865,N_13613);
or U19806 (N_19806,N_10654,N_10007);
and U19807 (N_19807,N_13103,N_13530);
nor U19808 (N_19808,N_13840,N_11852);
nor U19809 (N_19809,N_14232,N_10141);
or U19810 (N_19810,N_11026,N_13485);
and U19811 (N_19811,N_12213,N_13028);
and U19812 (N_19812,N_11709,N_10822);
nor U19813 (N_19813,N_13108,N_10099);
nor U19814 (N_19814,N_11300,N_10146);
nor U19815 (N_19815,N_10564,N_11944);
nor U19816 (N_19816,N_11569,N_12212);
and U19817 (N_19817,N_14448,N_10400);
nand U19818 (N_19818,N_10050,N_11618);
nor U19819 (N_19819,N_11026,N_11312);
xor U19820 (N_19820,N_10274,N_14688);
and U19821 (N_19821,N_13372,N_10034);
xor U19822 (N_19822,N_13285,N_10961);
nor U19823 (N_19823,N_12452,N_13300);
nand U19824 (N_19824,N_10496,N_10211);
xor U19825 (N_19825,N_11187,N_12777);
nand U19826 (N_19826,N_13241,N_10641);
and U19827 (N_19827,N_12894,N_12940);
or U19828 (N_19828,N_10753,N_11261);
nand U19829 (N_19829,N_10557,N_13734);
nor U19830 (N_19830,N_13813,N_10500);
or U19831 (N_19831,N_13886,N_13044);
xor U19832 (N_19832,N_10976,N_13732);
and U19833 (N_19833,N_13728,N_13751);
nand U19834 (N_19834,N_14578,N_10393);
xor U19835 (N_19835,N_14688,N_11985);
xnor U19836 (N_19836,N_13136,N_13154);
and U19837 (N_19837,N_13216,N_14341);
nor U19838 (N_19838,N_10951,N_12324);
and U19839 (N_19839,N_11631,N_10260);
or U19840 (N_19840,N_10527,N_13316);
or U19841 (N_19841,N_13415,N_14878);
and U19842 (N_19842,N_11996,N_10418);
nand U19843 (N_19843,N_12175,N_12299);
or U19844 (N_19844,N_13411,N_10710);
nand U19845 (N_19845,N_11889,N_10452);
nor U19846 (N_19846,N_14262,N_12548);
and U19847 (N_19847,N_10885,N_11012);
nor U19848 (N_19848,N_13491,N_14907);
and U19849 (N_19849,N_12821,N_10400);
nand U19850 (N_19850,N_11937,N_11328);
nor U19851 (N_19851,N_13975,N_10018);
nand U19852 (N_19852,N_12380,N_12740);
or U19853 (N_19853,N_14805,N_10268);
and U19854 (N_19854,N_13089,N_12244);
nor U19855 (N_19855,N_14224,N_11378);
nand U19856 (N_19856,N_11350,N_14782);
xnor U19857 (N_19857,N_10246,N_14626);
and U19858 (N_19858,N_13621,N_13767);
or U19859 (N_19859,N_12423,N_13096);
nand U19860 (N_19860,N_10883,N_12446);
nand U19861 (N_19861,N_11009,N_11246);
and U19862 (N_19862,N_12512,N_12174);
and U19863 (N_19863,N_13947,N_14003);
nor U19864 (N_19864,N_13470,N_13613);
and U19865 (N_19865,N_11909,N_11766);
or U19866 (N_19866,N_12869,N_11204);
or U19867 (N_19867,N_11525,N_12033);
nor U19868 (N_19868,N_14957,N_10761);
nor U19869 (N_19869,N_12772,N_14008);
nand U19870 (N_19870,N_14039,N_14810);
nor U19871 (N_19871,N_11157,N_12111);
or U19872 (N_19872,N_14154,N_13682);
nand U19873 (N_19873,N_13434,N_10605);
nand U19874 (N_19874,N_12518,N_12593);
nor U19875 (N_19875,N_12349,N_10714);
or U19876 (N_19876,N_11604,N_14999);
xnor U19877 (N_19877,N_12239,N_11870);
or U19878 (N_19878,N_10389,N_12078);
nand U19879 (N_19879,N_12110,N_10010);
and U19880 (N_19880,N_10040,N_10310);
nand U19881 (N_19881,N_14627,N_12949);
or U19882 (N_19882,N_10896,N_10689);
or U19883 (N_19883,N_13054,N_13248);
nand U19884 (N_19884,N_11380,N_14374);
xor U19885 (N_19885,N_14635,N_13863);
nand U19886 (N_19886,N_11206,N_12075);
xor U19887 (N_19887,N_11608,N_11808);
and U19888 (N_19888,N_14934,N_12025);
nor U19889 (N_19889,N_14387,N_13354);
nand U19890 (N_19890,N_14541,N_14389);
nor U19891 (N_19891,N_11135,N_10342);
and U19892 (N_19892,N_13866,N_14572);
or U19893 (N_19893,N_13535,N_10927);
nand U19894 (N_19894,N_11815,N_12532);
and U19895 (N_19895,N_12297,N_14302);
or U19896 (N_19896,N_14310,N_10212);
xnor U19897 (N_19897,N_14756,N_10187);
and U19898 (N_19898,N_12627,N_14684);
nand U19899 (N_19899,N_12813,N_11347);
and U19900 (N_19900,N_13033,N_11376);
xor U19901 (N_19901,N_14927,N_13805);
and U19902 (N_19902,N_10335,N_11940);
or U19903 (N_19903,N_13874,N_10598);
nand U19904 (N_19904,N_12407,N_10356);
nand U19905 (N_19905,N_11117,N_11529);
and U19906 (N_19906,N_10304,N_10904);
nand U19907 (N_19907,N_12607,N_10815);
nand U19908 (N_19908,N_11599,N_14546);
nor U19909 (N_19909,N_11866,N_10109);
and U19910 (N_19910,N_13017,N_14159);
or U19911 (N_19911,N_14332,N_11037);
nor U19912 (N_19912,N_10223,N_12695);
or U19913 (N_19913,N_14382,N_10669);
and U19914 (N_19914,N_13584,N_11446);
nand U19915 (N_19915,N_13747,N_10144);
nand U19916 (N_19916,N_11527,N_13998);
or U19917 (N_19917,N_14839,N_11524);
or U19918 (N_19918,N_13675,N_11362);
or U19919 (N_19919,N_12148,N_12832);
and U19920 (N_19920,N_10257,N_14192);
xor U19921 (N_19921,N_10557,N_14264);
or U19922 (N_19922,N_14665,N_10778);
and U19923 (N_19923,N_13659,N_13260);
or U19924 (N_19924,N_12850,N_12979);
or U19925 (N_19925,N_10477,N_10602);
and U19926 (N_19926,N_12754,N_12273);
and U19927 (N_19927,N_11630,N_10247);
nand U19928 (N_19928,N_14054,N_10700);
or U19929 (N_19929,N_11623,N_10866);
nor U19930 (N_19930,N_10296,N_11012);
nand U19931 (N_19931,N_11467,N_10022);
nor U19932 (N_19932,N_13224,N_14084);
nand U19933 (N_19933,N_13479,N_12957);
or U19934 (N_19934,N_14214,N_11105);
or U19935 (N_19935,N_10423,N_12530);
or U19936 (N_19936,N_14765,N_13539);
xnor U19937 (N_19937,N_10599,N_14272);
nor U19938 (N_19938,N_13429,N_13976);
or U19939 (N_19939,N_10631,N_14139);
and U19940 (N_19940,N_13136,N_11625);
xnor U19941 (N_19941,N_13361,N_10922);
nand U19942 (N_19942,N_11774,N_10948);
nor U19943 (N_19943,N_11415,N_13110);
or U19944 (N_19944,N_12512,N_13739);
and U19945 (N_19945,N_13606,N_12854);
and U19946 (N_19946,N_13535,N_12860);
or U19947 (N_19947,N_14905,N_13729);
nor U19948 (N_19948,N_11481,N_13355);
or U19949 (N_19949,N_14960,N_11759);
or U19950 (N_19950,N_10406,N_12233);
nor U19951 (N_19951,N_11223,N_10959);
nor U19952 (N_19952,N_11474,N_10284);
xnor U19953 (N_19953,N_10122,N_10942);
nand U19954 (N_19954,N_14102,N_12089);
and U19955 (N_19955,N_14017,N_12931);
xor U19956 (N_19956,N_12533,N_13370);
and U19957 (N_19957,N_13232,N_14236);
or U19958 (N_19958,N_10926,N_10424);
and U19959 (N_19959,N_13509,N_10498);
nand U19960 (N_19960,N_10893,N_11261);
or U19961 (N_19961,N_11558,N_12693);
and U19962 (N_19962,N_12694,N_13303);
xnor U19963 (N_19963,N_12336,N_11180);
and U19964 (N_19964,N_11510,N_11199);
or U19965 (N_19965,N_11668,N_10991);
nand U19966 (N_19966,N_14721,N_10096);
nor U19967 (N_19967,N_14048,N_14109);
or U19968 (N_19968,N_10057,N_10719);
or U19969 (N_19969,N_11557,N_11205);
xnor U19970 (N_19970,N_11825,N_13632);
and U19971 (N_19971,N_13039,N_11543);
nor U19972 (N_19972,N_12151,N_13515);
nand U19973 (N_19973,N_12135,N_10265);
xnor U19974 (N_19974,N_13482,N_11478);
nor U19975 (N_19975,N_12458,N_13419);
nand U19976 (N_19976,N_12089,N_11304);
nor U19977 (N_19977,N_13740,N_10856);
nand U19978 (N_19978,N_12192,N_14690);
nor U19979 (N_19979,N_11530,N_13727);
or U19980 (N_19980,N_14908,N_11664);
xor U19981 (N_19981,N_11207,N_13675);
xnor U19982 (N_19982,N_12368,N_12342);
nand U19983 (N_19983,N_13672,N_10359);
nor U19984 (N_19984,N_13007,N_12657);
xor U19985 (N_19985,N_14761,N_13553);
or U19986 (N_19986,N_12765,N_12017);
nor U19987 (N_19987,N_12807,N_14017);
nor U19988 (N_19988,N_14376,N_13688);
and U19989 (N_19989,N_10004,N_14565);
and U19990 (N_19990,N_11263,N_13911);
nor U19991 (N_19991,N_14966,N_13904);
nor U19992 (N_19992,N_12460,N_12027);
nor U19993 (N_19993,N_12358,N_11816);
nor U19994 (N_19994,N_12430,N_14576);
nand U19995 (N_19995,N_14485,N_12969);
nor U19996 (N_19996,N_10039,N_13866);
xor U19997 (N_19997,N_11992,N_10788);
and U19998 (N_19998,N_13505,N_10002);
or U19999 (N_19999,N_13783,N_13954);
and U20000 (N_20000,N_18680,N_16253);
or U20001 (N_20001,N_15438,N_16863);
and U20002 (N_20002,N_16040,N_15071);
and U20003 (N_20003,N_16114,N_17795);
or U20004 (N_20004,N_18960,N_18085);
nand U20005 (N_20005,N_19238,N_17310);
and U20006 (N_20006,N_18916,N_17863);
and U20007 (N_20007,N_17450,N_17134);
nor U20008 (N_20008,N_15934,N_19890);
or U20009 (N_20009,N_16617,N_19098);
or U20010 (N_20010,N_18641,N_16756);
nor U20011 (N_20011,N_18084,N_17517);
nor U20012 (N_20012,N_19863,N_18290);
and U20013 (N_20013,N_19386,N_19639);
nor U20014 (N_20014,N_16461,N_15311);
or U20015 (N_20015,N_15608,N_15022);
and U20016 (N_20016,N_18650,N_17510);
nor U20017 (N_20017,N_15764,N_19810);
or U20018 (N_20018,N_17504,N_19821);
or U20019 (N_20019,N_16249,N_19579);
or U20020 (N_20020,N_17708,N_19813);
nor U20021 (N_20021,N_15024,N_18675);
or U20022 (N_20022,N_15594,N_15807);
nor U20023 (N_20023,N_17165,N_18741);
xor U20024 (N_20024,N_19086,N_17571);
or U20025 (N_20025,N_17373,N_19219);
or U20026 (N_20026,N_18712,N_17952);
and U20027 (N_20027,N_16551,N_19176);
or U20028 (N_20028,N_19940,N_16886);
or U20029 (N_20029,N_18321,N_16592);
nor U20030 (N_20030,N_15339,N_16792);
nor U20031 (N_20031,N_18262,N_19405);
xnor U20032 (N_20032,N_17512,N_15372);
and U20033 (N_20033,N_16939,N_17545);
xnor U20034 (N_20034,N_17052,N_15785);
or U20035 (N_20035,N_19761,N_19433);
xnor U20036 (N_20036,N_17726,N_16810);
nor U20037 (N_20037,N_16423,N_19037);
nand U20038 (N_20038,N_17663,N_17765);
nor U20039 (N_20039,N_19335,N_18893);
or U20040 (N_20040,N_16187,N_16287);
nor U20041 (N_20041,N_16086,N_15383);
and U20042 (N_20042,N_15564,N_16010);
xor U20043 (N_20043,N_15911,N_15473);
nor U20044 (N_20044,N_16186,N_19828);
nor U20045 (N_20045,N_15512,N_16787);
and U20046 (N_20046,N_19731,N_15603);
nand U20047 (N_20047,N_18306,N_17573);
or U20048 (N_20048,N_15411,N_17791);
nor U20049 (N_20049,N_15454,N_18217);
or U20050 (N_20050,N_16550,N_18630);
nand U20051 (N_20051,N_18663,N_16830);
and U20052 (N_20052,N_15646,N_15283);
xor U20053 (N_20053,N_17930,N_17678);
or U20054 (N_20054,N_17948,N_17323);
and U20055 (N_20055,N_16754,N_18662);
nor U20056 (N_20056,N_17981,N_15441);
and U20057 (N_20057,N_19625,N_16682);
and U20058 (N_20058,N_19599,N_17018);
or U20059 (N_20059,N_19374,N_17520);
or U20060 (N_20060,N_16318,N_16215);
nor U20061 (N_20061,N_18905,N_16416);
or U20062 (N_20062,N_15139,N_18096);
and U20063 (N_20063,N_17226,N_17731);
nand U20064 (N_20064,N_18181,N_17409);
and U20065 (N_20065,N_18081,N_16957);
and U20066 (N_20066,N_16664,N_15795);
and U20067 (N_20067,N_16841,N_17536);
xnor U20068 (N_20068,N_17874,N_15824);
nand U20069 (N_20069,N_17271,N_17554);
nand U20070 (N_20070,N_17679,N_16130);
xor U20071 (N_20071,N_19048,N_16744);
nand U20072 (N_20072,N_15739,N_15984);
xor U20073 (N_20073,N_15137,N_16609);
nor U20074 (N_20074,N_19215,N_17438);
and U20075 (N_20075,N_17759,N_16731);
or U20076 (N_20076,N_18330,N_19224);
and U20077 (N_20077,N_16056,N_19907);
or U20078 (N_20078,N_18099,N_16614);
or U20079 (N_20079,N_17222,N_15029);
xnor U20080 (N_20080,N_16204,N_17137);
nand U20081 (N_20081,N_19920,N_16611);
or U20082 (N_20082,N_18428,N_15352);
nand U20083 (N_20083,N_16448,N_18487);
and U20084 (N_20084,N_18743,N_17652);
or U20085 (N_20085,N_19962,N_15002);
or U20086 (N_20086,N_16209,N_15213);
xnor U20087 (N_20087,N_19188,N_17811);
nor U20088 (N_20088,N_18431,N_17370);
nand U20089 (N_20089,N_17204,N_15691);
nor U20090 (N_20090,N_17102,N_18913);
or U20091 (N_20091,N_17000,N_16050);
and U20092 (N_20092,N_18086,N_18606);
and U20093 (N_20093,N_19118,N_16389);
and U20094 (N_20094,N_16049,N_18264);
nand U20095 (N_20095,N_19422,N_18579);
and U20096 (N_20096,N_15574,N_17586);
or U20097 (N_20097,N_17912,N_17774);
and U20098 (N_20098,N_17229,N_17243);
nor U20099 (N_20099,N_16161,N_16667);
and U20100 (N_20100,N_17164,N_18043);
and U20101 (N_20101,N_19269,N_18507);
xor U20102 (N_20102,N_16653,N_15910);
nor U20103 (N_20103,N_15282,N_16620);
nand U20104 (N_20104,N_17352,N_18398);
or U20105 (N_20105,N_18065,N_15370);
nor U20106 (N_20106,N_19420,N_15822);
or U20107 (N_20107,N_17939,N_16973);
nand U20108 (N_20108,N_19683,N_15222);
nand U20109 (N_20109,N_18826,N_16350);
nor U20110 (N_20110,N_16442,N_19152);
or U20111 (N_20111,N_16446,N_19008);
xnor U20112 (N_20112,N_18756,N_18496);
or U20113 (N_20113,N_15091,N_15456);
xor U20114 (N_20114,N_16746,N_19467);
nor U20115 (N_20115,N_16743,N_16352);
and U20116 (N_20116,N_19820,N_16066);
nor U20117 (N_20117,N_18400,N_19024);
nand U20118 (N_20118,N_15609,N_16391);
or U20119 (N_20119,N_19489,N_15647);
nor U20120 (N_20120,N_17387,N_16212);
nor U20121 (N_20121,N_18516,N_15044);
and U20122 (N_20122,N_19357,N_18774);
xor U20123 (N_20123,N_16177,N_16636);
nor U20124 (N_20124,N_19830,N_19363);
nand U20125 (N_20125,N_18036,N_18269);
xnor U20126 (N_20126,N_15099,N_16102);
and U20127 (N_20127,N_18145,N_15409);
and U20128 (N_20128,N_19979,N_17158);
xnor U20129 (N_20129,N_16349,N_18623);
and U20130 (N_20130,N_18563,N_15358);
or U20131 (N_20131,N_19040,N_18237);
or U20132 (N_20132,N_16474,N_16332);
nand U20133 (N_20133,N_16121,N_18955);
and U20134 (N_20134,N_19450,N_19802);
or U20135 (N_20135,N_15748,N_19703);
and U20136 (N_20136,N_16842,N_15871);
or U20137 (N_20137,N_18926,N_19619);
nand U20138 (N_20138,N_18986,N_16286);
nand U20139 (N_20139,N_19610,N_18188);
or U20140 (N_20140,N_17804,N_19513);
xor U20141 (N_20141,N_17183,N_16296);
nor U20142 (N_20142,N_16877,N_15868);
nor U20143 (N_20143,N_17544,N_18928);
and U20144 (N_20144,N_15809,N_15954);
or U20145 (N_20145,N_18862,N_17338);
and U20146 (N_20146,N_17268,N_16179);
nor U20147 (N_20147,N_19471,N_16910);
nand U20148 (N_20148,N_19894,N_18534);
and U20149 (N_20149,N_15017,N_18042);
and U20150 (N_20150,N_15964,N_16099);
nor U20151 (N_20151,N_16907,N_15280);
and U20152 (N_20152,N_18484,N_16689);
or U20153 (N_20153,N_17224,N_19137);
nor U20154 (N_20154,N_16971,N_18793);
nor U20155 (N_20155,N_15433,N_16678);
or U20156 (N_20156,N_19136,N_17088);
nor U20157 (N_20157,N_18608,N_17643);
nand U20158 (N_20158,N_18041,N_15472);
or U20159 (N_20159,N_15776,N_18551);
nor U20160 (N_20160,N_18707,N_17660);
and U20161 (N_20161,N_17128,N_17139);
nor U20162 (N_20162,N_19641,N_19502);
nor U20163 (N_20163,N_19538,N_17464);
and U20164 (N_20164,N_15787,N_16324);
or U20165 (N_20165,N_16206,N_15404);
and U20166 (N_20166,N_18929,N_15401);
xnor U20167 (N_20167,N_17314,N_19875);
nand U20168 (N_20168,N_15829,N_16726);
nand U20169 (N_20169,N_17262,N_18273);
nor U20170 (N_20170,N_19547,N_18722);
nand U20171 (N_20171,N_17069,N_17360);
nand U20172 (N_20172,N_18270,N_15162);
and U20173 (N_20173,N_17451,N_19418);
and U20174 (N_20174,N_19917,N_15183);
nand U20175 (N_20175,N_18508,N_15986);
and U20176 (N_20176,N_16955,N_18223);
nor U20177 (N_20177,N_17665,N_18346);
and U20178 (N_20178,N_16216,N_18512);
nor U20179 (N_20179,N_15123,N_18369);
nor U20180 (N_20180,N_16479,N_19303);
nor U20181 (N_20181,N_18985,N_16972);
and U20182 (N_20182,N_18934,N_18924);
nor U20183 (N_20183,N_17965,N_18192);
or U20184 (N_20184,N_16103,N_15212);
nor U20185 (N_20185,N_17127,N_18800);
and U20186 (N_20186,N_18925,N_16561);
and U20187 (N_20187,N_19464,N_19768);
nand U20188 (N_20188,N_15380,N_18874);
xor U20189 (N_20189,N_17294,N_18616);
nor U20190 (N_20190,N_17951,N_19580);
nand U20191 (N_20191,N_15168,N_18464);
and U20192 (N_20192,N_15593,N_19025);
nand U20193 (N_20193,N_18203,N_15346);
nor U20194 (N_20194,N_17032,N_15789);
nor U20195 (N_20195,N_17225,N_16931);
and U20196 (N_20196,N_17816,N_17682);
or U20197 (N_20197,N_19012,N_17973);
nand U20198 (N_20198,N_18936,N_17074);
nor U20199 (N_20199,N_15519,N_15520);
nand U20200 (N_20200,N_15988,N_16748);
or U20201 (N_20201,N_15649,N_15275);
or U20202 (N_20202,N_18678,N_18747);
and U20203 (N_20203,N_17133,N_16909);
and U20204 (N_20204,N_18975,N_15130);
xnor U20205 (N_20205,N_17239,N_16541);
nand U20206 (N_20206,N_19328,N_17447);
nand U20207 (N_20207,N_18331,N_16404);
or U20208 (N_20208,N_19292,N_18174);
and U20209 (N_20209,N_15354,N_18024);
and U20210 (N_20210,N_16856,N_15686);
nand U20211 (N_20211,N_15154,N_18129);
nor U20212 (N_20212,N_19426,N_18108);
nor U20213 (N_20213,N_17056,N_17602);
and U20214 (N_20214,N_17796,N_17515);
nand U20215 (N_20215,N_19986,N_17778);
nand U20216 (N_20216,N_16312,N_15299);
and U20217 (N_20217,N_18639,N_18821);
nand U20218 (N_20218,N_17532,N_17563);
nand U20219 (N_20219,N_15205,N_19101);
nand U20220 (N_20220,N_16127,N_16380);
or U20221 (N_20221,N_16301,N_18922);
and U20222 (N_20222,N_16284,N_19856);
and U20223 (N_20223,N_19053,N_18473);
xor U20224 (N_20224,N_15126,N_19373);
or U20225 (N_20225,N_19996,N_16426);
nor U20226 (N_20226,N_18293,N_16591);
or U20227 (N_20227,N_18419,N_18116);
xor U20228 (N_20228,N_19371,N_19428);
nand U20229 (N_20229,N_16872,N_17126);
nand U20230 (N_20230,N_16603,N_19209);
nor U20231 (N_20231,N_15478,N_18891);
nand U20232 (N_20232,N_17557,N_18555);
nand U20233 (N_20233,N_19337,N_16510);
nor U20234 (N_20234,N_16079,N_18144);
or U20235 (N_20235,N_19900,N_17347);
nor U20236 (N_20236,N_16623,N_18471);
xor U20237 (N_20237,N_19801,N_15716);
nand U20238 (N_20238,N_17689,N_17743);
nand U20239 (N_20239,N_16950,N_17711);
and U20240 (N_20240,N_18478,N_18133);
and U20241 (N_20241,N_17701,N_15669);
or U20242 (N_20242,N_15874,N_15150);
nand U20243 (N_20243,N_18648,N_18425);
or U20244 (N_20244,N_17328,N_15155);
nor U20245 (N_20245,N_16666,N_15962);
nand U20246 (N_20246,N_16697,N_18786);
nor U20247 (N_20247,N_19211,N_15706);
nor U20248 (N_20248,N_16208,N_18697);
xor U20249 (N_20249,N_16776,N_17704);
nor U20250 (N_20250,N_15684,N_19148);
nor U20251 (N_20251,N_15901,N_16741);
xor U20252 (N_20252,N_18577,N_16537);
xor U20253 (N_20253,N_17921,N_16245);
and U20254 (N_20254,N_19916,N_19249);
or U20255 (N_20255,N_17854,N_18586);
nand U20256 (N_20256,N_19793,N_15439);
and U20257 (N_20257,N_17090,N_15097);
xnor U20258 (N_20258,N_19491,N_16055);
nor U20259 (N_20259,N_18131,N_19628);
xor U20260 (N_20260,N_16037,N_19734);
or U20261 (N_20261,N_19779,N_19930);
and U20262 (N_20262,N_15942,N_15839);
nor U20263 (N_20263,N_16257,N_18114);
or U20264 (N_20264,N_17728,N_16393);
and U20265 (N_20265,N_19403,N_19861);
nand U20266 (N_20266,N_16871,N_19961);
nand U20267 (N_20267,N_15586,N_18613);
nand U20268 (N_20268,N_18128,N_19800);
xnor U20269 (N_20269,N_17480,N_17695);
nand U20270 (N_20270,N_19794,N_16912);
xnor U20271 (N_20271,N_18714,N_15843);
and U20272 (N_20272,N_16001,N_15307);
nand U20273 (N_20273,N_17214,N_15216);
nand U20274 (N_20274,N_15252,N_18629);
nand U20275 (N_20275,N_17024,N_18204);
or U20276 (N_20276,N_17266,N_15906);
nand U20277 (N_20277,N_15049,N_17505);
nand U20278 (N_20278,N_19702,N_15078);
nand U20279 (N_20279,N_18869,N_17861);
and U20280 (N_20280,N_15236,N_17206);
or U20281 (N_20281,N_15034,N_19095);
nor U20282 (N_20282,N_17657,N_15258);
or U20283 (N_20283,N_15577,N_15284);
or U20284 (N_20284,N_18255,N_19015);
nor U20285 (N_20285,N_19382,N_16076);
nand U20286 (N_20286,N_16095,N_16882);
xnor U20287 (N_20287,N_16725,N_17406);
or U20288 (N_20288,N_16235,N_15791);
or U20289 (N_20289,N_17500,N_19334);
nor U20290 (N_20290,N_16547,N_17369);
nor U20291 (N_20291,N_18618,N_17051);
nor U20292 (N_20292,N_19609,N_15194);
nor U20293 (N_20293,N_17430,N_15513);
and U20294 (N_20294,N_15994,N_15345);
nand U20295 (N_20295,N_17882,N_19031);
or U20296 (N_20296,N_17290,N_16749);
nand U20297 (N_20297,N_15715,N_18635);
nor U20298 (N_20298,N_18567,N_19327);
or U20299 (N_20299,N_16439,N_15929);
nand U20300 (N_20300,N_15769,N_18052);
or U20301 (N_20301,N_17197,N_19929);
nand U20302 (N_20302,N_18651,N_19096);
or U20303 (N_20303,N_18412,N_18783);
and U20304 (N_20304,N_17582,N_15443);
nor U20305 (N_20305,N_17255,N_19822);
nor U20306 (N_20306,N_19922,N_18920);
nor U20307 (N_20307,N_16498,N_19348);
or U20308 (N_20308,N_16896,N_19717);
nor U20309 (N_20309,N_17754,N_16964);
nor U20310 (N_20310,N_19921,N_17371);
and U20311 (N_20311,N_19169,N_15337);
xnor U20312 (N_20312,N_17730,N_19870);
and U20313 (N_20313,N_18225,N_15820);
nor U20314 (N_20314,N_17788,N_16714);
or U20315 (N_20315,N_15625,N_18860);
nor U20316 (N_20316,N_15459,N_19709);
nand U20317 (N_20317,N_18164,N_16906);
nand U20318 (N_20318,N_19562,N_17810);
xor U20319 (N_20319,N_16884,N_19959);
nand U20320 (N_20320,N_19675,N_18730);
or U20321 (N_20321,N_15878,N_19362);
nor U20322 (N_20322,N_19985,N_19456);
or U20323 (N_20323,N_15886,N_19650);
nand U20324 (N_20324,N_18620,N_19265);
xnor U20325 (N_20325,N_15487,N_17291);
nor U20326 (N_20326,N_15344,N_16529);
and U20327 (N_20327,N_19868,N_18523);
or U20328 (N_20328,N_17633,N_19207);
or U20329 (N_20329,N_17471,N_15696);
nand U20330 (N_20330,N_17960,N_15595);
nor U20331 (N_20331,N_18206,N_17993);
nand U20332 (N_20332,N_15397,N_16963);
nand U20333 (N_20333,N_15885,N_17770);
nor U20334 (N_20334,N_15179,N_17168);
and U20335 (N_20335,N_17033,N_19558);
or U20336 (N_20336,N_19615,N_17876);
nand U20337 (N_20337,N_18360,N_18596);
nor U20338 (N_20338,N_16732,N_18978);
and U20339 (N_20339,N_18760,N_18900);
and U20340 (N_20340,N_16643,N_17866);
or U20341 (N_20341,N_19771,N_19640);
or U20342 (N_20342,N_15730,N_17160);
and U20343 (N_20343,N_16181,N_15614);
or U20344 (N_20344,N_17123,N_17455);
or U20345 (N_20345,N_17150,N_16915);
or U20346 (N_20346,N_15710,N_15494);
nor U20347 (N_20347,N_16961,N_17004);
xnor U20348 (N_20348,N_17762,N_18031);
or U20349 (N_20349,N_15548,N_19617);
nor U20350 (N_20350,N_16034,N_17267);
nand U20351 (N_20351,N_17681,N_16000);
and U20352 (N_20352,N_15979,N_15606);
nor U20353 (N_20353,N_19947,N_18113);
and U20354 (N_20354,N_18382,N_17961);
nand U20355 (N_20355,N_18526,N_18669);
or U20356 (N_20356,N_16951,N_19692);
or U20357 (N_20357,N_18836,N_17926);
nor U20358 (N_20358,N_17490,N_16779);
nor U20359 (N_20359,N_19919,N_18310);
nor U20360 (N_20360,N_17814,N_18418);
xnor U20361 (N_20361,N_17379,N_15991);
nor U20362 (N_20362,N_15491,N_18448);
nor U20363 (N_20363,N_18311,N_15961);
and U20364 (N_20364,N_18820,N_15160);
and U20365 (N_20365,N_18040,N_19147);
or U20366 (N_20366,N_15766,N_18530);
or U20367 (N_20367,N_18137,N_17182);
and U20368 (N_20368,N_19622,N_17924);
nor U20369 (N_20369,N_16256,N_17333);
nor U20370 (N_20370,N_15151,N_16460);
xnor U20371 (N_20371,N_17015,N_17629);
xor U20372 (N_20372,N_16451,N_17761);
and U20373 (N_20373,N_18091,N_18120);
nor U20374 (N_20374,N_18536,N_16713);
or U20375 (N_20375,N_16342,N_18658);
and U20376 (N_20376,N_19333,N_19054);
nand U20377 (N_20377,N_15127,N_19448);
nand U20378 (N_20378,N_16465,N_19993);
xnor U20379 (N_20379,N_17990,N_17121);
xor U20380 (N_20380,N_15622,N_15356);
nor U20381 (N_20381,N_17440,N_19604);
nand U20382 (N_20382,N_17446,N_17215);
nand U20383 (N_20383,N_16226,N_16337);
xor U20384 (N_20384,N_17299,N_16969);
nand U20385 (N_20385,N_17170,N_17149);
nor U20386 (N_20386,N_19708,N_18199);
nor U20387 (N_20387,N_17035,N_19026);
and U20388 (N_20388,N_17188,N_16456);
or U20389 (N_20389,N_19595,N_18570);
nand U20390 (N_20390,N_19281,N_18778);
nand U20391 (N_20391,N_17145,N_15845);
nand U20392 (N_20392,N_17390,N_19546);
or U20393 (N_20393,N_19023,N_18685);
or U20394 (N_20394,N_16525,N_15321);
nand U20395 (N_20395,N_19463,N_18767);
nor U20396 (N_20396,N_17334,N_19700);
xnor U20397 (N_20397,N_15529,N_18395);
nor U20398 (N_20398,N_17904,N_16579);
nand U20399 (N_20399,N_19988,N_17664);
nand U20400 (N_20400,N_15110,N_16976);
and U20401 (N_20401,N_18763,N_15814);
nand U20402 (N_20402,N_18068,N_16429);
or U20403 (N_20403,N_18894,N_16003);
or U20404 (N_20404,N_19258,N_16436);
and U20405 (N_20405,N_16897,N_19059);
nor U20406 (N_20406,N_16853,N_17624);
and U20407 (N_20407,N_16953,N_15825);
and U20408 (N_20408,N_19107,N_18194);
and U20409 (N_20409,N_17671,N_17254);
nor U20410 (N_20410,N_19998,N_16230);
nand U20411 (N_20411,N_17097,N_17933);
nor U20412 (N_20412,N_17906,N_19946);
nand U20413 (N_20413,N_19738,N_16220);
nor U20414 (N_20414,N_17666,N_17959);
or U20415 (N_20415,N_17400,N_19166);
nand U20416 (N_20416,N_17306,N_18885);
or U20417 (N_20417,N_15448,N_17099);
and U20418 (N_20418,N_16699,N_19378);
nand U20419 (N_20419,N_16017,N_16967);
nor U20420 (N_20420,N_16098,N_17292);
and U20421 (N_20421,N_19069,N_16402);
nor U20422 (N_20422,N_19311,N_16300);
nor U20423 (N_20423,N_16934,N_16126);
nor U20424 (N_20424,N_16918,N_18598);
nor U20425 (N_20425,N_19637,N_19085);
and U20426 (N_20426,N_15800,N_15481);
nor U20427 (N_20427,N_15140,N_18098);
or U20428 (N_20428,N_16762,N_16885);
nor U20429 (N_20429,N_18968,N_18033);
nor U20430 (N_20430,N_15077,N_15844);
and U20431 (N_20431,N_16539,N_16149);
or U20432 (N_20432,N_16310,N_16362);
nand U20433 (N_20433,N_15920,N_16100);
nor U20434 (N_20434,N_17079,N_18316);
nor U20435 (N_20435,N_16061,N_16813);
or U20436 (N_20436,N_19174,N_15932);
and U20437 (N_20437,N_16588,N_16587);
and U20438 (N_20438,N_19056,N_18969);
or U20439 (N_20439,N_15281,N_19424);
or U20440 (N_20440,N_18835,N_17011);
nand U20441 (N_20441,N_16077,N_15772);
nor U20442 (N_20442,N_19545,N_18766);
xnor U20443 (N_20443,N_19079,N_17862);
and U20444 (N_20444,N_15249,N_16309);
and U20445 (N_20445,N_19742,N_18132);
nand U20446 (N_20446,N_19100,N_15851);
nor U20447 (N_20447,N_18365,N_19167);
nand U20448 (N_20448,N_15734,N_16693);
and U20449 (N_20449,N_15195,N_15161);
nand U20450 (N_20450,N_16238,N_19648);
or U20451 (N_20451,N_19255,N_18148);
nand U20452 (N_20452,N_18983,N_17697);
and U20453 (N_20453,N_15200,N_19182);
nand U20454 (N_20454,N_17417,N_18657);
nand U20455 (N_20455,N_17136,N_18610);
xor U20456 (N_20456,N_19193,N_19787);
and U20457 (N_20457,N_15244,N_18519);
nor U20458 (N_20458,N_18037,N_15351);
nand U20459 (N_20459,N_19361,N_17949);
nand U20460 (N_20460,N_19872,N_19543);
and U20461 (N_20461,N_17095,N_18938);
and U20462 (N_20462,N_19780,N_16926);
and U20463 (N_20463,N_15571,N_18724);
xor U20464 (N_20464,N_19831,N_15660);
nand U20465 (N_20465,N_19298,N_19050);
or U20466 (N_20466,N_15938,N_17955);
and U20467 (N_20467,N_19388,N_17138);
xor U20468 (N_20468,N_18472,N_19633);
nand U20469 (N_20469,N_18621,N_16033);
or U20470 (N_20470,N_18073,N_17055);
nor U20471 (N_20471,N_17424,N_19932);
or U20472 (N_20472,N_18720,N_19105);
nor U20473 (N_20473,N_16428,N_15550);
or U20474 (N_20474,N_16685,N_16109);
and U20475 (N_20475,N_16190,N_15523);
nor U20476 (N_20476,N_18443,N_18304);
xnor U20477 (N_20477,N_18397,N_15483);
xor U20478 (N_20478,N_17231,N_18465);
and U20479 (N_20479,N_19485,N_16839);
and U20480 (N_20480,N_19091,N_19377);
nand U20481 (N_20481,N_16785,N_19351);
and U20482 (N_20482,N_19161,N_19419);
and U20483 (N_20483,N_16798,N_15642);
or U20484 (N_20484,N_17783,N_19829);
xor U20485 (N_20485,N_17166,N_16512);
nand U20486 (N_20486,N_18529,N_19482);
nand U20487 (N_20487,N_19751,N_16898);
and U20488 (N_20488,N_15663,N_15267);
and U20489 (N_20489,N_19109,N_19332);
and U20490 (N_20490,N_18965,N_18746);
or U20491 (N_20491,N_19807,N_19329);
nor U20492 (N_20492,N_18261,N_17800);
nor U20493 (N_20493,N_19286,N_17997);
and U20494 (N_20494,N_16684,N_16517);
nor U20495 (N_20495,N_17491,N_15969);
or U20496 (N_20496,N_15892,N_17572);
or U20497 (N_20497,N_17321,N_17392);
or U20498 (N_20498,N_17014,N_15304);
and U20499 (N_20499,N_16409,N_15653);
or U20500 (N_20500,N_18542,N_15723);
nor U20501 (N_20501,N_16879,N_17481);
nand U20502 (N_20502,N_15418,N_18326);
or U20503 (N_20503,N_16306,N_16170);
xnor U20504 (N_20504,N_16467,N_15621);
nand U20505 (N_20505,N_15361,N_19819);
nand U20506 (N_20506,N_16608,N_19505);
and U20507 (N_20507,N_16093,N_17489);
or U20508 (N_20508,N_17896,N_17120);
and U20509 (N_20509,N_19789,N_15040);
and U20510 (N_20510,N_17460,N_15579);
nor U20511 (N_20511,N_15475,N_17767);
or U20512 (N_20512,N_16998,N_16760);
or U20513 (N_20513,N_19898,N_16155);
nor U20514 (N_20514,N_18322,N_16530);
xor U20515 (N_20515,N_19066,N_17036);
nor U20516 (N_20516,N_15793,N_18334);
nand U20517 (N_20517,N_15309,N_19613);
xnor U20518 (N_20518,N_17881,N_16084);
nand U20519 (N_20519,N_18661,N_15832);
nor U20520 (N_20520,N_18653,N_16786);
or U20521 (N_20521,N_16736,N_17022);
or U20522 (N_20522,N_15872,N_19150);
and U20523 (N_20523,N_15864,N_15303);
nor U20524 (N_20524,N_15292,N_15098);
nand U20525 (N_20525,N_17620,N_19564);
nor U20526 (N_20526,N_17203,N_19171);
nor U20527 (N_20527,N_16979,N_18353);
nor U20528 (N_20528,N_19847,N_16029);
and U20529 (N_20529,N_16606,N_18539);
and U20530 (N_20530,N_15084,N_17642);
nand U20531 (N_20531,N_15956,N_19237);
or U20532 (N_20532,N_17698,N_19933);
xnor U20533 (N_20533,N_18672,N_19638);
nor U20534 (N_20534,N_17928,N_19969);
nor U20535 (N_20535,N_19806,N_19210);
and U20536 (N_20536,N_17116,N_16106);
xor U20537 (N_20537,N_15350,N_19094);
nor U20538 (N_20538,N_16015,N_15186);
and U20539 (N_20539,N_19839,N_17122);
and U20540 (N_20540,N_17172,N_15322);
nand U20541 (N_20541,N_15582,N_15502);
nand U20542 (N_20542,N_15514,N_19304);
and U20543 (N_20543,N_18125,N_15738);
and U20544 (N_20544,N_17901,N_18066);
nand U20545 (N_20545,N_15985,N_16665);
and U20546 (N_20546,N_17335,N_16582);
nand U20547 (N_20547,N_17175,N_15695);
and U20548 (N_20548,N_15143,N_16662);
or U20549 (N_20549,N_18176,N_15288);
nor U20550 (N_20550,N_15987,N_15101);
or U20551 (N_20551,N_15899,N_17974);
nand U20552 (N_20552,N_16691,N_15315);
or U20553 (N_20553,N_15405,N_19439);
and U20554 (N_20554,N_19088,N_18294);
and U20555 (N_20555,N_15215,N_16956);
xnor U20556 (N_20556,N_17821,N_15256);
nand U20557 (N_20557,N_19125,N_17162);
nor U20558 (N_20558,N_19022,N_15152);
nand U20559 (N_20559,N_16980,N_18340);
or U20560 (N_20560,N_18328,N_19203);
nor U20561 (N_20561,N_16395,N_17385);
or U20562 (N_20562,N_17274,N_18158);
nor U20563 (N_20563,N_17411,N_15308);
nand U20564 (N_20564,N_19438,N_17105);
or U20565 (N_20565,N_17897,N_18357);
nand U20566 (N_20566,N_15341,N_18488);
or U20567 (N_20567,N_15955,N_19285);
nand U20568 (N_20568,N_16900,N_17826);
and U20569 (N_20569,N_19989,N_16021);
or U20570 (N_20570,N_16970,N_15270);
xnor U20571 (N_20571,N_16648,N_19866);
or U20572 (N_20572,N_18286,N_17546);
and U20573 (N_20573,N_16695,N_15014);
nand U20574 (N_20574,N_19122,N_15254);
nand U20575 (N_20575,N_18350,N_16729);
nor U20576 (N_20576,N_19090,N_16073);
nand U20577 (N_20577,N_17819,N_15963);
nand U20578 (N_20578,N_18455,N_18638);
nand U20579 (N_20579,N_19753,N_15941);
nor U20580 (N_20580,N_19507,N_16925);
nand U20581 (N_20581,N_17540,N_18141);
and U20582 (N_20582,N_18106,N_17789);
and U20583 (N_20583,N_16009,N_17478);
and U20584 (N_20584,N_16765,N_19585);
or U20585 (N_20585,N_15705,N_17048);
or U20586 (N_20586,N_16346,N_18414);
nor U20587 (N_20587,N_18585,N_19607);
xor U20588 (N_20588,N_18959,N_17300);
nand U20589 (N_20589,N_15238,N_17736);
or U20590 (N_20590,N_15768,N_19896);
nor U20591 (N_20591,N_17850,N_17604);
nor U20592 (N_20592,N_15879,N_15265);
nand U20593 (N_20593,N_17601,N_16861);
nor U20594 (N_20594,N_18706,N_19559);
nand U20595 (N_20595,N_15497,N_18583);
or U20596 (N_20596,N_16457,N_15960);
or U20597 (N_20597,N_16433,N_18146);
and U20598 (N_20598,N_16158,N_15816);
nor U20599 (N_20599,N_19548,N_15767);
and U20600 (N_20600,N_15980,N_16661);
nor U20601 (N_20601,N_15336,N_15020);
nor U20602 (N_20602,N_19886,N_19719);
and U20603 (N_20603,N_15469,N_19528);
and U20604 (N_20604,N_17030,N_18553);
and U20605 (N_20605,N_15403,N_16089);
nand U20606 (N_20606,N_18560,N_19903);
nor U20607 (N_20607,N_17848,N_19712);
or U20608 (N_20608,N_19437,N_16398);
nand U20609 (N_20609,N_19733,N_16947);
and U20610 (N_20610,N_17258,N_16070);
or U20611 (N_20611,N_18368,N_18196);
nor U20612 (N_20612,N_18126,N_19116);
nor U20613 (N_20613,N_17967,N_17198);
nand U20614 (N_20614,N_18918,N_16891);
nor U20615 (N_20615,N_17616,N_17673);
nand U20616 (N_20616,N_18160,N_17516);
and U20617 (N_20617,N_18233,N_19632);
nand U20618 (N_20618,N_19765,N_15096);
nand U20619 (N_20619,N_17298,N_15692);
nor U20620 (N_20620,N_17538,N_19033);
or U20621 (N_20621,N_19676,N_15070);
nor U20622 (N_20622,N_15210,N_16974);
or U20623 (N_20623,N_17191,N_17005);
nand U20624 (N_20624,N_15721,N_17787);
xnor U20625 (N_20625,N_16355,N_15794);
and U20626 (N_20626,N_19356,N_15480);
and U20627 (N_20627,N_19696,N_15717);
nand U20628 (N_20628,N_18263,N_19657);
or U20629 (N_20629,N_18424,N_18640);
or U20630 (N_20630,N_19966,N_19112);
and U20631 (N_20631,N_15854,N_17644);
and U20632 (N_20632,N_15652,N_16983);
xor U20633 (N_20633,N_16986,N_19379);
or U20634 (N_20634,N_15719,N_18260);
or U20635 (N_20635,N_18297,N_16225);
or U20636 (N_20636,N_15615,N_16039);
nor U20637 (N_20637,N_18045,N_16977);
nand U20638 (N_20638,N_17146,N_16219);
nor U20639 (N_20639,N_18665,N_17742);
or U20640 (N_20640,N_17931,N_17972);
or U20641 (N_20641,N_19612,N_17234);
and U20642 (N_20642,N_18361,N_17688);
and U20643 (N_20643,N_15619,N_18387);
nand U20644 (N_20644,N_19194,N_16605);
and U20645 (N_20645,N_15778,N_19741);
or U20646 (N_20646,N_17610,N_18094);
nor U20647 (N_20647,N_19243,N_19525);
and U20648 (N_20648,N_19710,N_17257);
and U20649 (N_20649,N_18168,N_19257);
nand U20650 (N_20650,N_17457,N_19178);
nor U20651 (N_20651,N_17724,N_17991);
nor U20652 (N_20652,N_19200,N_18951);
nand U20653 (N_20653,N_18870,N_16458);
and U20654 (N_20654,N_16718,N_17154);
nor U20655 (N_20655,N_15944,N_15058);
or U20656 (N_20656,N_17043,N_19837);
or U20657 (N_20657,N_18213,N_15326);
or U20658 (N_20658,N_16311,N_19248);
or U20659 (N_20659,N_17521,N_18319);
nor U20660 (N_20660,N_15940,N_16651);
xor U20661 (N_20661,N_15442,N_18899);
and U20662 (N_20662,N_19895,N_18725);
nand U20663 (N_20663,N_19749,N_15664);
nor U20664 (N_20664,N_17625,N_15041);
or U20665 (N_20665,N_19421,N_17284);
or U20666 (N_20666,N_17468,N_16595);
or U20667 (N_20667,N_18679,N_17838);
nand U20668 (N_20668,N_16329,N_15959);
nor U20669 (N_20669,N_15516,N_17727);
nand U20670 (N_20670,N_15109,N_19783);
or U20671 (N_20671,N_17979,N_15273);
nor U20672 (N_20672,N_18284,N_18505);
and U20673 (N_20673,N_19451,N_19699);
nand U20674 (N_20674,N_17776,N_19244);
nand U20675 (N_20675,N_17556,N_15509);
nor U20676 (N_20676,N_15263,N_19208);
or U20677 (N_20677,N_19729,N_15763);
nor U20678 (N_20678,N_19982,N_15325);
nand U20679 (N_20679,N_15575,N_17445);
nor U20680 (N_20680,N_15422,N_17944);
nor U20681 (N_20681,N_16672,N_17525);
nand U20682 (N_20682,N_15501,N_15209);
nand U20683 (N_20683,N_15460,N_16988);
and U20684 (N_20684,N_18761,N_16727);
or U20685 (N_20685,N_17087,N_15461);
or U20686 (N_20686,N_16113,N_16316);
or U20687 (N_20687,N_15290,N_19713);
and U20688 (N_20688,N_17593,N_19106);
nand U20689 (N_20689,N_17089,N_18420);
or U20690 (N_20690,N_19720,N_15072);
or U20691 (N_20691,N_19019,N_17713);
or U20692 (N_20692,N_17617,N_17608);
nand U20693 (N_20693,N_17712,N_15743);
and U20694 (N_20694,N_18504,N_17180);
nand U20695 (N_20695,N_17063,N_19995);
xnor U20696 (N_20696,N_15367,N_16940);
nand U20697 (N_20697,N_18147,N_18710);
or U20698 (N_20698,N_17046,N_19556);
xnor U20699 (N_20699,N_18824,N_18587);
and U20700 (N_20700,N_18102,N_18327);
or U20701 (N_20701,N_19515,N_19314);
nand U20702 (N_20702,N_16107,N_15784);
and U20703 (N_20703,N_18789,N_15266);
nand U20704 (N_20704,N_19569,N_17235);
or U20705 (N_20705,N_17053,N_17768);
and U20706 (N_20706,N_15122,N_19796);
nor U20707 (N_20707,N_16088,N_17322);
nor U20708 (N_20708,N_15765,N_18709);
or U20709 (N_20709,N_16405,N_18376);
or U20710 (N_20710,N_16562,N_17715);
and U20711 (N_20711,N_16450,N_19232);
nor U20712 (N_20712,N_19146,N_15038);
nor U20713 (N_20713,N_15952,N_16984);
or U20714 (N_20714,N_17739,N_19576);
xor U20715 (N_20715,N_18642,N_17858);
and U20716 (N_20716,N_19554,N_19519);
or U20717 (N_20717,N_16567,N_16356);
or U20718 (N_20718,N_19750,N_18251);
nand U20719 (N_20719,N_16738,N_19956);
nor U20720 (N_20720,N_19039,N_18363);
nor U20721 (N_20721,N_19473,N_18333);
or U20722 (N_20722,N_15223,N_16232);
xor U20723 (N_20723,N_18892,N_15505);
nand U20724 (N_20724,N_17619,N_15635);
xnor U20725 (N_20725,N_15206,N_16348);
and U20726 (N_20726,N_17890,N_16873);
nor U20727 (N_20727,N_18035,N_17662);
and U20728 (N_20728,N_17110,N_16002);
and U20729 (N_20729,N_19010,N_16011);
nand U20730 (N_20730,N_17331,N_19359);
nor U20731 (N_20731,N_18528,N_15108);
nand U20732 (N_20732,N_16014,N_18480);
or U20733 (N_20733,N_16519,N_19411);
nor U20734 (N_20734,N_19511,N_18970);
nor U20735 (N_20735,N_15668,N_17067);
or U20736 (N_20736,N_17330,N_19394);
xor U20737 (N_20737,N_15602,N_18942);
and U20738 (N_20738,N_15801,N_16270);
or U20739 (N_20739,N_17156,N_19384);
nor U20740 (N_20740,N_19756,N_17710);
nand U20741 (N_20741,N_15826,N_16092);
nand U20742 (N_20742,N_19603,N_19656);
and U20743 (N_20743,N_18385,N_16004);
or U20744 (N_20744,N_17236,N_18019);
and U20745 (N_20745,N_16484,N_16927);
nor U20746 (N_20746,N_19488,N_16619);
and U20747 (N_20747,N_19187,N_16777);
nor U20748 (N_20748,N_17092,N_17777);
or U20749 (N_20749,N_19301,N_15751);
and U20750 (N_20750,N_15371,N_15170);
nor U20751 (N_20751,N_15873,N_15187);
or U20752 (N_20752,N_16314,N_17509);
and U20753 (N_20753,N_17059,N_18552);
xnor U20754 (N_20754,N_18212,N_18868);
and U20755 (N_20755,N_16213,N_17355);
or U20756 (N_20756,N_18535,N_15157);
xor U20757 (N_20757,N_18476,N_19693);
or U20758 (N_20758,N_15408,N_19385);
and U20759 (N_20759,N_15918,N_18486);
or U20760 (N_20760,N_16764,N_15102);
or U20761 (N_20761,N_15016,N_19732);
nor U20762 (N_20762,N_19140,N_16440);
and U20763 (N_20763,N_15390,N_18185);
and U20764 (N_20764,N_16162,N_15803);
or U20765 (N_20765,N_18386,N_15667);
nand U20766 (N_20766,N_17252,N_16180);
nor U20767 (N_20767,N_15035,N_17118);
or U20768 (N_20768,N_16870,N_18711);
nand U20769 (N_20769,N_15611,N_17817);
nor U20770 (N_20770,N_17220,N_15399);
or U20771 (N_20771,N_16470,N_19695);
nand U20772 (N_20772,N_18879,N_17587);
nand U20773 (N_20773,N_16452,N_15148);
and U20774 (N_20774,N_16799,N_16293);
nand U20775 (N_20775,N_18351,N_19721);
nand U20776 (N_20776,N_15627,N_18556);
and U20777 (N_20777,N_19626,N_18812);
and U20778 (N_20778,N_18044,N_17435);
or U20779 (N_20779,N_19774,N_15375);
and U20780 (N_20780,N_15055,N_18025);
xnor U20781 (N_20781,N_15111,N_19972);
nor U20782 (N_20782,N_17132,N_18450);
and U20783 (N_20783,N_17281,N_19276);
or U20784 (N_20784,N_19191,N_19880);
and U20785 (N_20785,N_19017,N_15722);
nand U20786 (N_20786,N_18544,N_19724);
nand U20787 (N_20787,N_15493,N_19992);
or U20788 (N_20788,N_17757,N_18161);
nand U20789 (N_20789,N_19389,N_16464);
and U20790 (N_20790,N_17606,N_16938);
and U20791 (N_20791,N_19991,N_18243);
nor U20792 (N_20792,N_18461,N_19372);
nor U20793 (N_20793,N_15400,N_17834);
and U20794 (N_20794,N_18004,N_17627);
and U20795 (N_20795,N_17113,N_18378);
or U20796 (N_20796,N_15207,N_15488);
and U20797 (N_20797,N_15957,N_15939);
or U20798 (N_20798,N_17605,N_15009);
or U20799 (N_20799,N_19815,N_16434);
and U20800 (N_20800,N_15420,N_16146);
and U20801 (N_20801,N_15930,N_18447);
or U20802 (N_20802,N_15347,N_15530);
nand U20803 (N_20803,N_15232,N_19006);
xnor U20804 (N_20804,N_15255,N_17288);
nor U20805 (N_20805,N_16740,N_15432);
nor U20806 (N_20806,N_17978,N_17607);
or U20807 (N_20807,N_17856,N_18917);
or U20808 (N_20808,N_15164,N_16968);
nand U20809 (N_20809,N_19943,N_16205);
or U20810 (N_20810,N_19951,N_19914);
and U20811 (N_20811,N_16097,N_16432);
and U20812 (N_20812,N_19246,N_15189);
or U20813 (N_20813,N_19518,N_18005);
nor U20814 (N_20814,N_19493,N_16246);
nor U20815 (N_20815,N_16602,N_16991);
and U20816 (N_20816,N_19857,N_17522);
nand U20817 (N_20817,N_18693,N_16819);
xor U20818 (N_20818,N_19465,N_16472);
nand U20819 (N_20819,N_18582,N_15132);
nor U20820 (N_20820,N_15135,N_15553);
nor U20821 (N_20821,N_19684,N_18274);
or U20822 (N_20822,N_15543,N_15128);
or U20823 (N_20823,N_18105,N_18953);
and U20824 (N_20824,N_17007,N_16793);
nand U20825 (N_20825,N_19883,N_15975);
nor U20826 (N_20826,N_16679,N_19858);
nor U20827 (N_20827,N_17064,N_18142);
nand U20828 (N_20828,N_15467,N_17167);
and U20829 (N_20829,N_16370,N_19784);
or U20830 (N_20830,N_15417,N_18371);
or U20831 (N_20831,N_18628,N_17880);
nor U20832 (N_20832,N_16308,N_15891);
nand U20833 (N_20833,N_19646,N_17382);
nor U20834 (N_20834,N_16717,N_17669);
nand U20835 (N_20835,N_17583,N_15393);
nor U20836 (N_20836,N_18758,N_16942);
nor U20837 (N_20837,N_18354,N_16396);
and U20838 (N_20838,N_17383,N_18887);
nand U20839 (N_20839,N_19413,N_17687);
nand U20840 (N_20840,N_15711,N_18175);
or U20841 (N_20841,N_18490,N_15633);
nand U20842 (N_20842,N_16237,N_15704);
or U20843 (N_20843,N_16868,N_16901);
nand U20844 (N_20844,N_16486,N_18057);
nor U20845 (N_20845,N_15201,N_18877);
nor U20846 (N_20846,N_15757,N_18816);
and U20847 (N_20847,N_19621,N_16482);
nand U20848 (N_20848,N_16200,N_17612);
xnor U20849 (N_20849,N_18046,N_15269);
nor U20850 (N_20850,N_19487,N_18100);
and U20851 (N_20851,N_19375,N_19655);
and U20852 (N_20852,N_16832,N_16557);
nand U20853 (N_20853,N_19542,N_16524);
or U20854 (N_20854,N_17705,N_18878);
nor U20855 (N_20855,N_19740,N_16090);
nand U20856 (N_20856,N_17456,N_18935);
and U20857 (N_20857,N_15641,N_19936);
nand U20858 (N_20858,N_18103,N_15701);
nor U20859 (N_20859,N_17251,N_17081);
nand U20860 (N_20860,N_16357,N_19414);
or U20861 (N_20861,N_17529,N_18191);
and U20862 (N_20862,N_15850,N_18362);
nor U20863 (N_20863,N_17507,N_19715);
nand U20864 (N_20864,N_18339,N_15289);
xor U20865 (N_20865,N_15217,N_19701);
nor U20866 (N_20866,N_18941,N_18002);
and U20867 (N_20867,N_17391,N_18633);
and U20868 (N_20868,N_19845,N_17094);
and U20869 (N_20869,N_18292,N_17772);
xnor U20870 (N_20870,N_15247,N_19408);
nor U20871 (N_20871,N_17524,N_16132);
or U20872 (N_20872,N_15921,N_16295);
nor U20873 (N_20873,N_18254,N_18201);
or U20874 (N_20874,N_15792,N_19674);
and U20875 (N_20875,N_16586,N_16944);
or U20876 (N_20876,N_18107,N_18998);
nand U20877 (N_20877,N_19353,N_18165);
nor U20878 (N_20878,N_18817,N_15394);
xor U20879 (N_20879,N_17148,N_15902);
xnor U20880 (N_20880,N_15596,N_15694);
or U20881 (N_20881,N_19905,N_17551);
or U20882 (N_20882,N_15522,N_16548);
nor U20883 (N_20883,N_18518,N_17835);
and U20884 (N_20884,N_17913,N_16721);
nor U20885 (N_20885,N_19233,N_18000);
nand U20886 (N_20886,N_15999,N_15802);
or U20887 (N_20887,N_16171,N_15949);
or U20888 (N_20888,N_17101,N_17658);
nor U20889 (N_20889,N_19429,N_16327);
nand U20890 (N_20890,N_18423,N_18838);
nand U20891 (N_20891,N_16616,N_18940);
and U20892 (N_20892,N_18394,N_18485);
or U20893 (N_20893,N_17824,N_16641);
or U20894 (N_20894,N_17564,N_15852);
nor U20895 (N_20895,N_15391,N_16599);
nand U20896 (N_20896,N_19111,N_17362);
xnor U20897 (N_20897,N_17591,N_18828);
and U20898 (N_20898,N_16027,N_19397);
and U20899 (N_20899,N_18847,N_17117);
nand U20900 (N_20900,N_15895,N_19261);
or U20901 (N_20901,N_19901,N_19591);
and U20902 (N_20902,N_15486,N_16920);
or U20903 (N_20903,N_17549,N_17327);
or U20904 (N_20904,N_18803,N_15771);
nor U20905 (N_20905,N_16453,N_19347);
nor U20906 (N_20906,N_19283,N_15585);
and U20907 (N_20907,N_15534,N_16053);
or U20908 (N_20908,N_18895,N_16822);
or U20909 (N_20909,N_19611,N_17781);
and U20910 (N_20910,N_18749,N_15492);
and U20911 (N_20911,N_18110,N_18857);
or U20912 (N_20912,N_16706,N_19221);
nand U20913 (N_20913,N_18063,N_16783);
and U20914 (N_20914,N_16185,N_18704);
and U20915 (N_20915,N_19062,N_17983);
or U20916 (N_20916,N_17621,N_19275);
nor U20917 (N_20917,N_17336,N_15047);
xnor U20918 (N_20918,N_16996,N_17922);
nand U20919 (N_20919,N_15359,N_19352);
xnor U20920 (N_20920,N_15638,N_16198);
and U20921 (N_20921,N_19234,N_17269);
nand U20922 (N_20922,N_15342,N_17654);
and U20923 (N_20923,N_18776,N_15348);
nand U20924 (N_20924,N_16573,N_17169);
or U20925 (N_20925,N_15384,N_15970);
xor U20926 (N_20926,N_15707,N_17875);
nor U20927 (N_20927,N_18705,N_16271);
and U20928 (N_20928,N_19367,N_15798);
and U20929 (N_20929,N_19181,N_15278);
or U20930 (N_20930,N_16129,N_15214);
and U20931 (N_20931,N_15262,N_19259);
nand U20932 (N_20932,N_17441,N_17994);
xnor U20933 (N_20933,N_17326,N_17230);
nor U20934 (N_20934,N_19672,N_18492);
or U20935 (N_20935,N_17432,N_18982);
nand U20936 (N_20936,N_16794,N_19496);
nor U20937 (N_20937,N_17107,N_18309);
nor U20938 (N_20938,N_17891,N_16892);
or U20939 (N_20939,N_15752,N_18688);
nand U20940 (N_20940,N_15218,N_15665);
or U20941 (N_20941,N_18660,N_15312);
or U20942 (N_20942,N_18830,N_17414);
or U20943 (N_20943,N_16292,N_16993);
xor U20944 (N_20944,N_17636,N_15082);
nor U20945 (N_20945,N_17820,N_16640);
xor U20946 (N_20946,N_17753,N_15376);
or U20947 (N_20947,N_17833,N_15012);
nand U20948 (N_20948,N_18216,N_15729);
xnor U20949 (N_20949,N_17803,N_16902);
nor U20950 (N_20950,N_18061,N_15357);
nor U20951 (N_20951,N_16251,N_16507);
nor U20952 (N_20952,N_16378,N_15679);
and U20953 (N_20953,N_18849,N_18522);
or U20954 (N_20954,N_17155,N_18984);
or U20955 (N_20955,N_15755,N_19679);
xnor U20956 (N_20956,N_15662,N_18180);
xor U20957 (N_20957,N_17256,N_18547);
or U20958 (N_20958,N_15051,N_16600);
xnor U20959 (N_20959,N_19381,N_17575);
nor U20960 (N_20960,N_17041,N_15366);
xor U20961 (N_20961,N_18396,N_15515);
or U20962 (N_20962,N_17109,N_19536);
and U20963 (N_20963,N_18258,N_18202);
nand U20964 (N_20964,N_17301,N_15640);
nor U20965 (N_20965,N_18564,N_15294);
xor U20966 (N_20966,N_15453,N_16742);
nor U20967 (N_20967,N_17295,N_19075);
and U20968 (N_20968,N_15607,N_15181);
and U20969 (N_20969,N_19902,N_16656);
nand U20970 (N_20970,N_17119,N_15449);
and U20971 (N_20971,N_15656,N_15300);
xnor U20972 (N_20972,N_15117,N_19472);
or U20973 (N_20973,N_18977,N_17205);
nor U20974 (N_20974,N_19173,N_16800);
xor U20975 (N_20975,N_16737,N_18433);
or U20976 (N_20976,N_19874,N_19336);
and U20977 (N_20977,N_18289,N_15907);
or U20978 (N_20978,N_15786,N_19583);
nor U20979 (N_20979,N_18479,N_19268);
xnor U20980 (N_20980,N_19436,N_15887);
and U20981 (N_20981,N_18475,N_17395);
or U20982 (N_20982,N_16739,N_15849);
nand U20983 (N_20983,N_19670,N_16500);
and U20984 (N_20984,N_18762,N_16770);
or U20985 (N_20985,N_17050,N_18430);
or U20986 (N_20986,N_17384,N_17958);
nor U20987 (N_20987,N_17552,N_17068);
and U20988 (N_20988,N_15735,N_17233);
nand U20989 (N_20989,N_19577,N_15295);
or U20990 (N_20990,N_17893,N_18546);
nor U20991 (N_20991,N_18592,N_17935);
and U20992 (N_20992,N_17925,N_15759);
nor U20993 (N_20993,N_18375,N_18440);
and U20994 (N_20994,N_18402,N_17207);
nand U20995 (N_20995,N_18072,N_15427);
or U20996 (N_20996,N_15306,N_18445);
nor U20997 (N_20997,N_18342,N_19160);
nor U20998 (N_20998,N_17238,N_18080);
xnor U20999 (N_20999,N_16366,N_15681);
xnor U21000 (N_21000,N_16921,N_18364);
or U21001 (N_21001,N_19299,N_19454);
nand U21002 (N_21002,N_15718,N_15225);
xor U21003 (N_21003,N_17929,N_17364);
nand U21004 (N_21004,N_17272,N_18790);
nor U21005 (N_21005,N_15720,N_18858);
nor U21006 (N_21006,N_15203,N_18796);
and U21007 (N_21007,N_15982,N_17954);
nor U21008 (N_21008,N_18332,N_15587);
and U21009 (N_21009,N_16790,N_18622);
nand U21010 (N_21010,N_18604,N_19470);
and U21011 (N_21011,N_16922,N_19522);
nor U21012 (N_21012,N_19478,N_19910);
or U21013 (N_21013,N_15863,N_19020);
or U21014 (N_21014,N_15027,N_18077);
or U21015 (N_21015,N_15458,N_15589);
nand U21016 (N_21016,N_16914,N_19506);
nand U21017 (N_21017,N_18503,N_18624);
nor U21018 (N_21018,N_18314,N_17723);
or U21019 (N_21019,N_19434,N_18345);
or U21020 (N_21020,N_18531,N_17685);
nand U21021 (N_21021,N_15118,N_17999);
nand U21022 (N_21022,N_17569,N_16285);
xnor U21023 (N_21023,N_19401,N_18200);
nand U21024 (N_21024,N_19202,N_17171);
nand U21025 (N_21025,N_19341,N_16865);
nand U21026 (N_21026,N_18909,N_19097);
nor U21027 (N_21027,N_16379,N_19747);
nor U21028 (N_21028,N_16607,N_18915);
or U21029 (N_21029,N_15966,N_18449);
nor U21030 (N_21030,N_16532,N_18923);
and U21031 (N_21031,N_17309,N_19325);
nand U21032 (N_21032,N_18715,N_19654);
nor U21033 (N_21033,N_16064,N_18023);
nand U21034 (N_21034,N_18244,N_15323);
or U21035 (N_21035,N_17375,N_19773);
nand U21036 (N_21036,N_16668,N_16376);
nor U21037 (N_21037,N_19805,N_19596);
nor U21038 (N_21038,N_17111,N_18966);
nand U21039 (N_21039,N_19290,N_17860);
xnor U21040 (N_21040,N_16990,N_16307);
xnor U21041 (N_21041,N_16552,N_15010);
nand U21042 (N_21042,N_15060,N_19263);
and U21043 (N_21043,N_16854,N_15972);
or U21044 (N_21044,N_18318,N_19157);
nand U21045 (N_21045,N_19214,N_18139);
nand U21046 (N_21046,N_15057,N_15463);
nand U21047 (N_21047,N_18525,N_15841);
nor U21048 (N_21048,N_16240,N_16490);
and U21049 (N_21049,N_17054,N_18121);
and U21050 (N_21050,N_19184,N_19462);
nand U21051 (N_21051,N_19581,N_16060);
nor U21052 (N_21052,N_16193,N_17286);
and U21053 (N_21053,N_19404,N_18337);
and U21054 (N_21054,N_17058,N_17070);
nand U21055 (N_21055,N_17579,N_17399);
xor U21056 (N_21056,N_17147,N_16645);
and U21057 (N_21057,N_16598,N_16394);
and U21058 (N_21058,N_15623,N_15220);
nand U21059 (N_21059,N_16435,N_18236);
nand U21060 (N_21060,N_16932,N_15993);
or U21061 (N_21061,N_16159,N_17574);
or U21062 (N_21062,N_16101,N_16593);
nand U21063 (N_21063,N_19293,N_16509);
nand U21064 (N_21064,N_15019,N_16710);
or U21065 (N_21065,N_19748,N_17844);
and U21066 (N_21066,N_18205,N_18901);
nor U21067 (N_21067,N_17434,N_15833);
or U21068 (N_21068,N_17407,N_18676);
nor U21069 (N_21069,N_16545,N_15746);
or U21070 (N_21070,N_15661,N_18238);
nor U21071 (N_21071,N_16046,N_16085);
nor U21072 (N_21072,N_19058,N_17847);
and U21073 (N_21073,N_15296,N_17802);
xnor U21074 (N_21074,N_18482,N_16811);
nor U21075 (N_21075,N_17638,N_16043);
or U21076 (N_21076,N_17280,N_18843);
nand U21077 (N_21077,N_18457,N_17332);
nor U21078 (N_21078,N_17899,N_16410);
nor U21079 (N_21079,N_19534,N_18415);
xnor U21080 (N_21080,N_16228,N_17790);
and U21081 (N_21081,N_17427,N_15338);
and U21082 (N_21082,N_15678,N_17603);
or U21083 (N_21083,N_19446,N_18446);
nand U21084 (N_21084,N_16852,N_15452);
nor U21085 (N_21085,N_18028,N_15810);
nor U21086 (N_21086,N_16893,N_15912);
and U21087 (N_21087,N_15484,N_19659);
and U21088 (N_21088,N_19521,N_18392);
nand U21089 (N_21089,N_15182,N_16128);
xor U21090 (N_21090,N_18198,N_16504);
nor U21091 (N_21091,N_18348,N_19009);
nor U21092 (N_21092,N_16576,N_17210);
and U21093 (N_21093,N_19253,N_18173);
nor U21094 (N_21094,N_18580,N_16020);
nand U21095 (N_21095,N_15107,N_19954);
and U21096 (N_21096,N_15659,N_15882);
nor U21097 (N_21097,N_15597,N_19406);
nand U21098 (N_21098,N_16274,N_18226);
and U21099 (N_21099,N_18881,N_16688);
xor U21100 (N_21100,N_17717,N_15699);
and U21101 (N_21101,N_18358,N_19036);
and U21102 (N_21102,N_15645,N_15556);
nor U21103 (N_21103,N_19977,N_16628);
or U21104 (N_21104,N_17216,N_19677);
nand U21105 (N_21105,N_15889,N_17246);
nor U21106 (N_21106,N_19963,N_18576);
nor U21107 (N_21107,N_18325,N_15369);
nand U21108 (N_21108,N_16642,N_15134);
nand U21109 (N_21109,N_17813,N_16157);
nand U21110 (N_21110,N_15120,N_17872);
xnor U21111 (N_21111,N_16372,N_17771);
and U21112 (N_21112,N_17047,N_19881);
nor U21113 (N_21113,N_18003,N_17547);
nand U21114 (N_21114,N_16803,N_17454);
or U21115 (N_21115,N_15353,N_16140);
or U21116 (N_21116,N_19313,N_16758);
or U21117 (N_21117,N_19909,N_19736);
nand U21118 (N_21118,N_15568,N_17350);
and U21119 (N_21119,N_18250,N_18429);
or U21120 (N_21120,N_15819,N_18561);
xor U21121 (N_21121,N_17096,N_18690);
or U21122 (N_21122,N_17245,N_17289);
nand U21123 (N_21123,N_17600,N_17415);
or U21124 (N_21124,N_18593,N_16502);
nor U21125 (N_21125,N_18381,N_17729);
nor U21126 (N_21126,N_15450,N_16188);
xor U21127 (N_21127,N_15431,N_16222);
or U21128 (N_21128,N_16297,N_19119);
nand U21129 (N_21129,N_17115,N_16791);
or U21130 (N_21130,N_16650,N_19163);
nand U21131 (N_21131,N_19461,N_18597);
or U21132 (N_21132,N_19279,N_16836);
and U21133 (N_21133,N_17885,N_18018);
nand U21134 (N_21134,N_15797,N_15011);
xor U21135 (N_21135,N_19737,N_18054);
nor U21136 (N_21136,N_15429,N_18012);
nor U21137 (N_21137,N_17648,N_15781);
nor U21138 (N_21138,N_17003,N_19971);
xor U21139 (N_21139,N_18831,N_15243);
xnor U21140 (N_21140,N_16277,N_17805);
and U21141 (N_21141,N_17469,N_15092);
xor U21142 (N_21142,N_16334,N_18751);
nor U21143 (N_21143,N_16276,N_16554);
nor U21144 (N_21144,N_19846,N_16449);
nor U21145 (N_21145,N_16150,N_15913);
nor U21146 (N_21146,N_16397,N_17916);
or U21147 (N_21147,N_15430,N_19274);
nor U21148 (N_21148,N_15651,N_19230);
nor U21149 (N_21149,N_19592,N_15790);
nand U21150 (N_21150,N_15498,N_17502);
xor U21151 (N_21151,N_15043,N_16473);
xor U21152 (N_21152,N_16163,N_16686);
nor U21153 (N_21153,N_15318,N_18632);
and U21154 (N_21154,N_19206,N_17348);
and U21155 (N_21155,N_18166,N_19808);
xor U21156 (N_21156,N_18300,N_18249);
and U21157 (N_21157,N_19678,N_16735);
nand U21158 (N_21158,N_18034,N_15447);
or U21159 (N_21159,N_19500,N_19767);
nand U21160 (N_21160,N_16131,N_18341);
nand U21161 (N_21161,N_15893,N_15693);
xor U21162 (N_21162,N_15570,N_15629);
nand U21163 (N_21163,N_18875,N_15094);
or U21164 (N_21164,N_18716,N_18976);
nor U21165 (N_21165,N_15334,N_19124);
nand U21166 (N_21166,N_16183,N_18296);
nor U21167 (N_21167,N_19447,N_18861);
nand U21168 (N_21168,N_19795,N_15758);
and U21169 (N_21169,N_18143,N_18463);
nor U21170 (N_21170,N_16048,N_18728);
nand U21171 (N_21171,N_18271,N_19938);
nor U21172 (N_21172,N_18265,N_18647);
nand U21173 (N_21173,N_17060,N_18218);
nand U21174 (N_21174,N_18569,N_15144);
and U21175 (N_21175,N_19266,N_16824);
nand U21176 (N_21176,N_19572,N_16818);
nand U21177 (N_21177,N_16958,N_19885);
nor U21178 (N_21178,N_17100,N_16597);
and U21179 (N_21179,N_18873,N_15248);
and U21180 (N_21180,N_15046,N_18154);
nand U21181 (N_21181,N_15500,N_17153);
xnor U21182 (N_21182,N_19185,N_19860);
and U21183 (N_21183,N_19754,N_15875);
nor U21184 (N_21184,N_18557,N_15688);
xor U21185 (N_21185,N_15698,N_15731);
or U21186 (N_21186,N_16444,N_19142);
nor U21187 (N_21187,N_18695,N_19840);
nand U21188 (N_21188,N_15834,N_16420);
and U21189 (N_21189,N_19778,N_17526);
xnor U21190 (N_21190,N_15917,N_18007);
xnor U21191 (N_21191,N_16847,N_19871);
nand U21192 (N_21192,N_17686,N_19046);
or U21193 (N_21193,N_16759,N_18193);
or U21194 (N_21194,N_17356,N_17349);
and U21195 (N_21195,N_19387,N_16982);
or U21196 (N_21196,N_19175,N_16025);
and U21197 (N_21197,N_18117,N_17232);
nor U21198 (N_21198,N_15045,N_15846);
nand U21199 (N_21199,N_16248,N_15451);
nand U21200 (N_21200,N_19571,N_17589);
xor U21201 (N_21201,N_16564,N_16054);
and U21202 (N_21202,N_15971,N_15286);
nand U21203 (N_21203,N_16328,N_16629);
nor U21204 (N_21204,N_16821,N_19594);
and U21205 (N_21205,N_16058,N_19994);
xor U21206 (N_21206,N_18666,N_18514);
or U21207 (N_21207,N_15812,N_17676);
and U21208 (N_21208,N_19509,N_19691);
and U21209 (N_21209,N_18702,N_19222);
xor U21210 (N_21210,N_16401,N_16166);
or U21211 (N_21211,N_16438,N_17213);
nand U21212 (N_21212,N_19550,N_18056);
and U21213 (N_21213,N_19063,N_16326);
or U21214 (N_21214,N_16626,N_19688);
and U21215 (N_21215,N_19034,N_15613);
nor U21216 (N_21216,N_17822,N_15683);
nand U21217 (N_21217,N_19172,N_19980);
and U21218 (N_21218,N_17260,N_19516);
or U21219 (N_21219,N_19380,N_15173);
nor U21220 (N_21220,N_19041,N_17702);
nor U21221 (N_21221,N_17886,N_19110);
xnor U21222 (N_21222,N_17186,N_19126);
nand U21223 (N_21223,N_17313,N_17934);
xnor U21224 (N_21224,N_17859,N_16138);
and U21225 (N_21225,N_19772,N_19824);
xnor U21226 (N_21226,N_16203,N_16639);
and U21227 (N_21227,N_18854,N_16577);
and U21228 (N_21228,N_17038,N_18060);
nor U21229 (N_21229,N_15230,N_17910);
or U21230 (N_21230,N_16634,N_17488);
and U21231 (N_21231,N_16696,N_17285);
nand U21232 (N_21232,N_15796,N_19143);
or U21233 (N_21233,N_17534,N_15624);
xnor U21234 (N_21234,N_17523,N_17539);
and U21235 (N_21235,N_18127,N_19681);
nor U21236 (N_21236,N_19782,N_17372);
nand U21237 (N_21237,N_18997,N_18744);
nand U21238 (N_21238,N_18171,N_19089);
and U21239 (N_21239,N_17263,N_18652);
nor U21240 (N_21240,N_18851,N_15204);
nor U21241 (N_21241,N_19345,N_15774);
nand U21242 (N_21242,N_17264,N_18483);
and U21243 (N_21243,N_19631,N_17966);
nor U21244 (N_21244,N_17410,N_19052);
nor U21245 (N_21245,N_19060,N_18509);
nand U21246 (N_21246,N_16514,N_16336);
nand U21247 (N_21247,N_18474,N_19931);
nor U21248 (N_21248,N_17413,N_16338);
or U21249 (N_21249,N_19080,N_19867);
nand U21250 (N_21250,N_19851,N_15410);
nand U21251 (N_21251,N_18787,N_19117);
nand U21252 (N_21252,N_19164,N_15555);
xnor U21253 (N_21253,N_19553,N_17192);
nor U21254 (N_21254,N_18090,N_19555);
nor U21255 (N_21255,N_18152,N_17738);
nor U21256 (N_21256,N_15156,N_19934);
nand U21257 (N_21257,N_17690,N_19159);
xor U21258 (N_21258,N_18527,N_19882);
xnor U21259 (N_21259,N_16807,N_19355);
or U21260 (N_21260,N_19130,N_17684);
and U21261 (N_21261,N_19376,N_15324);
xnor U21262 (N_21262,N_17404,N_18089);
and U21263 (N_21263,N_19974,N_19662);
nor U21264 (N_21264,N_15026,N_18432);
nand U21265 (N_21265,N_15241,N_16078);
xnor U21266 (N_21266,N_15657,N_18119);
and U21267 (N_21267,N_17537,N_17363);
and U21268 (N_21268,N_19177,N_17010);
nand U21269 (N_21269,N_19312,N_19658);
xnor U21270 (N_21270,N_18303,N_17645);
or U21271 (N_21271,N_19643,N_18886);
nor U21272 (N_21272,N_19145,N_16304);
and U21273 (N_21273,N_19809,N_16223);
nor U21274 (N_21274,N_19770,N_17066);
xnor U21275 (N_21275,N_19197,N_18845);
nor U21276 (N_21276,N_15310,N_18183);
nor U21277 (N_21277,N_19412,N_17075);
and U21278 (N_21278,N_19315,N_18684);
or U21279 (N_21279,N_19671,N_18609);
nand U21280 (N_21280,N_15581,N_18591);
or U21281 (N_21281,N_17718,N_19635);
nand U21282 (N_21282,N_15702,N_16526);
or U21283 (N_21283,N_19155,N_19955);
nand U21284 (N_21284,N_16864,N_18852);
and U21285 (N_21285,N_15246,N_16437);
or U21286 (N_21286,N_17325,N_16618);
nor U21287 (N_21287,N_17980,N_16867);
or U21288 (N_21288,N_15386,N_18298);
nor U21289 (N_21289,N_18278,N_19814);
or U21290 (N_21290,N_17623,N_19370);
xnor U21291 (N_21291,N_19494,N_18466);
or U21292 (N_21292,N_17227,N_19844);
nor U21293 (N_21293,N_16513,N_16387);
xor U21294 (N_21294,N_16382,N_18022);
nor U21295 (N_21295,N_18987,N_18155);
and U21296 (N_21296,N_19330,N_15036);
xor U21297 (N_21297,N_15178,N_15567);
nor U21298 (N_21298,N_15740,N_17378);
nor U21299 (N_21299,N_16894,N_16330);
nand U21300 (N_21300,N_18912,N_16859);
and U21301 (N_21301,N_18442,N_15539);
nand U21302 (N_21302,N_15544,N_19151);
or U21303 (N_21303,N_18156,N_17827);
nand U21304 (N_21304,N_15167,N_16041);
nand U21305 (N_21305,N_18619,N_15425);
or U21306 (N_21306,N_16383,N_17784);
nor U21307 (N_21307,N_19132,N_15590);
nand U21308 (N_21308,N_19575,N_18750);
and U21309 (N_21309,N_18841,N_17706);
and U21310 (N_21310,N_16817,N_19180);
or U21311 (N_21311,N_17228,N_18979);
nand U21312 (N_21312,N_15566,N_15436);
xnor U21313 (N_21313,N_15015,N_18867);
and U21314 (N_21314,N_18062,N_19444);
nor U21315 (N_21315,N_15297,N_18545);
nor U21316 (N_21316,N_16369,N_15532);
nand U21317 (N_21317,N_15005,N_19698);
or U21318 (N_21318,N_15783,N_18130);
nor U21319 (N_21319,N_15507,N_15565);
nor U21320 (N_21320,N_18823,N_15842);
nand U21321 (N_21321,N_17157,N_16747);
nor U21322 (N_21322,N_15229,N_19442);
or U21323 (N_21323,N_16627,N_16072);
xor U21324 (N_21324,N_16298,N_16267);
nor U21325 (N_21325,N_17595,N_15021);
nor U21326 (N_21326,N_15142,N_17769);
or U21327 (N_21327,N_18521,N_17940);
nand U21328 (N_21328,N_16480,N_18871);
nor U21329 (N_21329,N_17247,N_19527);
or U21330 (N_21330,N_18259,N_18839);
nor U21331 (N_21331,N_18764,N_19544);
nand U21332 (N_21332,N_18543,N_17773);
nand U21333 (N_21333,N_16063,N_15227);
and U21334 (N_21334,N_17530,N_19510);
and U21335 (N_21335,N_18093,N_15329);
nor U21336 (N_21336,N_18307,N_17809);
and U21337 (N_21337,N_19804,N_19899);
nand U21338 (N_21338,N_15428,N_17042);
and U21339 (N_21339,N_17248,N_19342);
and U21340 (N_21340,N_16838,N_18459);
xnor U21341 (N_21341,N_16199,N_19791);
nand U21342 (N_21342,N_16663,N_15175);
nor U21343 (N_21343,N_19590,N_17140);
nor U21344 (N_21344,N_15989,N_18439);
and U21345 (N_21345,N_17151,N_19714);
and U21346 (N_21346,N_16904,N_18973);
nand U21347 (N_21347,N_16361,N_19305);
nor U21348 (N_21348,N_19192,N_15388);
nand U21349 (N_21349,N_16018,N_18379);
or U21350 (N_21350,N_18742,N_17202);
or U21351 (N_21351,N_17946,N_16323);
and U21352 (N_21352,N_15032,N_17659);
and U21353 (N_21353,N_15086,N_17677);
nand U21354 (N_21354,N_18426,N_17836);
xnor U21355 (N_21355,N_15632,N_19912);
nand U21356 (N_21356,N_19131,N_17031);
and U21357 (N_21357,N_18727,N_18510);
and U21358 (N_21358,N_16069,N_17745);
nand U21359 (N_21359,N_17026,N_18752);
and U21360 (N_21360,N_18568,N_19623);
nor U21361 (N_21361,N_17631,N_16890);
or U21362 (N_21362,N_18323,N_19229);
nand U21363 (N_21363,N_16734,N_16943);
or U21364 (N_21364,N_16124,N_19668);
and U21365 (N_21365,N_19460,N_17473);
or U21366 (N_21366,N_15905,N_19597);
and U21367 (N_21367,N_15184,N_18308);
and U21368 (N_21368,N_17982,N_16196);
nor U21369 (N_21369,N_19490,N_15504);
and U21370 (N_21370,N_16903,N_19790);
and U21371 (N_21371,N_16281,N_18087);
and U21372 (N_21372,N_16506,N_17756);
and U21373 (N_21373,N_19120,N_17458);
nor U21374 (N_21374,N_19213,N_15499);
nand U21375 (N_21375,N_15482,N_17439);
nand U21376 (N_21376,N_17592,N_18734);
and U21377 (N_21377,N_15916,N_15676);
or U21378 (N_21378,N_16520,N_18095);
nor U21379 (N_21379,N_16630,N_17452);
or U21380 (N_21380,N_19165,N_19318);
nand U21381 (N_21381,N_18367,N_17792);
nand U21382 (N_21382,N_19973,N_18388);
or U21383 (N_21383,N_16546,N_19786);
and U21384 (N_21384,N_18159,N_18413);
nand U21385 (N_21385,N_16962,N_17029);
and U21386 (N_21386,N_15037,N_19114);
nand U21387 (N_21387,N_18427,N_18458);
nor U21388 (N_21388,N_19523,N_19825);
or U21389 (N_21389,N_16026,N_19660);
nor U21390 (N_21390,N_17311,N_15489);
nor U21391 (N_21391,N_16141,N_15328);
nand U21392 (N_21392,N_19254,N_19884);
xor U21393 (N_21393,N_19766,N_16543);
or U21394 (N_21394,N_19073,N_16125);
and U21395 (N_21395,N_18540,N_19326);
and U21396 (N_21396,N_17535,N_15202);
or U21397 (N_21397,N_16533,N_15251);
nor U21398 (N_21398,N_19570,N_19044);
or U21399 (N_21399,N_19587,N_18015);
nor U21400 (N_21400,N_16981,N_15136);
nand U21401 (N_21401,N_18897,N_15511);
and U21402 (N_21402,N_15407,N_16916);
and U21403 (N_21403,N_16911,N_18001);
nor U21404 (N_21404,N_19399,N_19686);
xnor U21405 (N_21405,N_18962,N_18211);
or U21406 (N_21406,N_16260,N_17221);
xor U21407 (N_21407,N_15747,N_16094);
nand U21408 (N_21408,N_15639,N_18383);
and U21409 (N_21409,N_15908,N_16647);
nor U21410 (N_21410,N_18994,N_16283);
nor U21411 (N_21411,N_17108,N_15847);
nor U21412 (N_21412,N_18021,N_15990);
nor U21413 (N_21413,N_16876,N_19302);
or U21414 (N_21414,N_16655,N_18729);
nor U21415 (N_21415,N_17217,N_16143);
or U21416 (N_21416,N_19944,N_17869);
nor U21417 (N_21417,N_19849,N_16515);
nand U21418 (N_21418,N_18636,N_18305);
and U21419 (N_21419,N_16621,N_16521);
and U21420 (N_21420,N_18390,N_15476);
nand U21421 (N_21421,N_19503,N_16364);
nor U21422 (N_21422,N_17419,N_16949);
xnor U21423 (N_21423,N_18682,N_18335);
or U21424 (N_21424,N_16844,N_16294);
nand U21425 (N_21425,N_19323,N_19666);
or U21426 (N_21426,N_17733,N_18078);
nor U21427 (N_21427,N_15285,N_15062);
nand U21428 (N_21428,N_18071,N_16221);
and U21429 (N_21429,N_19149,N_16574);
and U21430 (N_21430,N_17420,N_19480);
and U21431 (N_21431,N_18315,N_18374);
or U21432 (N_21432,N_15066,N_19217);
xor U21433 (N_21433,N_18380,N_17195);
and U21434 (N_21434,N_16834,N_15395);
and U21435 (N_21435,N_16711,N_17237);
nor U21436 (N_21436,N_18842,N_17436);
nor U21437 (N_21437,N_18153,N_19764);
nand U21438 (N_21438,N_16067,N_17428);
nand U21439 (N_21439,N_16359,N_16707);
xor U21440 (N_21440,N_17312,N_15373);
and U21441 (N_21441,N_18898,N_17316);
or U21442 (N_21442,N_19497,N_17588);
and U21443 (N_21443,N_17998,N_16145);
or U21444 (N_21444,N_16469,N_19297);
nand U21445 (N_21445,N_19728,N_16511);
and U21446 (N_21446,N_17040,N_17072);
and U21447 (N_21447,N_15006,N_16837);
and U21448 (N_21448,N_17849,N_15105);
nand U21449 (N_21449,N_17433,N_16989);
xor U21450 (N_21450,N_18691,N_18805);
and U21451 (N_21451,N_17477,N_15733);
and U21452 (N_21452,N_17173,N_16826);
or U21453 (N_21453,N_18232,N_19321);
or U21454 (N_21454,N_18195,N_15116);
nand U21455 (N_21455,N_18882,N_17125);
nand U21456 (N_21456,N_15806,N_19727);
or U21457 (N_21457,N_19081,N_18735);
or U21458 (N_21458,N_19289,N_15457);
or U21459 (N_21459,N_15048,N_16895);
and U21460 (N_21460,N_19826,N_15714);
or U21461 (N_21461,N_15750,N_18122);
nand U21462 (N_21462,N_15379,N_16692);
nand U21463 (N_21463,N_18853,N_16182);
and U21464 (N_21464,N_17580,N_17672);
xnor U21465 (N_21465,N_19360,N_17193);
nand U21466 (N_21466,N_17506,N_16139);
nor U21467 (N_21467,N_17577,N_19799);
xnor U21468 (N_21468,N_15535,N_17720);
nor U21469 (N_21469,N_17818,N_16805);
and U21470 (N_21470,N_18588,N_16368);
xnor U21471 (N_21471,N_15946,N_15415);
nor U21472 (N_21472,N_17907,N_19560);
nand U21473 (N_21473,N_19068,N_17649);
nor U21474 (N_21474,N_18104,N_18088);
nor U21475 (N_21475,N_16772,N_18670);
and U21476 (N_21476,N_16241,N_17968);
or U21477 (N_21477,N_16224,N_19369);
nor U21478 (N_21478,N_16268,N_16771);
xnor U21479 (N_21479,N_18366,N_18958);
and U21480 (N_21480,N_17374,N_16173);
nor U21481 (N_21481,N_16261,N_15967);
nor U21482 (N_21482,N_16007,N_17798);
nor U21483 (N_21483,N_15250,N_18837);
and U21484 (N_21484,N_18441,N_17293);
nor U21485 (N_21485,N_17466,N_19958);
xnor U21486 (N_21486,N_19231,N_15628);
nor U21487 (N_21487,N_19445,N_18772);
or U21488 (N_21488,N_16160,N_15199);
and U21489 (N_21489,N_15172,N_19832);
and U21490 (N_21490,N_19945,N_17315);
nor U21491 (N_21491,N_19526,N_17656);
or U21492 (N_21492,N_16358,N_16715);
or U21493 (N_21493,N_18497,N_16411);
or U21494 (N_21494,N_16167,N_18956);
and U21495 (N_21495,N_16108,N_15276);
or U21496 (N_21496,N_17297,N_16933);
and U21497 (N_21497,N_18157,N_15305);
xor U21498 (N_21498,N_15419,N_16135);
or U21499 (N_21499,N_17344,N_17218);
or U21500 (N_21500,N_19201,N_16936);
nor U21501 (N_21501,N_19300,N_19873);
or U21502 (N_21502,N_19354,N_19968);
nand U21503 (N_21503,N_18190,N_19529);
nand U21504 (N_21504,N_19324,N_15104);
nor U21505 (N_21505,N_19262,N_19453);
and U21506 (N_21506,N_17780,N_16303);
and U21507 (N_21507,N_15933,N_18075);
nor U21508 (N_21508,N_19074,N_16443);
nand U21509 (N_21509,N_18178,N_17970);
nor U21510 (N_21510,N_16536,N_16412);
and U21511 (N_21511,N_18538,N_15059);
nor U21512 (N_21512,N_18162,N_19183);
nor U21513 (N_21513,N_16848,N_19001);
or U21514 (N_21514,N_17986,N_15039);
nor U21515 (N_21515,N_17086,N_16363);
nand U21516 (N_21516,N_16365,N_17812);
and U21517 (N_21517,N_16508,N_18014);
and U21518 (N_21518,N_15228,N_18694);
nand U21519 (N_21519,N_17276,N_18301);
nor U21520 (N_21520,N_17421,N_17590);
nor U21521 (N_21521,N_18452,N_15935);
or U21522 (N_21522,N_15245,N_17527);
or U21523 (N_21523,N_18489,N_15112);
xnor U21524 (N_21524,N_18069,N_19449);
and U21525 (N_21525,N_18801,N_18981);
or U21526 (N_21526,N_18498,N_19964);
nor U21527 (N_21527,N_15837,N_17305);
xor U21528 (N_21528,N_18699,N_17422);
nand U21529 (N_21529,N_18453,N_17570);
nor U21530 (N_21530,N_18625,N_19532);
or U21531 (N_21531,N_17932,N_19043);
xnor U21532 (N_21532,N_15065,N_17212);
nand U21533 (N_21533,N_19665,N_19927);
and U21534 (N_21534,N_18295,N_19011);
nor U21535 (N_21535,N_18524,N_19236);
nor U21536 (N_21536,N_15090,N_19440);
xor U21537 (N_21537,N_16147,N_16210);
or U21538 (N_21538,N_15185,N_15259);
or U21539 (N_21539,N_18500,N_17962);
xnor U21540 (N_21540,N_16006,N_19077);
and U21541 (N_21541,N_16505,N_15068);
nor U21542 (N_21542,N_19199,N_15630);
and U21543 (N_21543,N_15079,N_19064);
or U21544 (N_21544,N_15508,N_16322);
nand U21545 (N_21545,N_16110,N_17542);
nor U21546 (N_21546,N_17025,N_15159);
or U21547 (N_21547,N_15612,N_16846);
and U21548 (N_21548,N_16559,N_17852);
nand U21549 (N_21549,N_16683,N_17129);
nor U21550 (N_21550,N_18995,N_15008);
nand U21551 (N_21551,N_16769,N_17832);
or U21552 (N_21552,N_18584,N_19409);
or U21553 (N_21553,N_15004,N_18773);
and U21554 (N_21554,N_16466,N_19735);
nand U21555 (N_21555,N_15552,N_18177);
nand U21556 (N_21556,N_15007,N_15301);
or U21557 (N_21557,N_15559,N_15387);
and U21558 (N_21558,N_18410,N_15927);
xnor U21559 (N_21559,N_19084,N_19435);
or U21560 (N_21560,N_15277,N_17845);
nor U21561 (N_21561,N_15948,N_15685);
and U21562 (N_21562,N_15053,N_15392);
xor U21563 (N_21563,N_17920,N_18930);
xnor U21564 (N_21564,N_15856,N_15145);
or U21565 (N_21565,N_15030,N_19812);
xnor U21566 (N_21566,N_19295,N_17303);
or U21567 (N_21567,N_18214,N_18248);
nand U21568 (N_21568,N_18723,N_18187);
or U21569 (N_21569,N_18280,N_16493);
xor U21570 (N_21570,N_16660,N_16494);
and U21571 (N_21571,N_19014,N_18257);
or U21572 (N_21572,N_18317,N_15293);
nand U21573 (N_21573,N_18602,N_19935);
nand U21574 (N_21574,N_17553,N_17797);
nor U21575 (N_21575,N_16899,N_15188);
nand U21576 (N_21576,N_15580,N_15421);
nor U21577 (N_21577,N_17495,N_16254);
and U21578 (N_21578,N_16151,N_16945);
nor U21579 (N_21579,N_16252,N_16768);
and U21580 (N_21580,N_17365,N_19614);
nor U21581 (N_21581,N_16485,N_17749);
or U21582 (N_21582,N_16860,N_15904);
and U21583 (N_21583,N_17278,N_16814);
nor U21584 (N_21584,N_17200,N_18276);
nor U21585 (N_21585,N_15536,N_17461);
and U21586 (N_21586,N_19153,N_16455);
and U21587 (N_21587,N_17721,N_19055);
or U21588 (N_21588,N_15211,N_17104);
nand U21589 (N_21589,N_16201,N_18506);
and U21590 (N_21590,N_17950,N_15465);
and U21591 (N_21591,N_15713,N_15708);
nand U21592 (N_21592,N_17357,N_16802);
or U21593 (N_21593,N_17799,N_15601);
and U21594 (N_21594,N_16673,N_15368);
and U21595 (N_21595,N_17159,N_18677);
nand U21596 (N_21596,N_15226,N_18434);
or U21597 (N_21597,N_15340,N_17057);
and U21598 (N_21598,N_18914,N_18907);
and U21599 (N_21599,N_15521,N_17273);
nand U21600 (N_21600,N_15978,N_17584);
nor U21601 (N_21601,N_15830,N_15818);
and U21602 (N_21602,N_16612,N_17562);
and U21603 (N_21603,N_16462,N_18903);
and U21604 (N_21604,N_15637,N_17794);
xnor U21605 (N_21605,N_19838,N_16289);
nor U21606 (N_21606,N_16137,N_17287);
nand U21607 (N_21607,N_15332,N_18058);
or U21608 (N_21608,N_17696,N_15671);
or U21609 (N_21609,N_18813,N_18501);
and U21610 (N_21610,N_15365,N_15518);
nand U21611 (N_21611,N_17719,N_16833);
or U21612 (N_21612,N_18209,N_18689);
and U21613 (N_21613,N_19777,N_18614);
nor U21614 (N_21614,N_15853,N_17339);
or U21615 (N_21615,N_15389,N_16136);
nor U21616 (N_21616,N_17519,N_17453);
nor U21617 (N_21617,N_19245,N_17651);
or U21618 (N_21618,N_17637,N_19339);
xnor U21619 (N_21619,N_19083,N_19392);
and U21620 (N_21620,N_19739,N_16775);
nor U21621 (N_21621,N_19627,N_16534);
nor U21622 (N_21622,N_19047,N_19280);
and U21623 (N_21623,N_16789,N_18313);
or U21624 (N_21624,N_19976,N_16445);
nand U21625 (N_21625,N_19170,N_19457);
nor U21626 (N_21626,N_19102,N_19198);
xor U21627 (N_21627,N_15883,N_19620);
xor U21628 (N_21628,N_19904,N_18559);
xnor U21629 (N_21629,N_18511,N_17639);
nand U21630 (N_21630,N_16258,N_16279);
and U21631 (N_21631,N_19495,N_19950);
or U21632 (N_21632,N_18123,N_16763);
nand U21633 (N_21633,N_16275,N_16291);
or U21634 (N_21634,N_16148,N_17044);
nand U21635 (N_21635,N_18902,N_15925);
xnor U21636 (N_21636,N_15424,N_17494);
or U21637 (N_21637,N_18355,N_18407);
and U21638 (N_21638,N_15726,N_18782);
nand U21639 (N_21639,N_15081,N_15001);
xnor U21640 (N_21640,N_16408,N_17062);
nand U21641 (N_21641,N_17985,N_19349);
nand U21642 (N_21642,N_15741,N_15050);
and U21643 (N_21643,N_16476,N_18932);
or U21644 (N_21644,N_17740,N_18896);
xnor U21645 (N_21645,N_19417,N_17479);
and U21646 (N_21646,N_18287,N_19716);
nor U21647 (N_21647,N_16930,N_15914);
and U21648 (N_21648,N_19129,N_18771);
nand U21649 (N_21649,N_19541,N_19319);
nand U21650 (N_21650,N_15541,N_19606);
xnor U21651 (N_21651,N_16057,N_18320);
xor U21652 (N_21652,N_18683,N_16635);
xnor U21653 (N_21653,N_19888,N_18589);
and U21654 (N_21654,N_17911,N_15859);
nand U21655 (N_21655,N_17006,N_19358);
and U21656 (N_21656,N_16570,N_16499);
and U21657 (N_21657,N_19196,N_17977);
nor U21658 (N_21658,N_18572,N_17873);
nand U21659 (N_21659,N_17661,N_19618);
nand U21660 (N_21660,N_16496,N_19535);
and U21661 (N_21661,N_16468,N_16975);
xnor U21662 (N_21662,N_18356,N_16266);
nand U21663 (N_21663,N_17091,N_15147);
or U21664 (N_21664,N_18565,N_15561);
xnor U21665 (N_21665,N_18186,N_15076);
or U21666 (N_21666,N_19984,N_18435);
nand U21667 (N_21667,N_17947,N_18267);
and U21668 (N_21668,N_16999,N_17628);
xnor U21669 (N_21669,N_16610,N_17296);
nand U21670 (N_21670,N_15067,N_18006);
xnor U21671 (N_21671,N_15973,N_18948);
nand U21672 (N_21672,N_19540,N_19983);
and U21673 (N_21673,N_17864,N_18468);
nor U21674 (N_21674,N_18208,N_19427);
and U21675 (N_21675,N_16835,N_16024);
and U21676 (N_21676,N_19135,N_16071);
or U21677 (N_21677,N_15677,N_17448);
xnor U21678 (N_21678,N_18844,N_16489);
nand U21679 (N_21679,N_15725,N_18607);
nor U21680 (N_21680,N_18737,N_16812);
or U21681 (N_21681,N_18169,N_17442);
nor U21682 (N_21682,N_16825,N_18224);
or U21683 (N_21683,N_16540,N_19792);
nor U21684 (N_21684,N_19520,N_17431);
or U21685 (N_21685,N_18347,N_19864);
nand U21686 (N_21686,N_19769,N_19410);
or U21687 (N_21687,N_17599,N_19697);
nand U21688 (N_21688,N_15138,N_18027);
or U21689 (N_21689,N_18736,N_17449);
and U21690 (N_21690,N_17163,N_18548);
nor U21691 (N_21691,N_19390,N_17443);
nor U21692 (N_21692,N_17883,N_17747);
and U21693 (N_21693,N_19029,N_19763);
and U21694 (N_21694,N_17402,N_18646);
nand U21695 (N_21695,N_15414,N_17189);
nor U21696 (N_21696,N_17843,N_19999);
nand U21697 (N_21697,N_18469,N_19997);
xnor U21698 (N_21698,N_15054,N_16016);
and U21699 (N_21699,N_19441,N_18302);
nand U21700 (N_21700,N_19291,N_17020);
and U21701 (N_21701,N_16351,N_16154);
nand U21702 (N_21702,N_18937,N_18795);
and U21703 (N_21703,N_17548,N_17640);
and U21704 (N_21704,N_15680,N_16596);
nor U21705 (N_21705,N_19758,N_15997);
or U21706 (N_21706,N_18745,N_15923);
nor U21707 (N_21707,N_16840,N_16516);
and U21708 (N_21708,N_19514,N_18999);
nand U21709 (N_21709,N_19752,N_16827);
xnor U21710 (N_21710,N_18352,N_17351);
nor U21711 (N_21711,N_19070,N_18566);
xnor U21712 (N_21712,N_16264,N_18227);
nor U21713 (N_21713,N_18291,N_16594);
or U21714 (N_21714,N_16008,N_19455);
nand U21715 (N_21715,N_16556,N_16823);
nor U21716 (N_21716,N_18732,N_18819);
or U21717 (N_21717,N_19531,N_17752);
and U21718 (N_21718,N_16414,N_15644);
nand U21719 (N_21719,N_19486,N_16421);
nor U21720 (N_21720,N_17199,N_16463);
nor U21721 (N_21721,N_17131,N_18032);
xor U21722 (N_21722,N_19139,N_19918);
nor U21723 (N_21723,N_15287,N_17987);
nand U21724 (N_21724,N_17851,N_16888);
and U21725 (N_21725,N_15584,N_15745);
nor U21726 (N_21726,N_16288,N_19264);
nor U21727 (N_21727,N_15355,N_17211);
and U21728 (N_21728,N_16035,N_17734);
or U21729 (N_21729,N_17130,N_18408);
xor U21730 (N_21730,N_15666,N_19115);
xnor U21731 (N_21731,N_19072,N_15234);
and U21732 (N_21732,N_16415,N_15291);
nand U21733 (N_21733,N_19990,N_18950);
and U21734 (N_21734,N_17037,N_18686);
nor U21735 (N_21735,N_17611,N_17541);
nor U21736 (N_21736,N_17012,N_17963);
nand U21737 (N_21737,N_19760,N_15069);
nor U21738 (N_21738,N_18111,N_18615);
xor U21739 (N_21739,N_18404,N_16302);
nand U21740 (N_21740,N_18017,N_16340);
nor U21741 (N_21741,N_16808,N_15426);
or U21742 (N_21742,N_15855,N_18239);
and U21743 (N_21743,N_19744,N_15866);
or U21744 (N_21744,N_18671,N_17779);
and U21745 (N_21745,N_17401,N_17302);
nor U21746 (N_21746,N_19092,N_17317);
xnor U21747 (N_21747,N_16820,N_17867);
nand U21748 (N_21748,N_15828,N_18738);
or U21749 (N_21749,N_18974,N_15823);
xnor U21750 (N_21750,N_19551,N_16935);
nand U21751 (N_21751,N_15313,N_16087);
or U21752 (N_21752,N_15398,N_18039);
and U21753 (N_21753,N_15636,N_16431);
or U21754 (N_21754,N_17008,N_16104);
and U21755 (N_21755,N_15468,N_19568);
nor U21756 (N_21756,N_19949,N_15274);
and U21757 (N_21757,N_15943,N_16580);
or U21758 (N_21758,N_17576,N_17828);
and U21759 (N_21759,N_17039,N_16454);
xor U21760 (N_21760,N_19704,N_17744);
and U21761 (N_21761,N_16044,N_16236);
or U21762 (N_21762,N_18020,N_16344);
xnor U21763 (N_21763,N_17114,N_18791);
xor U21764 (N_21764,N_17242,N_17408);
xor U21765 (N_21765,N_15261,N_19270);
and U21766 (N_21766,N_15115,N_15437);
nand U21767 (N_21767,N_17013,N_16675);
nor U21768 (N_21768,N_16385,N_17368);
nor U21769 (N_21769,N_15233,N_16806);
and U21770 (N_21770,N_19924,N_19817);
or U21771 (N_21771,N_16374,N_15074);
or U21772 (N_21772,N_19007,N_18097);
or U21773 (N_21773,N_17614,N_17124);
nand U21774 (N_21774,N_17377,N_15936);
nor U21775 (N_21775,N_18645,N_16217);
or U21776 (N_21776,N_19803,N_17511);
nand U21777 (N_21777,N_16702,N_16527);
nor U21778 (N_21778,N_19843,N_17514);
or U21779 (N_21779,N_19913,N_18634);
or U21780 (N_21780,N_18189,N_16377);
nand U21781 (N_21781,N_16780,N_15727);
or U21782 (N_21782,N_19365,N_17343);
xnor U21783 (N_21783,N_16631,N_18207);
or U21784 (N_21784,N_16239,N_16845);
nand U21785 (N_21785,N_15177,N_19049);
or U21786 (N_21786,N_18574,N_15171);
nor U21787 (N_21787,N_17184,N_15782);
xnor U21788 (N_21788,N_18904,N_15703);
nor U21789 (N_21789,N_19878,N_17641);
and U21790 (N_21790,N_17380,N_15562);
or U21791 (N_21791,N_15922,N_18687);
and U21792 (N_21792,N_17045,N_18554);
and U21793 (N_21793,N_19915,N_18784);
nor U21794 (N_21794,N_19273,N_17879);
and U21795 (N_21795,N_16831,N_16544);
nand U21796 (N_21796,N_19726,N_18436);
nand U21797 (N_21797,N_19552,N_15600);
or U21798 (N_21798,N_16441,N_15506);
nand U21799 (N_21799,N_15479,N_17106);
or U21800 (N_21800,N_18884,N_16153);
and U21801 (N_21801,N_18668,N_16866);
or U21802 (N_21802,N_15761,N_17975);
nand U21803 (N_21803,N_15945,N_17622);
xnor U21804 (N_21804,N_17178,N_19908);
and U21805 (N_21805,N_18856,N_18016);
nor U21806 (N_21806,N_19530,N_16889);
xor U21807 (N_21807,N_15327,N_18692);
or U21808 (N_21808,N_17393,N_19757);
xnor U21809 (N_21809,N_17398,N_15003);
and U21810 (N_21810,N_17353,N_16422);
nor U21811 (N_21811,N_17187,N_19651);
and U21812 (N_21812,N_19539,N_16475);
nand U21813 (N_21813,N_16722,N_16858);
nor U21814 (N_21814,N_16234,N_16030);
or U21815 (N_21815,N_19396,N_16753);
and U21816 (N_21816,N_15349,N_18182);
xnor U21817 (N_21817,N_19076,N_19466);
xor U21818 (N_21818,N_19458,N_17396);
xnor U21819 (N_21819,N_15557,N_15770);
and U21820 (N_21820,N_15762,N_17560);
nand U21821 (N_21821,N_17249,N_19630);
nand U21822 (N_21822,N_19239,N_15056);
nand U21823 (N_21823,N_19316,N_15018);
or U21824 (N_21824,N_16565,N_17943);
nand U21825 (N_21825,N_19690,N_18074);
nand U21826 (N_21826,N_15528,N_17751);
nand U21827 (N_21827,N_15525,N_16960);
xnor U21828 (N_21828,N_18972,N_18241);
nor U21829 (N_21829,N_17470,N_17760);
or U21830 (N_21830,N_17016,N_18416);
xnor U21831 (N_21831,N_18467,N_15083);
nand U21832 (N_21832,N_18864,N_18573);
or U21833 (N_21833,N_19123,N_16112);
and U21834 (N_21834,N_16575,N_18834);
or U21835 (N_21835,N_15114,N_15158);
xor U21836 (N_21836,N_19957,N_18859);
nand U21837 (N_21837,N_17842,N_16581);
and U21838 (N_21838,N_18810,N_15298);
or U21839 (N_21839,N_18863,N_15648);
and U21840 (N_21840,N_15598,N_16719);
or U21841 (N_21841,N_17714,N_18499);
nand U21842 (N_21842,N_17518,N_18399);
nor U21843 (N_21843,N_17181,N_17764);
or U21844 (N_21844,N_19647,N_15888);
or U21845 (N_21845,N_17634,N_17493);
or U21846 (N_21846,N_18659,N_15377);
and U21847 (N_21847,N_16701,N_19593);
nor U21848 (N_21848,N_19869,N_15867);
and U21849 (N_21849,N_17177,N_19524);
nand U21850 (N_21850,N_17275,N_19517);
nand U21851 (N_21851,N_19492,N_18581);
nand U21852 (N_21852,N_18654,N_19252);
nor U21853 (N_21853,N_16189,N_15113);
xor U21854 (N_21854,N_19216,N_19827);
xnor U21855 (N_21855,N_18719,N_19939);
xnor U21856 (N_21856,N_19294,N_18644);
nor U21857 (N_21857,N_18136,N_18405);
nor U21858 (N_21858,N_19016,N_16728);
nor U21859 (N_21859,N_16558,N_15813);
nor U21860 (N_21860,N_18417,N_18228);
and U21861 (N_21861,N_17855,N_19889);
nor U21862 (N_21862,N_18541,N_16031);
or U21863 (N_21863,N_17806,N_18285);
nor U21864 (N_21864,N_17732,N_18532);
nor U21865 (N_21865,N_16501,N_15928);
and U21866 (N_21866,N_17261,N_16815);
or U21867 (N_21867,N_16211,N_15865);
and U21868 (N_21868,N_17837,N_17892);
and U21869 (N_21869,N_18409,N_15095);
or U21870 (N_21870,N_18210,N_16954);
nand U21871 (N_21871,N_18883,N_15896);
nor U21872 (N_21872,N_15756,N_18957);
nor U21873 (N_21873,N_17801,N_19600);
or U21874 (N_21874,N_16849,N_18558);
nand U21875 (N_21875,N_19928,N_16528);
nand U21876 (N_21876,N_17485,N_18708);
and U21877 (N_21877,N_15995,N_17884);
or U21878 (N_21878,N_19241,N_17632);
nand U21879 (N_21879,N_16553,N_17937);
nor U21880 (N_21880,N_17775,N_16178);
xnor U21881 (N_21881,N_19430,N_15827);
nor U21882 (N_21882,N_17080,N_16341);
or U21883 (N_21883,N_15817,N_15221);
nor U21884 (N_21884,N_19484,N_16492);
nand U21885 (N_21885,N_15821,N_15440);
nand U21886 (N_21886,N_15242,N_16005);
nand U21887 (N_21887,N_15495,N_19680);
and U21888 (N_21888,N_17065,N_18804);
nand U21889 (N_21889,N_19661,N_18848);
or U21890 (N_21890,N_19468,N_15279);
nor U21891 (N_21891,N_18030,N_15196);
and U21892 (N_21892,N_17635,N_15804);
and U21893 (N_21893,N_15654,N_15658);
or U21894 (N_21894,N_16065,N_15381);
nand U21895 (N_21895,N_16804,N_18667);
or U21896 (N_21896,N_19818,N_16367);
and U21897 (N_21897,N_16400,N_15413);
nand U21898 (N_21898,N_17346,N_18549);
nor U21899 (N_21899,N_19664,N_15176);
nand U21900 (N_21900,N_17426,N_17437);
and U21901 (N_21901,N_17895,N_19481);
and U21902 (N_21902,N_15149,N_17902);
nor U21903 (N_21903,N_18491,N_17988);
nand U21904 (N_21904,N_18799,N_19887);
nand U21905 (N_21905,N_19346,N_18612);
and U21906 (N_21906,N_17467,N_18513);
and U21907 (N_21907,N_16569,N_17021);
xnor U21908 (N_21908,N_17498,N_16013);
xor U21909 (N_21909,N_16869,N_16850);
and U21910 (N_21910,N_15235,N_15087);
nor U21911 (N_21911,N_16913,N_19189);
or U21912 (N_21912,N_17244,N_16115);
or U21913 (N_21913,N_15926,N_18256);
or U21914 (N_21914,N_17462,N_16373);
or U21915 (N_21915,N_17613,N_15996);
nor U21916 (N_21916,N_17971,N_16995);
or U21917 (N_21917,N_19853,N_17329);
and U21918 (N_21918,N_18406,N_17581);
and U21919 (N_21919,N_16096,N_18140);
nand U21920 (N_21920,N_17240,N_15697);
nand U21921 (N_21921,N_16012,N_16331);
or U21922 (N_21922,N_15237,N_18338);
nand U21923 (N_21923,N_19948,N_18637);
or U21924 (N_21924,N_19477,N_15333);
nand U21925 (N_21925,N_16724,N_19942);
nand U21926 (N_21926,N_16585,N_16720);
xnor U21927 (N_21927,N_15897,N_18393);
nor U21928 (N_21928,N_18242,N_16674);
xor U21929 (N_21929,N_15588,N_17646);
xnor U21930 (N_21930,N_15146,N_17917);
or U21931 (N_21931,N_19223,N_16774);
nand U21932 (N_21932,N_16680,N_18921);
or U21933 (N_21933,N_16447,N_15977);
nor U21934 (N_21934,N_19652,N_15165);
or U21935 (N_21935,N_17459,N_17358);
and U21936 (N_21936,N_17566,N_18832);
and U21937 (N_21937,N_16111,N_19911);
or U21938 (N_21938,N_19865,N_18083);
or U21939 (N_21939,N_19891,N_15533);
and U21940 (N_21940,N_15208,N_19310);
or U21941 (N_21941,N_15073,N_18989);
or U21942 (N_21942,N_18595,N_15931);
nand U21943 (N_21943,N_16320,N_18411);
and U21944 (N_21944,N_19498,N_19104);
nand U21945 (N_21945,N_16315,N_18008);
xor U21946 (N_21946,N_19103,N_15924);
nor U21947 (N_21947,N_16299,N_18220);
xor U21948 (N_21948,N_19296,N_15712);
nor U21949 (N_21949,N_16142,N_18600);
nand U21950 (N_21950,N_16250,N_18757);
nand U21951 (N_21951,N_19893,N_17909);
nor U21952 (N_21952,N_16325,N_17735);
xnor U21953 (N_21953,N_17865,N_15540);
nor U21954 (N_21954,N_15560,N_19366);
nand U21955 (N_21955,N_19602,N_17900);
or U21956 (N_21956,N_16709,N_15272);
nand U21957 (N_21957,N_19923,N_16197);
nand U21958 (N_21958,N_16946,N_19027);
and U21959 (N_21959,N_17841,N_19673);
and U21960 (N_21960,N_17655,N_17561);
or U21961 (N_21961,N_17103,N_16152);
and U21962 (N_21962,N_16038,N_15788);
nand U21963 (N_21963,N_18064,N_16062);
nand U21964 (N_21964,N_15958,N_15103);
nand U21965 (N_21965,N_16227,N_18945);
or U21966 (N_21966,N_17598,N_19848);
nor U21967 (N_21967,N_15573,N_16156);
nor U21968 (N_21968,N_19051,N_16247);
or U21969 (N_21969,N_18163,N_19035);
xor U21970 (N_21970,N_19138,N_16700);
or U21971 (N_21971,N_16386,N_18717);
xor U21972 (N_21972,N_16563,N_16589);
or U21973 (N_21973,N_19616,N_16795);
nor U21974 (N_21974,N_16133,N_19850);
and U21975 (N_21975,N_18403,N_17984);
and U21976 (N_21976,N_15268,N_17829);
and U21977 (N_21977,N_19636,N_17194);
nand U21978 (N_21978,N_16347,N_17693);
or U21979 (N_21979,N_19879,N_19667);
or U21980 (N_21980,N_17497,N_15919);
nor U21981 (N_21981,N_16966,N_16272);
or U21982 (N_21982,N_17956,N_18197);
and U21983 (N_21983,N_17938,N_16418);
and U21984 (N_21984,N_15382,N_19168);
nor U21985 (N_21985,N_18768,N_19533);
xnor U21986 (N_21986,N_19338,N_17870);
or U21987 (N_21987,N_16390,N_18754);
nand U21988 (N_21988,N_18780,N_18890);
nand U21989 (N_21989,N_16192,N_18806);
or U21990 (N_21990,N_16333,N_17320);
and U21991 (N_21991,N_16184,N_19045);
nor U21992 (N_21992,N_17630,N_17142);
or U21993 (N_21993,N_17253,N_17381);
nand U21994 (N_21994,N_19967,N_16273);
and U21995 (N_21995,N_17763,N_16169);
nand U21996 (N_21996,N_19797,N_18343);
nand U21997 (N_21997,N_17176,N_16497);
nand U21998 (N_21998,N_17201,N_18247);
nand U21999 (N_21999,N_17416,N_15569);
and U22000 (N_22000,N_16231,N_18880);
xor U22001 (N_22001,N_15385,N_19057);
and U22002 (N_22002,N_18359,N_17340);
and U22003 (N_22003,N_19842,N_17750);
nor U22004 (N_22004,N_19228,N_17887);
nand U22005 (N_22005,N_19624,N_15363);
or U22006 (N_22006,N_18785,N_15174);
nand U22007 (N_22007,N_15271,N_17342);
or U22008 (N_22008,N_19608,N_15900);
xnor U22009 (N_22009,N_18971,N_15517);
nand U22010 (N_22010,N_18814,N_19582);
nor U22011 (N_22011,N_16280,N_18170);
nor U22012 (N_22012,N_16105,N_18324);
and U22013 (N_22013,N_17009,N_15023);
or U22014 (N_22014,N_15862,N_15682);
nor U22015 (N_22015,N_17389,N_18571);
nor U22016 (N_22016,N_15838,N_18336);
nand U22017 (N_22017,N_16233,N_16491);
or U22018 (N_22018,N_15835,N_17746);
nor U22019 (N_22019,N_19431,N_18050);
nor U22020 (N_22020,N_18594,N_17823);
nor U22021 (N_22021,N_16531,N_17953);
nand U22022 (N_22022,N_16074,N_18109);
nor U22023 (N_22023,N_16255,N_19508);
nand U22024 (N_22024,N_16290,N_17425);
nand U22025 (N_22025,N_17304,N_16649);
and U22026 (N_22026,N_17017,N_16730);
nor U22027 (N_22027,N_18627,N_19499);
or U22028 (N_22028,N_19762,N_15124);
nor U22029 (N_22029,N_19965,N_17444);
xor U22030 (N_22030,N_18477,N_16406);
nand U22031 (N_22031,N_16045,N_16978);
xor U22032 (N_22032,N_15362,N_17366);
nand U22033 (N_22033,N_18993,N_18515);
nor U22034 (N_22034,N_19834,N_19859);
or U22035 (N_22035,N_16878,N_17996);
nor U22036 (N_22036,N_18740,N_17028);
nor U22037 (N_22037,N_17002,N_19452);
and U22038 (N_22038,N_17135,N_15974);
nor U22039 (N_22039,N_18721,N_15634);
or U22040 (N_22040,N_18067,N_17927);
xnor U22041 (N_22041,N_16413,N_15153);
nand U22042 (N_22042,N_19469,N_18550);
or U22043 (N_22043,N_18038,N_18344);
and U22044 (N_22044,N_16175,N_16243);
nand U22045 (N_22045,N_18655,N_19383);
xor U22046 (N_22046,N_15549,N_15239);
and U22047 (N_22047,N_19584,N_19687);
xor U22048 (N_22048,N_16483,N_18739);
xor U22049 (N_22049,N_19287,N_15316);
and U22050 (N_22050,N_15319,N_17830);
and U22051 (N_22051,N_16164,N_15724);
nor U22052 (N_22052,N_19288,N_15510);
or U22053 (N_22053,N_15546,N_17568);
or U22054 (N_22054,N_15808,N_17474);
xor U22055 (N_22055,N_19835,N_16637);
nor U22056 (N_22056,N_16671,N_19925);
or U22057 (N_22057,N_17650,N_18770);
or U22058 (N_22058,N_15180,N_17208);
and U22059 (N_22059,N_19416,N_19250);
and U22060 (N_22060,N_16773,N_17386);
nand U22061 (N_22061,N_18235,N_19195);
or U22062 (N_22062,N_18933,N_19730);
nor U22063 (N_22063,N_16118,N_17082);
or U22064 (N_22064,N_16471,N_16477);
xnor U22065 (N_22065,N_16503,N_18822);
or U22066 (N_22066,N_15650,N_16880);
or U22067 (N_22067,N_18222,N_18456);
nand U22068 (N_22068,N_15709,N_15224);
xor U22069 (N_22069,N_19156,N_19350);
and U22070 (N_22070,N_19395,N_18377);
nand U22071 (N_22071,N_15396,N_19645);
nor U22072 (N_22072,N_19271,N_17223);
nor U22073 (N_22073,N_15890,N_17919);
nand U22074 (N_22074,N_17905,N_18079);
nand U22075 (N_22075,N_17492,N_18990);
nor U22076 (N_22076,N_19256,N_19755);
nor U22077 (N_22077,N_15558,N_16207);
nand U22078 (N_22078,N_16997,N_19785);
and U22079 (N_22079,N_16047,N_16937);
or U22080 (N_22080,N_17668,N_15042);
or U22081 (N_22081,N_15617,N_16625);
or U22082 (N_22082,N_15538,N_18949);
and U22083 (N_22083,N_15848,N_16687);
and U22084 (N_22084,N_19746,N_19306);
or U22085 (N_22085,N_17034,N_16994);
nor U22086 (N_22086,N_19393,N_15526);
nor U22087 (N_22087,N_18070,N_16042);
or U22088 (N_22088,N_17482,N_16119);
nor U22089 (N_22089,N_16908,N_18943);
and U22090 (N_22090,N_18268,N_19689);
nor U22091 (N_22091,N_15572,N_15675);
and U22092 (N_22092,N_18946,N_18794);
nor U22093 (N_22093,N_16343,N_16755);
nor U22094 (N_22094,N_19003,N_18462);
and U22095 (N_22095,N_17992,N_17359);
nand U22096 (N_22096,N_19941,N_18372);
xnor U22097 (N_22097,N_16887,N_16929);
nand U22098 (N_22098,N_18246,N_17001);
and U22099 (N_22099,N_18275,N_16941);
nor U22100 (N_22100,N_19653,N_16952);
nand U22101 (N_22101,N_16081,N_16624);
and U22102 (N_22102,N_17319,N_19629);
nor U22103 (N_22103,N_15728,N_19067);
or U22104 (N_22104,N_16924,N_17250);
and U22105 (N_22105,N_17265,N_18010);
nand U22106 (N_22106,N_16375,N_19694);
nand U22107 (N_22107,N_18026,N_19320);
and U22108 (N_22108,N_16174,N_18454);
nand U22109 (N_22109,N_17807,N_16229);
or U22110 (N_22110,N_19186,N_15616);
or U22111 (N_22111,N_16766,N_18815);
or U22112 (N_22112,N_19432,N_15496);
or U22113 (N_22113,N_15799,N_16784);
and U22114 (N_22114,N_15775,N_17868);
nor U22115 (N_22115,N_16905,N_16478);
xor U22116 (N_22116,N_17403,N_15474);
and U22117 (N_22117,N_16761,N_16427);
and U22118 (N_22118,N_17675,N_16828);
nand U22119 (N_22119,N_19601,N_18059);
nand U22120 (N_22120,N_18931,N_16032);
and U22121 (N_22121,N_18798,N_15674);
nor U22122 (N_22122,N_18952,N_16875);
xnor U22123 (N_22123,N_18349,N_17914);
xnor U22124 (N_22124,N_16917,N_19981);
nand U22125 (N_22125,N_18939,N_15025);
nand U22126 (N_22126,N_17597,N_15687);
or U22127 (N_22127,N_15257,N_18151);
nand U22128 (N_22128,N_18134,N_17674);
nand U22129 (N_22129,N_17513,N_15412);
and U22130 (N_22130,N_16403,N_19561);
and U22131 (N_22131,N_15626,N_15870);
nor U22132 (N_22132,N_16068,N_19952);
nand U22133 (N_22133,N_17465,N_19978);
nor U22134 (N_22134,N_15840,N_16028);
and U22135 (N_22135,N_16165,N_18631);
xor U22136 (N_22136,N_16959,N_18470);
xor U22137 (N_22137,N_19005,N_18495);
nor U22138 (N_22138,N_17112,N_15106);
nand U22139 (N_22139,N_16075,N_16657);
nor U22140 (N_22140,N_17093,N_19398);
nand U22141 (N_22141,N_19642,N_17839);
or U22142 (N_22142,N_19154,N_18421);
nand U22143 (N_22143,N_16788,N_16681);
and U22144 (N_22144,N_19705,N_18696);
or U22145 (N_22145,N_15836,N_16319);
and U22146 (N_22146,N_18603,N_19368);
or U22147 (N_22147,N_19573,N_16459);
nor U22148 (N_22148,N_16654,N_15364);
xnor U22149 (N_22149,N_18231,N_18288);
nor U22150 (N_22150,N_15192,N_15537);
and U22151 (N_22151,N_18329,N_19141);
nand U22152 (N_22152,N_15779,N_18906);
xor U22153 (N_22153,N_16116,N_18947);
nor U22154 (N_22154,N_19970,N_16371);
nor U22155 (N_22155,N_19218,N_18048);
or U22156 (N_22156,N_19586,N_15302);
and U22157 (N_22157,N_16313,N_15992);
nor U22158 (N_22158,N_18533,N_15485);
and U22159 (N_22159,N_17700,N_18888);
nand U22160 (N_22160,N_19605,N_18245);
nor U22161 (N_22161,N_17496,N_18954);
and U22162 (N_22162,N_16542,N_19190);
and U22163 (N_22163,N_15089,N_17670);
or U22164 (N_22164,N_17241,N_19400);
xor U22165 (N_22165,N_18272,N_16669);
nor U22166 (N_22166,N_19578,N_15876);
or U22167 (N_22167,N_19877,N_19113);
nand U22168 (N_22168,N_17412,N_17259);
nand U22169 (N_22169,N_16134,N_19479);
nand U22170 (N_22170,N_17283,N_16195);
or U22171 (N_22171,N_18092,N_17324);
and U22172 (N_22172,N_18537,N_17846);
and U22173 (N_22173,N_16353,N_18765);
and U22174 (N_22174,N_15869,N_15434);
nand U22175 (N_22175,N_18703,N_19669);
nand U22176 (N_22176,N_15605,N_15965);
and U22177 (N_22177,N_17085,N_16555);
nor U22178 (N_22178,N_19892,N_17618);
nor U22179 (N_22179,N_16801,N_15950);
nor U22180 (N_22180,N_19278,N_18283);
and U22181 (N_22181,N_16992,N_15075);
and U22182 (N_22182,N_17915,N_18855);
nand U22183 (N_22183,N_15028,N_18460);
or U22184 (N_22184,N_18866,N_19277);
nand U22185 (N_22185,N_16259,N_17282);
and U22186 (N_22186,N_19282,N_17898);
xnor U22187 (N_22187,N_18219,N_15524);
or U22188 (N_22188,N_16923,N_19000);
nand U22189 (N_22189,N_17853,N_16694);
or U22190 (N_22190,N_16948,N_15471);
or U22191 (N_22191,N_19876,N_17475);
xor U22192 (N_22192,N_16752,N_17196);
and U22193 (N_22193,N_17503,N_17683);
or U22194 (N_22194,N_17903,N_18731);
nand U22195 (N_22195,N_19975,N_18047);
and U22196 (N_22196,N_16321,N_15983);
nor U22197 (N_22197,N_15857,N_15700);
xor U22198 (N_22198,N_18517,N_15610);
nand U22199 (N_22199,N_15780,N_15462);
and U22200 (N_22200,N_16218,N_19906);
nand U22201 (N_22201,N_19204,N_15503);
nand U22202 (N_22202,N_16244,N_17078);
or U22203 (N_22203,N_18493,N_16305);
xnor U22204 (N_22204,N_19862,N_17908);
and U22205 (N_22205,N_18135,N_18575);
nor U22206 (N_22206,N_16560,N_18726);
or U22207 (N_22207,N_16676,N_18282);
xor U22208 (N_22208,N_16424,N_19926);
xnor U22209 (N_22209,N_15455,N_15416);
and U22210 (N_22210,N_18277,N_17555);
or U22211 (N_22211,N_16928,N_18617);
xnor U22212 (N_22212,N_19212,N_19402);
or U22213 (N_22213,N_15670,N_17061);
xnor U22214 (N_22214,N_16857,N_16535);
or U22215 (N_22215,N_18865,N_19788);
or U22216 (N_22216,N_15231,N_18605);
nor U22217 (N_22217,N_16407,N_16123);
or U22218 (N_22218,N_17871,N_17667);
nor U22219 (N_22219,N_17361,N_16269);
nor U22220 (N_22220,N_18049,N_18802);
nor U22221 (N_22221,N_18370,N_16425);
nor U22222 (N_22222,N_16384,N_17185);
or U22223 (N_22223,N_19002,N_15877);
nor U22224 (N_22224,N_18281,N_19317);
and U22225 (N_22225,N_17073,N_18919);
and U22226 (N_22226,N_16566,N_15064);
and U22227 (N_22227,N_15937,N_17691);
and U22228 (N_22228,N_18451,N_18649);
xnor U22229 (N_22229,N_17083,N_15737);
and U22230 (N_22230,N_17528,N_19512);
nand U22231 (N_22231,N_16987,N_16712);
or U22232 (N_22232,N_15133,N_19307);
and U22233 (N_22233,N_15061,N_16658);
or U22234 (N_22234,N_16809,N_18681);
xor U22235 (N_22235,N_15880,N_15777);
xor U22236 (N_22236,N_17388,N_16782);
or U22237 (N_22237,N_17429,N_17709);
and U22238 (N_22238,N_16677,N_15881);
nor U22239 (N_22239,N_16335,N_15805);
nor U22240 (N_22240,N_15749,N_18011);
nand U22241 (N_22241,N_19205,N_16778);
nor U22242 (N_22242,N_19391,N_16392);
or U22243 (N_22243,N_15141,N_18988);
nor U22244 (N_22244,N_19483,N_15563);
nor U22245 (N_22245,N_18437,N_17936);
nand U22246 (N_22246,N_18753,N_15402);
or U22247 (N_22247,N_16622,N_15773);
nand U22248 (N_22248,N_18184,N_15554);
or U22249 (N_22249,N_15253,N_15673);
nand U22250 (N_22250,N_18013,N_15976);
or U22251 (N_22251,N_17889,N_15689);
nand U22252 (N_22252,N_17722,N_17472);
nand U22253 (N_22253,N_19443,N_17694);
nand U22254 (N_22254,N_16144,N_18438);
xnor U22255 (N_22255,N_16052,N_16985);
and U22256 (N_22256,N_18827,N_16091);
and U22257 (N_22257,N_17476,N_15190);
or U22258 (N_22258,N_17957,N_19854);
or U22259 (N_22259,N_19158,N_18389);
xor U22260 (N_22260,N_17766,N_15732);
and U22261 (N_22261,N_19557,N_15331);
or U22262 (N_22262,N_15374,N_15578);
xor U22263 (N_22263,N_17071,N_17337);
or U22264 (N_22264,N_16855,N_15631);
nor U22265 (N_22265,N_19644,N_16265);
and U22266 (N_22266,N_18700,N_18112);
nor U22267 (N_22267,N_17463,N_16083);
nand U22268 (N_22268,N_15088,N_17345);
and U22269 (N_22269,N_17558,N_15063);
nor U22270 (N_22270,N_18167,N_17486);
nor U22271 (N_22271,N_18124,N_15858);
nand U22272 (N_22272,N_16843,N_19549);
or U22273 (N_22273,N_18118,N_18833);
and U22274 (N_22274,N_17815,N_16757);
or U22275 (N_22275,N_18029,N_18590);
nor U22276 (N_22276,N_19099,N_15620);
nand U22277 (N_22277,N_16263,N_17840);
nor U22278 (N_22278,N_17367,N_16829);
and U22279 (N_22279,N_17918,N_16242);
and U22280 (N_22280,N_15470,N_18115);
or U22281 (N_22281,N_15981,N_19108);
nand U22282 (N_22282,N_19759,N_19574);
nor U22283 (N_22283,N_15193,N_17594);
xnor U22284 (N_22284,N_18138,N_16633);
and U22285 (N_22285,N_19953,N_18967);
and U22286 (N_22286,N_18076,N_18980);
and U22287 (N_22287,N_16751,N_16601);
and U22288 (N_22288,N_16523,N_18055);
or U22289 (N_22289,N_17615,N_15240);
and U22290 (N_22290,N_19476,N_19566);
or U22291 (N_22291,N_18829,N_19722);
nor U22292 (N_22292,N_19649,N_15219);
or U22293 (N_22293,N_17023,N_19032);
nand U22294 (N_22294,N_17737,N_17174);
nor U22295 (N_22295,N_17533,N_19021);
nor U22296 (N_22296,N_16051,N_17219);
or U22297 (N_22297,N_15915,N_15903);
nor U22298 (N_22298,N_19937,N_16708);
xor U22299 (N_22299,N_19987,N_18444);
nand U22300 (N_22300,N_15166,N_19423);
or U22301 (N_22301,N_17354,N_19272);
or U22302 (N_22302,N_18009,N_17405);
nand U22303 (N_22303,N_15320,N_17483);
and U22304 (N_22304,N_16723,N_17487);
xor U22305 (N_22305,N_19816,N_15197);
and U22306 (N_22306,N_18809,N_19343);
or U22307 (N_22307,N_19501,N_15464);
and U22308 (N_22308,N_18101,N_19781);
and U22309 (N_22309,N_17945,N_19504);
nand U22310 (N_22310,N_15119,N_17209);
nand U22311 (N_22311,N_19425,N_16345);
xnor U22312 (N_22312,N_18961,N_15477);
and U22313 (N_22313,N_18944,N_17499);
xor U22314 (N_22314,N_16082,N_17831);
and U22315 (N_22315,N_16481,N_19071);
or U22316 (N_22316,N_18149,N_15811);
xor U22317 (N_22317,N_16522,N_18312);
nor U22318 (N_22318,N_18818,N_16278);
or U22319 (N_22319,N_19004,N_15547);
xnor U22320 (N_22320,N_19162,N_19588);
and U22321 (N_22321,N_17877,N_16690);
and U22322 (N_22322,N_18992,N_17565);
nor U22323 (N_22323,N_19475,N_18229);
or U22324 (N_22324,N_18769,N_17725);
or U22325 (N_22325,N_19018,N_15861);
and U22326 (N_22326,N_19242,N_16036);
or U22327 (N_22327,N_19240,N_18578);
nand U22328 (N_22328,N_17942,N_16354);
nor U22329 (N_22329,N_17585,N_16767);
nand U22330 (N_22330,N_16883,N_15335);
or U22331 (N_22331,N_19711,N_18082);
and U22332 (N_22332,N_17423,N_18872);
or U22333 (N_22333,N_17508,N_17308);
nand U22334 (N_22334,N_16176,N_15947);
nor U22335 (N_22335,N_15736,N_17703);
and U22336 (N_22336,N_18401,N_16019);
nand U22337 (N_22337,N_16568,N_17653);
and U22338 (N_22338,N_15466,N_19775);
or U22339 (N_22339,N_16652,N_17152);
nand U22340 (N_22340,N_19340,N_18266);
or U22341 (N_22341,N_17785,N_19251);
and U22342 (N_22342,N_18889,N_18996);
or U22343 (N_22343,N_19634,N_18850);
and U22344 (N_22344,N_15360,N_15490);
or U22345 (N_22345,N_19220,N_15264);
or U22346 (N_22346,N_18221,N_18748);
nand U22347 (N_22347,N_17989,N_16080);
or U22348 (N_22348,N_15343,N_15951);
or U22349 (N_22349,N_19235,N_18755);
xor U22350 (N_22350,N_17976,N_16571);
nand U22351 (N_22351,N_19030,N_15884);
or U22352 (N_22352,N_16583,N_17394);
and U22353 (N_22353,N_17084,N_19028);
and U22354 (N_22354,N_18391,N_16388);
nand U22355 (N_22355,N_19725,N_18481);
and U22356 (N_22356,N_16578,N_17190);
nor U22357 (N_22357,N_19682,N_16584);
xor U22358 (N_22358,N_19144,N_18230);
and U22359 (N_22359,N_15260,N_17141);
nor U22360 (N_22360,N_15898,N_15542);
xnor U22361 (N_22361,N_19723,N_19459);
nor U22362 (N_22362,N_15191,N_16646);
or U22363 (N_22363,N_16495,N_19897);
or U22364 (N_22364,N_18781,N_18601);
nand U22365 (N_22365,N_17825,N_16705);
and U22366 (N_22366,N_19706,N_16360);
nand U22367 (N_22367,N_17418,N_16604);
or U22368 (N_22368,N_19565,N_15033);
nor U22369 (N_22369,N_17307,N_17559);
nand U22370 (N_22370,N_19811,N_17748);
and U22371 (N_22371,N_19474,N_19344);
nor U22372 (N_22372,N_17341,N_18991);
xor U22373 (N_22373,N_16168,N_19407);
or U22374 (N_22374,N_18797,N_18053);
nand U22375 (N_22375,N_18656,N_17894);
xnor U22376 (N_22376,N_19960,N_16417);
or U22377 (N_22377,N_15446,N_19598);
nor U22378 (N_22378,N_16194,N_19537);
xnor U22379 (N_22379,N_17279,N_15052);
nor U22380 (N_22380,N_16488,N_15000);
or U22381 (N_22381,N_15753,N_17578);
and U22382 (N_22382,N_17626,N_18664);
or U22383 (N_22383,N_19087,N_15655);
nor U22384 (N_22384,N_15131,N_17144);
and U22385 (N_22385,N_16202,N_16117);
or U22386 (N_22386,N_16733,N_16191);
and U22387 (N_22387,N_18775,N_16670);
xnor U22388 (N_22388,N_18215,N_16644);
or U22389 (N_22389,N_15163,N_18808);
or U22390 (N_22390,N_18172,N_18179);
nor U22391 (N_22391,N_16704,N_19663);
nand U22392 (N_22392,N_16549,N_17567);
nand U22393 (N_22393,N_16381,N_18253);
xnor U22394 (N_22394,N_17596,N_15031);
nor U22395 (N_22395,N_19179,N_18643);
nand U22396 (N_22396,N_16339,N_19267);
nor U22397 (N_22397,N_18927,N_15968);
and U22398 (N_22398,N_18910,N_17755);
nor U22399 (N_22399,N_15527,N_17888);
nor U22400 (N_22400,N_17270,N_18911);
and U22401 (N_22401,N_19833,N_16122);
or U22402 (N_22402,N_16816,N_15330);
and U22403 (N_22403,N_19225,N_15080);
and U22404 (N_22404,N_17501,N_17995);
nor U22405 (N_22405,N_17793,N_15406);
nand U22406 (N_22406,N_19284,N_15690);
xor U22407 (N_22407,N_15604,N_16874);
nor U22408 (N_22408,N_16262,N_18718);
and U22409 (N_22409,N_18673,N_18252);
or U22410 (N_22410,N_17857,N_16282);
nand U22411 (N_22411,N_15576,N_15169);
xnor U22412 (N_22412,N_15672,N_18674);
xnor U22413 (N_22413,N_17049,N_17098);
or U22414 (N_22414,N_16613,N_18713);
nand U22415 (N_22415,N_16862,N_16750);
or U22416 (N_22416,N_18373,N_18840);
nand U22417 (N_22417,N_16638,N_16487);
xor U22418 (N_22418,N_16797,N_17318);
or U22419 (N_22419,N_16572,N_17019);
or U22420 (N_22420,N_17707,N_18733);
and U22421 (N_22421,N_17878,N_15378);
nor U22422 (N_22422,N_17716,N_18384);
nand U22423 (N_22423,N_16919,N_17397);
xnor U22424 (N_22424,N_18825,N_16538);
nor U22425 (N_22425,N_15643,N_17543);
or U22426 (N_22426,N_15129,N_16698);
or U22427 (N_22427,N_16615,N_19745);
or U22428 (N_22428,N_18279,N_18626);
nand U22429 (N_22429,N_18779,N_19013);
xor U22430 (N_22430,N_16851,N_17964);
or U22431 (N_22431,N_18422,N_18150);
and U22432 (N_22432,N_18234,N_16796);
or U22433 (N_22433,N_15583,N_19309);
nand U22434 (N_22434,N_18502,N_17808);
and U22435 (N_22435,N_19823,N_16059);
nand U22436 (N_22436,N_16022,N_19227);
nand U22437 (N_22437,N_19836,N_19134);
or U22438 (N_22438,N_18792,N_15317);
or U22439 (N_22439,N_19415,N_15100);
xor U22440 (N_22440,N_15013,N_17692);
xor U22441 (N_22441,N_19061,N_16716);
nand U22442 (N_22442,N_15085,N_15545);
or U22443 (N_22443,N_18051,N_16120);
nand U22444 (N_22444,N_19743,N_15754);
and U22445 (N_22445,N_18562,N_17143);
nor U22446 (N_22446,N_18701,N_15760);
xnor U22447 (N_22447,N_15314,N_19563);
or U22448 (N_22448,N_18964,N_17076);
nor U22449 (N_22449,N_15592,N_18846);
nand U22450 (N_22450,N_17484,N_16023);
nand U22451 (N_22451,N_17376,N_17550);
xnor U22452 (N_22452,N_15121,N_17647);
nor U22453 (N_22453,N_19567,N_15435);
nand U22454 (N_22454,N_17179,N_18599);
or U22455 (N_22455,N_15894,N_19322);
or U22456 (N_22456,N_15953,N_16590);
nor U22457 (N_22457,N_17969,N_17609);
and U22458 (N_22458,N_18759,N_19776);
nand U22459 (N_22459,N_19852,N_19065);
or U22460 (N_22460,N_15093,N_15445);
or U22461 (N_22461,N_18299,N_17786);
or U22462 (N_22462,N_15444,N_19133);
nand U22463 (N_22463,N_15198,N_17027);
xnor U22464 (N_22464,N_19331,N_19685);
or U22465 (N_22465,N_19226,N_16703);
xnor U22466 (N_22466,N_16317,N_19308);
and U22467 (N_22467,N_19078,N_17758);
nor U22468 (N_22468,N_15744,N_18240);
or U22469 (N_22469,N_16430,N_19855);
nand U22470 (N_22470,N_18520,N_19841);
nand U22471 (N_22471,N_18876,N_15831);
nand U22472 (N_22472,N_19589,N_19121);
nand U22473 (N_22473,N_19364,N_17741);
or U22474 (N_22474,N_19128,N_17161);
nand U22475 (N_22475,N_19127,N_16518);
xnor U22476 (N_22476,N_15591,N_17680);
xor U22477 (N_22477,N_15125,N_19718);
or U22478 (N_22478,N_16214,N_15551);
nand U22479 (N_22479,N_18908,N_19042);
nor U22480 (N_22480,N_19038,N_17531);
xnor U22481 (N_22481,N_16659,N_19707);
nor U22482 (N_22482,N_16632,N_18807);
and U22483 (N_22483,N_16881,N_15423);
nand U22484 (N_22484,N_16172,N_15909);
nand U22485 (N_22485,N_19247,N_16745);
nor U22486 (N_22486,N_15860,N_15742);
nor U22487 (N_22487,N_17077,N_17923);
or U22488 (N_22488,N_18788,N_18963);
or U22489 (N_22489,N_15618,N_17782);
and U22490 (N_22490,N_18494,N_18698);
nand U22491 (N_22491,N_16399,N_18777);
nor U22492 (N_22492,N_19082,N_15599);
or U22493 (N_22493,N_17941,N_18811);
and U22494 (N_22494,N_18611,N_15815);
or U22495 (N_22495,N_16419,N_16965);
and U22496 (N_22496,N_17277,N_19093);
nand U22497 (N_22497,N_15998,N_19798);
nor U22498 (N_22498,N_15531,N_19260);
and U22499 (N_22499,N_17699,N_16781);
xnor U22500 (N_22500,N_19337,N_18211);
or U22501 (N_22501,N_16252,N_15730);
and U22502 (N_22502,N_16228,N_16320);
nor U22503 (N_22503,N_19829,N_16843);
nor U22504 (N_22504,N_18672,N_19203);
xnor U22505 (N_22505,N_19173,N_18609);
or U22506 (N_22506,N_16189,N_16784);
nor U22507 (N_22507,N_19383,N_18925);
or U22508 (N_22508,N_19162,N_16531);
nor U22509 (N_22509,N_15545,N_18381);
and U22510 (N_22510,N_17131,N_15572);
or U22511 (N_22511,N_18076,N_18663);
nor U22512 (N_22512,N_18977,N_15351);
xor U22513 (N_22513,N_16130,N_18472);
or U22514 (N_22514,N_17612,N_16223);
nor U22515 (N_22515,N_15435,N_16730);
nor U22516 (N_22516,N_19239,N_19553);
or U22517 (N_22517,N_18614,N_15517);
and U22518 (N_22518,N_19599,N_18924);
nand U22519 (N_22519,N_16866,N_19979);
nand U22520 (N_22520,N_15550,N_16736);
nor U22521 (N_22521,N_17235,N_19146);
nand U22522 (N_22522,N_15901,N_19345);
or U22523 (N_22523,N_19626,N_17242);
or U22524 (N_22524,N_17493,N_19061);
and U22525 (N_22525,N_17816,N_17101);
or U22526 (N_22526,N_19915,N_19771);
nor U22527 (N_22527,N_18623,N_17042);
nor U22528 (N_22528,N_15037,N_18136);
nand U22529 (N_22529,N_18786,N_17985);
nor U22530 (N_22530,N_18505,N_16723);
nor U22531 (N_22531,N_18458,N_19344);
nor U22532 (N_22532,N_15820,N_16633);
nor U22533 (N_22533,N_19143,N_16183);
nor U22534 (N_22534,N_16730,N_19928);
and U22535 (N_22535,N_16341,N_18520);
nand U22536 (N_22536,N_19566,N_19326);
xnor U22537 (N_22537,N_16513,N_19635);
and U22538 (N_22538,N_19814,N_15838);
xnor U22539 (N_22539,N_19122,N_16677);
nor U22540 (N_22540,N_15524,N_18026);
nand U22541 (N_22541,N_19278,N_16643);
and U22542 (N_22542,N_16661,N_18212);
nand U22543 (N_22543,N_16051,N_16232);
and U22544 (N_22544,N_16260,N_18541);
or U22545 (N_22545,N_16795,N_15671);
and U22546 (N_22546,N_18469,N_18868);
or U22547 (N_22547,N_16226,N_17823);
nor U22548 (N_22548,N_19967,N_17666);
xor U22549 (N_22549,N_18818,N_17870);
or U22550 (N_22550,N_19043,N_19095);
nand U22551 (N_22551,N_19973,N_17743);
nand U22552 (N_22552,N_16712,N_17198);
nand U22553 (N_22553,N_16692,N_16930);
nand U22554 (N_22554,N_17269,N_19470);
and U22555 (N_22555,N_18187,N_19840);
and U22556 (N_22556,N_16535,N_18977);
or U22557 (N_22557,N_16171,N_19224);
or U22558 (N_22558,N_15269,N_16753);
nand U22559 (N_22559,N_17982,N_18455);
nor U22560 (N_22560,N_17862,N_15847);
nor U22561 (N_22561,N_18208,N_17723);
and U22562 (N_22562,N_19348,N_19155);
nand U22563 (N_22563,N_16265,N_18236);
or U22564 (N_22564,N_17006,N_19745);
and U22565 (N_22565,N_18533,N_19667);
or U22566 (N_22566,N_19656,N_15894);
xor U22567 (N_22567,N_18562,N_18615);
nor U22568 (N_22568,N_18672,N_19456);
nand U22569 (N_22569,N_15875,N_15024);
or U22570 (N_22570,N_17611,N_19302);
nand U22571 (N_22571,N_17643,N_17918);
nand U22572 (N_22572,N_17430,N_16914);
or U22573 (N_22573,N_19712,N_17043);
nor U22574 (N_22574,N_19736,N_15662);
nor U22575 (N_22575,N_18590,N_16948);
or U22576 (N_22576,N_17659,N_17055);
or U22577 (N_22577,N_16321,N_16324);
or U22578 (N_22578,N_17024,N_19757);
nor U22579 (N_22579,N_18723,N_16439);
nor U22580 (N_22580,N_19369,N_18960);
and U22581 (N_22581,N_17799,N_17764);
and U22582 (N_22582,N_19298,N_15023);
nand U22583 (N_22583,N_15168,N_16102);
nor U22584 (N_22584,N_19877,N_18828);
and U22585 (N_22585,N_17191,N_19197);
nor U22586 (N_22586,N_19944,N_15043);
nor U22587 (N_22587,N_16401,N_19757);
nand U22588 (N_22588,N_16734,N_18544);
nor U22589 (N_22589,N_15258,N_15948);
or U22590 (N_22590,N_18758,N_19402);
or U22591 (N_22591,N_19784,N_19844);
or U22592 (N_22592,N_18539,N_15321);
or U22593 (N_22593,N_17986,N_18831);
nor U22594 (N_22594,N_18755,N_15564);
or U22595 (N_22595,N_15404,N_19254);
or U22596 (N_22596,N_19211,N_18375);
or U22597 (N_22597,N_19290,N_18201);
and U22598 (N_22598,N_16210,N_16764);
or U22599 (N_22599,N_16146,N_18126);
or U22600 (N_22600,N_18121,N_17026);
nand U22601 (N_22601,N_17700,N_15926);
nor U22602 (N_22602,N_19949,N_17874);
xnor U22603 (N_22603,N_18883,N_18010);
nand U22604 (N_22604,N_17862,N_18530);
nor U22605 (N_22605,N_18932,N_17981);
nand U22606 (N_22606,N_18332,N_18207);
or U22607 (N_22607,N_18474,N_18163);
or U22608 (N_22608,N_19354,N_19011);
or U22609 (N_22609,N_15073,N_19836);
and U22610 (N_22610,N_18220,N_19604);
or U22611 (N_22611,N_17457,N_19517);
nor U22612 (N_22612,N_17872,N_17217);
and U22613 (N_22613,N_19131,N_15075);
nand U22614 (N_22614,N_17358,N_19462);
and U22615 (N_22615,N_19841,N_18291);
and U22616 (N_22616,N_16047,N_17193);
or U22617 (N_22617,N_16827,N_17079);
and U22618 (N_22618,N_15009,N_18124);
nor U22619 (N_22619,N_17426,N_16845);
and U22620 (N_22620,N_19152,N_15687);
or U22621 (N_22621,N_15921,N_18044);
xor U22622 (N_22622,N_16939,N_18072);
or U22623 (N_22623,N_16374,N_16027);
or U22624 (N_22624,N_15325,N_15706);
and U22625 (N_22625,N_19921,N_18660);
or U22626 (N_22626,N_16677,N_17073);
and U22627 (N_22627,N_15908,N_15635);
xnor U22628 (N_22628,N_17268,N_16918);
and U22629 (N_22629,N_18788,N_18317);
or U22630 (N_22630,N_18411,N_17681);
and U22631 (N_22631,N_19765,N_18060);
nor U22632 (N_22632,N_19864,N_16527);
xnor U22633 (N_22633,N_17548,N_17078);
nor U22634 (N_22634,N_16114,N_18440);
and U22635 (N_22635,N_17099,N_15357);
or U22636 (N_22636,N_15492,N_17498);
or U22637 (N_22637,N_19242,N_16525);
xnor U22638 (N_22638,N_18015,N_16879);
nor U22639 (N_22639,N_15455,N_18591);
and U22640 (N_22640,N_19933,N_16360);
nor U22641 (N_22641,N_18825,N_19745);
xnor U22642 (N_22642,N_15384,N_15807);
nand U22643 (N_22643,N_16083,N_15584);
or U22644 (N_22644,N_15558,N_16094);
nand U22645 (N_22645,N_17165,N_15470);
or U22646 (N_22646,N_16361,N_17568);
or U22647 (N_22647,N_18610,N_17243);
or U22648 (N_22648,N_16149,N_17749);
nor U22649 (N_22649,N_18801,N_19813);
or U22650 (N_22650,N_18174,N_15471);
nand U22651 (N_22651,N_19004,N_15481);
nand U22652 (N_22652,N_17531,N_18988);
xor U22653 (N_22653,N_19046,N_17489);
and U22654 (N_22654,N_15447,N_18283);
and U22655 (N_22655,N_17683,N_19698);
or U22656 (N_22656,N_15013,N_15305);
or U22657 (N_22657,N_15326,N_18657);
nand U22658 (N_22658,N_16866,N_17153);
and U22659 (N_22659,N_15386,N_19184);
xnor U22660 (N_22660,N_17468,N_17460);
nand U22661 (N_22661,N_16892,N_19391);
or U22662 (N_22662,N_15228,N_15732);
and U22663 (N_22663,N_18330,N_17060);
nand U22664 (N_22664,N_19861,N_19056);
and U22665 (N_22665,N_19373,N_18121);
xor U22666 (N_22666,N_15414,N_16625);
or U22667 (N_22667,N_16369,N_18907);
xnor U22668 (N_22668,N_15988,N_19731);
nand U22669 (N_22669,N_16904,N_19930);
xor U22670 (N_22670,N_15237,N_17095);
or U22671 (N_22671,N_16212,N_16188);
nand U22672 (N_22672,N_17686,N_16300);
or U22673 (N_22673,N_18454,N_16904);
or U22674 (N_22674,N_17658,N_15970);
nor U22675 (N_22675,N_18597,N_18357);
nor U22676 (N_22676,N_18256,N_18985);
and U22677 (N_22677,N_18941,N_18947);
or U22678 (N_22678,N_19579,N_15405);
nand U22679 (N_22679,N_18439,N_19654);
nand U22680 (N_22680,N_16197,N_15723);
nand U22681 (N_22681,N_15957,N_18671);
or U22682 (N_22682,N_19132,N_16003);
or U22683 (N_22683,N_18805,N_17686);
or U22684 (N_22684,N_15161,N_17056);
or U22685 (N_22685,N_16762,N_16951);
nor U22686 (N_22686,N_18786,N_18747);
nor U22687 (N_22687,N_18170,N_16101);
xor U22688 (N_22688,N_16139,N_15484);
nor U22689 (N_22689,N_17876,N_18591);
or U22690 (N_22690,N_19977,N_18821);
or U22691 (N_22691,N_16332,N_17223);
and U22692 (N_22692,N_16409,N_17252);
or U22693 (N_22693,N_18215,N_16079);
nor U22694 (N_22694,N_16354,N_19699);
and U22695 (N_22695,N_17015,N_17691);
and U22696 (N_22696,N_18648,N_17995);
nand U22697 (N_22697,N_15508,N_18972);
or U22698 (N_22698,N_15778,N_16477);
xor U22699 (N_22699,N_19358,N_18405);
or U22700 (N_22700,N_19707,N_17796);
xor U22701 (N_22701,N_15379,N_17249);
or U22702 (N_22702,N_19854,N_17500);
nand U22703 (N_22703,N_16344,N_18403);
and U22704 (N_22704,N_19932,N_17974);
or U22705 (N_22705,N_18920,N_15326);
nor U22706 (N_22706,N_19662,N_16822);
nand U22707 (N_22707,N_15976,N_18150);
nor U22708 (N_22708,N_19887,N_19592);
or U22709 (N_22709,N_19586,N_18624);
nand U22710 (N_22710,N_19939,N_17943);
or U22711 (N_22711,N_16758,N_16117);
xnor U22712 (N_22712,N_17103,N_19584);
or U22713 (N_22713,N_15386,N_19609);
nor U22714 (N_22714,N_19630,N_16403);
nor U22715 (N_22715,N_18440,N_17008);
nor U22716 (N_22716,N_17224,N_16591);
nor U22717 (N_22717,N_19239,N_18426);
and U22718 (N_22718,N_16176,N_16345);
nand U22719 (N_22719,N_16980,N_18915);
or U22720 (N_22720,N_17051,N_15381);
or U22721 (N_22721,N_16399,N_19757);
and U22722 (N_22722,N_18668,N_16502);
or U22723 (N_22723,N_18703,N_18925);
and U22724 (N_22724,N_15490,N_19920);
or U22725 (N_22725,N_15889,N_16573);
or U22726 (N_22726,N_16419,N_15074);
or U22727 (N_22727,N_17628,N_19038);
nand U22728 (N_22728,N_19586,N_15238);
xor U22729 (N_22729,N_15086,N_18284);
nand U22730 (N_22730,N_15089,N_19434);
and U22731 (N_22731,N_15823,N_17224);
and U22732 (N_22732,N_16798,N_15738);
and U22733 (N_22733,N_16523,N_19375);
nor U22734 (N_22734,N_15633,N_15419);
or U22735 (N_22735,N_16633,N_16007);
nor U22736 (N_22736,N_17606,N_17081);
or U22737 (N_22737,N_19768,N_15289);
or U22738 (N_22738,N_18211,N_15123);
and U22739 (N_22739,N_17784,N_19797);
and U22740 (N_22740,N_19813,N_17911);
or U22741 (N_22741,N_17732,N_15790);
or U22742 (N_22742,N_16003,N_15352);
and U22743 (N_22743,N_19625,N_15244);
nand U22744 (N_22744,N_17797,N_16622);
nand U22745 (N_22745,N_15193,N_19116);
nand U22746 (N_22746,N_18807,N_16192);
and U22747 (N_22747,N_15435,N_16298);
or U22748 (N_22748,N_17158,N_17698);
or U22749 (N_22749,N_18431,N_19366);
and U22750 (N_22750,N_19175,N_15055);
nor U22751 (N_22751,N_15029,N_19979);
or U22752 (N_22752,N_18027,N_18902);
and U22753 (N_22753,N_19499,N_19200);
and U22754 (N_22754,N_19628,N_17778);
nand U22755 (N_22755,N_16250,N_16637);
or U22756 (N_22756,N_18388,N_15392);
or U22757 (N_22757,N_15981,N_16900);
nand U22758 (N_22758,N_18370,N_17958);
nor U22759 (N_22759,N_19690,N_17032);
nor U22760 (N_22760,N_19453,N_15546);
nor U22761 (N_22761,N_19232,N_15937);
or U22762 (N_22762,N_15441,N_19533);
nand U22763 (N_22763,N_15708,N_18966);
or U22764 (N_22764,N_17200,N_17575);
and U22765 (N_22765,N_18589,N_17072);
nor U22766 (N_22766,N_16460,N_15975);
nand U22767 (N_22767,N_17384,N_18421);
and U22768 (N_22768,N_17493,N_16316);
and U22769 (N_22769,N_19539,N_19722);
nand U22770 (N_22770,N_16412,N_17872);
nor U22771 (N_22771,N_15099,N_16697);
nand U22772 (N_22772,N_19146,N_18999);
nor U22773 (N_22773,N_17741,N_17980);
nor U22774 (N_22774,N_17686,N_19750);
or U22775 (N_22775,N_18171,N_18502);
nand U22776 (N_22776,N_18115,N_15486);
or U22777 (N_22777,N_18314,N_19686);
or U22778 (N_22778,N_18792,N_18086);
and U22779 (N_22779,N_19646,N_18017);
and U22780 (N_22780,N_19413,N_15627);
nor U22781 (N_22781,N_17967,N_15486);
and U22782 (N_22782,N_17659,N_17526);
nor U22783 (N_22783,N_19075,N_15748);
or U22784 (N_22784,N_18687,N_15425);
nor U22785 (N_22785,N_19815,N_15092);
or U22786 (N_22786,N_19605,N_19713);
xnor U22787 (N_22787,N_16675,N_16672);
nor U22788 (N_22788,N_15963,N_18406);
and U22789 (N_22789,N_16603,N_17335);
nor U22790 (N_22790,N_15593,N_17245);
nand U22791 (N_22791,N_17433,N_19044);
or U22792 (N_22792,N_15980,N_15078);
and U22793 (N_22793,N_17321,N_19461);
nor U22794 (N_22794,N_19102,N_18090);
nor U22795 (N_22795,N_15191,N_16119);
and U22796 (N_22796,N_16013,N_15287);
and U22797 (N_22797,N_16529,N_15475);
or U22798 (N_22798,N_17488,N_17565);
nor U22799 (N_22799,N_15115,N_18983);
or U22800 (N_22800,N_19089,N_19691);
nor U22801 (N_22801,N_17981,N_16313);
or U22802 (N_22802,N_17769,N_19563);
or U22803 (N_22803,N_16992,N_16553);
or U22804 (N_22804,N_19562,N_18211);
and U22805 (N_22805,N_17033,N_16905);
and U22806 (N_22806,N_18609,N_15942);
and U22807 (N_22807,N_18208,N_15881);
and U22808 (N_22808,N_15556,N_15050);
nor U22809 (N_22809,N_17749,N_18935);
nand U22810 (N_22810,N_17026,N_15869);
or U22811 (N_22811,N_16810,N_17408);
nand U22812 (N_22812,N_15251,N_15591);
and U22813 (N_22813,N_16836,N_19731);
or U22814 (N_22814,N_18273,N_16174);
nor U22815 (N_22815,N_18323,N_17007);
or U22816 (N_22816,N_15514,N_17198);
nor U22817 (N_22817,N_19311,N_18713);
or U22818 (N_22818,N_18171,N_18735);
nand U22819 (N_22819,N_16753,N_19426);
nand U22820 (N_22820,N_18932,N_15200);
and U22821 (N_22821,N_16496,N_15200);
xor U22822 (N_22822,N_18810,N_19901);
nand U22823 (N_22823,N_18463,N_16324);
nand U22824 (N_22824,N_19679,N_15497);
and U22825 (N_22825,N_19328,N_17106);
nor U22826 (N_22826,N_18345,N_17750);
nand U22827 (N_22827,N_17878,N_19087);
nor U22828 (N_22828,N_18427,N_17473);
xor U22829 (N_22829,N_15156,N_17114);
nand U22830 (N_22830,N_16322,N_17121);
or U22831 (N_22831,N_15493,N_18707);
nor U22832 (N_22832,N_19170,N_18027);
and U22833 (N_22833,N_18505,N_16114);
or U22834 (N_22834,N_19187,N_15486);
nor U22835 (N_22835,N_18031,N_16855);
nand U22836 (N_22836,N_15392,N_18426);
nand U22837 (N_22837,N_18341,N_16210);
or U22838 (N_22838,N_16286,N_18133);
and U22839 (N_22839,N_17912,N_16843);
and U22840 (N_22840,N_19082,N_19006);
and U22841 (N_22841,N_18566,N_16550);
nor U22842 (N_22842,N_19436,N_19174);
or U22843 (N_22843,N_16901,N_15952);
and U22844 (N_22844,N_19327,N_17906);
or U22845 (N_22845,N_15699,N_16524);
nor U22846 (N_22846,N_19847,N_19978);
or U22847 (N_22847,N_16202,N_19391);
or U22848 (N_22848,N_17720,N_17677);
nor U22849 (N_22849,N_19863,N_19914);
and U22850 (N_22850,N_18100,N_16751);
and U22851 (N_22851,N_15243,N_17569);
and U22852 (N_22852,N_18775,N_15273);
nor U22853 (N_22853,N_18607,N_16927);
and U22854 (N_22854,N_17509,N_16517);
and U22855 (N_22855,N_15898,N_18332);
and U22856 (N_22856,N_16996,N_17595);
nor U22857 (N_22857,N_15475,N_19571);
or U22858 (N_22858,N_15784,N_16324);
nand U22859 (N_22859,N_16944,N_15803);
nand U22860 (N_22860,N_16390,N_15918);
and U22861 (N_22861,N_19093,N_19289);
nor U22862 (N_22862,N_17857,N_17378);
nand U22863 (N_22863,N_19831,N_16877);
and U22864 (N_22864,N_15747,N_19128);
and U22865 (N_22865,N_15513,N_17026);
nand U22866 (N_22866,N_19649,N_18565);
nor U22867 (N_22867,N_18334,N_15432);
nand U22868 (N_22868,N_17226,N_18517);
nor U22869 (N_22869,N_17702,N_19991);
and U22870 (N_22870,N_16986,N_15723);
and U22871 (N_22871,N_19948,N_18877);
and U22872 (N_22872,N_16592,N_18101);
or U22873 (N_22873,N_19004,N_15258);
and U22874 (N_22874,N_19777,N_17185);
or U22875 (N_22875,N_18556,N_15456);
and U22876 (N_22876,N_15989,N_15764);
nand U22877 (N_22877,N_16000,N_17449);
nand U22878 (N_22878,N_18419,N_19720);
xnor U22879 (N_22879,N_16979,N_18763);
or U22880 (N_22880,N_19236,N_16755);
or U22881 (N_22881,N_17711,N_18635);
or U22882 (N_22882,N_19308,N_18372);
nand U22883 (N_22883,N_19400,N_17580);
nand U22884 (N_22884,N_18051,N_19037);
nand U22885 (N_22885,N_15564,N_18292);
and U22886 (N_22886,N_18780,N_16590);
xnor U22887 (N_22887,N_16184,N_16194);
or U22888 (N_22888,N_17074,N_16120);
and U22889 (N_22889,N_19271,N_19591);
nor U22890 (N_22890,N_18228,N_15847);
or U22891 (N_22891,N_16387,N_18361);
and U22892 (N_22892,N_16434,N_18320);
or U22893 (N_22893,N_17456,N_15843);
nand U22894 (N_22894,N_19661,N_17275);
nor U22895 (N_22895,N_15762,N_19512);
or U22896 (N_22896,N_18187,N_17882);
nor U22897 (N_22897,N_15495,N_17406);
nand U22898 (N_22898,N_18834,N_19836);
nor U22899 (N_22899,N_18943,N_15586);
or U22900 (N_22900,N_18621,N_18755);
nand U22901 (N_22901,N_19885,N_16322);
and U22902 (N_22902,N_17912,N_16011);
nand U22903 (N_22903,N_18947,N_19591);
and U22904 (N_22904,N_15954,N_19850);
nand U22905 (N_22905,N_16951,N_17759);
nor U22906 (N_22906,N_17309,N_16103);
or U22907 (N_22907,N_15792,N_17869);
and U22908 (N_22908,N_19125,N_16056);
and U22909 (N_22909,N_16154,N_15234);
nor U22910 (N_22910,N_16597,N_17708);
and U22911 (N_22911,N_19510,N_17816);
nand U22912 (N_22912,N_19814,N_18811);
nand U22913 (N_22913,N_16952,N_15120);
nor U22914 (N_22914,N_18185,N_17301);
nor U22915 (N_22915,N_18264,N_19900);
nand U22916 (N_22916,N_19739,N_17192);
nor U22917 (N_22917,N_18758,N_18258);
xnor U22918 (N_22918,N_17564,N_18618);
nand U22919 (N_22919,N_19762,N_16232);
or U22920 (N_22920,N_18587,N_17519);
nor U22921 (N_22921,N_17595,N_18436);
or U22922 (N_22922,N_15971,N_18371);
and U22923 (N_22923,N_19926,N_15947);
and U22924 (N_22924,N_18524,N_19655);
and U22925 (N_22925,N_18536,N_17049);
nor U22926 (N_22926,N_15841,N_19837);
nor U22927 (N_22927,N_18336,N_16420);
and U22928 (N_22928,N_18991,N_18670);
nand U22929 (N_22929,N_15174,N_19090);
nand U22930 (N_22930,N_19479,N_19798);
and U22931 (N_22931,N_16016,N_17494);
nand U22932 (N_22932,N_17705,N_17784);
nand U22933 (N_22933,N_18295,N_18318);
and U22934 (N_22934,N_17466,N_15089);
nor U22935 (N_22935,N_16244,N_17511);
nor U22936 (N_22936,N_18729,N_16381);
and U22937 (N_22937,N_15548,N_19465);
and U22938 (N_22938,N_18706,N_16262);
nand U22939 (N_22939,N_17343,N_16508);
xnor U22940 (N_22940,N_19634,N_18431);
nor U22941 (N_22941,N_17766,N_18421);
and U22942 (N_22942,N_19076,N_19112);
and U22943 (N_22943,N_18994,N_17047);
or U22944 (N_22944,N_19908,N_17243);
or U22945 (N_22945,N_17991,N_19861);
and U22946 (N_22946,N_17812,N_18783);
nand U22947 (N_22947,N_16970,N_18937);
or U22948 (N_22948,N_16849,N_16999);
or U22949 (N_22949,N_16531,N_15523);
and U22950 (N_22950,N_17399,N_19388);
and U22951 (N_22951,N_18941,N_19931);
or U22952 (N_22952,N_17785,N_18308);
nand U22953 (N_22953,N_18283,N_18722);
nand U22954 (N_22954,N_16204,N_16590);
or U22955 (N_22955,N_15530,N_18954);
or U22956 (N_22956,N_15300,N_18734);
nor U22957 (N_22957,N_17790,N_18530);
nor U22958 (N_22958,N_17308,N_15698);
nand U22959 (N_22959,N_16661,N_19926);
and U22960 (N_22960,N_17675,N_16063);
and U22961 (N_22961,N_19671,N_18498);
xor U22962 (N_22962,N_16052,N_17163);
nand U22963 (N_22963,N_18528,N_18062);
nand U22964 (N_22964,N_17140,N_17711);
or U22965 (N_22965,N_15240,N_15694);
nor U22966 (N_22966,N_17538,N_16904);
and U22967 (N_22967,N_19291,N_16745);
xor U22968 (N_22968,N_18879,N_16366);
nor U22969 (N_22969,N_18847,N_17000);
and U22970 (N_22970,N_18266,N_15715);
nor U22971 (N_22971,N_19066,N_16914);
or U22972 (N_22972,N_16622,N_19296);
and U22973 (N_22973,N_18014,N_15473);
nand U22974 (N_22974,N_15644,N_15733);
or U22975 (N_22975,N_17709,N_15245);
and U22976 (N_22976,N_19772,N_18478);
nand U22977 (N_22977,N_16992,N_18206);
nor U22978 (N_22978,N_16670,N_15145);
or U22979 (N_22979,N_16424,N_15654);
and U22980 (N_22980,N_19550,N_17318);
nand U22981 (N_22981,N_15200,N_15440);
nand U22982 (N_22982,N_16410,N_16498);
nor U22983 (N_22983,N_18687,N_17470);
or U22984 (N_22984,N_16191,N_19979);
nand U22985 (N_22985,N_17245,N_19175);
or U22986 (N_22986,N_17723,N_18416);
nand U22987 (N_22987,N_15038,N_19954);
nand U22988 (N_22988,N_16515,N_18381);
nand U22989 (N_22989,N_16293,N_17565);
or U22990 (N_22990,N_15985,N_17322);
nor U22991 (N_22991,N_18061,N_17115);
and U22992 (N_22992,N_15570,N_18034);
and U22993 (N_22993,N_19733,N_15489);
nand U22994 (N_22994,N_17559,N_16528);
nand U22995 (N_22995,N_16379,N_16415);
nor U22996 (N_22996,N_15944,N_19805);
and U22997 (N_22997,N_15013,N_19554);
and U22998 (N_22998,N_19014,N_18705);
nand U22999 (N_22999,N_17558,N_16241);
and U23000 (N_23000,N_19262,N_15189);
nand U23001 (N_23001,N_15110,N_15544);
nand U23002 (N_23002,N_18668,N_18786);
nor U23003 (N_23003,N_16049,N_15248);
or U23004 (N_23004,N_19974,N_17570);
xor U23005 (N_23005,N_18431,N_15011);
nand U23006 (N_23006,N_16410,N_16097);
nor U23007 (N_23007,N_16021,N_15873);
or U23008 (N_23008,N_18762,N_15790);
or U23009 (N_23009,N_17519,N_18432);
nand U23010 (N_23010,N_19141,N_17766);
and U23011 (N_23011,N_18834,N_19570);
and U23012 (N_23012,N_18917,N_16083);
nor U23013 (N_23013,N_16418,N_15036);
and U23014 (N_23014,N_18937,N_16713);
and U23015 (N_23015,N_15722,N_16929);
or U23016 (N_23016,N_18768,N_18503);
and U23017 (N_23017,N_16156,N_18452);
or U23018 (N_23018,N_15611,N_15535);
nor U23019 (N_23019,N_19970,N_17106);
or U23020 (N_23020,N_15296,N_19956);
and U23021 (N_23021,N_16467,N_18223);
nor U23022 (N_23022,N_15070,N_16374);
or U23023 (N_23023,N_19724,N_16531);
or U23024 (N_23024,N_17410,N_19142);
nand U23025 (N_23025,N_19271,N_16768);
nand U23026 (N_23026,N_15395,N_19056);
and U23027 (N_23027,N_15151,N_18287);
or U23028 (N_23028,N_19896,N_16902);
and U23029 (N_23029,N_19550,N_15259);
nand U23030 (N_23030,N_17684,N_19511);
or U23031 (N_23031,N_18908,N_17037);
nor U23032 (N_23032,N_16589,N_16901);
and U23033 (N_23033,N_17566,N_16762);
nand U23034 (N_23034,N_16541,N_15166);
and U23035 (N_23035,N_17830,N_17411);
nand U23036 (N_23036,N_15697,N_19099);
or U23037 (N_23037,N_19741,N_15680);
and U23038 (N_23038,N_19990,N_18051);
xnor U23039 (N_23039,N_15300,N_15055);
nand U23040 (N_23040,N_18746,N_18697);
nor U23041 (N_23041,N_18929,N_17217);
nor U23042 (N_23042,N_19453,N_17434);
or U23043 (N_23043,N_15650,N_19754);
nor U23044 (N_23044,N_17450,N_17143);
and U23045 (N_23045,N_17288,N_18852);
or U23046 (N_23046,N_18571,N_17382);
nand U23047 (N_23047,N_19169,N_17065);
or U23048 (N_23048,N_15654,N_15208);
nand U23049 (N_23049,N_15721,N_17081);
nor U23050 (N_23050,N_19252,N_19328);
nor U23051 (N_23051,N_15096,N_18056);
and U23052 (N_23052,N_15124,N_15365);
and U23053 (N_23053,N_16703,N_18208);
and U23054 (N_23054,N_16950,N_15297);
xor U23055 (N_23055,N_17214,N_19966);
xnor U23056 (N_23056,N_18767,N_16483);
nand U23057 (N_23057,N_16737,N_16702);
nor U23058 (N_23058,N_15850,N_18582);
nor U23059 (N_23059,N_19643,N_19754);
and U23060 (N_23060,N_15397,N_15722);
and U23061 (N_23061,N_15182,N_15024);
nor U23062 (N_23062,N_17985,N_19396);
nor U23063 (N_23063,N_18338,N_15269);
nand U23064 (N_23064,N_16786,N_15848);
nor U23065 (N_23065,N_15785,N_16850);
xor U23066 (N_23066,N_18214,N_15218);
nand U23067 (N_23067,N_15871,N_17444);
nor U23068 (N_23068,N_18191,N_16132);
nor U23069 (N_23069,N_15358,N_18079);
or U23070 (N_23070,N_15752,N_18559);
or U23071 (N_23071,N_18382,N_19066);
and U23072 (N_23072,N_18545,N_18623);
xnor U23073 (N_23073,N_17498,N_19716);
or U23074 (N_23074,N_17930,N_15766);
and U23075 (N_23075,N_18988,N_16443);
or U23076 (N_23076,N_15469,N_18064);
or U23077 (N_23077,N_19278,N_17026);
nor U23078 (N_23078,N_19659,N_16213);
nand U23079 (N_23079,N_19182,N_17794);
and U23080 (N_23080,N_17019,N_17342);
nand U23081 (N_23081,N_17015,N_17165);
or U23082 (N_23082,N_19030,N_19594);
and U23083 (N_23083,N_16509,N_17923);
nand U23084 (N_23084,N_19239,N_19786);
nand U23085 (N_23085,N_19554,N_18463);
and U23086 (N_23086,N_18906,N_16804);
nor U23087 (N_23087,N_16894,N_15554);
and U23088 (N_23088,N_15851,N_17156);
xor U23089 (N_23089,N_15682,N_18982);
and U23090 (N_23090,N_16473,N_17284);
or U23091 (N_23091,N_18041,N_18645);
nand U23092 (N_23092,N_16273,N_16047);
and U23093 (N_23093,N_18575,N_17222);
and U23094 (N_23094,N_17403,N_15134);
and U23095 (N_23095,N_16616,N_16288);
and U23096 (N_23096,N_19264,N_19328);
and U23097 (N_23097,N_18451,N_15522);
nand U23098 (N_23098,N_16550,N_15746);
nand U23099 (N_23099,N_19999,N_17380);
and U23100 (N_23100,N_17722,N_19760);
and U23101 (N_23101,N_15541,N_15895);
nand U23102 (N_23102,N_19970,N_17672);
nor U23103 (N_23103,N_19349,N_16043);
nor U23104 (N_23104,N_16914,N_19312);
xnor U23105 (N_23105,N_19823,N_19717);
nor U23106 (N_23106,N_17679,N_17331);
and U23107 (N_23107,N_18277,N_17385);
nor U23108 (N_23108,N_18577,N_17943);
nand U23109 (N_23109,N_19700,N_17533);
xnor U23110 (N_23110,N_16754,N_16275);
nor U23111 (N_23111,N_15442,N_15906);
nor U23112 (N_23112,N_19625,N_18277);
nand U23113 (N_23113,N_17134,N_18471);
or U23114 (N_23114,N_18147,N_15850);
or U23115 (N_23115,N_19551,N_19806);
xnor U23116 (N_23116,N_16348,N_19756);
xor U23117 (N_23117,N_19343,N_17924);
nand U23118 (N_23118,N_17187,N_17647);
nand U23119 (N_23119,N_17357,N_19448);
nor U23120 (N_23120,N_17401,N_19361);
and U23121 (N_23121,N_16146,N_16573);
or U23122 (N_23122,N_18000,N_18892);
or U23123 (N_23123,N_18209,N_15721);
or U23124 (N_23124,N_19108,N_16654);
nand U23125 (N_23125,N_19679,N_16642);
nor U23126 (N_23126,N_17544,N_17296);
or U23127 (N_23127,N_16607,N_16107);
xor U23128 (N_23128,N_17792,N_15393);
xor U23129 (N_23129,N_17652,N_17655);
or U23130 (N_23130,N_19307,N_17670);
and U23131 (N_23131,N_15383,N_16008);
nand U23132 (N_23132,N_18157,N_18165);
nor U23133 (N_23133,N_17489,N_18605);
and U23134 (N_23134,N_19384,N_17628);
nand U23135 (N_23135,N_15667,N_19377);
nor U23136 (N_23136,N_15233,N_18636);
nand U23137 (N_23137,N_18528,N_18413);
and U23138 (N_23138,N_16933,N_15933);
or U23139 (N_23139,N_18239,N_19215);
or U23140 (N_23140,N_15013,N_15597);
xor U23141 (N_23141,N_16719,N_16586);
and U23142 (N_23142,N_16325,N_17952);
and U23143 (N_23143,N_15218,N_16055);
nand U23144 (N_23144,N_18681,N_16130);
and U23145 (N_23145,N_16901,N_19857);
nand U23146 (N_23146,N_17235,N_16515);
nand U23147 (N_23147,N_19395,N_15560);
nand U23148 (N_23148,N_19847,N_17460);
and U23149 (N_23149,N_15909,N_18224);
and U23150 (N_23150,N_16141,N_17954);
nand U23151 (N_23151,N_18372,N_17591);
and U23152 (N_23152,N_15250,N_19045);
nand U23153 (N_23153,N_17651,N_16751);
and U23154 (N_23154,N_16699,N_17556);
xor U23155 (N_23155,N_16261,N_15805);
and U23156 (N_23156,N_17510,N_17762);
xnor U23157 (N_23157,N_15271,N_17228);
or U23158 (N_23158,N_19266,N_15624);
or U23159 (N_23159,N_15171,N_15728);
and U23160 (N_23160,N_16975,N_19711);
xnor U23161 (N_23161,N_16980,N_18516);
nand U23162 (N_23162,N_18381,N_19353);
nand U23163 (N_23163,N_15885,N_15706);
or U23164 (N_23164,N_19746,N_19930);
nand U23165 (N_23165,N_17166,N_19510);
nor U23166 (N_23166,N_16216,N_18324);
nand U23167 (N_23167,N_16694,N_17860);
nor U23168 (N_23168,N_17774,N_16603);
or U23169 (N_23169,N_17796,N_15813);
nor U23170 (N_23170,N_19244,N_19866);
nor U23171 (N_23171,N_19619,N_18798);
and U23172 (N_23172,N_19211,N_18650);
or U23173 (N_23173,N_18788,N_15178);
and U23174 (N_23174,N_16587,N_17337);
nor U23175 (N_23175,N_15930,N_19607);
and U23176 (N_23176,N_17943,N_18395);
or U23177 (N_23177,N_15695,N_16368);
nor U23178 (N_23178,N_16458,N_16080);
and U23179 (N_23179,N_17354,N_15110);
and U23180 (N_23180,N_16382,N_19965);
nor U23181 (N_23181,N_15283,N_15904);
nor U23182 (N_23182,N_19971,N_16702);
or U23183 (N_23183,N_16283,N_15897);
nand U23184 (N_23184,N_17134,N_15307);
nor U23185 (N_23185,N_17519,N_18253);
or U23186 (N_23186,N_16946,N_17408);
nand U23187 (N_23187,N_15380,N_19934);
nor U23188 (N_23188,N_15216,N_18743);
or U23189 (N_23189,N_15074,N_19235);
or U23190 (N_23190,N_15793,N_16868);
and U23191 (N_23191,N_15743,N_18214);
nor U23192 (N_23192,N_16873,N_16368);
and U23193 (N_23193,N_19422,N_17082);
and U23194 (N_23194,N_17401,N_18469);
xnor U23195 (N_23195,N_17750,N_17269);
and U23196 (N_23196,N_15543,N_15513);
or U23197 (N_23197,N_15310,N_15280);
and U23198 (N_23198,N_19934,N_18468);
xnor U23199 (N_23199,N_18351,N_18998);
nor U23200 (N_23200,N_19877,N_18077);
nor U23201 (N_23201,N_18173,N_18106);
nand U23202 (N_23202,N_17060,N_17308);
or U23203 (N_23203,N_18079,N_17767);
or U23204 (N_23204,N_18407,N_17774);
nor U23205 (N_23205,N_17194,N_15746);
and U23206 (N_23206,N_17969,N_18030);
nor U23207 (N_23207,N_19973,N_18361);
and U23208 (N_23208,N_15038,N_19874);
or U23209 (N_23209,N_17806,N_19279);
nand U23210 (N_23210,N_17800,N_18861);
xor U23211 (N_23211,N_16475,N_16095);
and U23212 (N_23212,N_17547,N_17083);
or U23213 (N_23213,N_19438,N_16879);
and U23214 (N_23214,N_17322,N_15475);
nand U23215 (N_23215,N_19762,N_17844);
xor U23216 (N_23216,N_15653,N_19759);
nor U23217 (N_23217,N_19407,N_18216);
nor U23218 (N_23218,N_18540,N_19889);
and U23219 (N_23219,N_15986,N_19013);
nand U23220 (N_23220,N_15518,N_17587);
nor U23221 (N_23221,N_15889,N_19032);
or U23222 (N_23222,N_15493,N_15968);
nand U23223 (N_23223,N_18884,N_19505);
or U23224 (N_23224,N_19848,N_18568);
or U23225 (N_23225,N_17196,N_18096);
and U23226 (N_23226,N_16718,N_19945);
nand U23227 (N_23227,N_17597,N_17606);
and U23228 (N_23228,N_17913,N_15175);
xor U23229 (N_23229,N_17881,N_16689);
nand U23230 (N_23230,N_19745,N_17823);
and U23231 (N_23231,N_19288,N_18170);
nand U23232 (N_23232,N_18156,N_19821);
and U23233 (N_23233,N_17910,N_16349);
and U23234 (N_23234,N_16376,N_15631);
nand U23235 (N_23235,N_17076,N_16341);
nor U23236 (N_23236,N_17679,N_19217);
nor U23237 (N_23237,N_16749,N_19187);
and U23238 (N_23238,N_17758,N_16719);
or U23239 (N_23239,N_18781,N_17172);
and U23240 (N_23240,N_16153,N_15621);
nor U23241 (N_23241,N_18574,N_15783);
or U23242 (N_23242,N_15319,N_16982);
or U23243 (N_23243,N_16569,N_15084);
nor U23244 (N_23244,N_17408,N_18676);
xnor U23245 (N_23245,N_15770,N_17627);
or U23246 (N_23246,N_17947,N_15004);
nand U23247 (N_23247,N_16370,N_19135);
or U23248 (N_23248,N_18818,N_15946);
xor U23249 (N_23249,N_18582,N_19638);
nand U23250 (N_23250,N_18269,N_17759);
or U23251 (N_23251,N_17437,N_15579);
or U23252 (N_23252,N_16753,N_18773);
xor U23253 (N_23253,N_15463,N_19218);
and U23254 (N_23254,N_17629,N_19752);
and U23255 (N_23255,N_17280,N_19121);
xnor U23256 (N_23256,N_15574,N_15788);
or U23257 (N_23257,N_16917,N_19095);
nor U23258 (N_23258,N_19808,N_19371);
or U23259 (N_23259,N_18634,N_19804);
and U23260 (N_23260,N_18691,N_19472);
or U23261 (N_23261,N_18637,N_16657);
or U23262 (N_23262,N_18168,N_16238);
nand U23263 (N_23263,N_19445,N_19261);
nor U23264 (N_23264,N_19725,N_16902);
nor U23265 (N_23265,N_16534,N_15043);
nand U23266 (N_23266,N_15812,N_19213);
nor U23267 (N_23267,N_19949,N_19057);
xor U23268 (N_23268,N_17245,N_15922);
or U23269 (N_23269,N_15086,N_15646);
nor U23270 (N_23270,N_15013,N_16426);
nand U23271 (N_23271,N_18324,N_15471);
nand U23272 (N_23272,N_17592,N_16437);
nand U23273 (N_23273,N_19643,N_18728);
nor U23274 (N_23274,N_19623,N_17496);
or U23275 (N_23275,N_19824,N_15048);
nor U23276 (N_23276,N_16635,N_17505);
nand U23277 (N_23277,N_19554,N_17566);
xor U23278 (N_23278,N_17991,N_17054);
nand U23279 (N_23279,N_17157,N_18588);
xor U23280 (N_23280,N_19298,N_17807);
or U23281 (N_23281,N_19354,N_16252);
nand U23282 (N_23282,N_17546,N_16884);
nor U23283 (N_23283,N_17646,N_18876);
nor U23284 (N_23284,N_15082,N_17046);
nor U23285 (N_23285,N_18259,N_17046);
nand U23286 (N_23286,N_18044,N_15661);
xnor U23287 (N_23287,N_17951,N_17936);
nor U23288 (N_23288,N_18538,N_17207);
xnor U23289 (N_23289,N_16004,N_17054);
nor U23290 (N_23290,N_16594,N_15050);
nand U23291 (N_23291,N_15799,N_15495);
nand U23292 (N_23292,N_17419,N_17502);
or U23293 (N_23293,N_16707,N_19395);
xor U23294 (N_23294,N_17091,N_17563);
nor U23295 (N_23295,N_19003,N_19207);
xnor U23296 (N_23296,N_17582,N_19829);
or U23297 (N_23297,N_19732,N_17884);
or U23298 (N_23298,N_15126,N_15751);
xnor U23299 (N_23299,N_15644,N_18373);
nand U23300 (N_23300,N_16588,N_17444);
and U23301 (N_23301,N_16135,N_15186);
nand U23302 (N_23302,N_18902,N_17903);
or U23303 (N_23303,N_18753,N_19837);
nor U23304 (N_23304,N_15884,N_17995);
and U23305 (N_23305,N_18107,N_17037);
or U23306 (N_23306,N_16554,N_19644);
and U23307 (N_23307,N_19267,N_16541);
or U23308 (N_23308,N_19530,N_18119);
and U23309 (N_23309,N_19862,N_17399);
nand U23310 (N_23310,N_17707,N_15073);
or U23311 (N_23311,N_18667,N_16264);
and U23312 (N_23312,N_19415,N_19134);
nor U23313 (N_23313,N_16980,N_17788);
nor U23314 (N_23314,N_16194,N_17980);
and U23315 (N_23315,N_16920,N_16535);
or U23316 (N_23316,N_16935,N_19941);
nor U23317 (N_23317,N_17870,N_16247);
or U23318 (N_23318,N_16057,N_16113);
nor U23319 (N_23319,N_17076,N_17798);
xor U23320 (N_23320,N_15422,N_18670);
or U23321 (N_23321,N_16647,N_17293);
nand U23322 (N_23322,N_15499,N_18794);
or U23323 (N_23323,N_17869,N_15823);
or U23324 (N_23324,N_15822,N_17880);
nor U23325 (N_23325,N_19787,N_17043);
and U23326 (N_23326,N_17392,N_18039);
or U23327 (N_23327,N_16562,N_19397);
nor U23328 (N_23328,N_16310,N_15192);
nor U23329 (N_23329,N_18552,N_19379);
xnor U23330 (N_23330,N_19281,N_15753);
or U23331 (N_23331,N_15068,N_15890);
nor U23332 (N_23332,N_19268,N_15248);
nand U23333 (N_23333,N_18657,N_17364);
or U23334 (N_23334,N_19438,N_19032);
nand U23335 (N_23335,N_15748,N_19604);
or U23336 (N_23336,N_18561,N_18027);
or U23337 (N_23337,N_16688,N_17130);
or U23338 (N_23338,N_18432,N_17638);
nand U23339 (N_23339,N_15586,N_15701);
and U23340 (N_23340,N_15018,N_16089);
xnor U23341 (N_23341,N_19048,N_18109);
nor U23342 (N_23342,N_18772,N_17933);
xor U23343 (N_23343,N_15366,N_15791);
or U23344 (N_23344,N_18003,N_17235);
and U23345 (N_23345,N_15513,N_18398);
and U23346 (N_23346,N_19982,N_15622);
and U23347 (N_23347,N_16986,N_17025);
nor U23348 (N_23348,N_18805,N_17254);
xnor U23349 (N_23349,N_16349,N_18157);
or U23350 (N_23350,N_17310,N_18818);
nor U23351 (N_23351,N_18363,N_18195);
or U23352 (N_23352,N_18210,N_18473);
or U23353 (N_23353,N_18306,N_17996);
nand U23354 (N_23354,N_19763,N_16068);
xor U23355 (N_23355,N_18777,N_15829);
xnor U23356 (N_23356,N_15473,N_19653);
and U23357 (N_23357,N_16150,N_18260);
or U23358 (N_23358,N_16142,N_17603);
or U23359 (N_23359,N_18835,N_15478);
nor U23360 (N_23360,N_17902,N_17681);
nand U23361 (N_23361,N_19310,N_16123);
nor U23362 (N_23362,N_17140,N_17404);
and U23363 (N_23363,N_15951,N_19146);
nor U23364 (N_23364,N_15805,N_15316);
xor U23365 (N_23365,N_16177,N_16520);
nand U23366 (N_23366,N_18914,N_19226);
and U23367 (N_23367,N_19623,N_15635);
nand U23368 (N_23368,N_17335,N_17187);
xor U23369 (N_23369,N_15984,N_18218);
nor U23370 (N_23370,N_19748,N_16298);
and U23371 (N_23371,N_17129,N_16975);
or U23372 (N_23372,N_19418,N_15509);
nand U23373 (N_23373,N_16208,N_16533);
xnor U23374 (N_23374,N_17642,N_16119);
or U23375 (N_23375,N_19162,N_17204);
or U23376 (N_23376,N_16430,N_18766);
or U23377 (N_23377,N_17914,N_16912);
nand U23378 (N_23378,N_17234,N_16675);
nor U23379 (N_23379,N_18009,N_19248);
and U23380 (N_23380,N_19354,N_18637);
xnor U23381 (N_23381,N_16353,N_17369);
xor U23382 (N_23382,N_19684,N_19620);
nand U23383 (N_23383,N_17668,N_15405);
xor U23384 (N_23384,N_17576,N_19156);
nor U23385 (N_23385,N_16803,N_16509);
nand U23386 (N_23386,N_19858,N_18183);
or U23387 (N_23387,N_17369,N_16678);
or U23388 (N_23388,N_16797,N_16795);
nand U23389 (N_23389,N_16342,N_17809);
and U23390 (N_23390,N_17192,N_18318);
or U23391 (N_23391,N_19234,N_19421);
or U23392 (N_23392,N_18530,N_18896);
xnor U23393 (N_23393,N_19603,N_16227);
or U23394 (N_23394,N_17055,N_19282);
xnor U23395 (N_23395,N_19474,N_17012);
or U23396 (N_23396,N_18488,N_18778);
xnor U23397 (N_23397,N_15544,N_16625);
xor U23398 (N_23398,N_19566,N_18929);
and U23399 (N_23399,N_15916,N_18593);
xnor U23400 (N_23400,N_15445,N_17047);
nor U23401 (N_23401,N_15178,N_19299);
and U23402 (N_23402,N_18170,N_19975);
or U23403 (N_23403,N_17450,N_19754);
or U23404 (N_23404,N_15127,N_15881);
nand U23405 (N_23405,N_16548,N_18856);
xor U23406 (N_23406,N_17325,N_18368);
nand U23407 (N_23407,N_19459,N_17336);
and U23408 (N_23408,N_17119,N_15026);
xnor U23409 (N_23409,N_16381,N_15259);
and U23410 (N_23410,N_16339,N_19801);
nand U23411 (N_23411,N_17190,N_19523);
nor U23412 (N_23412,N_15620,N_17970);
nand U23413 (N_23413,N_15489,N_19478);
nand U23414 (N_23414,N_18229,N_19899);
nor U23415 (N_23415,N_15764,N_15678);
and U23416 (N_23416,N_18002,N_19092);
or U23417 (N_23417,N_18930,N_15485);
and U23418 (N_23418,N_16817,N_15708);
nor U23419 (N_23419,N_15486,N_16014);
and U23420 (N_23420,N_19825,N_16118);
nor U23421 (N_23421,N_15439,N_18089);
nor U23422 (N_23422,N_19916,N_16244);
or U23423 (N_23423,N_16254,N_19425);
xor U23424 (N_23424,N_16332,N_19848);
nor U23425 (N_23425,N_15076,N_16977);
and U23426 (N_23426,N_16546,N_17446);
or U23427 (N_23427,N_17696,N_15458);
or U23428 (N_23428,N_18723,N_16703);
nor U23429 (N_23429,N_18847,N_18474);
and U23430 (N_23430,N_19670,N_17389);
nor U23431 (N_23431,N_17088,N_17354);
xnor U23432 (N_23432,N_19533,N_16116);
and U23433 (N_23433,N_16937,N_15032);
and U23434 (N_23434,N_16836,N_18445);
xnor U23435 (N_23435,N_17595,N_15979);
and U23436 (N_23436,N_17169,N_15921);
xnor U23437 (N_23437,N_15035,N_18851);
or U23438 (N_23438,N_17103,N_15994);
nor U23439 (N_23439,N_15122,N_16349);
or U23440 (N_23440,N_18044,N_18009);
nor U23441 (N_23441,N_15519,N_16342);
and U23442 (N_23442,N_17912,N_19790);
and U23443 (N_23443,N_18143,N_18941);
xnor U23444 (N_23444,N_16606,N_15778);
nor U23445 (N_23445,N_16636,N_19264);
or U23446 (N_23446,N_15590,N_19187);
nor U23447 (N_23447,N_15367,N_19494);
nor U23448 (N_23448,N_18681,N_16014);
or U23449 (N_23449,N_16873,N_18218);
or U23450 (N_23450,N_19111,N_18124);
nand U23451 (N_23451,N_16713,N_15310);
and U23452 (N_23452,N_18332,N_17393);
nor U23453 (N_23453,N_17143,N_17292);
nand U23454 (N_23454,N_16055,N_18471);
nand U23455 (N_23455,N_16966,N_15326);
nor U23456 (N_23456,N_18926,N_15691);
nor U23457 (N_23457,N_18513,N_19920);
nor U23458 (N_23458,N_19765,N_16023);
nand U23459 (N_23459,N_17123,N_18057);
nand U23460 (N_23460,N_17730,N_19167);
nor U23461 (N_23461,N_19687,N_19974);
or U23462 (N_23462,N_19058,N_15524);
and U23463 (N_23463,N_17434,N_19404);
nand U23464 (N_23464,N_18953,N_17179);
and U23465 (N_23465,N_16383,N_19609);
or U23466 (N_23466,N_17863,N_18271);
xor U23467 (N_23467,N_18186,N_15188);
or U23468 (N_23468,N_18969,N_18067);
nor U23469 (N_23469,N_18883,N_18470);
nor U23470 (N_23470,N_18433,N_15743);
nand U23471 (N_23471,N_18749,N_18260);
or U23472 (N_23472,N_18501,N_19192);
nor U23473 (N_23473,N_15735,N_17721);
or U23474 (N_23474,N_19770,N_18808);
and U23475 (N_23475,N_17558,N_18989);
nor U23476 (N_23476,N_15954,N_19569);
nand U23477 (N_23477,N_18136,N_18661);
nand U23478 (N_23478,N_16275,N_16042);
nor U23479 (N_23479,N_16301,N_16198);
nor U23480 (N_23480,N_16192,N_15684);
xnor U23481 (N_23481,N_15004,N_18548);
and U23482 (N_23482,N_17470,N_16189);
nor U23483 (N_23483,N_15727,N_19985);
and U23484 (N_23484,N_17533,N_16026);
and U23485 (N_23485,N_17442,N_18641);
or U23486 (N_23486,N_18015,N_19677);
nand U23487 (N_23487,N_16501,N_17186);
or U23488 (N_23488,N_19053,N_15868);
or U23489 (N_23489,N_18808,N_15195);
nor U23490 (N_23490,N_18161,N_16186);
or U23491 (N_23491,N_18014,N_19143);
xor U23492 (N_23492,N_17662,N_17792);
nand U23493 (N_23493,N_17942,N_15283);
nand U23494 (N_23494,N_15503,N_17957);
nand U23495 (N_23495,N_17110,N_15029);
nand U23496 (N_23496,N_15982,N_15505);
or U23497 (N_23497,N_15474,N_19644);
or U23498 (N_23498,N_16982,N_15740);
nand U23499 (N_23499,N_16062,N_15126);
or U23500 (N_23500,N_17510,N_19066);
nand U23501 (N_23501,N_15086,N_17207);
nor U23502 (N_23502,N_18123,N_17403);
or U23503 (N_23503,N_19381,N_18994);
xnor U23504 (N_23504,N_17286,N_19239);
or U23505 (N_23505,N_19440,N_15290);
or U23506 (N_23506,N_19046,N_17052);
xor U23507 (N_23507,N_16066,N_19109);
nor U23508 (N_23508,N_19082,N_19206);
and U23509 (N_23509,N_18283,N_15865);
nand U23510 (N_23510,N_17527,N_18367);
nor U23511 (N_23511,N_16497,N_19594);
nor U23512 (N_23512,N_18293,N_18434);
nand U23513 (N_23513,N_19765,N_15080);
nand U23514 (N_23514,N_15720,N_16344);
nand U23515 (N_23515,N_18248,N_19943);
nand U23516 (N_23516,N_18181,N_19328);
and U23517 (N_23517,N_19031,N_18499);
nor U23518 (N_23518,N_18558,N_15371);
nor U23519 (N_23519,N_18104,N_18820);
or U23520 (N_23520,N_17872,N_15518);
nand U23521 (N_23521,N_17162,N_17009);
nor U23522 (N_23522,N_18304,N_17060);
nand U23523 (N_23523,N_16997,N_17286);
nor U23524 (N_23524,N_18481,N_15460);
nor U23525 (N_23525,N_18230,N_15231);
and U23526 (N_23526,N_16862,N_17399);
or U23527 (N_23527,N_19862,N_16200);
and U23528 (N_23528,N_19402,N_18266);
nand U23529 (N_23529,N_16408,N_16776);
nand U23530 (N_23530,N_18475,N_18708);
or U23531 (N_23531,N_17368,N_18740);
or U23532 (N_23532,N_16714,N_19030);
nand U23533 (N_23533,N_15161,N_18148);
nand U23534 (N_23534,N_18586,N_19567);
nand U23535 (N_23535,N_19931,N_16763);
xor U23536 (N_23536,N_15002,N_19296);
and U23537 (N_23537,N_18801,N_17063);
xor U23538 (N_23538,N_15225,N_18567);
and U23539 (N_23539,N_18359,N_15348);
or U23540 (N_23540,N_19910,N_16907);
and U23541 (N_23541,N_15520,N_15757);
nand U23542 (N_23542,N_16691,N_15939);
xor U23543 (N_23543,N_17219,N_19352);
xor U23544 (N_23544,N_18396,N_16672);
xnor U23545 (N_23545,N_18384,N_16175);
or U23546 (N_23546,N_18580,N_16732);
or U23547 (N_23547,N_18831,N_15751);
nor U23548 (N_23548,N_19540,N_17817);
nand U23549 (N_23549,N_18575,N_19056);
nor U23550 (N_23550,N_17569,N_17119);
nand U23551 (N_23551,N_18045,N_15661);
or U23552 (N_23552,N_16697,N_17803);
xor U23553 (N_23553,N_18227,N_17884);
xnor U23554 (N_23554,N_16024,N_16272);
nand U23555 (N_23555,N_16526,N_17289);
nor U23556 (N_23556,N_17756,N_19726);
or U23557 (N_23557,N_18992,N_16085);
nand U23558 (N_23558,N_16642,N_15244);
and U23559 (N_23559,N_15008,N_18436);
and U23560 (N_23560,N_15074,N_19906);
or U23561 (N_23561,N_15127,N_15913);
nor U23562 (N_23562,N_19051,N_18954);
and U23563 (N_23563,N_18486,N_19264);
and U23564 (N_23564,N_17556,N_19266);
nor U23565 (N_23565,N_17818,N_18076);
nor U23566 (N_23566,N_18572,N_18994);
or U23567 (N_23567,N_19582,N_16669);
xnor U23568 (N_23568,N_18840,N_16461);
or U23569 (N_23569,N_18586,N_19214);
nor U23570 (N_23570,N_19712,N_17331);
nor U23571 (N_23571,N_16017,N_16145);
and U23572 (N_23572,N_15520,N_17441);
nand U23573 (N_23573,N_15050,N_19866);
nor U23574 (N_23574,N_19399,N_19169);
nor U23575 (N_23575,N_16825,N_16646);
or U23576 (N_23576,N_15102,N_18460);
and U23577 (N_23577,N_17704,N_19486);
and U23578 (N_23578,N_15984,N_18930);
nor U23579 (N_23579,N_19628,N_16126);
and U23580 (N_23580,N_19887,N_15034);
or U23581 (N_23581,N_18656,N_16860);
xnor U23582 (N_23582,N_15790,N_19957);
or U23583 (N_23583,N_15666,N_15293);
and U23584 (N_23584,N_15232,N_16916);
nand U23585 (N_23585,N_16443,N_17342);
or U23586 (N_23586,N_15424,N_15953);
or U23587 (N_23587,N_19943,N_15385);
nor U23588 (N_23588,N_18655,N_17519);
nor U23589 (N_23589,N_18771,N_19569);
and U23590 (N_23590,N_19600,N_19703);
nand U23591 (N_23591,N_18935,N_16714);
nor U23592 (N_23592,N_19876,N_15187);
or U23593 (N_23593,N_19219,N_16656);
and U23594 (N_23594,N_19244,N_19705);
xor U23595 (N_23595,N_15343,N_19245);
nor U23596 (N_23596,N_18402,N_15212);
or U23597 (N_23597,N_17384,N_15043);
or U23598 (N_23598,N_15497,N_16180);
xor U23599 (N_23599,N_15392,N_19846);
nor U23600 (N_23600,N_17722,N_16175);
or U23601 (N_23601,N_15670,N_18340);
or U23602 (N_23602,N_16454,N_16217);
and U23603 (N_23603,N_19853,N_18401);
and U23604 (N_23604,N_15955,N_15095);
xor U23605 (N_23605,N_18677,N_18927);
or U23606 (N_23606,N_18641,N_15528);
or U23607 (N_23607,N_19200,N_17129);
xnor U23608 (N_23608,N_19750,N_15106);
and U23609 (N_23609,N_15257,N_15110);
or U23610 (N_23610,N_18027,N_17975);
xor U23611 (N_23611,N_18610,N_18193);
and U23612 (N_23612,N_17788,N_19830);
nand U23613 (N_23613,N_15884,N_15616);
and U23614 (N_23614,N_19123,N_18995);
xnor U23615 (N_23615,N_15970,N_16767);
and U23616 (N_23616,N_17101,N_16091);
nand U23617 (N_23617,N_19609,N_15867);
nor U23618 (N_23618,N_17056,N_16683);
nand U23619 (N_23619,N_19326,N_16238);
and U23620 (N_23620,N_15989,N_15385);
and U23621 (N_23621,N_19438,N_17362);
nand U23622 (N_23622,N_17648,N_15040);
and U23623 (N_23623,N_15864,N_19152);
nor U23624 (N_23624,N_15908,N_15039);
xor U23625 (N_23625,N_15947,N_17013);
or U23626 (N_23626,N_16171,N_19805);
or U23627 (N_23627,N_18565,N_16978);
xnor U23628 (N_23628,N_18147,N_16555);
nand U23629 (N_23629,N_17031,N_19326);
or U23630 (N_23630,N_17699,N_16967);
nor U23631 (N_23631,N_19748,N_15728);
nand U23632 (N_23632,N_15835,N_15609);
and U23633 (N_23633,N_17445,N_17126);
xnor U23634 (N_23634,N_18762,N_19238);
xnor U23635 (N_23635,N_17040,N_17045);
nand U23636 (N_23636,N_16619,N_19900);
or U23637 (N_23637,N_16397,N_15997);
and U23638 (N_23638,N_18508,N_17320);
and U23639 (N_23639,N_16061,N_19056);
and U23640 (N_23640,N_16341,N_18029);
and U23641 (N_23641,N_17572,N_19470);
or U23642 (N_23642,N_16820,N_15815);
xnor U23643 (N_23643,N_17353,N_15850);
or U23644 (N_23644,N_19047,N_18375);
xor U23645 (N_23645,N_19267,N_16324);
and U23646 (N_23646,N_17804,N_15158);
nor U23647 (N_23647,N_18860,N_15348);
and U23648 (N_23648,N_16868,N_17598);
nor U23649 (N_23649,N_15095,N_16745);
or U23650 (N_23650,N_16537,N_16792);
xor U23651 (N_23651,N_19633,N_19973);
nor U23652 (N_23652,N_17253,N_15642);
and U23653 (N_23653,N_17860,N_19058);
nand U23654 (N_23654,N_15797,N_17807);
nand U23655 (N_23655,N_18411,N_17960);
nor U23656 (N_23656,N_18907,N_15653);
or U23657 (N_23657,N_19681,N_15495);
and U23658 (N_23658,N_19667,N_19073);
xor U23659 (N_23659,N_18200,N_17775);
nand U23660 (N_23660,N_18564,N_17882);
nor U23661 (N_23661,N_19259,N_19883);
and U23662 (N_23662,N_17469,N_18146);
xnor U23663 (N_23663,N_17322,N_17613);
nand U23664 (N_23664,N_17993,N_19425);
nand U23665 (N_23665,N_18327,N_19533);
nand U23666 (N_23666,N_17139,N_15013);
or U23667 (N_23667,N_19358,N_15475);
or U23668 (N_23668,N_18149,N_17230);
and U23669 (N_23669,N_16669,N_19130);
and U23670 (N_23670,N_17736,N_16501);
xnor U23671 (N_23671,N_15704,N_18055);
and U23672 (N_23672,N_19095,N_17680);
nor U23673 (N_23673,N_16261,N_16354);
or U23674 (N_23674,N_16677,N_16298);
nand U23675 (N_23675,N_18868,N_18730);
nand U23676 (N_23676,N_16095,N_17654);
nand U23677 (N_23677,N_18818,N_19953);
xor U23678 (N_23678,N_19957,N_18948);
or U23679 (N_23679,N_18798,N_19431);
or U23680 (N_23680,N_18243,N_17887);
or U23681 (N_23681,N_19204,N_17430);
nor U23682 (N_23682,N_15168,N_19823);
or U23683 (N_23683,N_17575,N_16453);
xor U23684 (N_23684,N_16281,N_18055);
or U23685 (N_23685,N_19684,N_15632);
or U23686 (N_23686,N_16425,N_15723);
and U23687 (N_23687,N_15143,N_15964);
and U23688 (N_23688,N_16566,N_15926);
and U23689 (N_23689,N_16263,N_17817);
or U23690 (N_23690,N_15574,N_15105);
or U23691 (N_23691,N_18349,N_18166);
or U23692 (N_23692,N_15450,N_19713);
nand U23693 (N_23693,N_17603,N_18107);
and U23694 (N_23694,N_15596,N_19702);
and U23695 (N_23695,N_19994,N_18492);
or U23696 (N_23696,N_16815,N_17927);
nor U23697 (N_23697,N_15417,N_19509);
nand U23698 (N_23698,N_17018,N_16838);
nor U23699 (N_23699,N_17878,N_17584);
and U23700 (N_23700,N_19673,N_15602);
or U23701 (N_23701,N_19631,N_18022);
or U23702 (N_23702,N_18901,N_15552);
nand U23703 (N_23703,N_15277,N_17654);
nand U23704 (N_23704,N_15230,N_19921);
nor U23705 (N_23705,N_15938,N_15516);
nand U23706 (N_23706,N_16122,N_18835);
xor U23707 (N_23707,N_19760,N_19030);
nand U23708 (N_23708,N_16841,N_18858);
nor U23709 (N_23709,N_16004,N_17122);
nand U23710 (N_23710,N_18647,N_17799);
nor U23711 (N_23711,N_16189,N_19508);
nor U23712 (N_23712,N_19615,N_18380);
and U23713 (N_23713,N_18449,N_16547);
nor U23714 (N_23714,N_15320,N_18693);
nand U23715 (N_23715,N_16169,N_17215);
nor U23716 (N_23716,N_16688,N_16278);
nor U23717 (N_23717,N_16096,N_15757);
nand U23718 (N_23718,N_19905,N_16162);
nand U23719 (N_23719,N_16830,N_19725);
and U23720 (N_23720,N_18588,N_17043);
and U23721 (N_23721,N_18856,N_18022);
xnor U23722 (N_23722,N_17701,N_19943);
and U23723 (N_23723,N_19611,N_18597);
nor U23724 (N_23724,N_18917,N_18688);
xor U23725 (N_23725,N_19402,N_15727);
nor U23726 (N_23726,N_17208,N_16834);
nand U23727 (N_23727,N_18744,N_17543);
nor U23728 (N_23728,N_15467,N_19034);
nand U23729 (N_23729,N_17463,N_16476);
nand U23730 (N_23730,N_19928,N_16086);
or U23731 (N_23731,N_18537,N_16564);
nand U23732 (N_23732,N_19871,N_15013);
and U23733 (N_23733,N_18494,N_16201);
or U23734 (N_23734,N_16705,N_15473);
xnor U23735 (N_23735,N_17529,N_18444);
nor U23736 (N_23736,N_16793,N_17282);
or U23737 (N_23737,N_16916,N_18225);
nor U23738 (N_23738,N_17865,N_17800);
or U23739 (N_23739,N_17467,N_17943);
nand U23740 (N_23740,N_16109,N_18568);
or U23741 (N_23741,N_17991,N_19366);
and U23742 (N_23742,N_15932,N_16269);
nor U23743 (N_23743,N_16472,N_18822);
and U23744 (N_23744,N_17659,N_17725);
nand U23745 (N_23745,N_18175,N_17042);
nor U23746 (N_23746,N_19384,N_15748);
nand U23747 (N_23747,N_15363,N_19374);
nor U23748 (N_23748,N_16250,N_17698);
nor U23749 (N_23749,N_16451,N_19070);
nor U23750 (N_23750,N_15579,N_19840);
and U23751 (N_23751,N_19919,N_15481);
nand U23752 (N_23752,N_17064,N_17840);
or U23753 (N_23753,N_18908,N_19084);
or U23754 (N_23754,N_16205,N_19318);
or U23755 (N_23755,N_17661,N_18089);
and U23756 (N_23756,N_17744,N_16994);
xor U23757 (N_23757,N_16609,N_16916);
nor U23758 (N_23758,N_18053,N_18192);
nand U23759 (N_23759,N_15559,N_17193);
or U23760 (N_23760,N_16835,N_17154);
nor U23761 (N_23761,N_16661,N_17426);
or U23762 (N_23762,N_16552,N_16693);
nand U23763 (N_23763,N_15302,N_16588);
nand U23764 (N_23764,N_18579,N_15010);
nor U23765 (N_23765,N_17621,N_15139);
xor U23766 (N_23766,N_16600,N_19216);
nor U23767 (N_23767,N_17292,N_15834);
or U23768 (N_23768,N_18075,N_16297);
and U23769 (N_23769,N_19889,N_19286);
or U23770 (N_23770,N_19121,N_17227);
nor U23771 (N_23771,N_15128,N_19831);
nand U23772 (N_23772,N_17030,N_17461);
and U23773 (N_23773,N_19559,N_17594);
xnor U23774 (N_23774,N_17217,N_17297);
or U23775 (N_23775,N_18782,N_16213);
xor U23776 (N_23776,N_18574,N_18597);
and U23777 (N_23777,N_15148,N_18828);
or U23778 (N_23778,N_16204,N_15863);
or U23779 (N_23779,N_16525,N_19784);
nor U23780 (N_23780,N_17336,N_16449);
nand U23781 (N_23781,N_17781,N_15516);
nand U23782 (N_23782,N_19174,N_19217);
nand U23783 (N_23783,N_18317,N_15485);
nand U23784 (N_23784,N_17181,N_18378);
and U23785 (N_23785,N_16328,N_16185);
xnor U23786 (N_23786,N_17071,N_18777);
nand U23787 (N_23787,N_18804,N_17956);
xnor U23788 (N_23788,N_18594,N_16954);
xnor U23789 (N_23789,N_19400,N_17642);
or U23790 (N_23790,N_18614,N_17513);
xnor U23791 (N_23791,N_15004,N_15415);
and U23792 (N_23792,N_19293,N_19442);
xor U23793 (N_23793,N_19474,N_18014);
nand U23794 (N_23794,N_19448,N_19690);
and U23795 (N_23795,N_16765,N_19562);
nor U23796 (N_23796,N_17092,N_15321);
xnor U23797 (N_23797,N_17381,N_17351);
nor U23798 (N_23798,N_15829,N_15516);
nand U23799 (N_23799,N_17193,N_19606);
nor U23800 (N_23800,N_18958,N_16994);
and U23801 (N_23801,N_18301,N_19568);
nand U23802 (N_23802,N_17233,N_19967);
xnor U23803 (N_23803,N_18727,N_16765);
nand U23804 (N_23804,N_15058,N_15183);
and U23805 (N_23805,N_19837,N_15378);
xnor U23806 (N_23806,N_16891,N_16602);
and U23807 (N_23807,N_16394,N_17003);
nor U23808 (N_23808,N_15695,N_15178);
nand U23809 (N_23809,N_16610,N_16644);
xnor U23810 (N_23810,N_15129,N_16562);
nand U23811 (N_23811,N_17561,N_17388);
nand U23812 (N_23812,N_15887,N_16935);
nor U23813 (N_23813,N_16359,N_16990);
nor U23814 (N_23814,N_17367,N_16808);
and U23815 (N_23815,N_18438,N_19545);
xor U23816 (N_23816,N_17126,N_16053);
nand U23817 (N_23817,N_15463,N_18614);
xor U23818 (N_23818,N_19017,N_18334);
nor U23819 (N_23819,N_19271,N_15677);
and U23820 (N_23820,N_16268,N_19919);
and U23821 (N_23821,N_17494,N_19665);
nor U23822 (N_23822,N_16422,N_15647);
and U23823 (N_23823,N_16823,N_15237);
nor U23824 (N_23824,N_15511,N_19483);
nand U23825 (N_23825,N_18280,N_15174);
and U23826 (N_23826,N_18275,N_19861);
or U23827 (N_23827,N_16532,N_16158);
nor U23828 (N_23828,N_18088,N_17995);
nand U23829 (N_23829,N_17852,N_19488);
or U23830 (N_23830,N_17623,N_18297);
and U23831 (N_23831,N_15098,N_16742);
nand U23832 (N_23832,N_16173,N_18122);
and U23833 (N_23833,N_19539,N_16675);
and U23834 (N_23834,N_19042,N_16289);
nand U23835 (N_23835,N_18664,N_19062);
or U23836 (N_23836,N_18744,N_15080);
nand U23837 (N_23837,N_16649,N_18242);
or U23838 (N_23838,N_19714,N_19254);
and U23839 (N_23839,N_18190,N_16075);
and U23840 (N_23840,N_18531,N_19426);
and U23841 (N_23841,N_17660,N_17912);
nor U23842 (N_23842,N_16782,N_16799);
and U23843 (N_23843,N_17588,N_19672);
and U23844 (N_23844,N_19958,N_19115);
nand U23845 (N_23845,N_15497,N_19366);
or U23846 (N_23846,N_17865,N_19964);
nor U23847 (N_23847,N_19995,N_19155);
nand U23848 (N_23848,N_15669,N_19003);
or U23849 (N_23849,N_17253,N_18938);
nor U23850 (N_23850,N_17888,N_18004);
nor U23851 (N_23851,N_15314,N_16186);
and U23852 (N_23852,N_19741,N_19715);
and U23853 (N_23853,N_16003,N_18041);
xnor U23854 (N_23854,N_17163,N_15802);
xnor U23855 (N_23855,N_16006,N_15128);
nor U23856 (N_23856,N_16115,N_19332);
and U23857 (N_23857,N_17168,N_17955);
nor U23858 (N_23858,N_17376,N_19308);
or U23859 (N_23859,N_17145,N_16708);
nor U23860 (N_23860,N_16499,N_17831);
nor U23861 (N_23861,N_17049,N_19529);
or U23862 (N_23862,N_18767,N_16001);
nor U23863 (N_23863,N_15515,N_15960);
nor U23864 (N_23864,N_18857,N_15894);
nand U23865 (N_23865,N_15993,N_19195);
or U23866 (N_23866,N_15489,N_18201);
and U23867 (N_23867,N_18055,N_17305);
or U23868 (N_23868,N_19124,N_17536);
nand U23869 (N_23869,N_18739,N_18067);
xor U23870 (N_23870,N_16927,N_17300);
nand U23871 (N_23871,N_17435,N_18434);
nand U23872 (N_23872,N_19567,N_17606);
and U23873 (N_23873,N_16382,N_19314);
nand U23874 (N_23874,N_18532,N_19357);
xnor U23875 (N_23875,N_16323,N_19548);
and U23876 (N_23876,N_16647,N_18798);
or U23877 (N_23877,N_15121,N_16681);
or U23878 (N_23878,N_19747,N_19595);
nor U23879 (N_23879,N_19797,N_18160);
nor U23880 (N_23880,N_15959,N_16815);
nor U23881 (N_23881,N_18682,N_17631);
and U23882 (N_23882,N_16685,N_16801);
xor U23883 (N_23883,N_15639,N_16510);
xor U23884 (N_23884,N_18319,N_19683);
and U23885 (N_23885,N_18704,N_18810);
nand U23886 (N_23886,N_16956,N_18528);
and U23887 (N_23887,N_17714,N_15449);
or U23888 (N_23888,N_16957,N_16093);
nand U23889 (N_23889,N_15338,N_15552);
and U23890 (N_23890,N_18377,N_16277);
or U23891 (N_23891,N_19677,N_15936);
nor U23892 (N_23892,N_15161,N_18098);
nor U23893 (N_23893,N_19480,N_17053);
and U23894 (N_23894,N_16777,N_15140);
nand U23895 (N_23895,N_15745,N_19258);
nor U23896 (N_23896,N_18301,N_16801);
nand U23897 (N_23897,N_19564,N_18437);
or U23898 (N_23898,N_17234,N_17183);
nand U23899 (N_23899,N_16204,N_17332);
and U23900 (N_23900,N_16659,N_17457);
nor U23901 (N_23901,N_17579,N_19331);
nor U23902 (N_23902,N_18775,N_16913);
nor U23903 (N_23903,N_19417,N_16669);
nor U23904 (N_23904,N_15649,N_16560);
xor U23905 (N_23905,N_18596,N_15624);
and U23906 (N_23906,N_16981,N_17236);
nor U23907 (N_23907,N_16744,N_18771);
nor U23908 (N_23908,N_19059,N_19462);
nor U23909 (N_23909,N_17293,N_17975);
nand U23910 (N_23910,N_18894,N_19001);
nand U23911 (N_23911,N_16727,N_16061);
and U23912 (N_23912,N_19548,N_18013);
nand U23913 (N_23913,N_17014,N_18184);
nand U23914 (N_23914,N_15094,N_17947);
nand U23915 (N_23915,N_17245,N_16659);
or U23916 (N_23916,N_17723,N_17715);
and U23917 (N_23917,N_16268,N_16132);
or U23918 (N_23918,N_19977,N_16026);
nor U23919 (N_23919,N_15855,N_17826);
xor U23920 (N_23920,N_17644,N_16679);
nor U23921 (N_23921,N_18810,N_18328);
nand U23922 (N_23922,N_19576,N_15222);
or U23923 (N_23923,N_19452,N_19430);
and U23924 (N_23924,N_15088,N_18419);
nand U23925 (N_23925,N_17136,N_16247);
nor U23926 (N_23926,N_18751,N_15842);
and U23927 (N_23927,N_17387,N_18032);
nand U23928 (N_23928,N_16686,N_18407);
nand U23929 (N_23929,N_18927,N_19657);
nand U23930 (N_23930,N_17562,N_15415);
or U23931 (N_23931,N_19206,N_18681);
and U23932 (N_23932,N_19019,N_18312);
and U23933 (N_23933,N_16356,N_16360);
and U23934 (N_23934,N_17445,N_17078);
nor U23935 (N_23935,N_16364,N_19836);
nand U23936 (N_23936,N_16052,N_16765);
and U23937 (N_23937,N_19545,N_15992);
and U23938 (N_23938,N_16280,N_17799);
nor U23939 (N_23939,N_17196,N_16424);
nor U23940 (N_23940,N_17540,N_16929);
and U23941 (N_23941,N_18884,N_19818);
or U23942 (N_23942,N_18273,N_18854);
nand U23943 (N_23943,N_19777,N_17841);
and U23944 (N_23944,N_16559,N_18703);
nand U23945 (N_23945,N_15398,N_16173);
xor U23946 (N_23946,N_19606,N_18521);
nand U23947 (N_23947,N_15620,N_17188);
and U23948 (N_23948,N_16942,N_18822);
and U23949 (N_23949,N_18471,N_16814);
nand U23950 (N_23950,N_17100,N_17013);
or U23951 (N_23951,N_16358,N_17562);
or U23952 (N_23952,N_16329,N_19902);
xor U23953 (N_23953,N_15528,N_15043);
xnor U23954 (N_23954,N_18375,N_18993);
xnor U23955 (N_23955,N_18388,N_18418);
or U23956 (N_23956,N_18732,N_18514);
and U23957 (N_23957,N_15759,N_15250);
nand U23958 (N_23958,N_18672,N_19662);
nand U23959 (N_23959,N_16616,N_15820);
nor U23960 (N_23960,N_15939,N_16664);
nor U23961 (N_23961,N_16871,N_16541);
or U23962 (N_23962,N_16128,N_15332);
nand U23963 (N_23963,N_18782,N_16426);
xnor U23964 (N_23964,N_17004,N_16287);
and U23965 (N_23965,N_19314,N_19853);
nand U23966 (N_23966,N_19482,N_17932);
nor U23967 (N_23967,N_16819,N_17539);
nor U23968 (N_23968,N_15286,N_19466);
nand U23969 (N_23969,N_17338,N_18103);
and U23970 (N_23970,N_18363,N_16248);
nand U23971 (N_23971,N_17168,N_15476);
xor U23972 (N_23972,N_17325,N_19672);
and U23973 (N_23973,N_15250,N_19936);
or U23974 (N_23974,N_17200,N_19274);
nand U23975 (N_23975,N_17917,N_16263);
or U23976 (N_23976,N_15365,N_19481);
xor U23977 (N_23977,N_18906,N_18336);
nor U23978 (N_23978,N_19546,N_19396);
nand U23979 (N_23979,N_16038,N_15999);
nor U23980 (N_23980,N_16271,N_16758);
xor U23981 (N_23981,N_17219,N_17134);
xor U23982 (N_23982,N_18310,N_17824);
nor U23983 (N_23983,N_18456,N_16906);
and U23984 (N_23984,N_16100,N_17174);
nand U23985 (N_23985,N_17581,N_18552);
nand U23986 (N_23986,N_16081,N_15241);
nand U23987 (N_23987,N_17379,N_17571);
and U23988 (N_23988,N_16590,N_19972);
and U23989 (N_23989,N_18042,N_16737);
or U23990 (N_23990,N_16266,N_15181);
xor U23991 (N_23991,N_16197,N_16743);
or U23992 (N_23992,N_17095,N_18698);
and U23993 (N_23993,N_18480,N_17922);
and U23994 (N_23994,N_16082,N_15116);
xor U23995 (N_23995,N_17693,N_17721);
nor U23996 (N_23996,N_15583,N_18622);
nand U23997 (N_23997,N_15678,N_17056);
nand U23998 (N_23998,N_16085,N_17017);
and U23999 (N_23999,N_17067,N_18383);
nand U24000 (N_24000,N_15220,N_17033);
nand U24001 (N_24001,N_18777,N_19993);
xnor U24002 (N_24002,N_15155,N_18572);
or U24003 (N_24003,N_18981,N_17456);
nand U24004 (N_24004,N_19060,N_17899);
and U24005 (N_24005,N_18940,N_18962);
or U24006 (N_24006,N_16729,N_15564);
nor U24007 (N_24007,N_19417,N_16909);
and U24008 (N_24008,N_17600,N_18196);
and U24009 (N_24009,N_16122,N_16602);
nor U24010 (N_24010,N_17301,N_15482);
or U24011 (N_24011,N_17024,N_18990);
nor U24012 (N_24012,N_18536,N_17499);
and U24013 (N_24013,N_17537,N_19249);
and U24014 (N_24014,N_15161,N_18877);
nor U24015 (N_24015,N_18754,N_18712);
xor U24016 (N_24016,N_17089,N_19132);
xnor U24017 (N_24017,N_17352,N_16493);
or U24018 (N_24018,N_15869,N_17095);
and U24019 (N_24019,N_19269,N_15094);
or U24020 (N_24020,N_17689,N_19201);
nor U24021 (N_24021,N_15599,N_19931);
xnor U24022 (N_24022,N_18747,N_18247);
nor U24023 (N_24023,N_17424,N_17560);
nand U24024 (N_24024,N_19918,N_18543);
or U24025 (N_24025,N_18935,N_18801);
xnor U24026 (N_24026,N_16603,N_15938);
nor U24027 (N_24027,N_19242,N_19060);
and U24028 (N_24028,N_15570,N_18804);
nor U24029 (N_24029,N_18392,N_18793);
and U24030 (N_24030,N_16355,N_17998);
nor U24031 (N_24031,N_19538,N_15367);
nand U24032 (N_24032,N_19117,N_18755);
and U24033 (N_24033,N_18925,N_19345);
nand U24034 (N_24034,N_17528,N_17089);
nor U24035 (N_24035,N_18745,N_18107);
and U24036 (N_24036,N_15650,N_16456);
or U24037 (N_24037,N_17399,N_17526);
xor U24038 (N_24038,N_19566,N_18908);
nand U24039 (N_24039,N_15171,N_18001);
nor U24040 (N_24040,N_15462,N_16063);
and U24041 (N_24041,N_15591,N_19682);
or U24042 (N_24042,N_15455,N_18616);
nor U24043 (N_24043,N_16805,N_16787);
or U24044 (N_24044,N_19645,N_18478);
and U24045 (N_24045,N_19423,N_17646);
nor U24046 (N_24046,N_17955,N_15882);
and U24047 (N_24047,N_15222,N_16435);
nand U24048 (N_24048,N_19367,N_17144);
nor U24049 (N_24049,N_16995,N_17412);
nor U24050 (N_24050,N_15064,N_18837);
and U24051 (N_24051,N_16187,N_15650);
and U24052 (N_24052,N_15467,N_15385);
nor U24053 (N_24053,N_15108,N_15511);
nor U24054 (N_24054,N_18119,N_17659);
nand U24055 (N_24055,N_19746,N_19777);
or U24056 (N_24056,N_18052,N_17658);
or U24057 (N_24057,N_19797,N_19677);
nor U24058 (N_24058,N_17509,N_16459);
or U24059 (N_24059,N_18902,N_15125);
and U24060 (N_24060,N_16049,N_15572);
nand U24061 (N_24061,N_19482,N_17727);
nor U24062 (N_24062,N_15684,N_15255);
or U24063 (N_24063,N_15702,N_16182);
nand U24064 (N_24064,N_16037,N_19697);
xor U24065 (N_24065,N_17270,N_16101);
and U24066 (N_24066,N_18330,N_18637);
and U24067 (N_24067,N_19266,N_19930);
xnor U24068 (N_24068,N_15208,N_19066);
or U24069 (N_24069,N_17735,N_18908);
nor U24070 (N_24070,N_18532,N_16636);
xnor U24071 (N_24071,N_15539,N_17914);
nor U24072 (N_24072,N_16226,N_17912);
and U24073 (N_24073,N_19702,N_19541);
nor U24074 (N_24074,N_17867,N_16190);
nand U24075 (N_24075,N_17955,N_16244);
nor U24076 (N_24076,N_19473,N_15197);
nor U24077 (N_24077,N_16790,N_15467);
or U24078 (N_24078,N_15802,N_19252);
nand U24079 (N_24079,N_18484,N_15957);
nor U24080 (N_24080,N_16333,N_15669);
nand U24081 (N_24081,N_19810,N_17691);
nor U24082 (N_24082,N_19016,N_16158);
nor U24083 (N_24083,N_19549,N_19350);
nor U24084 (N_24084,N_16818,N_19732);
or U24085 (N_24085,N_15070,N_16032);
nand U24086 (N_24086,N_18183,N_17625);
nand U24087 (N_24087,N_16713,N_15370);
xnor U24088 (N_24088,N_18979,N_18233);
nor U24089 (N_24089,N_17074,N_17087);
nand U24090 (N_24090,N_19214,N_15426);
and U24091 (N_24091,N_18308,N_18111);
or U24092 (N_24092,N_17679,N_15617);
nor U24093 (N_24093,N_19487,N_18490);
nand U24094 (N_24094,N_19624,N_18708);
nand U24095 (N_24095,N_15234,N_16786);
nor U24096 (N_24096,N_19802,N_17607);
or U24097 (N_24097,N_16542,N_18476);
or U24098 (N_24098,N_19424,N_17457);
and U24099 (N_24099,N_17602,N_17830);
nor U24100 (N_24100,N_17833,N_19846);
or U24101 (N_24101,N_15693,N_16673);
and U24102 (N_24102,N_15883,N_19437);
nand U24103 (N_24103,N_19665,N_16974);
and U24104 (N_24104,N_18841,N_18857);
nor U24105 (N_24105,N_18318,N_19077);
or U24106 (N_24106,N_19566,N_19036);
nor U24107 (N_24107,N_17396,N_16689);
or U24108 (N_24108,N_18142,N_17336);
or U24109 (N_24109,N_17104,N_19253);
or U24110 (N_24110,N_15679,N_15553);
xor U24111 (N_24111,N_16905,N_18220);
or U24112 (N_24112,N_15743,N_15336);
and U24113 (N_24113,N_19308,N_15738);
nand U24114 (N_24114,N_19823,N_16807);
nor U24115 (N_24115,N_17614,N_18694);
nand U24116 (N_24116,N_19369,N_16514);
nor U24117 (N_24117,N_19218,N_17455);
nand U24118 (N_24118,N_16973,N_18651);
nand U24119 (N_24119,N_18020,N_15855);
or U24120 (N_24120,N_17363,N_18464);
and U24121 (N_24121,N_15849,N_16841);
nor U24122 (N_24122,N_18133,N_18164);
nand U24123 (N_24123,N_15379,N_15447);
nor U24124 (N_24124,N_15429,N_16210);
nand U24125 (N_24125,N_16827,N_17384);
or U24126 (N_24126,N_18997,N_16719);
xnor U24127 (N_24127,N_17227,N_19143);
and U24128 (N_24128,N_16450,N_15510);
or U24129 (N_24129,N_19844,N_17037);
nand U24130 (N_24130,N_18043,N_15678);
nand U24131 (N_24131,N_16020,N_18046);
or U24132 (N_24132,N_18207,N_18050);
nor U24133 (N_24133,N_15380,N_19788);
nand U24134 (N_24134,N_19330,N_17605);
or U24135 (N_24135,N_17206,N_15775);
xnor U24136 (N_24136,N_19905,N_18942);
or U24137 (N_24137,N_18086,N_19146);
nand U24138 (N_24138,N_19017,N_16029);
or U24139 (N_24139,N_15996,N_16734);
nor U24140 (N_24140,N_15144,N_18417);
or U24141 (N_24141,N_19243,N_16892);
nor U24142 (N_24142,N_17548,N_15044);
nand U24143 (N_24143,N_19833,N_18955);
and U24144 (N_24144,N_15663,N_16619);
and U24145 (N_24145,N_16557,N_16568);
nand U24146 (N_24146,N_16186,N_18565);
or U24147 (N_24147,N_15195,N_18629);
nor U24148 (N_24148,N_15262,N_18978);
or U24149 (N_24149,N_18839,N_19806);
xnor U24150 (N_24150,N_17787,N_15850);
nor U24151 (N_24151,N_19167,N_16221);
nand U24152 (N_24152,N_16657,N_16679);
xnor U24153 (N_24153,N_17267,N_18944);
nor U24154 (N_24154,N_18925,N_16487);
or U24155 (N_24155,N_17051,N_19096);
nor U24156 (N_24156,N_17416,N_15679);
or U24157 (N_24157,N_16141,N_18501);
and U24158 (N_24158,N_15531,N_18367);
xnor U24159 (N_24159,N_16015,N_17093);
and U24160 (N_24160,N_15648,N_16270);
nor U24161 (N_24161,N_16940,N_19497);
and U24162 (N_24162,N_15190,N_15289);
nor U24163 (N_24163,N_19276,N_17563);
nand U24164 (N_24164,N_17964,N_17140);
xor U24165 (N_24165,N_17103,N_17148);
nor U24166 (N_24166,N_15812,N_18103);
or U24167 (N_24167,N_19095,N_15823);
or U24168 (N_24168,N_17102,N_16965);
nand U24169 (N_24169,N_17744,N_18858);
and U24170 (N_24170,N_18289,N_17445);
nor U24171 (N_24171,N_19213,N_17596);
xnor U24172 (N_24172,N_17995,N_18665);
and U24173 (N_24173,N_19454,N_15625);
nor U24174 (N_24174,N_18622,N_15786);
and U24175 (N_24175,N_15570,N_18942);
nor U24176 (N_24176,N_19078,N_18971);
or U24177 (N_24177,N_18286,N_18246);
nand U24178 (N_24178,N_19423,N_17107);
xor U24179 (N_24179,N_17982,N_16548);
nand U24180 (N_24180,N_15132,N_15675);
xnor U24181 (N_24181,N_17317,N_16248);
and U24182 (N_24182,N_16621,N_18527);
and U24183 (N_24183,N_17524,N_15812);
nand U24184 (N_24184,N_15379,N_15860);
or U24185 (N_24185,N_18502,N_16279);
nor U24186 (N_24186,N_15381,N_18157);
or U24187 (N_24187,N_15480,N_19764);
nand U24188 (N_24188,N_15658,N_17126);
or U24189 (N_24189,N_17266,N_15148);
and U24190 (N_24190,N_17832,N_16823);
nand U24191 (N_24191,N_15547,N_18933);
xnor U24192 (N_24192,N_18922,N_16679);
or U24193 (N_24193,N_19672,N_18150);
xor U24194 (N_24194,N_16859,N_17991);
and U24195 (N_24195,N_18956,N_16502);
or U24196 (N_24196,N_19175,N_18922);
nor U24197 (N_24197,N_16617,N_19965);
nor U24198 (N_24198,N_19494,N_19796);
or U24199 (N_24199,N_15808,N_15851);
and U24200 (N_24200,N_19333,N_15874);
and U24201 (N_24201,N_17994,N_16854);
nand U24202 (N_24202,N_16016,N_18212);
or U24203 (N_24203,N_15421,N_18720);
and U24204 (N_24204,N_16438,N_16218);
xor U24205 (N_24205,N_16251,N_15370);
nor U24206 (N_24206,N_17867,N_18347);
or U24207 (N_24207,N_15511,N_16459);
nor U24208 (N_24208,N_17954,N_17392);
nor U24209 (N_24209,N_18320,N_17887);
and U24210 (N_24210,N_19490,N_15303);
nand U24211 (N_24211,N_17753,N_16752);
nand U24212 (N_24212,N_16937,N_16447);
or U24213 (N_24213,N_18993,N_17546);
nor U24214 (N_24214,N_18848,N_17046);
and U24215 (N_24215,N_18466,N_19887);
nor U24216 (N_24216,N_17538,N_17061);
xnor U24217 (N_24217,N_17821,N_15761);
nor U24218 (N_24218,N_17702,N_19384);
xor U24219 (N_24219,N_16733,N_18820);
nor U24220 (N_24220,N_19072,N_19062);
nor U24221 (N_24221,N_15544,N_19064);
and U24222 (N_24222,N_16222,N_16517);
xor U24223 (N_24223,N_19945,N_17918);
xor U24224 (N_24224,N_17761,N_16467);
and U24225 (N_24225,N_17793,N_19667);
nor U24226 (N_24226,N_17988,N_16096);
nor U24227 (N_24227,N_16246,N_16155);
nand U24228 (N_24228,N_18630,N_18081);
nor U24229 (N_24229,N_18130,N_15476);
or U24230 (N_24230,N_15066,N_17680);
nand U24231 (N_24231,N_15129,N_18147);
nand U24232 (N_24232,N_15738,N_17580);
and U24233 (N_24233,N_19439,N_19858);
and U24234 (N_24234,N_19824,N_18861);
nor U24235 (N_24235,N_18183,N_15244);
nor U24236 (N_24236,N_16398,N_18322);
xor U24237 (N_24237,N_15466,N_17141);
nand U24238 (N_24238,N_19573,N_15117);
or U24239 (N_24239,N_18085,N_18238);
nor U24240 (N_24240,N_18651,N_15635);
nand U24241 (N_24241,N_17036,N_18502);
xnor U24242 (N_24242,N_19986,N_17655);
or U24243 (N_24243,N_17521,N_17360);
or U24244 (N_24244,N_16704,N_15107);
nand U24245 (N_24245,N_16209,N_15174);
nor U24246 (N_24246,N_19279,N_17987);
or U24247 (N_24247,N_15593,N_15267);
nand U24248 (N_24248,N_19102,N_19504);
or U24249 (N_24249,N_19512,N_17594);
nand U24250 (N_24250,N_17648,N_17384);
nand U24251 (N_24251,N_16266,N_16468);
or U24252 (N_24252,N_19919,N_16917);
and U24253 (N_24253,N_18310,N_18551);
and U24254 (N_24254,N_15964,N_18679);
or U24255 (N_24255,N_16759,N_16388);
and U24256 (N_24256,N_16143,N_16026);
nand U24257 (N_24257,N_16916,N_16095);
and U24258 (N_24258,N_15983,N_15971);
nor U24259 (N_24259,N_18531,N_18544);
xnor U24260 (N_24260,N_19488,N_19533);
nor U24261 (N_24261,N_16190,N_16567);
nand U24262 (N_24262,N_15401,N_19435);
xnor U24263 (N_24263,N_15808,N_19679);
and U24264 (N_24264,N_16532,N_15767);
or U24265 (N_24265,N_19838,N_15216);
nand U24266 (N_24266,N_18997,N_19421);
and U24267 (N_24267,N_18888,N_15453);
or U24268 (N_24268,N_16058,N_19587);
or U24269 (N_24269,N_15745,N_19758);
nand U24270 (N_24270,N_19651,N_18367);
and U24271 (N_24271,N_17967,N_17360);
and U24272 (N_24272,N_15838,N_19226);
or U24273 (N_24273,N_16310,N_17021);
and U24274 (N_24274,N_16980,N_15036);
or U24275 (N_24275,N_19062,N_18539);
and U24276 (N_24276,N_19896,N_15388);
xnor U24277 (N_24277,N_19769,N_17178);
and U24278 (N_24278,N_16572,N_16515);
xnor U24279 (N_24279,N_18917,N_15519);
and U24280 (N_24280,N_19761,N_17342);
and U24281 (N_24281,N_18027,N_19225);
nand U24282 (N_24282,N_17522,N_15059);
and U24283 (N_24283,N_15846,N_17354);
nand U24284 (N_24284,N_17727,N_17356);
nand U24285 (N_24285,N_16059,N_16790);
and U24286 (N_24286,N_15669,N_18418);
and U24287 (N_24287,N_19974,N_17476);
or U24288 (N_24288,N_15995,N_17158);
nand U24289 (N_24289,N_15792,N_19705);
xnor U24290 (N_24290,N_16190,N_19487);
xnor U24291 (N_24291,N_18816,N_15620);
nand U24292 (N_24292,N_16039,N_17555);
and U24293 (N_24293,N_17775,N_18347);
or U24294 (N_24294,N_18674,N_16288);
nand U24295 (N_24295,N_19699,N_19292);
or U24296 (N_24296,N_15080,N_16199);
or U24297 (N_24297,N_18748,N_17962);
nand U24298 (N_24298,N_17068,N_19837);
and U24299 (N_24299,N_18140,N_15030);
nand U24300 (N_24300,N_17716,N_18288);
nor U24301 (N_24301,N_17668,N_16005);
or U24302 (N_24302,N_17122,N_16705);
and U24303 (N_24303,N_16187,N_16968);
and U24304 (N_24304,N_18861,N_15749);
nand U24305 (N_24305,N_18559,N_15697);
nand U24306 (N_24306,N_15530,N_18253);
nor U24307 (N_24307,N_15039,N_19059);
and U24308 (N_24308,N_17881,N_16624);
nand U24309 (N_24309,N_15256,N_18980);
nor U24310 (N_24310,N_16925,N_15325);
nor U24311 (N_24311,N_18509,N_16494);
or U24312 (N_24312,N_16188,N_15953);
nor U24313 (N_24313,N_19273,N_18228);
nor U24314 (N_24314,N_18570,N_19373);
and U24315 (N_24315,N_18416,N_15810);
or U24316 (N_24316,N_18611,N_16014);
and U24317 (N_24317,N_15494,N_17604);
or U24318 (N_24318,N_15984,N_15667);
or U24319 (N_24319,N_18252,N_17362);
or U24320 (N_24320,N_18472,N_18230);
nor U24321 (N_24321,N_19941,N_19165);
xnor U24322 (N_24322,N_15208,N_16397);
and U24323 (N_24323,N_16845,N_15874);
and U24324 (N_24324,N_19340,N_19877);
nand U24325 (N_24325,N_16661,N_16194);
nand U24326 (N_24326,N_15568,N_16756);
or U24327 (N_24327,N_16209,N_17525);
xor U24328 (N_24328,N_17655,N_15522);
or U24329 (N_24329,N_15925,N_19151);
nor U24330 (N_24330,N_17903,N_17960);
nor U24331 (N_24331,N_18059,N_17839);
and U24332 (N_24332,N_19757,N_17608);
and U24333 (N_24333,N_19719,N_18379);
xnor U24334 (N_24334,N_19393,N_17334);
nor U24335 (N_24335,N_16384,N_15755);
nand U24336 (N_24336,N_17241,N_17074);
nand U24337 (N_24337,N_19172,N_17243);
nor U24338 (N_24338,N_15794,N_18769);
nor U24339 (N_24339,N_16815,N_15360);
and U24340 (N_24340,N_17048,N_15345);
nand U24341 (N_24341,N_15596,N_19278);
or U24342 (N_24342,N_16681,N_16356);
nor U24343 (N_24343,N_17309,N_16524);
nand U24344 (N_24344,N_16020,N_18427);
and U24345 (N_24345,N_17585,N_18021);
xor U24346 (N_24346,N_16341,N_16106);
nand U24347 (N_24347,N_19361,N_15431);
nor U24348 (N_24348,N_16298,N_15362);
or U24349 (N_24349,N_16977,N_18092);
xor U24350 (N_24350,N_15827,N_18096);
and U24351 (N_24351,N_15351,N_19688);
or U24352 (N_24352,N_16483,N_15922);
nor U24353 (N_24353,N_18846,N_19276);
and U24354 (N_24354,N_15035,N_19270);
or U24355 (N_24355,N_16705,N_16714);
nand U24356 (N_24356,N_19431,N_18080);
or U24357 (N_24357,N_16614,N_19487);
or U24358 (N_24358,N_16810,N_19949);
or U24359 (N_24359,N_15170,N_16318);
nand U24360 (N_24360,N_17875,N_17790);
xnor U24361 (N_24361,N_17305,N_15989);
or U24362 (N_24362,N_15972,N_18635);
nand U24363 (N_24363,N_19836,N_17692);
nor U24364 (N_24364,N_16171,N_15985);
and U24365 (N_24365,N_15942,N_19102);
nor U24366 (N_24366,N_15329,N_19353);
and U24367 (N_24367,N_18927,N_15644);
nand U24368 (N_24368,N_19915,N_19486);
and U24369 (N_24369,N_19593,N_18680);
xnor U24370 (N_24370,N_19631,N_15093);
xor U24371 (N_24371,N_15531,N_18380);
and U24372 (N_24372,N_19413,N_19698);
xor U24373 (N_24373,N_19830,N_16903);
nand U24374 (N_24374,N_16751,N_19444);
nor U24375 (N_24375,N_17253,N_17735);
nand U24376 (N_24376,N_19727,N_15867);
and U24377 (N_24377,N_19140,N_19973);
and U24378 (N_24378,N_18242,N_18357);
and U24379 (N_24379,N_15903,N_19743);
nor U24380 (N_24380,N_19202,N_15867);
and U24381 (N_24381,N_19920,N_17798);
nand U24382 (N_24382,N_15666,N_19070);
xnor U24383 (N_24383,N_15940,N_18021);
and U24384 (N_24384,N_19785,N_18221);
nand U24385 (N_24385,N_19390,N_15582);
nor U24386 (N_24386,N_15582,N_17289);
nand U24387 (N_24387,N_16590,N_19245);
and U24388 (N_24388,N_16824,N_19163);
nand U24389 (N_24389,N_17511,N_16332);
nand U24390 (N_24390,N_17721,N_19012);
nor U24391 (N_24391,N_16955,N_19165);
nor U24392 (N_24392,N_16770,N_17650);
nand U24393 (N_24393,N_17706,N_17920);
or U24394 (N_24394,N_19525,N_18142);
or U24395 (N_24395,N_17162,N_17736);
or U24396 (N_24396,N_19365,N_16745);
and U24397 (N_24397,N_17277,N_16578);
or U24398 (N_24398,N_15357,N_17101);
or U24399 (N_24399,N_17548,N_19695);
xnor U24400 (N_24400,N_15953,N_18778);
nand U24401 (N_24401,N_18059,N_17316);
nor U24402 (N_24402,N_15532,N_15917);
xor U24403 (N_24403,N_17418,N_17821);
nand U24404 (N_24404,N_16249,N_17651);
or U24405 (N_24405,N_16126,N_15052);
nor U24406 (N_24406,N_19576,N_16464);
or U24407 (N_24407,N_19178,N_15485);
and U24408 (N_24408,N_17390,N_19733);
nand U24409 (N_24409,N_17370,N_18812);
nand U24410 (N_24410,N_19293,N_19300);
and U24411 (N_24411,N_16858,N_15550);
nor U24412 (N_24412,N_15677,N_19723);
nand U24413 (N_24413,N_17546,N_15358);
nor U24414 (N_24414,N_19144,N_15195);
xnor U24415 (N_24415,N_18058,N_17282);
or U24416 (N_24416,N_19379,N_17493);
nor U24417 (N_24417,N_16124,N_18742);
or U24418 (N_24418,N_16219,N_16110);
nor U24419 (N_24419,N_19221,N_18006);
nand U24420 (N_24420,N_18957,N_15857);
or U24421 (N_24421,N_19584,N_15047);
or U24422 (N_24422,N_15507,N_15242);
nor U24423 (N_24423,N_19497,N_18205);
and U24424 (N_24424,N_19394,N_15062);
nand U24425 (N_24425,N_18407,N_16081);
nand U24426 (N_24426,N_16228,N_19979);
and U24427 (N_24427,N_16207,N_18387);
or U24428 (N_24428,N_15933,N_18044);
nor U24429 (N_24429,N_15252,N_17317);
and U24430 (N_24430,N_16067,N_15325);
nand U24431 (N_24431,N_19665,N_17198);
nand U24432 (N_24432,N_18476,N_17083);
or U24433 (N_24433,N_16446,N_17836);
nand U24434 (N_24434,N_16721,N_16777);
and U24435 (N_24435,N_18216,N_17181);
nor U24436 (N_24436,N_18255,N_16876);
nor U24437 (N_24437,N_16754,N_18377);
nand U24438 (N_24438,N_16926,N_19683);
nor U24439 (N_24439,N_19673,N_15558);
and U24440 (N_24440,N_15965,N_16256);
and U24441 (N_24441,N_19316,N_18861);
and U24442 (N_24442,N_18953,N_16500);
or U24443 (N_24443,N_15105,N_16116);
and U24444 (N_24444,N_18369,N_17385);
xnor U24445 (N_24445,N_17025,N_19486);
nor U24446 (N_24446,N_19705,N_18143);
nor U24447 (N_24447,N_18106,N_17350);
nand U24448 (N_24448,N_17910,N_17647);
nand U24449 (N_24449,N_17080,N_18792);
and U24450 (N_24450,N_15419,N_15599);
and U24451 (N_24451,N_16414,N_15195);
and U24452 (N_24452,N_17580,N_17244);
nand U24453 (N_24453,N_16885,N_17740);
and U24454 (N_24454,N_16309,N_16247);
nor U24455 (N_24455,N_18153,N_15790);
nand U24456 (N_24456,N_18682,N_19106);
nor U24457 (N_24457,N_16611,N_16739);
nor U24458 (N_24458,N_17993,N_17499);
or U24459 (N_24459,N_18028,N_15157);
xor U24460 (N_24460,N_19280,N_19662);
nand U24461 (N_24461,N_18443,N_17973);
nor U24462 (N_24462,N_16129,N_15590);
and U24463 (N_24463,N_16201,N_16567);
xnor U24464 (N_24464,N_15901,N_19327);
or U24465 (N_24465,N_19516,N_19562);
or U24466 (N_24466,N_17836,N_17087);
xor U24467 (N_24467,N_18424,N_19790);
nand U24468 (N_24468,N_16328,N_15113);
nor U24469 (N_24469,N_17088,N_15883);
or U24470 (N_24470,N_16354,N_17856);
and U24471 (N_24471,N_15700,N_18697);
nand U24472 (N_24472,N_19341,N_19088);
nor U24473 (N_24473,N_18768,N_18047);
nand U24474 (N_24474,N_15346,N_19205);
nor U24475 (N_24475,N_15752,N_15909);
xnor U24476 (N_24476,N_19780,N_16467);
nand U24477 (N_24477,N_17803,N_15338);
and U24478 (N_24478,N_16741,N_16982);
and U24479 (N_24479,N_16743,N_15414);
and U24480 (N_24480,N_16289,N_17802);
xnor U24481 (N_24481,N_18482,N_17644);
nand U24482 (N_24482,N_17719,N_16435);
or U24483 (N_24483,N_16241,N_19078);
or U24484 (N_24484,N_15515,N_19670);
nor U24485 (N_24485,N_15263,N_18043);
nand U24486 (N_24486,N_18318,N_19859);
and U24487 (N_24487,N_19226,N_16828);
or U24488 (N_24488,N_19160,N_15162);
nor U24489 (N_24489,N_16152,N_19388);
nor U24490 (N_24490,N_18594,N_17862);
nor U24491 (N_24491,N_16307,N_18663);
nand U24492 (N_24492,N_19901,N_17425);
or U24493 (N_24493,N_17779,N_15625);
nand U24494 (N_24494,N_16643,N_17175);
or U24495 (N_24495,N_16112,N_18768);
nor U24496 (N_24496,N_17048,N_16782);
and U24497 (N_24497,N_19279,N_16675);
and U24498 (N_24498,N_19982,N_17263);
or U24499 (N_24499,N_18528,N_19213);
nor U24500 (N_24500,N_16624,N_18750);
or U24501 (N_24501,N_19721,N_19988);
xnor U24502 (N_24502,N_17462,N_19871);
and U24503 (N_24503,N_18725,N_19725);
and U24504 (N_24504,N_16900,N_16075);
and U24505 (N_24505,N_15274,N_16659);
and U24506 (N_24506,N_16879,N_17188);
nand U24507 (N_24507,N_18502,N_16830);
or U24508 (N_24508,N_18427,N_17873);
and U24509 (N_24509,N_16475,N_16356);
xor U24510 (N_24510,N_16414,N_17139);
or U24511 (N_24511,N_15407,N_19069);
nand U24512 (N_24512,N_19002,N_19265);
nand U24513 (N_24513,N_18946,N_19083);
nor U24514 (N_24514,N_16916,N_19198);
and U24515 (N_24515,N_16122,N_18492);
or U24516 (N_24516,N_18432,N_19497);
and U24517 (N_24517,N_16083,N_16606);
nor U24518 (N_24518,N_16694,N_17600);
or U24519 (N_24519,N_19015,N_17573);
nor U24520 (N_24520,N_18441,N_15761);
and U24521 (N_24521,N_15654,N_18589);
nand U24522 (N_24522,N_16116,N_18993);
xnor U24523 (N_24523,N_16027,N_17740);
nand U24524 (N_24524,N_16453,N_16068);
nor U24525 (N_24525,N_16773,N_16867);
nor U24526 (N_24526,N_19205,N_15523);
and U24527 (N_24527,N_15822,N_16073);
nand U24528 (N_24528,N_15644,N_18409);
nor U24529 (N_24529,N_15398,N_15641);
nand U24530 (N_24530,N_17953,N_16060);
nand U24531 (N_24531,N_16386,N_15267);
xor U24532 (N_24532,N_15105,N_18861);
nand U24533 (N_24533,N_15742,N_19933);
xor U24534 (N_24534,N_19415,N_18133);
and U24535 (N_24535,N_17059,N_17290);
and U24536 (N_24536,N_19186,N_16231);
nand U24537 (N_24537,N_16570,N_16098);
nor U24538 (N_24538,N_15165,N_16489);
nand U24539 (N_24539,N_17430,N_15575);
and U24540 (N_24540,N_16706,N_16258);
and U24541 (N_24541,N_17101,N_15028);
nand U24542 (N_24542,N_15500,N_19476);
nand U24543 (N_24543,N_16221,N_17442);
nor U24544 (N_24544,N_18491,N_18740);
nand U24545 (N_24545,N_16842,N_16171);
nand U24546 (N_24546,N_15038,N_16925);
or U24547 (N_24547,N_15530,N_18451);
nand U24548 (N_24548,N_18931,N_19550);
nand U24549 (N_24549,N_18861,N_18549);
or U24550 (N_24550,N_18985,N_17276);
and U24551 (N_24551,N_17126,N_16906);
or U24552 (N_24552,N_17348,N_17482);
and U24553 (N_24553,N_15036,N_19263);
or U24554 (N_24554,N_19384,N_17007);
nand U24555 (N_24555,N_18442,N_19058);
nor U24556 (N_24556,N_16648,N_18008);
nand U24557 (N_24557,N_17587,N_19934);
nor U24558 (N_24558,N_16893,N_15365);
and U24559 (N_24559,N_19370,N_16810);
nor U24560 (N_24560,N_16326,N_19743);
or U24561 (N_24561,N_19714,N_18390);
nand U24562 (N_24562,N_18378,N_16925);
nor U24563 (N_24563,N_15270,N_15252);
and U24564 (N_24564,N_16160,N_19784);
or U24565 (N_24565,N_15947,N_19371);
and U24566 (N_24566,N_16440,N_19827);
nor U24567 (N_24567,N_15036,N_17239);
or U24568 (N_24568,N_17841,N_19045);
nand U24569 (N_24569,N_16773,N_18218);
or U24570 (N_24570,N_15723,N_19469);
xnor U24571 (N_24571,N_17652,N_19227);
and U24572 (N_24572,N_16939,N_15701);
xor U24573 (N_24573,N_19299,N_15169);
and U24574 (N_24574,N_15884,N_18020);
nand U24575 (N_24575,N_18462,N_18075);
nand U24576 (N_24576,N_19322,N_16055);
nand U24577 (N_24577,N_17492,N_16135);
or U24578 (N_24578,N_15726,N_19489);
nand U24579 (N_24579,N_18061,N_19001);
nand U24580 (N_24580,N_19895,N_16726);
nor U24581 (N_24581,N_17730,N_19275);
and U24582 (N_24582,N_17846,N_16872);
nor U24583 (N_24583,N_19334,N_17782);
nand U24584 (N_24584,N_19831,N_15171);
and U24585 (N_24585,N_16119,N_16210);
nand U24586 (N_24586,N_16039,N_15540);
or U24587 (N_24587,N_18789,N_16646);
or U24588 (N_24588,N_16799,N_15028);
nand U24589 (N_24589,N_18393,N_17079);
or U24590 (N_24590,N_16601,N_17971);
and U24591 (N_24591,N_19825,N_16827);
nor U24592 (N_24592,N_19297,N_19231);
nor U24593 (N_24593,N_18115,N_18683);
nand U24594 (N_24594,N_15501,N_15036);
and U24595 (N_24595,N_16151,N_18520);
nand U24596 (N_24596,N_15633,N_17689);
xnor U24597 (N_24597,N_17749,N_18851);
nor U24598 (N_24598,N_16055,N_15044);
nand U24599 (N_24599,N_18020,N_18853);
or U24600 (N_24600,N_18186,N_19684);
and U24601 (N_24601,N_16449,N_19135);
and U24602 (N_24602,N_18951,N_17585);
and U24603 (N_24603,N_15060,N_18644);
nor U24604 (N_24604,N_16155,N_18357);
nand U24605 (N_24605,N_18440,N_17326);
nand U24606 (N_24606,N_18725,N_18423);
or U24607 (N_24607,N_17743,N_19697);
or U24608 (N_24608,N_18295,N_18229);
and U24609 (N_24609,N_18465,N_19686);
nand U24610 (N_24610,N_16161,N_17204);
and U24611 (N_24611,N_18006,N_15455);
and U24612 (N_24612,N_18662,N_17915);
nand U24613 (N_24613,N_16282,N_18626);
nand U24614 (N_24614,N_18975,N_17827);
and U24615 (N_24615,N_19220,N_17963);
nand U24616 (N_24616,N_17115,N_19671);
and U24617 (N_24617,N_17281,N_15233);
nand U24618 (N_24618,N_17309,N_17567);
nand U24619 (N_24619,N_17114,N_15399);
xnor U24620 (N_24620,N_16687,N_18807);
nand U24621 (N_24621,N_16808,N_17730);
or U24622 (N_24622,N_15543,N_19973);
or U24623 (N_24623,N_17065,N_15497);
or U24624 (N_24624,N_19222,N_18040);
nor U24625 (N_24625,N_17268,N_18294);
xor U24626 (N_24626,N_19696,N_15928);
nor U24627 (N_24627,N_17970,N_19415);
and U24628 (N_24628,N_16340,N_19904);
or U24629 (N_24629,N_17382,N_19345);
nor U24630 (N_24630,N_16921,N_19633);
xnor U24631 (N_24631,N_19403,N_18580);
nand U24632 (N_24632,N_17030,N_15039);
xnor U24633 (N_24633,N_15546,N_18916);
nand U24634 (N_24634,N_15955,N_18350);
nor U24635 (N_24635,N_19447,N_15729);
or U24636 (N_24636,N_19531,N_15581);
nor U24637 (N_24637,N_16609,N_17928);
nand U24638 (N_24638,N_18190,N_16822);
or U24639 (N_24639,N_15198,N_16738);
nor U24640 (N_24640,N_19479,N_15090);
or U24641 (N_24641,N_19125,N_19802);
nor U24642 (N_24642,N_17130,N_19146);
and U24643 (N_24643,N_16312,N_15216);
and U24644 (N_24644,N_15952,N_16370);
and U24645 (N_24645,N_17315,N_15618);
xnor U24646 (N_24646,N_17015,N_16159);
nor U24647 (N_24647,N_16123,N_16432);
and U24648 (N_24648,N_16307,N_19149);
or U24649 (N_24649,N_16573,N_16316);
and U24650 (N_24650,N_15657,N_19822);
or U24651 (N_24651,N_17317,N_18621);
nor U24652 (N_24652,N_18659,N_18877);
or U24653 (N_24653,N_16837,N_19549);
or U24654 (N_24654,N_18160,N_16608);
or U24655 (N_24655,N_15419,N_15388);
and U24656 (N_24656,N_18248,N_19597);
and U24657 (N_24657,N_17340,N_19850);
or U24658 (N_24658,N_17150,N_15081);
or U24659 (N_24659,N_15625,N_15030);
xor U24660 (N_24660,N_19219,N_18483);
and U24661 (N_24661,N_18563,N_17933);
or U24662 (N_24662,N_16137,N_18500);
or U24663 (N_24663,N_17408,N_15830);
nor U24664 (N_24664,N_18354,N_15043);
or U24665 (N_24665,N_17599,N_16771);
nand U24666 (N_24666,N_16616,N_16218);
and U24667 (N_24667,N_19215,N_17467);
or U24668 (N_24668,N_18334,N_18949);
nor U24669 (N_24669,N_19487,N_15832);
xor U24670 (N_24670,N_16873,N_18633);
nor U24671 (N_24671,N_19496,N_19149);
or U24672 (N_24672,N_15959,N_17862);
or U24673 (N_24673,N_16632,N_18221);
nand U24674 (N_24674,N_19369,N_15913);
xnor U24675 (N_24675,N_19802,N_15100);
or U24676 (N_24676,N_18179,N_18313);
nand U24677 (N_24677,N_19572,N_19268);
and U24678 (N_24678,N_16383,N_16799);
nand U24679 (N_24679,N_18169,N_17873);
and U24680 (N_24680,N_19363,N_16408);
xnor U24681 (N_24681,N_15855,N_15206);
nor U24682 (N_24682,N_16026,N_16275);
and U24683 (N_24683,N_15946,N_19406);
xor U24684 (N_24684,N_19441,N_17332);
and U24685 (N_24685,N_15283,N_16128);
nand U24686 (N_24686,N_16639,N_18650);
nor U24687 (N_24687,N_17917,N_18896);
and U24688 (N_24688,N_17413,N_19310);
nand U24689 (N_24689,N_19307,N_16235);
nor U24690 (N_24690,N_16034,N_19709);
nand U24691 (N_24691,N_17208,N_19854);
nor U24692 (N_24692,N_16825,N_19902);
nand U24693 (N_24693,N_16334,N_17398);
nand U24694 (N_24694,N_19534,N_19581);
or U24695 (N_24695,N_17917,N_15221);
nand U24696 (N_24696,N_18165,N_18919);
nand U24697 (N_24697,N_19333,N_17613);
or U24698 (N_24698,N_18324,N_19073);
or U24699 (N_24699,N_19395,N_15758);
nand U24700 (N_24700,N_19969,N_17004);
and U24701 (N_24701,N_18890,N_17702);
nor U24702 (N_24702,N_17909,N_18835);
nor U24703 (N_24703,N_18809,N_15653);
and U24704 (N_24704,N_19365,N_18270);
or U24705 (N_24705,N_16515,N_15201);
or U24706 (N_24706,N_16511,N_15144);
or U24707 (N_24707,N_15396,N_19123);
and U24708 (N_24708,N_16179,N_15396);
nor U24709 (N_24709,N_19042,N_19673);
nand U24710 (N_24710,N_15225,N_16409);
nor U24711 (N_24711,N_15759,N_18873);
or U24712 (N_24712,N_16791,N_16192);
or U24713 (N_24713,N_18681,N_19827);
nand U24714 (N_24714,N_19256,N_16030);
and U24715 (N_24715,N_17881,N_18355);
or U24716 (N_24716,N_15260,N_15306);
nor U24717 (N_24717,N_19449,N_15002);
nand U24718 (N_24718,N_17553,N_18550);
nand U24719 (N_24719,N_17228,N_18013);
nor U24720 (N_24720,N_16556,N_16939);
nand U24721 (N_24721,N_15182,N_16789);
nor U24722 (N_24722,N_17090,N_16769);
xnor U24723 (N_24723,N_19230,N_15318);
and U24724 (N_24724,N_18959,N_18024);
xnor U24725 (N_24725,N_18439,N_18165);
nand U24726 (N_24726,N_19485,N_15527);
and U24727 (N_24727,N_17578,N_19624);
nor U24728 (N_24728,N_18202,N_16806);
nor U24729 (N_24729,N_16694,N_18652);
nor U24730 (N_24730,N_17107,N_16986);
or U24731 (N_24731,N_16232,N_19306);
nor U24732 (N_24732,N_17955,N_19345);
or U24733 (N_24733,N_18537,N_19067);
and U24734 (N_24734,N_15396,N_18953);
nor U24735 (N_24735,N_18702,N_19762);
or U24736 (N_24736,N_16013,N_18357);
or U24737 (N_24737,N_16195,N_18064);
and U24738 (N_24738,N_18504,N_18594);
nor U24739 (N_24739,N_16497,N_17682);
or U24740 (N_24740,N_18483,N_17651);
nor U24741 (N_24741,N_19438,N_18869);
nor U24742 (N_24742,N_18279,N_15281);
or U24743 (N_24743,N_19715,N_16693);
and U24744 (N_24744,N_15910,N_18069);
nor U24745 (N_24745,N_16448,N_17436);
nand U24746 (N_24746,N_19607,N_18377);
nand U24747 (N_24747,N_17612,N_19730);
nand U24748 (N_24748,N_16436,N_19575);
and U24749 (N_24749,N_16707,N_16451);
nor U24750 (N_24750,N_19860,N_15525);
nand U24751 (N_24751,N_17887,N_19986);
nand U24752 (N_24752,N_16197,N_16762);
nor U24753 (N_24753,N_19372,N_17783);
and U24754 (N_24754,N_15671,N_18859);
or U24755 (N_24755,N_19613,N_17839);
nor U24756 (N_24756,N_19244,N_17980);
and U24757 (N_24757,N_16736,N_15627);
nor U24758 (N_24758,N_19991,N_17664);
nor U24759 (N_24759,N_19420,N_16818);
nand U24760 (N_24760,N_18239,N_19841);
xor U24761 (N_24761,N_18445,N_19797);
nand U24762 (N_24762,N_18880,N_17661);
and U24763 (N_24763,N_19749,N_16132);
nor U24764 (N_24764,N_16999,N_17017);
or U24765 (N_24765,N_15638,N_16868);
nand U24766 (N_24766,N_16366,N_17479);
nand U24767 (N_24767,N_16148,N_19533);
or U24768 (N_24768,N_16691,N_18146);
or U24769 (N_24769,N_17334,N_16187);
nand U24770 (N_24770,N_16539,N_15418);
and U24771 (N_24771,N_17025,N_15755);
nor U24772 (N_24772,N_19304,N_16659);
nor U24773 (N_24773,N_15583,N_18319);
or U24774 (N_24774,N_16325,N_15487);
nand U24775 (N_24775,N_17729,N_19646);
or U24776 (N_24776,N_18759,N_19330);
or U24777 (N_24777,N_17726,N_16669);
nand U24778 (N_24778,N_18259,N_19121);
nor U24779 (N_24779,N_18543,N_16897);
nor U24780 (N_24780,N_17361,N_15142);
or U24781 (N_24781,N_15417,N_17002);
and U24782 (N_24782,N_17995,N_19858);
nand U24783 (N_24783,N_19270,N_18700);
or U24784 (N_24784,N_15094,N_17678);
and U24785 (N_24785,N_17168,N_16969);
or U24786 (N_24786,N_15710,N_18184);
and U24787 (N_24787,N_17054,N_16160);
and U24788 (N_24788,N_18394,N_17515);
or U24789 (N_24789,N_17073,N_18147);
nand U24790 (N_24790,N_18288,N_18828);
nor U24791 (N_24791,N_18761,N_16000);
xnor U24792 (N_24792,N_19896,N_16177);
nand U24793 (N_24793,N_15214,N_18170);
nand U24794 (N_24794,N_19070,N_19810);
and U24795 (N_24795,N_17362,N_15699);
nor U24796 (N_24796,N_15058,N_15483);
and U24797 (N_24797,N_16470,N_19236);
nor U24798 (N_24798,N_16195,N_15741);
nor U24799 (N_24799,N_15775,N_19917);
and U24800 (N_24800,N_16677,N_16900);
nand U24801 (N_24801,N_17013,N_16593);
nor U24802 (N_24802,N_19865,N_18000);
nor U24803 (N_24803,N_17259,N_18481);
nor U24804 (N_24804,N_15954,N_15950);
xnor U24805 (N_24805,N_17896,N_15124);
or U24806 (N_24806,N_16427,N_18959);
nor U24807 (N_24807,N_16476,N_19005);
nor U24808 (N_24808,N_15866,N_18895);
nor U24809 (N_24809,N_17035,N_16438);
nand U24810 (N_24810,N_15939,N_16526);
nand U24811 (N_24811,N_16413,N_16141);
or U24812 (N_24812,N_19637,N_17555);
and U24813 (N_24813,N_15499,N_16747);
xnor U24814 (N_24814,N_17568,N_16650);
or U24815 (N_24815,N_16942,N_19926);
xor U24816 (N_24816,N_19260,N_18188);
nand U24817 (N_24817,N_15402,N_19870);
nand U24818 (N_24818,N_15398,N_19731);
xnor U24819 (N_24819,N_17779,N_16230);
and U24820 (N_24820,N_15587,N_15206);
nor U24821 (N_24821,N_16911,N_16630);
and U24822 (N_24822,N_17885,N_15285);
and U24823 (N_24823,N_17661,N_17141);
xor U24824 (N_24824,N_18212,N_19964);
or U24825 (N_24825,N_17625,N_15493);
xnor U24826 (N_24826,N_15006,N_18426);
nor U24827 (N_24827,N_15148,N_16432);
or U24828 (N_24828,N_18390,N_18500);
nand U24829 (N_24829,N_17664,N_15684);
or U24830 (N_24830,N_19475,N_15497);
and U24831 (N_24831,N_15041,N_17207);
or U24832 (N_24832,N_18475,N_18889);
nand U24833 (N_24833,N_16334,N_17036);
nand U24834 (N_24834,N_18793,N_18454);
nor U24835 (N_24835,N_15207,N_19934);
nand U24836 (N_24836,N_18918,N_16122);
or U24837 (N_24837,N_18281,N_18053);
nand U24838 (N_24838,N_18656,N_18132);
and U24839 (N_24839,N_19904,N_18652);
and U24840 (N_24840,N_16044,N_16749);
nor U24841 (N_24841,N_17360,N_18659);
xor U24842 (N_24842,N_17503,N_15879);
and U24843 (N_24843,N_16094,N_19222);
and U24844 (N_24844,N_17238,N_19467);
nand U24845 (N_24845,N_17134,N_18851);
nor U24846 (N_24846,N_19754,N_15526);
nand U24847 (N_24847,N_15784,N_15628);
nor U24848 (N_24848,N_16232,N_18048);
and U24849 (N_24849,N_17647,N_17777);
or U24850 (N_24850,N_15401,N_17484);
nand U24851 (N_24851,N_15898,N_16262);
nor U24852 (N_24852,N_17516,N_19364);
or U24853 (N_24853,N_16459,N_16025);
nor U24854 (N_24854,N_18391,N_15704);
and U24855 (N_24855,N_18582,N_18082);
nand U24856 (N_24856,N_19162,N_17700);
or U24857 (N_24857,N_19312,N_16362);
and U24858 (N_24858,N_17835,N_15540);
or U24859 (N_24859,N_18877,N_15271);
nor U24860 (N_24860,N_19228,N_17411);
and U24861 (N_24861,N_18502,N_16546);
nand U24862 (N_24862,N_15435,N_18788);
and U24863 (N_24863,N_15515,N_17378);
or U24864 (N_24864,N_17371,N_19764);
nand U24865 (N_24865,N_19852,N_18962);
and U24866 (N_24866,N_15484,N_19968);
and U24867 (N_24867,N_18076,N_17377);
nor U24868 (N_24868,N_16908,N_16754);
and U24869 (N_24869,N_15073,N_19087);
and U24870 (N_24870,N_19426,N_19169);
nand U24871 (N_24871,N_19118,N_17893);
and U24872 (N_24872,N_19700,N_15367);
nand U24873 (N_24873,N_18952,N_16027);
and U24874 (N_24874,N_19287,N_18354);
nand U24875 (N_24875,N_18429,N_15020);
xor U24876 (N_24876,N_17507,N_16964);
and U24877 (N_24877,N_16771,N_18435);
xor U24878 (N_24878,N_19342,N_18566);
nor U24879 (N_24879,N_19958,N_17924);
nand U24880 (N_24880,N_17175,N_17418);
or U24881 (N_24881,N_19534,N_16960);
and U24882 (N_24882,N_17578,N_18678);
or U24883 (N_24883,N_17324,N_15159);
or U24884 (N_24884,N_17813,N_18615);
nor U24885 (N_24885,N_18218,N_19109);
and U24886 (N_24886,N_18756,N_17777);
and U24887 (N_24887,N_16707,N_17315);
xor U24888 (N_24888,N_16689,N_19479);
nand U24889 (N_24889,N_16341,N_19374);
and U24890 (N_24890,N_17420,N_16047);
nand U24891 (N_24891,N_16898,N_19297);
nor U24892 (N_24892,N_16025,N_18891);
nor U24893 (N_24893,N_17205,N_17969);
nor U24894 (N_24894,N_19099,N_18534);
or U24895 (N_24895,N_15189,N_18502);
nor U24896 (N_24896,N_16572,N_16827);
nor U24897 (N_24897,N_15556,N_16412);
or U24898 (N_24898,N_16999,N_18327);
nor U24899 (N_24899,N_19292,N_19775);
nor U24900 (N_24900,N_16795,N_16639);
nand U24901 (N_24901,N_15041,N_18723);
and U24902 (N_24902,N_15096,N_17780);
or U24903 (N_24903,N_19512,N_18162);
or U24904 (N_24904,N_19017,N_19961);
and U24905 (N_24905,N_16989,N_15516);
nor U24906 (N_24906,N_18475,N_17569);
and U24907 (N_24907,N_18459,N_18616);
nand U24908 (N_24908,N_15473,N_16951);
nor U24909 (N_24909,N_16975,N_17100);
or U24910 (N_24910,N_18564,N_17769);
or U24911 (N_24911,N_19057,N_15938);
and U24912 (N_24912,N_19209,N_15329);
nand U24913 (N_24913,N_18012,N_16088);
or U24914 (N_24914,N_18063,N_15438);
or U24915 (N_24915,N_15085,N_17776);
nor U24916 (N_24916,N_18179,N_19601);
or U24917 (N_24917,N_18381,N_16965);
or U24918 (N_24918,N_16811,N_18252);
and U24919 (N_24919,N_16388,N_15678);
nor U24920 (N_24920,N_19716,N_18379);
nand U24921 (N_24921,N_16555,N_18599);
and U24922 (N_24922,N_16394,N_18615);
nor U24923 (N_24923,N_18275,N_18454);
nor U24924 (N_24924,N_19050,N_17526);
and U24925 (N_24925,N_16509,N_18782);
xor U24926 (N_24926,N_19692,N_15976);
and U24927 (N_24927,N_16685,N_19690);
nor U24928 (N_24928,N_18200,N_15158);
or U24929 (N_24929,N_18014,N_19647);
or U24930 (N_24930,N_15585,N_17256);
nand U24931 (N_24931,N_18353,N_16728);
nand U24932 (N_24932,N_15699,N_17009);
nand U24933 (N_24933,N_17016,N_18842);
or U24934 (N_24934,N_15356,N_15121);
and U24935 (N_24935,N_18229,N_18642);
nand U24936 (N_24936,N_19805,N_15516);
nor U24937 (N_24937,N_15049,N_15361);
or U24938 (N_24938,N_19955,N_15444);
nor U24939 (N_24939,N_19321,N_19453);
nor U24940 (N_24940,N_17724,N_18698);
nand U24941 (N_24941,N_15247,N_17727);
or U24942 (N_24942,N_16867,N_15428);
nor U24943 (N_24943,N_17683,N_18253);
nor U24944 (N_24944,N_19027,N_17111);
nand U24945 (N_24945,N_15139,N_15930);
nand U24946 (N_24946,N_18069,N_17911);
and U24947 (N_24947,N_16110,N_17603);
nor U24948 (N_24948,N_15252,N_19705);
and U24949 (N_24949,N_19730,N_17281);
and U24950 (N_24950,N_15659,N_16118);
and U24951 (N_24951,N_17588,N_19294);
or U24952 (N_24952,N_18194,N_17832);
or U24953 (N_24953,N_17334,N_18797);
nand U24954 (N_24954,N_18004,N_18162);
and U24955 (N_24955,N_15784,N_16734);
and U24956 (N_24956,N_15380,N_16946);
nand U24957 (N_24957,N_19757,N_15405);
xor U24958 (N_24958,N_15940,N_15354);
and U24959 (N_24959,N_17031,N_17819);
xor U24960 (N_24960,N_16047,N_18030);
nand U24961 (N_24961,N_17625,N_16005);
xor U24962 (N_24962,N_17163,N_18369);
nor U24963 (N_24963,N_19898,N_18038);
nand U24964 (N_24964,N_16404,N_18005);
nor U24965 (N_24965,N_18558,N_19416);
nand U24966 (N_24966,N_19611,N_19599);
xor U24967 (N_24967,N_17402,N_18438);
and U24968 (N_24968,N_18671,N_15542);
nand U24969 (N_24969,N_15478,N_19098);
nand U24970 (N_24970,N_15382,N_15280);
or U24971 (N_24971,N_16690,N_16830);
and U24972 (N_24972,N_17992,N_15590);
nor U24973 (N_24973,N_18913,N_18082);
nand U24974 (N_24974,N_17220,N_15545);
nor U24975 (N_24975,N_18764,N_16373);
or U24976 (N_24976,N_18662,N_16989);
nand U24977 (N_24977,N_17580,N_19726);
nor U24978 (N_24978,N_16616,N_15275);
nand U24979 (N_24979,N_17210,N_16235);
nor U24980 (N_24980,N_18308,N_15887);
nor U24981 (N_24981,N_17817,N_15340);
nor U24982 (N_24982,N_16705,N_19730);
nor U24983 (N_24983,N_16098,N_16337);
and U24984 (N_24984,N_17969,N_15445);
nor U24985 (N_24985,N_15198,N_15110);
xor U24986 (N_24986,N_18305,N_19837);
nand U24987 (N_24987,N_15513,N_16932);
or U24988 (N_24988,N_18081,N_16240);
xnor U24989 (N_24989,N_15625,N_18959);
or U24990 (N_24990,N_16486,N_18284);
nand U24991 (N_24991,N_15816,N_16759);
nor U24992 (N_24992,N_18827,N_19460);
and U24993 (N_24993,N_17771,N_18450);
and U24994 (N_24994,N_16749,N_18324);
and U24995 (N_24995,N_18367,N_17080);
nand U24996 (N_24996,N_19191,N_18216);
xnor U24997 (N_24997,N_15595,N_16740);
and U24998 (N_24998,N_17299,N_18511);
and U24999 (N_24999,N_19700,N_15864);
nand U25000 (N_25000,N_24808,N_24472);
and U25001 (N_25001,N_24750,N_21557);
or U25002 (N_25002,N_22164,N_24674);
nand U25003 (N_25003,N_20885,N_22533);
xor U25004 (N_25004,N_21112,N_23856);
and U25005 (N_25005,N_21042,N_21723);
or U25006 (N_25006,N_23354,N_20327);
xor U25007 (N_25007,N_22731,N_21802);
or U25008 (N_25008,N_20160,N_22680);
xor U25009 (N_25009,N_20624,N_23003);
xnor U25010 (N_25010,N_23889,N_24470);
and U25011 (N_25011,N_23147,N_23995);
or U25012 (N_25012,N_22694,N_20292);
nand U25013 (N_25013,N_22967,N_22051);
nor U25014 (N_25014,N_20842,N_22188);
or U25015 (N_25015,N_22190,N_21067);
nor U25016 (N_25016,N_24943,N_20094);
nand U25017 (N_25017,N_24695,N_22564);
and U25018 (N_25018,N_24967,N_22722);
nor U25019 (N_25019,N_21263,N_24792);
and U25020 (N_25020,N_20429,N_24208);
nor U25021 (N_25021,N_20375,N_20305);
or U25022 (N_25022,N_21897,N_21334);
nand U25023 (N_25023,N_24198,N_21249);
nand U25024 (N_25024,N_22105,N_24909);
and U25025 (N_25025,N_23890,N_23182);
nand U25026 (N_25026,N_20574,N_20288);
or U25027 (N_25027,N_20706,N_20577);
nand U25028 (N_25028,N_24012,N_21383);
or U25029 (N_25029,N_22862,N_21725);
and U25030 (N_25030,N_23608,N_24798);
nor U25031 (N_25031,N_23069,N_23283);
or U25032 (N_25032,N_23959,N_24234);
or U25033 (N_25033,N_21553,N_21406);
nor U25034 (N_25034,N_24227,N_23242);
or U25035 (N_25035,N_20037,N_22588);
or U25036 (N_25036,N_21985,N_20588);
and U25037 (N_25037,N_24144,N_23037);
or U25038 (N_25038,N_20064,N_23979);
or U25039 (N_25039,N_20736,N_24989);
xnor U25040 (N_25040,N_21801,N_23462);
and U25041 (N_25041,N_20204,N_21963);
and U25042 (N_25042,N_23918,N_23797);
and U25043 (N_25043,N_22599,N_22992);
nor U25044 (N_25044,N_21767,N_20866);
or U25045 (N_25045,N_20622,N_20551);
or U25046 (N_25046,N_22393,N_24405);
and U25047 (N_25047,N_21135,N_20262);
and U25048 (N_25048,N_23595,N_23492);
nor U25049 (N_25049,N_23371,N_21501);
and U25050 (N_25050,N_21270,N_22450);
nor U25051 (N_25051,N_24069,N_20059);
and U25052 (N_25052,N_22742,N_20272);
nand U25053 (N_25053,N_23596,N_21799);
or U25054 (N_25054,N_23772,N_23113);
nor U25055 (N_25055,N_21336,N_24694);
xnor U25056 (N_25056,N_21573,N_23080);
nand U25057 (N_25057,N_21397,N_23920);
nor U25058 (N_25058,N_23620,N_21746);
nor U25059 (N_25059,N_23280,N_22635);
xor U25060 (N_25060,N_23142,N_21011);
nor U25061 (N_25061,N_21450,N_22598);
or U25062 (N_25062,N_20744,N_21264);
xor U25063 (N_25063,N_23038,N_23234);
and U25064 (N_25064,N_20694,N_22622);
nand U25065 (N_25065,N_22053,N_24457);
or U25066 (N_25066,N_20021,N_21398);
xor U25067 (N_25067,N_20854,N_24094);
nand U25068 (N_25068,N_23087,N_22295);
nor U25069 (N_25069,N_24669,N_24140);
nand U25070 (N_25070,N_24135,N_24035);
xor U25071 (N_25071,N_20106,N_23843);
xor U25072 (N_25072,N_20897,N_20374);
or U25073 (N_25073,N_22034,N_24038);
nand U25074 (N_25074,N_24788,N_22528);
or U25075 (N_25075,N_21731,N_24157);
and U25076 (N_25076,N_21295,N_22878);
and U25077 (N_25077,N_24848,N_22296);
nand U25078 (N_25078,N_24937,N_20643);
nand U25079 (N_25079,N_20584,N_20051);
xor U25080 (N_25080,N_21500,N_24718);
and U25081 (N_25081,N_21818,N_21100);
and U25082 (N_25082,N_21780,N_22741);
or U25083 (N_25083,N_23128,N_23413);
and U25084 (N_25084,N_24359,N_22601);
nor U25085 (N_25085,N_23955,N_20916);
nor U25086 (N_25086,N_23992,N_22559);
xor U25087 (N_25087,N_20162,N_23146);
nor U25088 (N_25088,N_22752,N_20930);
and U25089 (N_25089,N_21179,N_20118);
or U25090 (N_25090,N_24830,N_21838);
nand U25091 (N_25091,N_20027,N_21886);
or U25092 (N_25092,N_21856,N_22772);
nand U25093 (N_25093,N_21745,N_21621);
nand U25094 (N_25094,N_23335,N_21775);
and U25095 (N_25095,N_21662,N_20435);
and U25096 (N_25096,N_20926,N_23731);
and U25097 (N_25097,N_21638,N_21187);
and U25098 (N_25098,N_23961,N_22327);
nor U25099 (N_25099,N_22616,N_23163);
and U25100 (N_25100,N_20666,N_21485);
nor U25101 (N_25101,N_21438,N_20750);
and U25102 (N_25102,N_23686,N_23783);
nand U25103 (N_25103,N_20069,N_22416);
nand U25104 (N_25104,N_22836,N_22063);
xnor U25105 (N_25105,N_21456,N_23557);
or U25106 (N_25106,N_24620,N_24513);
xor U25107 (N_25107,N_20680,N_20806);
nor U25108 (N_25108,N_23839,N_22012);
or U25109 (N_25109,N_20674,N_24995);
and U25110 (N_25110,N_22541,N_20180);
and U25111 (N_25111,N_23018,N_21218);
or U25112 (N_25112,N_23135,N_20539);
nand U25113 (N_25113,N_24266,N_21589);
or U25114 (N_25114,N_21867,N_24195);
xnor U25115 (N_25115,N_20194,N_20918);
nor U25116 (N_25116,N_21722,N_24554);
xnor U25117 (N_25117,N_22817,N_21835);
or U25118 (N_25118,N_24782,N_21757);
or U25119 (N_25119,N_20271,N_24019);
nand U25120 (N_25120,N_21971,N_22434);
nand U25121 (N_25121,N_21462,N_24084);
and U25122 (N_25122,N_24889,N_22647);
nor U25123 (N_25123,N_21890,N_20083);
or U25124 (N_25124,N_22284,N_22766);
and U25125 (N_25125,N_23415,N_21453);
nand U25126 (N_25126,N_23987,N_22414);
nor U25127 (N_25127,N_24357,N_20815);
nand U25128 (N_25128,N_22511,N_22659);
nor U25129 (N_25129,N_21110,N_24903);
nand U25130 (N_25130,N_24600,N_22707);
nand U25131 (N_25131,N_20128,N_23793);
nand U25132 (N_25132,N_23359,N_23784);
xnor U25133 (N_25133,N_22687,N_23516);
or U25134 (N_25134,N_20058,N_20267);
nor U25135 (N_25135,N_21504,N_21093);
nand U25136 (N_25136,N_20936,N_24429);
nand U25137 (N_25137,N_22787,N_23118);
or U25138 (N_25138,N_24948,N_24957);
or U25139 (N_25139,N_22775,N_24459);
and U25140 (N_25140,N_22555,N_20260);
nor U25141 (N_25141,N_20434,N_24502);
nor U25142 (N_25142,N_20320,N_23198);
nor U25143 (N_25143,N_20682,N_20556);
and U25144 (N_25144,N_21498,N_21915);
and U25145 (N_25145,N_24749,N_23081);
nand U25146 (N_25146,N_22235,N_21178);
or U25147 (N_25147,N_24020,N_20036);
and U25148 (N_25148,N_21229,N_22308);
nor U25149 (N_25149,N_22663,N_24462);
nor U25150 (N_25150,N_21044,N_21900);
xnor U25151 (N_25151,N_21743,N_21477);
or U25152 (N_25152,N_21733,N_20505);
nand U25153 (N_25153,N_23704,N_22797);
xor U25154 (N_25154,N_21030,N_23877);
and U25155 (N_25155,N_23989,N_21469);
nand U25156 (N_25156,N_21926,N_23144);
or U25157 (N_25157,N_24703,N_21415);
or U25158 (N_25158,N_20686,N_22332);
or U25159 (N_25159,N_22170,N_23226);
nor U25160 (N_25160,N_23040,N_21108);
nor U25161 (N_25161,N_23327,N_20595);
xnor U25162 (N_25162,N_21858,N_21615);
nand U25163 (N_25163,N_23747,N_23068);
or U25164 (N_25164,N_21672,N_24833);
or U25165 (N_25165,N_22801,N_22789);
or U25166 (N_25166,N_23153,N_23716);
nand U25167 (N_25167,N_21717,N_21987);
or U25168 (N_25168,N_21774,N_23074);
nor U25169 (N_25169,N_22065,N_23973);
nor U25170 (N_25170,N_20544,N_22904);
and U25171 (N_25171,N_21523,N_22685);
nor U25172 (N_25172,N_22173,N_22861);
nand U25173 (N_25173,N_23493,N_21944);
xor U25174 (N_25174,N_23565,N_20486);
nand U25175 (N_25175,N_23116,N_21443);
and U25176 (N_25176,N_20931,N_23422);
and U25177 (N_25177,N_24872,N_22761);
or U25178 (N_25178,N_23237,N_20517);
nor U25179 (N_25179,N_22712,N_20279);
xor U25180 (N_25180,N_24315,N_20452);
nor U25181 (N_25181,N_20131,N_24886);
xor U25182 (N_25182,N_20770,N_24356);
xor U25183 (N_25183,N_23452,N_23501);
nand U25184 (N_25184,N_21982,N_20074);
nor U25185 (N_25185,N_21768,N_22197);
or U25186 (N_25186,N_23864,N_23336);
or U25187 (N_25187,N_20468,N_21511);
and U25188 (N_25188,N_23477,N_24192);
and U25189 (N_25189,N_23360,N_22859);
nand U25190 (N_25190,N_21430,N_20910);
or U25191 (N_25191,N_23795,N_23285);
and U25192 (N_25192,N_20711,N_21008);
and U25193 (N_25193,N_24021,N_21951);
nor U25194 (N_25194,N_20503,N_23779);
nand U25195 (N_25195,N_23088,N_23296);
nand U25196 (N_25196,N_24720,N_20585);
and U25197 (N_25197,N_22263,N_23152);
or U25198 (N_25198,N_20399,N_22944);
xnor U25199 (N_25199,N_23005,N_24312);
nor U25200 (N_25200,N_20309,N_21538);
nor U25201 (N_25201,N_22069,N_20735);
and U25202 (N_25202,N_24481,N_22786);
and U25203 (N_25203,N_22446,N_21822);
xnor U25204 (N_25204,N_22335,N_22668);
or U25205 (N_25205,N_22056,N_20566);
nand U25206 (N_25206,N_22782,N_21750);
nand U25207 (N_25207,N_24216,N_23885);
and U25208 (N_25208,N_20834,N_22223);
nor U25209 (N_25209,N_22358,N_22047);
and U25210 (N_25210,N_24221,N_22392);
nor U25211 (N_25211,N_23706,N_21842);
or U25212 (N_25212,N_21107,N_23337);
or U25213 (N_25213,N_20299,N_22273);
nand U25214 (N_25214,N_21947,N_22032);
nand U25215 (N_25215,N_23970,N_24278);
or U25216 (N_25216,N_22113,N_24797);
nand U25217 (N_25217,N_22045,N_21350);
or U25218 (N_25218,N_23489,N_22457);
nor U25219 (N_25219,N_24860,N_22409);
and U25220 (N_25220,N_20480,N_22042);
nor U25221 (N_25221,N_22341,N_23692);
nor U25222 (N_25222,N_22914,N_21751);
xor U25223 (N_25223,N_22426,N_21038);
or U25224 (N_25224,N_20779,N_21305);
nor U25225 (N_25225,N_23550,N_23913);
or U25226 (N_25226,N_23670,N_21661);
nor U25227 (N_25227,N_24888,N_22945);
nand U25228 (N_25228,N_22950,N_21075);
nand U25229 (N_25229,N_21645,N_20247);
or U25230 (N_25230,N_21316,N_20501);
and U25231 (N_25231,N_21091,N_22626);
and U25232 (N_25232,N_22571,N_24007);
or U25233 (N_25233,N_21495,N_22613);
nand U25234 (N_25234,N_24977,N_23494);
nor U25235 (N_25235,N_23714,N_23560);
and U25236 (N_25236,N_21377,N_24760);
xor U25237 (N_25237,N_20243,N_22200);
and U25238 (N_25238,N_20883,N_21676);
or U25239 (N_25239,N_21544,N_22675);
or U25240 (N_25240,N_24086,N_22184);
nand U25241 (N_25241,N_22812,N_24638);
nand U25242 (N_25242,N_24956,N_21532);
nand U25243 (N_25243,N_21126,N_20147);
or U25244 (N_25244,N_23257,N_24906);
nor U25245 (N_25245,N_21660,N_24257);
nand U25246 (N_25246,N_22863,N_21310);
and U25247 (N_25247,N_21580,N_24374);
nor U25248 (N_25248,N_24342,N_21476);
and U25249 (N_25249,N_22204,N_22606);
or U25250 (N_25250,N_23800,N_24656);
or U25251 (N_25251,N_23721,N_23181);
nor U25252 (N_25252,N_23259,N_21616);
or U25253 (N_25253,N_20889,N_23203);
and U25254 (N_25254,N_20870,N_22700);
nand U25255 (N_25255,N_20984,N_23591);
xnor U25256 (N_25256,N_21540,N_23936);
and U25257 (N_25257,N_21535,N_21781);
and U25258 (N_25258,N_21991,N_21988);
and U25259 (N_25259,N_20315,N_24183);
or U25260 (N_25260,N_21173,N_21932);
nand U25261 (N_25261,N_23272,N_20342);
nand U25262 (N_25262,N_21446,N_21650);
nor U25263 (N_25263,N_20265,N_20176);
nand U25264 (N_25264,N_20432,N_20905);
xnor U25265 (N_25265,N_21514,N_21211);
or U25266 (N_25266,N_21084,N_20678);
nand U25267 (N_25267,N_22552,N_24355);
nor U25268 (N_25268,N_21222,N_24509);
nand U25269 (N_25269,N_20290,N_24287);
nor U25270 (N_25270,N_20601,N_23654);
nor U25271 (N_25271,N_24096,N_22145);
xor U25272 (N_25272,N_21680,N_23625);
and U25273 (N_25273,N_21693,N_23490);
nand U25274 (N_25274,N_23811,N_23888);
nor U25275 (N_25275,N_22557,N_21833);
xor U25276 (N_25276,N_22514,N_24304);
or U25277 (N_25277,N_24139,N_20339);
nor U25278 (N_25278,N_22139,N_20990);
and U25279 (N_25279,N_22472,N_21040);
and U25280 (N_25280,N_21980,N_22444);
nand U25281 (N_25281,N_24710,N_22101);
and U25282 (N_25282,N_21828,N_21382);
nand U25283 (N_25283,N_23472,N_21655);
or U25284 (N_25284,N_22060,N_20301);
nand U25285 (N_25285,N_21508,N_20338);
nor U25286 (N_25286,N_21015,N_21132);
or U25287 (N_25287,N_20297,N_24521);
xnor U25288 (N_25288,N_21379,N_24577);
and U25289 (N_25289,N_24448,N_22739);
nand U25290 (N_25290,N_21512,N_22447);
or U25291 (N_25291,N_21527,N_23734);
nand U25292 (N_25292,N_22891,N_23943);
or U25293 (N_25293,N_24248,N_20580);
nor U25294 (N_25294,N_23394,N_22303);
and U25295 (N_25295,N_21599,N_24305);
or U25296 (N_25296,N_22664,N_21820);
nor U25297 (N_25297,N_20002,N_22090);
nand U25298 (N_25298,N_21570,N_20158);
nor U25299 (N_25299,N_21442,N_20859);
and U25300 (N_25300,N_21546,N_20394);
xnor U25301 (N_25301,N_22765,N_24874);
nand U25302 (N_25302,N_24325,N_20531);
or U25303 (N_25303,N_23642,N_20422);
or U25304 (N_25304,N_22109,N_22560);
and U25305 (N_25305,N_22026,N_22758);
nor U25306 (N_25306,N_24927,N_23491);
and U25307 (N_25307,N_20105,N_24804);
xor U25308 (N_25308,N_21274,N_20616);
nor U25309 (N_25309,N_22780,N_23180);
and U25310 (N_25310,N_24181,N_24009);
nand U25311 (N_25311,N_20203,N_20238);
and U25312 (N_25312,N_24911,N_23008);
xor U25313 (N_25313,N_21455,N_20634);
xnor U25314 (N_25314,N_22344,N_20372);
and U25315 (N_25315,N_20402,N_20075);
nor U25316 (N_25316,N_24384,N_24321);
xnor U25317 (N_25317,N_23053,N_23641);
nand U25318 (N_25318,N_20112,N_21291);
nand U25319 (N_25319,N_22144,N_23769);
and U25320 (N_25320,N_21646,N_24917);
xor U25321 (N_25321,N_20543,N_24487);
nor U25322 (N_25322,N_22316,N_20156);
xnor U25323 (N_25323,N_20840,N_20485);
and U25324 (N_25324,N_22381,N_22917);
or U25325 (N_25325,N_20438,N_23281);
and U25326 (N_25326,N_23112,N_23633);
and U25327 (N_25327,N_20475,N_20006);
nand U25328 (N_25328,N_21016,N_23511);
and U25329 (N_25329,N_24904,N_21425);
or U25330 (N_25330,N_21909,N_22259);
or U25331 (N_25331,N_20398,N_23695);
xnor U25332 (N_25332,N_21308,N_21513);
and U25333 (N_25333,N_20287,N_21727);
or U25334 (N_25334,N_24365,N_20157);
or U25335 (N_25335,N_23278,N_20691);
or U25336 (N_25336,N_22982,N_23759);
and U25337 (N_25337,N_23363,N_24857);
or U25338 (N_25338,N_23914,N_22075);
or U25339 (N_25339,N_21195,N_23332);
and U25340 (N_25340,N_22579,N_22994);
xnor U25341 (N_25341,N_24163,N_22007);
and U25342 (N_25342,N_20011,N_22238);
nand U25343 (N_25343,N_21841,N_22802);
and U25344 (N_25344,N_21868,N_22469);
nor U25345 (N_25345,N_22896,N_24178);
and U25346 (N_25346,N_21927,N_21470);
nand U25347 (N_25347,N_20071,N_24297);
nand U25348 (N_25348,N_22518,N_21635);
nand U25349 (N_25349,N_21748,N_23409);
nand U25350 (N_25350,N_22691,N_20166);
nand U25351 (N_25351,N_22875,N_21454);
nor U25352 (N_25352,N_22014,N_20135);
xnor U25353 (N_25353,N_20860,N_23323);
and U25354 (N_25354,N_20732,N_21531);
and U25355 (N_25355,N_20412,N_21332);
or U25356 (N_25356,N_23515,N_20082);
or U25357 (N_25357,N_21283,N_24252);
nor U25358 (N_25358,N_24476,N_20768);
and U25359 (N_25359,N_23200,N_20043);
or U25360 (N_25360,N_24166,N_24370);
nand U25361 (N_25361,N_21369,N_23300);
or U25362 (N_25362,N_20676,N_24465);
xnor U25363 (N_25363,N_24786,N_20762);
nand U25364 (N_25364,N_20519,N_23222);
xnor U25365 (N_25365,N_23372,N_24660);
nor U25366 (N_25366,N_20725,N_20641);
and U25367 (N_25367,N_23651,N_24998);
and U25368 (N_25368,N_23164,N_20276);
xor U25369 (N_25369,N_23276,N_22540);
nor U25370 (N_25370,N_24298,N_24002);
or U25371 (N_25371,N_24913,N_23166);
xor U25372 (N_25372,N_24552,N_21876);
nand U25373 (N_25373,N_21409,N_20258);
and U25374 (N_25374,N_22930,N_24489);
or U25375 (N_25375,N_22839,N_22454);
or U25376 (N_25376,N_21235,N_23626);
and U25377 (N_25377,N_24124,N_22121);
or U25378 (N_25378,N_22125,N_20314);
nor U25379 (N_25379,N_20493,N_20009);
and U25380 (N_25380,N_24576,N_20708);
or U25381 (N_25381,N_20555,N_23925);
xnor U25382 (N_25382,N_23937,N_21933);
nand U25383 (N_25383,N_22674,N_20459);
nor U25384 (N_25384,N_22634,N_22954);
nor U25385 (N_25385,N_21370,N_22777);
nor U25386 (N_25386,N_21564,N_23815);
xor U25387 (N_25387,N_21819,N_23674);
and U25388 (N_25388,N_20773,N_23831);
xor U25389 (N_25389,N_21879,N_22521);
nor U25390 (N_25390,N_20317,N_22157);
nor U25391 (N_25391,N_24033,N_20726);
or U25392 (N_25392,N_20192,N_23273);
nand U25393 (N_25393,N_22936,N_21471);
nor U25394 (N_25394,N_22743,N_21082);
xnor U25395 (N_25395,N_23917,N_23000);
and U25396 (N_25396,N_21236,N_24344);
xor U25397 (N_25397,N_23265,N_22881);
or U25398 (N_25398,N_23499,N_23046);
and U25399 (N_25399,N_22757,N_21797);
and U25400 (N_25400,N_20031,N_22401);
or U25401 (N_25401,N_20958,N_23867);
xnor U25402 (N_25402,N_20116,N_23509);
nand U25403 (N_25403,N_20099,N_21029);
and U25404 (N_25404,N_23423,N_24683);
and U25405 (N_25405,N_21254,N_22285);
and U25406 (N_25406,N_21571,N_20557);
nor U25407 (N_25407,N_22132,N_24188);
nand U25408 (N_25408,N_21266,N_21697);
nor U25409 (N_25409,N_22278,N_21167);
nand U25410 (N_25410,N_23878,N_21160);
or U25411 (N_25411,N_23709,N_22258);
nand U25412 (N_25412,N_23882,N_24551);
and U25413 (N_25413,N_24985,N_23282);
nand U25414 (N_25414,N_21541,N_23905);
nor U25415 (N_25415,N_24147,N_22079);
or U25416 (N_25416,N_20336,N_20609);
and U25417 (N_25417,N_24654,N_24867);
nor U25418 (N_25418,N_23397,N_22095);
nor U25419 (N_25419,N_22997,N_21039);
and U25420 (N_25420,N_24294,N_20964);
nor U25421 (N_25421,N_23441,N_20463);
nor U25422 (N_25422,N_21817,N_22404);
nand U25423 (N_25423,N_24882,N_20978);
nor U25424 (N_25424,N_23921,N_24617);
xor U25425 (N_25425,N_21217,N_20752);
or U25426 (N_25426,N_21681,N_20717);
or U25427 (N_25427,N_22181,N_22390);
and U25428 (N_25428,N_22524,N_22941);
nor U25429 (N_25429,N_23637,N_23115);
nand U25430 (N_25430,N_22440,N_24735);
nor U25431 (N_25431,N_21296,N_24256);
and U25432 (N_25432,N_21260,N_24742);
or U25433 (N_25433,N_22304,N_24547);
nor U25434 (N_25434,N_21782,N_23597);
or U25435 (N_25435,N_24719,N_24026);
xnor U25436 (N_25436,N_22895,N_22207);
nand U25437 (N_25437,N_22534,N_20410);
or U25438 (N_25438,N_24506,N_20256);
and U25439 (N_25439,N_24421,N_20291);
and U25440 (N_25440,N_22871,N_22495);
or U25441 (N_25441,N_20652,N_23542);
and U25442 (N_25442,N_23944,N_20396);
xnor U25443 (N_25443,N_21567,N_24326);
or U25444 (N_25444,N_22538,N_24066);
xor U25445 (N_25445,N_23322,N_21220);
or U25446 (N_25446,N_20344,N_24328);
nor U25447 (N_25447,N_23621,N_20513);
or U25448 (N_25448,N_24285,N_23151);
or U25449 (N_25449,N_20994,N_23435);
or U25450 (N_25450,N_22085,N_22709);
nor U25451 (N_25451,N_22467,N_22833);
or U25452 (N_25452,N_22522,N_24712);
nand U25453 (N_25453,N_20334,N_22435);
or U25454 (N_25454,N_23176,N_24402);
nor U25455 (N_25455,N_20115,N_21714);
or U25456 (N_25456,N_20799,N_22456);
and U25457 (N_25457,N_20951,N_24938);
or U25458 (N_25458,N_22856,N_20324);
or U25459 (N_25459,N_22824,N_22542);
xnor U25460 (N_25460,N_24338,N_23838);
or U25461 (N_25461,N_20259,N_24450);
xor U25462 (N_25462,N_24189,N_20619);
nand U25463 (N_25463,N_21068,N_20443);
nor U25464 (N_25464,N_23749,N_22030);
and U25465 (N_25465,N_24436,N_20545);
and U25466 (N_25466,N_23907,N_20030);
nand U25467 (N_25467,N_24350,N_21949);
xor U25468 (N_25468,N_21436,N_23975);
nand U25469 (N_25469,N_24032,N_22825);
nor U25470 (N_25470,N_24148,N_20350);
and U25471 (N_25471,N_20229,N_22239);
nand U25472 (N_25472,N_23603,N_21297);
and U25473 (N_25473,N_22214,N_20136);
nand U25474 (N_25474,N_23792,N_20662);
and U25475 (N_25475,N_22338,N_21278);
and U25476 (N_25476,N_23031,N_24934);
or U25477 (N_25477,N_22388,N_24564);
nand U25478 (N_25478,N_24884,N_21941);
nand U25479 (N_25479,N_22718,N_22064);
nor U25480 (N_25480,N_20241,N_22437);
or U25481 (N_25481,N_23999,N_22010);
nor U25482 (N_25482,N_24484,N_23931);
nor U25483 (N_25483,N_21989,N_21188);
and U25484 (N_25484,N_23904,N_24898);
nand U25485 (N_25485,N_22832,N_24275);
or U25486 (N_25486,N_20239,N_23352);
nor U25487 (N_25487,N_22888,N_24090);
xnor U25488 (N_25488,N_23810,N_24612);
and U25489 (N_25489,N_20386,N_22151);
nand U25490 (N_25490,N_24717,N_23030);
and U25491 (N_25491,N_22422,N_20949);
nand U25492 (N_25492,N_23589,N_24991);
nand U25493 (N_25493,N_20720,N_22880);
nand U25494 (N_25494,N_24052,N_21878);
and U25495 (N_25495,N_21507,N_24108);
nor U25496 (N_25496,N_21956,N_21489);
and U25497 (N_25497,N_24692,N_23440);
or U25498 (N_25498,N_24141,N_22903);
nand U25499 (N_25499,N_23240,N_21484);
nor U25500 (N_25500,N_23157,N_24925);
nor U25501 (N_25501,N_20472,N_22512);
nand U25502 (N_25502,N_24693,N_23712);
and U25503 (N_25503,N_23778,N_23017);
nor U25504 (N_25504,N_22412,N_21056);
nor U25505 (N_25505,N_20199,N_24268);
nand U25506 (N_25506,N_21996,N_21981);
xor U25507 (N_25507,N_24990,N_21806);
or U25508 (N_25508,N_23622,N_20182);
and U25509 (N_25509,N_24118,N_20492);
xnor U25510 (N_25510,N_24117,N_20117);
and U25511 (N_25511,N_21643,N_24228);
nor U25512 (N_25512,N_23884,N_22299);
and U25513 (N_25513,N_23250,N_23656);
xnor U25514 (N_25514,N_22037,N_23167);
xor U25515 (N_25515,N_22679,N_24153);
or U25516 (N_25516,N_21969,N_23400);
nand U25517 (N_25517,N_23924,N_21428);
nor U25518 (N_25518,N_23430,N_21911);
xor U25519 (N_25519,N_23184,N_23611);
or U25520 (N_25520,N_21275,N_24714);
or U25521 (N_25521,N_21123,N_24316);
or U25522 (N_25522,N_21788,N_24855);
nor U25523 (N_25523,N_22912,N_20347);
nor U25524 (N_25524,N_21130,N_21027);
nand U25525 (N_25525,N_24591,N_20010);
nor U25526 (N_25526,N_24615,N_23677);
or U25527 (N_25527,N_22172,N_22017);
nor U25528 (N_25528,N_22039,N_24779);
or U25529 (N_25529,N_20950,N_22291);
nor U25530 (N_25530,N_23404,N_23733);
or U25531 (N_25531,N_20923,N_24631);
or U25532 (N_25532,N_24605,N_23875);
and U25533 (N_25533,N_21063,N_21994);
nand U25534 (N_25534,N_23253,N_23421);
or U25535 (N_25535,N_21418,N_21881);
nand U25536 (N_25536,N_23015,N_22086);
and U25537 (N_25537,N_22206,N_22027);
and U25538 (N_25538,N_24527,N_22081);
and U25539 (N_25539,N_20185,N_21061);
nand U25540 (N_25540,N_24335,N_24277);
nand U25541 (N_25541,N_23393,N_23785);
or U25542 (N_25542,N_21482,N_23190);
nor U25543 (N_25543,N_22360,N_21057);
or U25544 (N_25544,N_24241,N_20201);
or U25545 (N_25545,N_22395,N_22166);
and U25546 (N_25546,N_20586,N_23034);
nand U25547 (N_25547,N_21948,N_24373);
or U25548 (N_25548,N_21059,N_20321);
nand U25549 (N_25549,N_20746,N_23236);
xnor U25550 (N_25550,N_20352,N_21182);
xnor U25551 (N_25551,N_21116,N_24048);
or U25552 (N_25552,N_24085,N_23739);
or U25553 (N_25553,N_22724,N_23358);
nor U25554 (N_25554,N_24361,N_22478);
or U25555 (N_25555,N_24924,N_23438);
nor U25556 (N_25556,N_22919,N_24469);
nand U25557 (N_25557,N_21776,N_20437);
and U25558 (N_25558,N_22792,N_20909);
and U25559 (N_25559,N_24736,N_22490);
and U25560 (N_25560,N_21997,N_22840);
or U25561 (N_25561,N_21137,N_22361);
nor U25562 (N_25562,N_22080,N_20046);
nand U25563 (N_25563,N_23583,N_21007);
nor U25564 (N_25564,N_22701,N_21707);
or U25565 (N_25565,N_20200,N_20389);
nor U25566 (N_25566,N_21268,N_22574);
and U25567 (N_25567,N_21323,N_20469);
nor U25568 (N_25568,N_22934,N_22355);
nor U25569 (N_25569,N_20822,N_21276);
or U25570 (N_25570,N_20563,N_24896);
nand U25571 (N_25571,N_23188,N_21639);
nor U25572 (N_25572,N_21018,N_24433);
xnor U25573 (N_25573,N_22900,N_24816);
nand U25574 (N_25574,N_22939,N_23449);
or U25575 (N_25575,N_23098,N_21753);
nor U25576 (N_25576,N_22357,N_20540);
or U25577 (N_25577,N_20390,N_24574);
nor U25578 (N_25578,N_21816,N_23083);
nor U25579 (N_25579,N_20677,N_23558);
nor U25580 (N_25580,N_24826,N_21921);
or U25581 (N_25581,N_24004,N_24819);
or U25582 (N_25582,N_24881,N_22067);
or U25583 (N_25583,N_21191,N_22644);
or U25584 (N_25584,N_24238,N_24870);
nand U25585 (N_25585,N_20535,N_24318);
nor U25586 (N_25586,N_21496,N_23262);
xor U25587 (N_25587,N_24423,N_21744);
nor U25588 (N_25588,N_22452,N_22494);
or U25589 (N_25589,N_22094,N_20364);
or U25590 (N_25590,N_24568,N_21562);
or U25591 (N_25591,N_20101,N_20568);
or U25592 (N_25592,N_20653,N_21486);
xor U25593 (N_25593,N_20733,N_23498);
and U25594 (N_25594,N_22572,N_23717);
nor U25595 (N_25595,N_21728,N_24150);
nor U25596 (N_25596,N_24877,N_24364);
nor U25597 (N_25597,N_23928,N_24636);
nand U25598 (N_25598,N_23871,N_24083);
xnor U25599 (N_25599,N_22177,N_20489);
and U25600 (N_25600,N_20683,N_23009);
nand U25601 (N_25601,N_21458,N_22046);
nor U25602 (N_25602,N_22191,N_23643);
nand U25603 (N_25603,N_22652,N_21036);
or U25604 (N_25604,N_22251,N_20847);
and U25605 (N_25605,N_21269,N_24396);
nor U25606 (N_25606,N_24151,N_20040);
and U25607 (N_25607,N_21355,N_24759);
xnor U25608 (N_25608,N_24045,N_22340);
xor U25609 (N_25609,N_24389,N_22376);
nor U25610 (N_25610,N_23659,N_20440);
nor U25611 (N_25611,N_22287,N_24313);
xor U25612 (N_25612,N_24001,N_21047);
xnor U25613 (N_25613,N_22972,N_22187);
nand U25614 (N_25614,N_22520,N_22868);
or U25615 (N_25615,N_20712,N_21373);
nor U25616 (N_25616,N_23343,N_21808);
nor U25617 (N_25617,N_24928,N_24665);
nor U25618 (N_25618,N_24825,N_20977);
or U25619 (N_25619,N_20629,N_24566);
and U25620 (N_25620,N_23102,N_20328);
nor U25621 (N_25621,N_20392,N_22485);
or U25622 (N_25622,N_23347,N_21559);
nand U25623 (N_25623,N_24801,N_24959);
nand U25624 (N_25624,N_20558,N_21691);
and U25625 (N_25625,N_20819,N_23531);
nand U25626 (N_25626,N_23630,N_20004);
xor U25627 (N_25627,N_20138,N_20329);
nand U25628 (N_25628,N_20604,N_22317);
and U25629 (N_25629,N_23101,N_21329);
xor U25630 (N_25630,N_21290,N_24171);
nand U25631 (N_25631,N_24603,N_22799);
or U25632 (N_25632,N_20227,N_24724);
or U25633 (N_25633,N_22302,N_24952);
or U25634 (N_25634,N_21338,N_23791);
nand U25635 (N_25635,N_22218,N_21863);
and U25636 (N_25636,N_23091,N_22893);
xor U25637 (N_25637,N_24134,N_22947);
xnor U25638 (N_25638,N_22654,N_21502);
nor U25639 (N_25639,N_20072,N_23892);
or U25640 (N_25640,N_20639,N_20388);
or U25641 (N_25641,N_22328,N_23544);
xor U25642 (N_25642,N_21081,N_21726);
and U25643 (N_25643,N_23817,N_24352);
and U25644 (N_25644,N_22441,N_21421);
nor U25645 (N_25645,N_20771,N_20831);
nor U25646 (N_25646,N_22174,N_22964);
or U25647 (N_25647,N_22165,N_24664);
xnor U25648 (N_25648,N_22676,N_20710);
or U25649 (N_25649,N_21433,N_20167);
or U25650 (N_25650,N_22953,N_20749);
xnor U25651 (N_25651,N_21395,N_22241);
and U25652 (N_25652,N_24900,N_23746);
xnor U25653 (N_25653,N_23865,N_24232);
xor U25654 (N_25654,N_20232,N_21023);
nand U25655 (N_25655,N_21537,N_20331);
nand U25656 (N_25656,N_21292,N_20022);
or U25657 (N_25657,N_21936,N_22369);
nand U25658 (N_25658,N_20471,N_20857);
nor U25659 (N_25659,N_23308,N_22536);
xnor U25660 (N_25660,N_22966,N_20792);
nand U25661 (N_25661,N_23958,N_21618);
or U25662 (N_25662,N_24976,N_21773);
xnor U25663 (N_25663,N_24109,N_24829);
or U25664 (N_25664,N_23260,N_22508);
xnor U25665 (N_25665,N_24293,N_23549);
or U25666 (N_25666,N_23700,N_22124);
or U25667 (N_25667,N_24260,N_21688);
xnor U25668 (N_25668,N_23060,N_24062);
nand U25669 (N_25669,N_24016,N_20920);
or U25670 (N_25670,N_20018,N_23495);
nand U25671 (N_25671,N_22107,N_20269);
and U25672 (N_25672,N_24916,N_23624);
and U25673 (N_25673,N_24968,N_22262);
or U25674 (N_25674,N_21550,N_21221);
nand U25675 (N_25675,N_21560,N_21597);
and U25676 (N_25676,N_23145,N_22897);
or U25677 (N_25677,N_23346,N_22725);
or U25678 (N_25678,N_20495,N_22929);
nor U25679 (N_25679,N_20441,N_24301);
xor U25680 (N_25680,N_23638,N_20126);
and U25681 (N_25681,N_24386,N_24725);
nand U25682 (N_25682,N_24213,N_22108);
or U25683 (N_25683,N_20536,N_21967);
or U25684 (N_25684,N_23279,N_24174);
xnor U25685 (N_25685,N_22847,N_21682);
nand U25686 (N_25686,N_21590,N_23392);
nor U25687 (N_25687,N_21124,N_23798);
xnor U25688 (N_25688,N_21186,N_22346);
nor U25689 (N_25689,N_21076,N_23103);
nor U25690 (N_25690,N_21674,N_24082);
or U25691 (N_25691,N_23255,N_21092);
nand U25692 (N_25692,N_20899,N_22209);
nor U25693 (N_25693,N_23428,N_20465);
nor U25694 (N_25694,N_22633,N_21313);
nand U25695 (N_25695,N_23807,N_22023);
and U25696 (N_25696,N_23715,N_22759);
and U25697 (N_25697,N_23160,N_23129);
nand U25698 (N_25698,N_20170,N_20210);
or U25699 (N_25699,N_23141,N_24836);
and U25700 (N_25700,N_23125,N_21247);
xor U25701 (N_25701,N_20943,N_20599);
and U25702 (N_25702,N_22918,N_22614);
nand U25703 (N_25703,N_22597,N_21586);
nand U25704 (N_25704,N_22623,N_20302);
xnor U25705 (N_25705,N_24049,N_24122);
nor U25706 (N_25706,N_20124,N_23459);
or U25707 (N_25707,N_20461,N_22257);
nand U25708 (N_25708,N_20985,N_21610);
nor U25709 (N_25709,N_24696,N_23664);
and U25710 (N_25710,N_24131,N_23427);
nor U25711 (N_25711,N_20196,N_23189);
nor U25712 (N_25712,N_23927,N_23019);
or U25713 (N_25713,N_22022,N_24563);
or U25714 (N_25714,N_22203,N_23929);
nor U25715 (N_25715,N_22098,N_21699);
xnor U25716 (N_25716,N_20479,N_21898);
or U25717 (N_25717,N_20612,N_21739);
nand U25718 (N_25718,N_20812,N_22461);
or U25719 (N_25719,N_23941,N_23614);
nor U25720 (N_25720,N_24922,N_20800);
nor U25721 (N_25721,N_21908,N_23095);
and U25722 (N_25722,N_21813,N_21020);
nor U25723 (N_25723,N_22199,N_23768);
nor U25724 (N_25724,N_23479,N_22306);
nor U25725 (N_25725,N_21902,N_23672);
xnor U25726 (N_25726,N_23598,N_21119);
or U25727 (N_25727,N_22215,N_20277);
nor U25728 (N_25728,N_22119,N_24835);
xor U25729 (N_25729,N_22048,N_23755);
nor U25730 (N_25730,N_20549,N_20382);
and U25731 (N_25731,N_23829,N_21893);
nand U25732 (N_25732,N_23305,N_20249);
nor U25733 (N_25733,N_21861,N_22590);
or U25734 (N_25734,N_20193,N_22816);
and U25735 (N_25735,N_20993,N_24524);
nand U25736 (N_25736,N_21777,N_21652);
nor U25737 (N_25737,N_20225,N_20451);
and U25738 (N_25738,N_22870,N_24056);
and U25739 (N_25739,N_20737,N_20945);
and U25740 (N_25740,N_20283,N_20025);
and U25741 (N_25741,N_20687,N_20991);
nand U25742 (N_25742,N_24962,N_20326);
or U25743 (N_25743,N_22504,N_21125);
nand U25744 (N_25744,N_23197,N_21793);
or U25745 (N_25745,N_22138,N_22201);
nor U25746 (N_25746,N_23123,N_22111);
or U25747 (N_25747,N_23874,N_21592);
xor U25748 (N_25748,N_23662,N_23667);
and U25749 (N_25749,N_22383,N_24587);
nand U25750 (N_25750,N_22353,N_23319);
nor U25751 (N_25751,N_24921,N_21390);
nor U25752 (N_25752,N_23602,N_24483);
and U25753 (N_25753,N_23130,N_22589);
nor U25754 (N_25754,N_24741,N_22049);
nor U25755 (N_25755,N_24961,N_22443);
nor U25756 (N_25756,N_20596,N_24346);
nand U25757 (N_25757,N_23020,N_22704);
and U25758 (N_25758,N_21631,N_24970);
nor U25759 (N_25759,N_21045,N_21491);
and U25760 (N_25760,N_20801,N_21961);
and U25761 (N_25761,N_23780,N_21299);
nor U25762 (N_25762,N_22270,N_22254);
xnor U25763 (N_25763,N_23632,N_22193);
nor U25764 (N_25764,N_23313,N_20803);
or U25765 (N_25765,N_20001,N_24348);
or U25766 (N_25766,N_20104,N_21174);
nand U25767 (N_25767,N_24112,N_23434);
nand U25768 (N_25768,N_21465,N_23541);
nor U25769 (N_25769,N_20174,N_23666);
xor U25770 (N_25770,N_23816,N_22043);
nor U25771 (N_25771,N_23334,N_24544);
nor U25772 (N_25772,N_21608,N_23788);
nand U25773 (N_25773,N_23230,N_23750);
and U25774 (N_25774,N_22147,N_24811);
and U25775 (N_25775,N_20383,N_21872);
and U25776 (N_25776,N_24107,N_21331);
nor U25777 (N_25777,N_23745,N_22835);
or U25778 (N_25778,N_20845,N_23683);
and U25779 (N_25779,N_24453,N_22320);
nor U25780 (N_25780,N_22421,N_20313);
nand U25781 (N_25781,N_24616,N_22993);
or U25782 (N_25782,N_24758,N_24091);
xnor U25783 (N_25783,N_23705,N_21457);
and U25784 (N_25784,N_23767,N_23437);
xnor U25785 (N_25785,N_23340,N_22318);
xor U25786 (N_25786,N_20355,N_21066);
nor U25787 (N_25787,N_22923,N_20895);
or U25788 (N_25788,N_20047,N_22503);
and U25789 (N_25789,N_24070,N_22509);
or U25790 (N_25790,N_22176,N_20095);
or U25791 (N_25791,N_24380,N_20730);
or U25792 (N_25792,N_24858,N_20790);
and U25793 (N_25793,N_24920,N_23513);
nor U25794 (N_25794,N_23376,N_23592);
xnor U25795 (N_25795,N_24607,N_23873);
nor U25796 (N_25796,N_23036,N_24838);
nor U25797 (N_25797,N_24649,N_21147);
nor U25798 (N_25798,N_20888,N_20962);
or U25799 (N_25799,N_21497,N_24497);
or U25800 (N_25800,N_22915,N_22650);
or U25801 (N_25801,N_21925,N_21686);
and U25802 (N_25802,N_23287,N_20638);
nand U25803 (N_25803,N_21238,N_23744);
nor U25804 (N_25804,N_21460,N_22087);
nor U25805 (N_25805,N_20380,N_23451);
nor U25806 (N_25806,N_23533,N_20019);
nor U25807 (N_25807,N_20722,N_21424);
xor U25808 (N_25808,N_21459,N_24642);
and U25809 (N_25809,N_20644,N_24785);
xnor U25810 (N_25810,N_20289,N_24733);
and U25811 (N_25811,N_24748,N_23827);
nor U25812 (N_25812,N_20791,N_23696);
or U25813 (N_25813,N_21918,N_22019);
or U25814 (N_25814,N_24068,N_21359);
nor U25815 (N_25815,N_23685,N_20965);
xor U25816 (N_25816,N_23284,N_20381);
or U25817 (N_25817,N_24367,N_24100);
xnor U25818 (N_25818,N_20924,N_20874);
nor U25819 (N_25819,N_23364,N_22247);
nand U25820 (N_25820,N_20727,N_24102);
nor U25821 (N_25821,N_24846,N_24199);
nor U25822 (N_25822,N_24914,N_20751);
nor U25823 (N_25823,N_22313,N_20523);
nand U25824 (N_25824,N_21342,N_23431);
nor U25825 (N_25825,N_20351,N_21322);
or U25826 (N_25826,N_21603,N_21328);
nand U25827 (N_25827,N_20405,N_23028);
and U25828 (N_25828,N_20255,N_24893);
nor U25829 (N_25829,N_22256,N_21128);
nand U25830 (N_25830,N_22820,N_22796);
or U25831 (N_25831,N_22627,N_21198);
or U25832 (N_25832,N_21611,N_24933);
nor U25833 (N_25833,N_23534,N_22883);
nor U25834 (N_25834,N_24639,N_21129);
xor U25835 (N_25835,N_24223,N_24400);
or U25836 (N_25836,N_23826,N_23966);
xnor U25837 (N_25837,N_20794,N_20606);
xor U25838 (N_25838,N_21293,N_23658);
nand U25839 (N_25839,N_20356,N_24013);
or U25840 (N_25840,N_21796,N_22280);
nor U25841 (N_25841,N_23840,N_23729);
xnor U25842 (N_25842,N_23934,N_24901);
and U25843 (N_25843,N_20917,N_22846);
or U25844 (N_25844,N_22153,N_21141);
nor U25845 (N_25845,N_22596,N_23245);
or U25846 (N_25846,N_24279,N_20378);
and U25847 (N_25847,N_24410,N_24686);
nor U25848 (N_25848,N_23218,N_21452);
and U25849 (N_25849,N_20642,N_24558);
and U25850 (N_25850,N_22311,N_23954);
nand U25851 (N_25851,N_20024,N_22767);
xnor U25852 (N_25852,N_21884,N_20760);
or U25853 (N_25853,N_20863,N_24869);
nor U25854 (N_25854,N_24358,N_21648);
nand U25855 (N_25855,N_22756,N_22260);
nor U25856 (N_25856,N_24701,N_22576);
or U25857 (N_25857,N_22008,N_24522);
xor U25858 (N_25858,N_22178,N_20598);
xor U25859 (N_25859,N_22002,N_24687);
xnor U25860 (N_25860,N_21964,N_22734);
nor U25861 (N_25861,N_20490,N_24875);
nand U25862 (N_25862,N_20772,N_23368);
xnor U25863 (N_25863,N_21159,N_23249);
and U25864 (N_25864,N_21569,N_22425);
and U25865 (N_25865,N_24030,N_22608);
and U25866 (N_25866,N_22882,N_20582);
xnor U25867 (N_25867,N_23316,N_24944);
nor U25868 (N_25868,N_20211,N_22300);
and U25869 (N_25869,N_22565,N_21755);
or U25870 (N_25870,N_23711,N_22637);
xnor U25871 (N_25871,N_23507,N_20955);
xor U25872 (N_25872,N_24800,N_21807);
nand U25873 (N_25873,N_24597,N_20957);
and U25874 (N_25874,N_22776,N_20922);
nand U25875 (N_25875,N_20763,N_24840);
nor U25876 (N_25876,N_24532,N_23953);
or U25877 (N_25877,N_22543,N_24265);
and U25878 (N_25878,N_21103,N_21656);
or U25879 (N_25879,N_21232,N_22690);
and U25880 (N_25880,N_24363,N_23497);
or U25881 (N_25881,N_23252,N_22815);
nor U25882 (N_25882,N_23764,N_21649);
nor U25883 (N_25883,N_24460,N_21547);
nor U25884 (N_25884,N_21852,N_23742);
nand U25885 (N_25885,N_24689,N_21365);
nor U25886 (N_25886,N_23474,N_24111);
nor U25887 (N_25887,N_23246,N_21765);
nand U25888 (N_25888,N_24780,N_23655);
xor U25889 (N_25889,N_21779,N_20705);
nor U25890 (N_25890,N_23628,N_23469);
nor U25891 (N_25891,N_21732,N_22484);
or U25892 (N_25892,N_23881,N_23475);
nor U25893 (N_25893,N_22243,N_22006);
xor U25894 (N_25894,N_21983,N_22805);
or U25895 (N_25895,N_23546,N_23381);
or U25896 (N_25896,N_21239,N_22656);
nor U25897 (N_25897,N_22058,N_22370);
and U25898 (N_25898,N_22442,N_21000);
or U25899 (N_25899,N_23782,N_21404);
xor U25900 (N_25900,N_23818,N_24087);
nor U25901 (N_25901,N_21598,N_23402);
or U25902 (N_25902,N_22523,N_23556);
and U25903 (N_25903,N_24403,N_21349);
nand U25904 (N_25904,N_21402,N_21156);
and U25905 (N_25905,N_22339,N_20731);
or U25906 (N_25906,N_23820,N_24789);
nand U25907 (N_25907,N_20921,N_24120);
or U25908 (N_25908,N_23395,N_21520);
nor U25909 (N_25909,N_24073,N_23195);
or U25910 (N_25910,N_21468,N_24817);
or U25911 (N_25911,N_22708,N_24653);
and U25912 (N_25912,N_24667,N_21347);
nand U25913 (N_25913,N_24569,N_20898);
and U25914 (N_25914,N_20467,N_24812);
and U25915 (N_25915,N_20188,N_21327);
and U25916 (N_25916,N_23736,N_22459);
nand U25917 (N_25917,N_20697,N_22729);
or U25918 (N_25918,N_20061,N_21975);
and U25919 (N_25919,N_23505,N_23199);
and U25920 (N_25920,N_20890,N_23370);
or U25921 (N_25921,N_21960,N_22645);
nand U25922 (N_25922,N_22334,N_20542);
nor U25923 (N_25923,N_23899,N_20828);
and U25924 (N_25924,N_23473,N_23812);
and U25925 (N_25925,N_22293,N_21420);
nor U25926 (N_25926,N_22092,N_24531);
nor U25927 (N_25927,N_20669,N_20120);
nand U25928 (N_25928,N_23618,N_20067);
xnor U25929 (N_25929,N_23669,N_21341);
nor U25930 (N_25930,N_22705,N_23012);
nand U25931 (N_25931,N_22884,N_23306);
or U25932 (N_25932,N_24890,N_20564);
nand U25933 (N_25933,N_21225,N_22500);
xor U25934 (N_25934,N_24892,N_24844);
nand U25935 (N_25935,N_24828,N_22077);
xnor U25936 (N_25936,N_21175,N_22229);
and U25937 (N_25937,N_20140,N_22429);
nand U25938 (N_25938,N_23389,N_22112);
or U25939 (N_25939,N_24739,N_22962);
or U25940 (N_25940,N_21240,N_20244);
xnor U25941 (N_25941,N_20632,N_22073);
nor U25942 (N_25942,N_20623,N_23708);
nor U25943 (N_25943,N_21405,N_20450);
or U25944 (N_25944,N_22368,N_22438);
nor U25945 (N_25945,N_21738,N_23926);
or U25946 (N_25946,N_24764,N_22431);
nor U25947 (N_25947,N_24093,N_24795);
and U25948 (N_25948,N_24501,N_20906);
xor U25949 (N_25949,N_24579,N_23120);
nor U25950 (N_25950,N_21945,N_22076);
nand U25951 (N_25951,N_22120,N_20307);
or U25952 (N_25952,N_21071,N_23356);
or U25953 (N_25953,N_21031,N_22771);
nand U25954 (N_25954,N_24666,N_20576);
nand U25955 (N_25955,N_21013,N_21843);
or U25956 (N_25956,N_24179,N_23814);
nand U25957 (N_25957,N_20893,N_22439);
or U25958 (N_25958,N_21846,N_20032);
or U25959 (N_25959,N_24332,N_20312);
and U25960 (N_25960,N_20003,N_23386);
or U25961 (N_25961,N_20470,N_20767);
nand U25962 (N_25962,N_23207,N_22349);
xor U25963 (N_25963,N_23328,N_22955);
or U25964 (N_25964,N_22956,N_22611);
and U25965 (N_25965,N_21234,N_21381);
nor U25966 (N_25966,N_20080,N_24856);
nand U25967 (N_25967,N_21475,N_20189);
nor U25968 (N_25968,N_22987,N_24503);
nor U25969 (N_25969,N_21834,N_21085);
or U25970 (N_25970,N_21563,N_20867);
nor U25971 (N_25971,N_20330,N_21215);
nand U25972 (N_25972,N_24394,N_23055);
nor U25973 (N_25973,N_23763,N_20323);
or U25974 (N_25974,N_21073,N_21677);
nand U25975 (N_25975,N_22501,N_23726);
or U25976 (N_25976,N_23148,N_21245);
or U25977 (N_25977,N_22730,N_24212);
and U25978 (N_25978,N_21367,N_21366);
nor U25979 (N_25979,N_22283,N_23379);
or U25980 (N_25980,N_23948,N_22544);
nand U25981 (N_25981,N_22916,N_21939);
and U25982 (N_25982,N_21172,N_20460);
nor U25983 (N_25983,N_23866,N_23923);
nor U25984 (N_25984,N_23244,N_22591);
xor U25985 (N_25985,N_22373,N_24236);
nand U25986 (N_25986,N_21380,N_24831);
and U25987 (N_25987,N_22136,N_24306);
and U25988 (N_25988,N_24142,N_21670);
and U25989 (N_25989,N_22803,N_22351);
or U25990 (N_25990,N_21798,N_23781);
nor U25991 (N_25991,N_22864,N_22532);
nor U25992 (N_25992,N_24539,N_21301);
nand U25993 (N_25993,N_22821,N_20190);
or U25994 (N_25994,N_24478,N_23671);
nand U25995 (N_25995,N_24965,N_21891);
nor U25996 (N_25996,N_20015,N_20298);
and U25997 (N_25997,N_24247,N_23317);
nand U25998 (N_25998,N_24243,N_23121);
or U25999 (N_25999,N_22502,N_23398);
or U26000 (N_26000,N_22604,N_21826);
or U26001 (N_26001,N_20026,N_23267);
or U26002 (N_26002,N_24923,N_24362);
xnor U26003 (N_26003,N_21653,N_20107);
or U26004 (N_26004,N_22746,N_24485);
nand U26005 (N_26005,N_24416,N_21393);
nor U26006 (N_26006,N_22359,N_22009);
and U26007 (N_26007,N_20520,N_21885);
xor U26008 (N_26008,N_23035,N_21480);
xnor U26009 (N_26009,N_24623,N_20952);
and U26010 (N_26010,N_24671,N_21561);
and U26011 (N_26011,N_24291,N_20657);
and U26012 (N_26012,N_21006,N_21472);
nor U26013 (N_26013,N_24392,N_21763);
and U26014 (N_26014,N_22096,N_20413);
or U26015 (N_26015,N_20497,N_22850);
nand U26016 (N_26016,N_23564,N_21715);
and U26017 (N_26017,N_22363,N_23476);
or U26018 (N_26018,N_21873,N_22482);
or U26019 (N_26019,N_21003,N_23694);
and U26020 (N_26020,N_24296,N_24550);
or U26021 (N_26021,N_24678,N_23418);
xor U26022 (N_26022,N_21977,N_21705);
nand U26023 (N_26023,N_21052,N_23374);
nor U26024 (N_26024,N_24110,N_23079);
xnor U26025 (N_26025,N_24618,N_20637);
or U26026 (N_26026,N_24964,N_22169);
or U26027 (N_26027,N_23590,N_21804);
nor U26028 (N_26028,N_24584,N_20122);
nor U26029 (N_26029,N_20774,N_24172);
xnor U26030 (N_26030,N_22653,N_24775);
and U26031 (N_26031,N_22933,N_23295);
and U26032 (N_26032,N_24590,N_21882);
nand U26033 (N_26033,N_24981,N_20416);
nor U26034 (N_26034,N_21166,N_23149);
nor U26035 (N_26035,N_24099,N_23223);
nor U26036 (N_26036,N_21241,N_20458);
xnor U26037 (N_26037,N_22628,N_23593);
nor U26038 (N_26038,N_24067,N_21086);
and U26039 (N_26039,N_24543,N_24437);
and U26040 (N_26040,N_22554,N_20590);
or U26041 (N_26041,N_21923,N_24207);
nand U26042 (N_26042,N_20944,N_24145);
nand U26043 (N_26043,N_20570,N_21284);
xnor U26044 (N_26044,N_23653,N_23991);
nand U26045 (N_26045,N_20278,N_24876);
or U26046 (N_26046,N_22684,N_23997);
or U26047 (N_26047,N_23178,N_23274);
nor U26048 (N_26048,N_23294,N_22516);
or U26049 (N_26049,N_24299,N_23224);
and U26050 (N_26050,N_24343,N_24963);
or U26051 (N_26051,N_22594,N_22242);
nor U26052 (N_26052,N_21488,N_20518);
nor U26053 (N_26053,N_20785,N_24634);
nand U26054 (N_26054,N_24598,N_24231);
or U26055 (N_26055,N_20377,N_24771);
or U26056 (N_26056,N_22736,N_22855);
and U26057 (N_26057,N_23893,N_23433);
and U26058 (N_26058,N_21698,N_23070);
nor U26059 (N_26059,N_24031,N_21094);
and U26060 (N_26060,N_21426,N_21671);
nor U26061 (N_26061,N_24814,N_24303);
nor U26062 (N_26062,N_24578,N_21766);
nor U26063 (N_26063,N_24619,N_22115);
nor U26064 (N_26064,N_22323,N_23001);
or U26065 (N_26065,N_20477,N_20139);
xnor U26066 (N_26066,N_24449,N_21972);
nor U26067 (N_26067,N_20125,N_23478);
nand U26068 (N_26068,N_24727,N_21026);
and U26069 (N_26069,N_22059,N_24613);
nor U26070 (N_26070,N_23536,N_23841);
nand U26071 (N_26071,N_21212,N_24681);
nor U26072 (N_26072,N_22636,N_20938);
nand U26073 (N_26073,N_22902,N_24704);
and U26074 (N_26074,N_20971,N_21943);
nor U26075 (N_26075,N_21242,N_23212);
nand U26076 (N_26076,N_22062,N_22935);
and U26077 (N_26077,N_22428,N_20756);
or U26078 (N_26078,N_23909,N_23813);
nor U26079 (N_26079,N_20939,N_20357);
and U26080 (N_26080,N_21593,N_24723);
or U26081 (N_26081,N_23661,N_21321);
nand U26082 (N_26082,N_23310,N_21683);
nor U26083 (N_26083,N_22991,N_24966);
and U26084 (N_26084,N_21702,N_20295);
nor U26085 (N_26085,N_21205,N_23106);
or U26086 (N_26086,N_22231,N_24728);
and U26087 (N_26087,N_23206,N_21929);
nand U26088 (N_26088,N_22468,N_22234);
nor U26089 (N_26089,N_23850,N_24589);
nor U26090 (N_26090,N_23289,N_24488);
or U26091 (N_26091,N_24036,N_24458);
xor U26092 (N_26092,N_22946,N_20538);
nand U26093 (N_26093,N_20723,N_20996);
nor U26094 (N_26094,N_23227,N_20186);
or U26095 (N_26095,N_20113,N_20894);
nand U26096 (N_26096,N_21493,N_24284);
or U26097 (N_26097,N_23539,N_22848);
xor U26098 (N_26098,N_22526,N_23663);
and U26099 (N_26099,N_21785,N_23110);
nor U26100 (N_26100,N_23933,N_21001);
nand U26101 (N_26101,N_20856,N_24106);
and U26102 (N_26102,N_23969,N_24322);
and U26103 (N_26103,N_21140,N_24397);
nor U26104 (N_26104,N_21168,N_24428);
and U26105 (N_26105,N_20237,N_20625);
and U26106 (N_26106,N_23916,N_24424);
nor U26107 (N_26107,N_20308,N_21669);
or U26108 (N_26108,N_21298,N_20788);
nand U26109 (N_26109,N_20960,N_21089);
and U26110 (N_26110,N_20005,N_24517);
xnor U26111 (N_26111,N_23728,N_21791);
xnor U26112 (N_26112,N_20533,N_24121);
nand U26113 (N_26113,N_21708,N_20420);
and U26114 (N_26114,N_20583,N_24769);
or U26115 (N_26115,N_21267,N_23822);
or U26116 (N_26116,N_21970,N_24581);
nor U26117 (N_26117,N_23872,N_22717);
nor U26118 (N_26118,N_24494,N_21543);
and U26119 (N_26119,N_22783,N_21077);
or U26120 (N_26120,N_24887,N_20363);
or U26121 (N_26121,N_23023,N_22130);
nand U26122 (N_26122,N_22312,N_22114);
nor U26123 (N_26123,N_21043,N_24273);
and U26124 (N_26124,N_22814,N_23568);
nand U26125 (N_26125,N_20028,N_21214);
or U26126 (N_26126,N_23540,N_20172);
xor U26127 (N_26127,N_24160,N_21004);
xnor U26128 (N_26128,N_23127,N_20636);
and U26129 (N_26129,N_22553,N_21104);
or U26130 (N_26130,N_24203,N_20483);
and U26131 (N_26131,N_22586,N_22703);
nand U26132 (N_26132,N_21333,N_23172);
nand U26133 (N_26133,N_21049,N_20060);
or U26134 (N_26134,N_21694,N_22948);
or U26135 (N_26135,N_22253,N_20742);
xor U26136 (N_26136,N_20833,N_22593);
or U26137 (N_26137,N_24077,N_20293);
nor U26138 (N_26138,N_20466,N_20482);
nand U26139 (N_26139,N_22099,N_21651);
xor U26140 (N_26140,N_20304,N_21106);
nand U26141 (N_26141,N_21330,N_22549);
nor U26142 (N_26142,N_21887,N_23801);
nand U26143 (N_26143,N_23737,N_24773);
or U26144 (N_26144,N_23612,N_24064);
or U26145 (N_26145,N_23131,N_24327);
and U26146 (N_26146,N_21864,N_20152);
or U26147 (N_26147,N_24595,N_24039);
or U26148 (N_26148,N_23776,N_22269);
nor U26149 (N_26149,N_23819,N_21992);
nand U26150 (N_26150,N_21017,N_20218);
and U26151 (N_26151,N_23514,N_21658);
or U26152 (N_26152,N_22890,N_23117);
nand U26153 (N_26153,N_24435,N_24180);
nor U26154 (N_26154,N_23174,N_22931);
and U26155 (N_26155,N_22506,N_21552);
nand U26156 (N_26156,N_20611,N_21870);
xnor U26157 (N_26157,N_21888,N_23471);
and U26158 (N_26158,N_23229,N_20510);
and U26159 (N_26159,N_20695,N_21180);
nand U26160 (N_26160,N_24377,N_22362);
or U26161 (N_26161,N_21901,N_21312);
or U26162 (N_26162,N_21087,N_21427);
and U26163 (N_26163,N_23631,N_24596);
and U26164 (N_26164,N_20765,N_21622);
or U26165 (N_26165,N_24209,N_20979);
nor U26166 (N_26166,N_20325,N_21111);
or U26167 (N_26167,N_21064,N_22582);
xor U26168 (N_26168,N_23580,N_21318);
or U26169 (N_26169,N_21630,N_23484);
nand U26170 (N_26170,N_23901,N_23794);
or U26171 (N_26171,N_21832,N_20811);
or U26172 (N_26172,N_23623,N_24430);
nand U26173 (N_26173,N_20212,N_24280);
or U26174 (N_26174,N_21620,N_24580);
nor U26175 (N_26175,N_23506,N_24908);
and U26176 (N_26176,N_23660,N_24625);
and U26177 (N_26177,N_20353,N_22005);
and U26178 (N_26178,N_20456,N_22330);
or U26179 (N_26179,N_21524,N_24926);
or U26180 (N_26180,N_21659,N_24594);
and U26181 (N_26181,N_21582,N_20581);
or U26182 (N_26182,N_22055,N_24471);
or U26183 (N_26183,N_22211,N_24330);
nand U26184 (N_26184,N_23520,N_24133);
nor U26185 (N_26185,N_24983,N_21233);
nor U26186 (N_26186,N_24010,N_20281);
nor U26187 (N_26187,N_23851,N_20049);
nor U26188 (N_26188,N_22969,N_20068);
nand U26189 (N_26189,N_21314,N_24820);
and U26190 (N_26190,N_22754,N_22609);
nand U26191 (N_26191,N_24177,N_24224);
and U26192 (N_26192,N_21736,N_22938);
nor U26193 (N_26193,N_23613,N_20780);
nor U26194 (N_26194,N_23179,N_23562);
and U26195 (N_26195,N_21619,N_21810);
nor U26196 (N_26196,N_22535,N_21815);
xnor U26197 (N_26197,N_23984,N_21522);
nand U26198 (N_26198,N_20053,N_20436);
nor U26199 (N_26199,N_20620,N_23802);
nand U26200 (N_26200,N_22298,N_23942);
nor U26201 (N_26201,N_20793,N_22451);
xor U26202 (N_26202,N_20795,N_20361);
and U26203 (N_26203,N_22054,N_24593);
xor U26204 (N_26204,N_24652,N_21022);
nor U26205 (N_26205,N_24744,N_23241);
and U26206 (N_26206,N_22723,N_21530);
nand U26207 (N_26207,N_23935,N_22768);
and U26208 (N_26208,N_24015,N_23271);
and U26209 (N_26209,N_24553,N_24984);
or U26210 (N_26210,N_24951,N_24661);
or U26211 (N_26211,N_23140,N_24218);
nor U26212 (N_26212,N_21678,N_23054);
or U26213 (N_26213,N_24899,N_24536);
nor U26214 (N_26214,N_21673,N_20371);
nor U26215 (N_26215,N_21399,N_20896);
nor U26216 (N_26216,N_24684,N_20852);
nor U26217 (N_26217,N_22585,N_21311);
or U26218 (N_26218,N_23187,N_24978);
nand U26219 (N_26219,N_20150,N_23073);
and U26220 (N_26220,N_20618,N_22906);
nand U26221 (N_26221,N_21675,N_21251);
nand U26222 (N_26222,N_21578,N_23169);
or U26223 (N_26223,N_23578,N_23021);
xor U26224 (N_26224,N_24037,N_21772);
xor U26225 (N_26225,N_24190,N_21362);
nor U26226 (N_26226,N_20989,N_24525);
or U26227 (N_26227,N_24510,N_20119);
xor U26228 (N_26228,N_22760,N_24393);
or U26229 (N_26229,N_24173,N_24385);
or U26230 (N_26230,N_23466,N_22785);
and U26231 (N_26231,N_22264,N_24507);
nand U26232 (N_26232,N_23635,N_20228);
and U26233 (N_26233,N_24088,N_22464);
or U26234 (N_26234,N_22545,N_21246);
or U26235 (N_26235,N_24401,N_22949);
or U26236 (N_26236,N_23806,N_22237);
and U26237 (N_26237,N_24210,N_24399);
and U26238 (N_26238,N_21394,N_21375);
nor U26239 (N_26239,N_23601,N_20655);
and U26240 (N_26240,N_20617,N_22336);
or U26241 (N_26241,N_21721,N_24611);
and U26242 (N_26242,N_22610,N_21474);
nor U26243 (N_26243,N_21642,N_24975);
nand U26244 (N_26244,N_21494,N_23825);
or U26245 (N_26245,N_24557,N_23485);
xnor U26246 (N_26246,N_24229,N_20242);
or U26247 (N_26247,N_24309,N_20953);
and U26248 (N_26248,N_20310,N_23693);
or U26249 (N_26249,N_20679,N_24953);
nor U26250 (N_26250,N_20709,N_22322);
nor U26251 (N_26251,N_21795,N_24853);
xnor U26252 (N_26252,N_20575,N_24709);
or U26253 (N_26253,N_24604,N_23504);
or U26254 (N_26254,N_20164,N_21216);
or U26255 (N_26255,N_23041,N_23304);
nand U26256 (N_26256,N_21197,N_24650);
or U26257 (N_26257,N_21935,N_24905);
or U26258 (N_26258,N_24535,N_21432);
nor U26259 (N_26259,N_20901,N_23447);
or U26260 (N_26260,N_23455,N_22809);
or U26261 (N_26261,N_22089,N_20488);
or U26262 (N_26262,N_20640,N_22103);
nor U26263 (N_26263,N_20769,N_20035);
nand U26264 (N_26264,N_21102,N_22577);
and U26265 (N_26265,N_23365,N_21138);
or U26266 (N_26266,N_22252,N_21171);
nor U26267 (N_26267,N_23338,N_22657);
or U26268 (N_26268,N_24381,N_23453);
nor U26269 (N_26269,N_23107,N_24137);
and U26270 (N_26270,N_22297,N_21814);
nand U26271 (N_26271,N_21515,N_23170);
nand U26272 (N_26272,N_20230,N_23446);
nor U26273 (N_26273,N_22849,N_21423);
nor U26274 (N_26274,N_20233,N_24512);
or U26275 (N_26275,N_20663,N_24753);
nor U26276 (N_26276,N_24690,N_24734);
nand U26277 (N_26277,N_21444,N_21934);
nand U26278 (N_26278,N_24894,N_21230);
nand U26279 (N_26279,N_23834,N_22873);
nand U26280 (N_26280,N_22678,N_23976);
and U26281 (N_26281,N_23962,N_23738);
and U26282 (N_26282,N_20935,N_22530);
xnor U26283 (N_26283,N_23486,N_21185);
xor U26284 (N_26284,N_22646,N_24292);
or U26285 (N_26285,N_23436,N_20614);
or U26286 (N_26286,N_23085,N_20499);
or U26287 (N_26287,N_23870,N_21021);
nand U26288 (N_26288,N_24477,N_23114);
or U26289 (N_26289,N_24076,N_20173);
or U26290 (N_26290,N_24565,N_23261);
xor U26291 (N_26291,N_24994,N_24055);
xor U26292 (N_26292,N_23998,N_20660);
nor U26293 (N_26293,N_21131,N_21903);
and U26294 (N_26294,N_21306,N_23220);
nand U26295 (N_26295,N_20569,N_20285);
nor U26296 (N_26296,N_20587,N_24463);
nand U26297 (N_26297,N_23719,N_22122);
and U26298 (N_26298,N_21170,N_24702);
nand U26299 (N_26299,N_23457,N_23947);
nor U26300 (N_26300,N_24713,N_20729);
nand U26301 (N_26301,N_21505,N_20716);
or U26302 (N_26302,N_24645,N_24841);
nand U26303 (N_26303,N_20473,N_21120);
and U26304 (N_26304,N_24662,N_23842);
nor U26305 (N_26305,N_20251,N_23450);
or U26306 (N_26306,N_23657,N_21984);
nor U26307 (N_26307,N_24822,N_24349);
xor U26308 (N_26308,N_23911,N_23248);
xnor U26309 (N_26309,N_24176,N_21255);
and U26310 (N_26310,N_22845,N_22394);
nand U26311 (N_26311,N_20217,N_23845);
xor U26312 (N_26312,N_22137,N_22093);
nand U26313 (N_26313,N_24440,N_21074);
and U26314 (N_26314,N_21352,N_20528);
nand U26315 (N_26315,N_21759,N_20146);
xor U26316 (N_26316,N_22568,N_20098);
and U26317 (N_26317,N_20358,N_21701);
nor U26318 (N_26318,N_20448,N_23465);
nor U26319 (N_26319,N_22641,N_22838);
nor U26320 (N_26320,N_20127,N_21163);
nand U26321 (N_26321,N_21320,N_22314);
nor U26322 (N_26322,N_20073,N_20048);
nor U26323 (N_26323,N_20967,N_21827);
xnor U26324 (N_26324,N_24371,N_21360);
nand U26325 (N_26325,N_20444,N_20696);
nor U26326 (N_26326,N_20547,N_20385);
nand U26327 (N_26327,N_24295,N_24794);
nor U26328 (N_26328,N_20565,N_22872);
or U26329 (N_26329,N_24159,N_20559);
or U26330 (N_26330,N_21952,N_22764);
or U26331 (N_26331,N_23062,N_23077);
or U26332 (N_26332,N_23275,N_20861);
or U26333 (N_26333,N_21962,N_23057);
and U26334 (N_26334,N_22837,N_22279);
and U26335 (N_26335,N_23682,N_24422);
or U26336 (N_26336,N_20484,N_21326);
nor U26337 (N_26337,N_21032,N_23990);
xnor U26338 (N_26338,N_20805,N_20561);
or U26339 (N_26339,N_23766,N_24763);
nor U26340 (N_26340,N_24054,N_23754);
xnor U26341 (N_26341,N_24651,N_21735);
or U26342 (N_26342,N_23243,N_23312);
and U26343 (N_26343,N_21830,N_22379);
and U26344 (N_26344,N_20245,N_23897);
or U26345 (N_26345,N_23824,N_22853);
nor U26346 (N_26346,N_21155,N_20912);
or U26347 (N_26347,N_21466,N_24187);
nor U26348 (N_26348,N_22224,N_23133);
and U26349 (N_26349,N_20552,N_24561);
nand U26350 (N_26350,N_20907,N_22141);
xnor U26351 (N_26351,N_24439,N_21549);
and U26352 (N_26352,N_23771,N_24796);
and U26353 (N_26353,N_20439,N_24799);
nor U26354 (N_26354,N_23254,N_20215);
or U26355 (N_26355,N_23898,N_24126);
nor U26356 (N_26356,N_22088,N_21875);
nand U26357 (N_26357,N_20600,N_23143);
or U26358 (N_26358,N_22276,N_23978);
nand U26359 (N_26359,N_20699,N_23239);
nor U26360 (N_26360,N_24340,N_21231);
nor U26361 (N_26361,N_22963,N_22958);
or U26362 (N_26362,N_24182,N_21441);
or U26363 (N_26363,N_23910,N_20515);
or U26364 (N_26364,N_22706,N_20808);
xnor U26365 (N_26365,N_23981,N_22788);
and U26366 (N_26366,N_23576,N_22894);
nor U26367 (N_26367,N_24395,N_20948);
nand U26368 (N_26368,N_24747,N_24336);
xnor U26369 (N_26369,N_23293,N_22629);
and U26370 (N_26370,N_20880,N_22460);
nand U26371 (N_26371,N_22831,N_20891);
and U26372 (N_26372,N_20980,N_20478);
and U26373 (N_26373,N_24699,N_24376);
or U26374 (N_26374,N_22640,N_20703);
or U26375 (N_26375,N_23579,N_22551);
nand U26376 (N_26376,N_23385,N_21809);
nor U26377 (N_26377,N_22372,N_24233);
or U26378 (N_26378,N_24345,N_23880);
or U26379 (N_26379,N_20319,N_20100);
or U26380 (N_26380,N_24490,N_23836);
and U26381 (N_26381,N_21417,N_24143);
nand U26382 (N_26382,N_23770,N_22714);
nand U26383 (N_26383,N_20810,N_24454);
and U26384 (N_26384,N_24046,N_23508);
nand U26385 (N_26385,N_20650,N_21287);
xor U26386 (N_26386,N_23828,N_21692);
nor U26387 (N_26387,N_21946,N_22928);
nor U26388 (N_26388,N_20915,N_24847);
and U26389 (N_26389,N_24300,N_21968);
nor U26390 (N_26390,N_23341,N_22097);
or U26391 (N_26391,N_23634,N_20747);
nor U26392 (N_26392,N_24075,N_22507);
nor U26393 (N_26393,N_22885,N_22481);
or U26394 (N_26394,N_21289,N_20151);
and U26395 (N_26395,N_24206,N_22569);
xor U26396 (N_26396,N_22580,N_21262);
nand U26397 (N_26397,N_22436,N_20739);
or U26398 (N_26398,N_22216,N_23215);
and U26399 (N_26399,N_23646,N_20474);
nor U26400 (N_26400,N_20872,N_21595);
xnor U26401 (N_26401,N_20903,N_22998);
or U26402 (N_26402,N_21142,N_21069);
nand U26403 (N_26403,N_20670,N_24168);
and U26404 (N_26404,N_23420,N_22877);
xor U26405 (N_26405,N_22794,N_24716);
or U26406 (N_26406,N_20578,N_24691);
nor U26407 (N_26407,N_21904,N_22852);
and U26408 (N_26408,N_23980,N_22649);
nand U26409 (N_26409,N_24711,N_21109);
nor U26410 (N_26410,N_22267,N_23461);
or U26411 (N_26411,N_22402,N_22603);
and U26412 (N_26412,N_23411,N_23311);
nand U26413 (N_26413,N_22294,N_23773);
or U26414 (N_26414,N_24314,N_23318);
or U26415 (N_26415,N_24572,N_21865);
nand U26416 (N_26416,N_24810,N_24935);
xor U26417 (N_26417,N_21461,N_22688);
and U26418 (N_26418,N_24802,N_23382);
and U26419 (N_26419,N_23859,N_23235);
nand U26420 (N_26420,N_23903,N_24546);
nand U26421 (N_26421,N_22116,N_23524);
nor U26422 (N_26422,N_21525,N_24185);
or U26423 (N_26423,N_21361,N_20165);
nor U26424 (N_26424,N_21574,N_21358);
and U26425 (N_26425,N_20209,N_21575);
or U26426 (N_26426,N_23727,N_21437);
nor U26427 (N_26427,N_21193,N_24941);
and U26428 (N_26428,N_23681,N_24254);
nand U26429 (N_26429,N_21401,N_22740);
nand U26430 (N_26430,N_23481,N_24319);
nand U26431 (N_26431,N_22942,N_22118);
xor U26432 (N_26432,N_22382,N_23443);
nor U26433 (N_26433,N_20216,N_24184);
and U26434 (N_26434,N_23680,N_23426);
nand U26435 (N_26435,N_24672,N_24730);
or U26436 (N_26436,N_23853,N_21919);
nor U26437 (N_26437,N_23315,N_22683);
nand U26438 (N_26438,N_21473,N_23269);
and U26439 (N_26439,N_23314,N_22185);
nand U26440 (N_26440,N_20675,N_23126);
and U26441 (N_26441,N_20873,N_24511);
nand U26442 (N_26442,N_23138,N_23830);
or U26443 (N_26443,N_23887,N_21754);
or U26444 (N_26444,N_22970,N_20266);
nand U26445 (N_26445,N_20254,N_22405);
or U26446 (N_26446,N_24824,N_22031);
nor U26447 (N_26447,N_24014,N_24222);
and U26448 (N_26448,N_22748,N_24575);
nor U26449 (N_26449,N_24929,N_22658);
and U26450 (N_26450,N_20956,N_21849);
nor U26451 (N_26451,N_24573,N_22035);
xor U26452 (N_26452,N_20008,N_22830);
and U26453 (N_26453,N_24999,N_24482);
nor U26454 (N_26454,N_21542,N_24058);
or U26455 (N_26455,N_23503,N_24155);
and U26456 (N_26456,N_21695,N_20701);
or U26457 (N_26457,N_21627,N_20376);
nand U26458 (N_26458,N_23383,N_23399);
nor U26459 (N_26459,N_20627,N_21192);
nor U26460 (N_26460,N_23225,N_22371);
or U26461 (N_26461,N_20830,N_22749);
and U26462 (N_26462,N_20603,N_22061);
and U26463 (N_26463,N_21280,N_24288);
nor U26464 (N_26464,N_23752,N_23741);
or U26465 (N_26465,N_21786,N_20685);
or U26466 (N_26466,N_21737,N_20970);
nor U26467 (N_26467,N_23968,N_21199);
nor U26468 (N_26468,N_21378,N_24545);
or U26469 (N_26469,N_24496,N_20114);
or U26470 (N_26470,N_20654,N_20044);
nor U26471 (N_26471,N_23977,N_22305);
nor U26472 (N_26472,N_21154,N_23210);
nor U26473 (N_26473,N_24697,N_20400);
and U26474 (N_26474,N_22727,N_23288);
or U26475 (N_26475,N_23339,N_20205);
and U26476 (N_26476,N_24034,N_22672);
and U26477 (N_26477,N_22733,N_24582);
and U26478 (N_26478,N_21041,N_24089);
and U26479 (N_26479,N_23753,N_22989);
nor U26480 (N_26480,N_24323,N_21055);
or U26481 (N_26481,N_20649,N_24104);
nor U26482 (N_26482,N_23432,N_20231);
nand U26483 (N_26483,N_22671,N_23460);
or U26484 (N_26484,N_20681,N_21761);
or U26485 (N_26485,N_24467,N_20961);
or U26486 (N_26486,N_21958,N_24648);
or U26487 (N_26487,N_20220,N_22040);
or U26488 (N_26488,N_21149,N_24382);
or U26489 (N_26489,N_23707,N_20090);
and U26490 (N_26490,N_22149,N_22750);
nor U26491 (N_26491,N_21568,N_20234);
and U26492 (N_26492,N_20550,N_20748);
nor U26493 (N_26493,N_23161,N_24194);
or U26494 (N_26494,N_24079,N_24432);
or U26495 (N_26495,N_23684,N_21954);
nand U26496 (N_26496,N_22348,N_23535);
nand U26497 (N_26497,N_22486,N_23648);
or U26498 (N_26498,N_23482,N_22841);
nor U26499 (N_26499,N_21411,N_24806);
nand U26500 (N_26500,N_21896,N_24602);
or U26501 (N_26501,N_22162,N_21526);
nand U26502 (N_26502,N_20145,N_22910);
nor U26503 (N_26503,N_22648,N_20573);
and U26504 (N_26504,N_21805,N_21758);
nor U26505 (N_26505,N_23616,N_20171);
or U26506 (N_26506,N_20507,N_20741);
and U26507 (N_26507,N_23345,N_22025);
nor U26508 (N_26508,N_20275,N_21910);
nor U26509 (N_26509,N_24562,N_21566);
and U26510 (N_26510,N_22366,N_20969);
nand U26511 (N_26511,N_22625,N_23640);
or U26512 (N_26512,N_24834,N_23604);
nand U26513 (N_26513,N_20121,N_20252);
and U26514 (N_26514,N_22167,N_24974);
xor U26515 (N_26515,N_23331,N_24907);
and U26516 (N_26516,N_20224,N_24599);
and U26517 (N_26517,N_23543,N_20264);
and U26518 (N_26518,N_22630,N_24271);
and U26519 (N_26519,N_23586,N_22670);
or U26520 (N_26520,N_21286,N_22537);
or U26521 (N_26521,N_21133,N_21844);
and U26522 (N_26522,N_21528,N_21957);
or U26523 (N_26523,N_22798,N_20816);
and U26524 (N_26524,N_24262,N_22292);
and U26525 (N_26525,N_21148,N_24390);
nand U26526 (N_26526,N_24426,N_20431);
and U26527 (N_26527,N_22222,N_20525);
nor U26528 (N_26528,N_24862,N_20879);
or U26529 (N_26529,N_20878,N_21204);
nor U26530 (N_26530,N_23996,N_24784);
or U26531 (N_26531,N_24737,N_24170);
nor U26532 (N_26532,N_21228,N_24969);
and U26533 (N_26533,N_22396,N_23644);
nand U26534 (N_26534,N_21724,N_22567);
nand U26535 (N_26535,N_23456,N_22981);
or U26536 (N_26536,N_22004,N_23058);
xor U26537 (N_26537,N_22738,N_23277);
or U26538 (N_26538,N_21410,N_22186);
and U26539 (N_26539,N_21194,N_24000);
and U26540 (N_26540,N_24540,N_21623);
xor U26541 (N_26541,N_22829,N_21577);
and U26542 (N_26542,N_24211,N_22665);
or U26543 (N_26543,N_21033,N_24731);
nand U26544 (N_26544,N_22556,N_21388);
nor U26545 (N_26545,N_22236,N_21257);
nor U26546 (N_26546,N_22926,N_23202);
and U26547 (N_26547,N_21337,N_24629);
nor U26548 (N_26548,N_20088,N_21990);
or U26549 (N_26549,N_22117,N_21265);
nand U26550 (N_26550,N_24193,N_21899);
and U26551 (N_26551,N_22011,N_21503);
nor U26552 (N_26552,N_23645,N_23002);
or U26553 (N_26553,N_22354,N_23026);
and U26554 (N_26554,N_24251,N_22104);
nor U26555 (N_26555,N_22710,N_20494);
or U26556 (N_26556,N_21354,N_24354);
xnor U26557 (N_26557,N_21277,N_23787);
nor U26558 (N_26558,N_20524,N_23159);
or U26559 (N_26559,N_23424,N_22790);
or U26560 (N_26560,N_22726,N_24992);
and U26561 (N_26561,N_23108,N_22505);
nor U26562 (N_26562,N_21587,N_22192);
and U26563 (N_26563,N_23732,N_23488);
nand U26564 (N_26564,N_22497,N_20081);
nor U26565 (N_26565,N_23765,N_20261);
nand U26566 (N_26566,N_22643,N_23532);
and U26567 (N_26567,N_24017,N_22696);
nor U26568 (N_26568,N_21050,N_21999);
and U26569 (N_26569,N_21176,N_22488);
nor U26570 (N_26570,N_22550,N_23701);
nand U26571 (N_26571,N_22407,N_23004);
or U26572 (N_26572,N_23963,N_23740);
or U26573 (N_26573,N_24726,N_21713);
or U26574 (N_26574,N_22282,N_20063);
and U26575 (N_26575,N_24095,N_23519);
nand U26576 (N_26576,N_22531,N_22033);
and U26577 (N_26577,N_23668,N_24871);
xor U26578 (N_26578,N_21364,N_23938);
and U26579 (N_26579,N_24411,N_22205);
xor U26580 (N_26580,N_24526,N_20875);
and U26581 (N_26581,N_20621,N_21099);
or U26582 (N_26582,N_23703,N_24883);
or U26583 (N_26583,N_21351,N_23326);
nor U26584 (N_26584,N_22128,N_24125);
or U26585 (N_26585,N_21243,N_21206);
nor U26586 (N_26586,N_23649,N_24761);
or U26587 (N_26587,N_23016,N_21848);
and U26588 (N_26588,N_23629,N_21521);
and U26589 (N_26589,N_23192,N_22288);
nand U26590 (N_26590,N_23193,N_21930);
and U26591 (N_26591,N_22978,N_23567);
nor U26592 (N_26592,N_22102,N_20370);
and U26593 (N_26593,N_22003,N_20346);
or U26594 (N_26594,N_24398,N_23177);
or U26595 (N_26595,N_20038,N_24754);
nand U26596 (N_26596,N_23930,N_21710);
nor U26597 (N_26597,N_22265,N_20183);
nor U26598 (N_26598,N_22310,N_23173);
nand U26599 (N_26599,N_21591,N_23886);
and U26600 (N_26600,N_24885,N_20714);
nand U26601 (N_26601,N_22721,N_24530);
nor U26602 (N_26602,N_23718,N_23089);
nand U26603 (N_26603,N_21509,N_22711);
xor U26604 (N_26604,N_21604,N_23523);
or U26605 (N_26605,N_23518,N_20191);
nand U26606 (N_26606,N_21709,N_22150);
nand U26607 (N_26607,N_24982,N_21812);
nor U26608 (N_26608,N_20526,N_24541);
nor U26609 (N_26609,N_23268,N_21034);
or U26610 (N_26610,N_21860,N_21237);
xnor U26611 (N_26611,N_22385,N_20849);
nand U26612 (N_26612,N_21483,N_23571);
nor U26613 (N_26613,N_22965,N_21153);
nor U26614 (N_26614,N_20825,N_22333);
xnor U26615 (N_26615,N_23652,N_23757);
nor U26616 (N_26616,N_24383,N_23067);
nor U26617 (N_26617,N_20671,N_23774);
nand U26618 (N_26618,N_24622,N_21729);
nand U26619 (N_26619,N_22879,N_20175);
or U26620 (N_26620,N_24097,N_24438);
and U26621 (N_26621,N_21654,N_22168);
nor U26622 (N_26622,N_22990,N_24025);
or U26623 (N_26623,N_24290,N_24447);
and U26624 (N_26624,N_22901,N_20824);
xor U26625 (N_26625,N_20442,N_21617);
nor U26626 (N_26626,N_22106,N_20414);
or U26627 (N_26627,N_20521,N_24538);
and U26628 (N_26628,N_24646,N_22052);
and U26629 (N_26629,N_23796,N_22100);
nor U26630 (N_26630,N_23584,N_22400);
nor U26631 (N_26631,N_20631,N_20415);
nand U26632 (N_26632,N_20079,N_22971);
nand U26633 (N_26633,N_24570,N_24473);
nor U26634 (N_26634,N_23391,N_22024);
nor U26635 (N_26635,N_22631,N_20384);
or U26636 (N_26636,N_24258,N_24269);
and U26637 (N_26637,N_23104,N_23971);
nor U26638 (N_26638,N_20981,N_20608);
and U26639 (N_26639,N_23932,N_20719);
or U26640 (N_26640,N_22819,N_23994);
or U26641 (N_26641,N_20871,N_23799);
nor U26642 (N_26642,N_20844,N_20821);
nand U26643 (N_26643,N_23521,N_22584);
xor U26644 (N_26644,N_20197,N_24225);
and U26645 (N_26645,N_24777,N_22375);
or U26646 (N_26646,N_23673,N_24774);
or U26647 (N_26647,N_21190,N_23512);
and U26648 (N_26648,N_24621,N_23247);
xor U26649 (N_26649,N_23569,N_23093);
and U26650 (N_26650,N_24950,N_24676);
or U26651 (N_26651,N_22466,N_22498);
nor U26652 (N_26652,N_22655,N_20758);
nand U26653 (N_26653,N_21953,N_20421);
nand U26654 (N_26654,N_23350,N_24931);
nor U26655 (N_26655,N_23214,N_23863);
nor U26656 (N_26656,N_24368,N_21857);
or U26657 (N_26657,N_23679,N_20925);
or U26658 (N_26658,N_23688,N_20572);
and U26659 (N_26659,N_20934,N_23264);
nand U26660 (N_26660,N_22575,N_20077);
or U26661 (N_26661,N_20397,N_20270);
nor U26662 (N_26662,N_24637,N_23879);
nand U26663 (N_26663,N_22857,N_23900);
or U26664 (N_26664,N_21177,N_21626);
nand U26665 (N_26665,N_21749,N_21386);
or U26666 (N_26666,N_20837,N_22563);
nor U26667 (N_26667,N_20594,N_23105);
nor U26668 (N_26668,N_21348,N_24839);
and U26669 (N_26669,N_21226,N_22876);
or U26670 (N_26670,N_24705,N_24320);
or U26671 (N_26671,N_21596,N_24047);
nand U26672 (N_26672,N_22078,N_24311);
or U26673 (N_26673,N_22163,N_20076);
nand U26674 (N_26674,N_21208,N_22865);
xor U26675 (N_26675,N_21938,N_23751);
xor U26676 (N_26676,N_20428,N_24065);
and U26677 (N_26677,N_20963,N_24842);
and U26678 (N_26678,N_24879,N_22066);
nand U26679 (N_26679,N_23906,N_24415);
and U26680 (N_26680,N_24283,N_21624);
and U26681 (N_26681,N_20560,N_21224);
nor U26682 (N_26682,N_22959,N_23165);
and U26683 (N_26683,N_24101,N_20700);
and U26684 (N_26684,N_22719,N_20992);
and U26685 (N_26685,N_20130,N_20820);
or U26686 (N_26686,N_20693,N_23291);
nor U26687 (N_26687,N_22615,N_21127);
nor U26688 (N_26688,N_20928,N_22922);
or U26689 (N_26689,N_24516,N_21207);
and U26690 (N_26690,N_24729,N_21200);
nor U26691 (N_26691,N_23993,N_20959);
or U26692 (N_26692,N_24161,N_21942);
and U26693 (N_26693,N_24334,N_23047);
nor U26694 (N_26694,N_23458,N_20827);
nor U26695 (N_26695,N_21636,N_22386);
or U26696 (N_26696,N_20141,N_24827);
nand U26697 (N_26697,N_20607,N_21628);
nor U26698 (N_26698,N_22143,N_22716);
xor U26699 (N_26699,N_20062,N_23725);
nor U26700 (N_26700,N_24215,N_22110);
or U26701 (N_26701,N_22927,N_24523);
nand U26702 (N_26702,N_20932,N_22695);
or U26703 (N_26703,N_20362,N_23480);
nand U26704 (N_26704,N_20511,N_21028);
or U26705 (N_26705,N_22561,N_20345);
and U26706 (N_26706,N_23075,N_22578);
or U26707 (N_26707,N_23676,N_23231);
nor U26708 (N_26708,N_24529,N_22778);
or U26709 (N_26709,N_24708,N_21640);
nand U26710 (N_26710,N_21973,N_22745);
or U26711 (N_26711,N_24105,N_22182);
nor U26712 (N_26712,N_24845,N_20411);
xor U26713 (N_26713,N_21053,N_24006);
nor U26714 (N_26714,N_20836,N_22720);
nand U26715 (N_26715,N_22976,N_20571);
and U26716 (N_26716,N_23290,N_23647);
or U26717 (N_26717,N_24466,N_23429);
or U26718 (N_26718,N_22208,N_22587);
nor U26719 (N_26719,N_24752,N_23946);
or U26720 (N_26720,N_21851,N_22477);
and U26721 (N_26721,N_22179,N_24196);
and U26722 (N_26722,N_24427,N_24116);
and U26723 (N_26723,N_21403,N_24980);
nor U26724 (N_26724,N_20333,N_24003);
xor U26725 (N_26725,N_24762,N_22356);
and U26726 (N_26726,N_20491,N_21600);
nor U26727 (N_26727,N_20610,N_23760);
and U26728 (N_26728,N_21279,N_24767);
nand U26729 (N_26729,N_23587,N_22681);
xor U26730 (N_26730,N_20633,N_22480);
and U26731 (N_26731,N_22909,N_22083);
and U26732 (N_26732,N_21445,N_24919);
nor U26733 (N_26733,N_24861,N_21309);
nand U26734 (N_26734,N_22984,N_22248);
and U26735 (N_26735,N_22301,N_22519);
nor U26736 (N_26736,N_23256,N_20656);
nand U26737 (N_26737,N_24624,N_23270);
or U26738 (N_26738,N_24051,N_20848);
nand U26739 (N_26739,N_22558,N_21790);
or U26740 (N_26740,N_22377,N_20379);
or U26741 (N_26741,N_21258,N_20446);
or U26742 (N_26742,N_20797,N_24912);
xor U26743 (N_26743,N_21009,N_22463);
xor U26744 (N_26744,N_21613,N_21734);
xor U26745 (N_26745,N_23150,N_22213);
nand U26746 (N_26746,N_24337,N_24668);
xor U26747 (N_26747,N_21062,N_22324);
and U26748 (N_26748,N_23297,N_23617);
nor U26749 (N_26749,N_23092,N_23844);
or U26750 (N_26750,N_21519,N_24866);
nand U26751 (N_26751,N_23333,N_24479);
xnor U26752 (N_26752,N_23574,N_20947);
nor U26753 (N_26753,N_20672,N_23403);
or U26754 (N_26754,N_21219,N_22347);
and U26755 (N_26755,N_24244,N_20645);
xnor U26756 (N_26756,N_21914,N_20408);
or U26757 (N_26757,N_21979,N_23320);
nand U26758 (N_26758,N_21335,N_24132);
or U26759 (N_26759,N_22082,N_20927);
and U26760 (N_26760,N_24255,N_21303);
nand U26761 (N_26761,N_20504,N_21002);
or U26762 (N_26762,N_23786,N_22581);
nand U26763 (N_26763,N_20109,N_21407);
nand U26764 (N_26764,N_23043,N_24679);
nor U26765 (N_26765,N_23124,N_21256);
nand U26766 (N_26766,N_23299,N_22423);
nand U26767 (N_26767,N_21181,N_24770);
xor U26768 (N_26768,N_20096,N_22465);
or U26769 (N_26769,N_23762,N_24005);
and U26770 (N_26770,N_20754,N_22084);
or U26771 (N_26771,N_20427,N_22548);
or U26772 (N_26772,N_22755,N_24863);
xnor U26773 (N_26773,N_23405,N_21866);
and U26774 (N_26774,N_23949,N_20407);
and U26775 (N_26775,N_23868,N_21429);
or U26776 (N_26776,N_22448,N_22397);
nand U26777 (N_26777,N_24214,N_21467);
nor U26778 (N_26778,N_24169,N_22321);
and U26779 (N_26779,N_23952,N_23367);
and U26780 (N_26780,N_21529,N_24443);
and U26781 (N_26781,N_22715,N_22476);
and U26782 (N_26782,N_23378,N_20250);
nor U26783 (N_26783,N_23132,N_24263);
or U26784 (N_26784,N_20029,N_20850);
nor U26785 (N_26785,N_21090,N_24369);
and U26786 (N_26786,N_24732,N_21769);
nand U26787 (N_26787,N_22249,N_23939);
or U26788 (N_26788,N_20123,N_24130);
xor U26789 (N_26789,N_22018,N_22791);
and U26790 (N_26790,N_21317,N_20343);
xor U26791 (N_26791,N_21451,N_21993);
nor U26792 (N_26792,N_24074,N_22529);
or U26793 (N_26793,N_20911,N_24803);
nand U26794 (N_26794,N_22389,N_21431);
nor U26795 (N_26795,N_20946,N_23554);
and U26796 (N_26796,N_20904,N_22148);
xor U26797 (N_26797,N_22513,N_22908);
nand U26798 (N_26798,N_22268,N_24738);
nand U26799 (N_26799,N_23605,N_22044);
nand U26800 (N_26800,N_21005,N_24351);
nand U26801 (N_26801,N_20529,N_21594);
or U26802 (N_26802,N_21189,N_22041);
nor U26803 (N_26803,N_21340,N_24688);
or U26804 (N_26804,N_22146,N_23216);
or U26805 (N_26805,N_24955,N_24499);
or U26806 (N_26806,N_20016,N_20476);
xor U26807 (N_26807,N_21492,N_22290);
nand U26808 (N_26808,N_21464,N_20206);
nand U26809 (N_26809,N_24136,N_24419);
nor U26810 (N_26810,N_20368,N_23090);
xor U26811 (N_26811,N_22374,N_22378);
xor U26812 (N_26812,N_22432,N_23321);
and U26813 (N_26813,N_20129,N_22133);
and U26814 (N_26814,N_23722,N_24864);
and U26815 (N_26815,N_22272,N_22212);
nand U26816 (N_26816,N_22029,N_21854);
xor U26817 (N_26817,N_24627,N_24022);
and U26818 (N_26818,N_20527,N_23575);
and U26819 (N_26819,N_21741,N_21169);
xnor U26820 (N_26820,N_23487,N_21244);
nor U26821 (N_26821,N_21101,N_21372);
or U26822 (N_26822,N_23059,N_23154);
and U26823 (N_26823,N_20862,N_20995);
or U26824 (N_26824,N_23029,N_22747);
nor U26825 (N_26825,N_24407,N_24226);
nand U26826 (N_26826,N_21663,N_22573);
xnor U26827 (N_26827,N_20704,N_23084);
or U26828 (N_26828,N_20784,N_22911);
or U26829 (N_26829,N_20591,N_22140);
xor U26830 (N_26830,N_24444,N_21012);
nor U26831 (N_26831,N_23171,N_24452);
or U26832 (N_26832,N_24746,N_20023);
xnor U26833 (N_26833,N_23156,N_20508);
nand U26834 (N_26834,N_22667,N_20715);
nand U26835 (N_26835,N_23951,N_20688);
and U26836 (N_26836,N_21548,N_23960);
nand U26837 (N_26837,N_24201,N_20718);
or U26838 (N_26838,N_23467,N_22618);
and U26839 (N_26839,N_24441,N_23076);
nor U26840 (N_26840,N_20728,N_23837);
and U26841 (N_26841,N_21282,N_24204);
and U26842 (N_26842,N_20103,N_23538);
nand U26843 (N_26843,N_23032,N_22924);
nand U26844 (N_26844,N_20335,N_20786);
or U26845 (N_26845,N_22898,N_21847);
and U26846 (N_26846,N_24024,N_20102);
nor U26847 (N_26847,N_24468,N_20221);
nand U26848 (N_26848,N_22319,N_20798);
and U26849 (N_26849,N_21440,N_22806);
or U26850 (N_26850,N_23442,N_23406);
and U26851 (N_26851,N_23330,N_23724);
or U26852 (N_26852,N_21151,N_24442);
nor U26853 (N_26853,N_22387,N_22843);
nor U26854 (N_26854,N_20738,N_20303);
and U26855 (N_26855,N_20365,N_22430);
nor U26856 (N_26856,N_21892,N_24149);
nor U26857 (N_26857,N_22230,N_20858);
xor U26858 (N_26858,N_21213,N_22013);
nor U26859 (N_26859,N_21307,N_24272);
nand U26860 (N_26860,N_20013,N_23832);
nor U26861 (N_26861,N_22642,N_23099);
or U26862 (N_26862,N_23194,N_22475);
or U26863 (N_26863,N_24408,N_21325);
xnor U26864 (N_26864,N_22364,N_22232);
xor U26865 (N_26865,N_21614,N_24113);
xor U26866 (N_26866,N_23238,N_24954);
nor U26867 (N_26867,N_20039,N_24504);
nand U26868 (N_26868,N_22155,N_20481);
or U26869 (N_26869,N_23027,N_23588);
nor U26870 (N_26870,N_20567,N_20142);
and U26871 (N_26871,N_22999,N_24880);
and U26872 (N_26872,N_20787,N_23251);
nor U26873 (N_26873,N_21536,N_23155);
and U26874 (N_26874,N_24420,N_22975);
and U26875 (N_26875,N_23353,N_21690);
and U26876 (N_26876,N_20987,N_22818);
nor U26877 (N_26877,N_23061,N_20087);
nand U26878 (N_26878,N_23219,N_22698);
nor U26879 (N_26879,N_23957,N_20110);
or U26880 (N_26880,N_24682,N_23748);
nor U26881 (N_26881,N_24308,N_23302);
and U26882 (N_26882,N_22899,N_22403);
nand U26883 (N_26883,N_22449,N_23344);
or U26884 (N_26884,N_21752,N_21824);
xnor U26885 (N_26885,N_22473,N_21162);
or U26886 (N_26886,N_22417,N_23720);
nor U26887 (N_26887,N_22325,N_21391);
and U26888 (N_26888,N_20690,N_24282);
and U26889 (N_26889,N_23500,N_23369);
nor U26890 (N_26890,N_24772,N_21606);
nand U26891 (N_26891,N_21764,N_22474);
or U26892 (N_26892,N_22479,N_20707);
and U26893 (N_26893,N_21581,N_23854);
or U26894 (N_26894,N_22813,N_22424);
or U26895 (N_26895,N_20667,N_23548);
and U26896 (N_26896,N_22961,N_23039);
nor U26897 (N_26897,N_21533,N_22602);
nand U26898 (N_26898,N_24755,N_21855);
nor U26899 (N_26899,N_23050,N_22413);
nand U26900 (N_26900,N_21647,N_24434);
nand U26901 (N_26901,N_20941,N_20184);
nand U26902 (N_26902,N_24643,N_22517);
nand U26903 (N_26903,N_20698,N_23883);
and U26904 (N_26904,N_22826,N_21339);
nand U26905 (N_26905,N_24677,N_22867);
xor U26906 (N_26906,N_21689,N_21770);
nor U26907 (N_26907,N_24757,N_23064);
and U26908 (N_26908,N_20684,N_20133);
or U26909 (N_26909,N_24787,N_24843);
and U26910 (N_26910,N_23697,N_23373);
or U26911 (N_26911,N_22822,N_21478);
or U26912 (N_26912,N_22281,N_23522);
and U26913 (N_26913,N_20153,N_24823);
and U26914 (N_26914,N_21998,N_23387);
nor U26915 (N_26915,N_22920,N_23407);
and U26916 (N_26916,N_20318,N_22770);
nor U26917 (N_26917,N_24537,N_20084);
nor U26918 (N_26918,N_21408,N_23362);
nor U26919 (N_26919,N_24486,N_22986);
nand U26920 (N_26920,N_21080,N_23158);
and U26921 (N_26921,N_22126,N_20919);
nor U26922 (N_26922,N_21794,N_20274);
or U26923 (N_26923,N_24063,N_23552);
or U26924 (N_26924,N_22607,N_23698);
nand U26925 (N_26925,N_21161,N_23530);
and U26926 (N_26926,N_21684,N_20839);
nor U26927 (N_26927,N_21632,N_24267);
nor U26928 (N_26928,N_23201,N_24464);
and U26929 (N_26929,N_23204,N_20433);
nand U26930 (N_26930,N_21019,N_23384);
nand U26931 (N_26931,N_21088,N_20589);
nor U26932 (N_26932,N_24445,N_22713);
or U26933 (N_26933,N_21097,N_23066);
or U26934 (N_26934,N_21853,N_21657);
and U26935 (N_26935,N_20219,N_24072);
or U26936 (N_26936,N_24372,N_24519);
or U26937 (N_26937,N_22496,N_24807);
and U26938 (N_26938,N_23577,N_23417);
or U26939 (N_26939,N_23390,N_22666);
nand U26940 (N_26940,N_23790,N_24412);
or U26941 (N_26941,N_20514,N_20391);
and U26942 (N_26942,N_23525,N_21014);
nand U26943 (N_26943,N_24940,N_20213);
nor U26944 (N_26944,N_22399,N_23594);
nor U26945 (N_26945,N_22195,N_23301);
or U26946 (N_26946,N_24897,N_20914);
nand U26947 (N_26947,N_22245,N_20349);
nand U26948 (N_26948,N_22233,N_24353);
and U26949 (N_26949,N_23342,N_24707);
or U26950 (N_26950,N_24202,N_20134);
nor U26951 (N_26951,N_24548,N_23388);
nand U26952 (N_26952,N_22940,N_23221);
and U26953 (N_26953,N_21771,N_22028);
and U26954 (N_26954,N_23049,N_20056);
nand U26955 (N_26955,N_22995,N_24781);
nand U26956 (N_26956,N_20579,N_24766);
or U26957 (N_26957,N_21916,N_24958);
nor U26958 (N_26958,N_24560,N_24307);
nor U26959 (N_26959,N_23857,N_24317);
and U26960 (N_26960,N_21051,N_20359);
nor U26961 (N_26961,N_24505,N_23122);
and U26962 (N_26962,N_23266,N_24854);
or U26963 (N_26963,N_22343,N_22617);
or U26964 (N_26964,N_24286,N_20042);
nand U26965 (N_26965,N_23573,N_24078);
nand U26966 (N_26966,N_22331,N_21113);
and U26967 (N_26967,N_21760,N_23361);
nand U26968 (N_26968,N_24071,N_22673);
nor U26969 (N_26969,N_22038,N_20778);
or U26970 (N_26970,N_21637,N_23175);
nand U26971 (N_26971,N_23743,N_23408);
nor U26972 (N_26972,N_21025,N_24751);
or U26973 (N_26973,N_22844,N_24670);
nor U26974 (N_26974,N_23526,N_23470);
or U26975 (N_26975,N_20496,N_21435);
nand U26976 (N_26976,N_24500,N_22737);
or U26977 (N_26977,N_23183,N_21937);
or U26978 (N_26978,N_23048,N_22887);
nand U26979 (N_26979,N_23849,N_22142);
nand U26980 (N_26980,N_22735,N_23985);
nor U26981 (N_26981,N_24790,N_23425);
or U26982 (N_26982,N_22250,N_23439);
nand U26983 (N_26983,N_23445,N_22974);
nand U26984 (N_26984,N_21271,N_21315);
nor U26985 (N_26985,N_20108,N_24146);
or U26986 (N_26986,N_24859,N_20395);
nand U26987 (N_26987,N_21730,N_23619);
nand U26988 (N_26988,N_20988,N_23528);
nor U26989 (N_26989,N_20393,N_23044);
and U26990 (N_26990,N_22510,N_20974);
or U26991 (N_26991,N_20530,N_20306);
or U26992 (N_26992,N_21490,N_21821);
nor U26993 (N_26993,N_24237,N_22329);
nor U26994 (N_26994,N_20886,N_21703);
and U26995 (N_26995,N_20367,N_22228);
nor U26996 (N_26996,N_22219,N_21095);
nand U26997 (N_26997,N_22937,N_20807);
and U26998 (N_26998,N_22869,N_24945);
or U26999 (N_26999,N_24972,N_20942);
nand U27000 (N_27000,N_23071,N_21152);
nor U27001 (N_27001,N_23858,N_24815);
and U27002 (N_27002,N_24455,N_21905);
nor U27003 (N_27003,N_23228,N_20613);
nand U27004 (N_27004,N_20776,N_20417);
or U27005 (N_27005,N_21778,N_20500);
nand U27006 (N_27006,N_20713,N_20253);
and U27007 (N_27007,N_24302,N_21565);
nor U27008 (N_27008,N_24028,N_21940);
xor U27009 (N_27009,N_24023,N_24528);
xnor U27010 (N_27010,N_20913,N_22921);
or U27011 (N_27011,N_22492,N_24246);
nor U27012 (N_27012,N_20541,N_20868);
nand U27013 (N_27013,N_24567,N_24175);
xor U27014 (N_27014,N_23349,N_22307);
and U27015 (N_27015,N_21416,N_23876);
xor U27016 (N_27016,N_20502,N_21955);
nand U27017 (N_27017,N_21196,N_23974);
and U27018 (N_27018,N_21602,N_24235);
xor U27019 (N_27019,N_20777,N_20972);
and U27020 (N_27020,N_21294,N_23599);
and U27021 (N_27021,N_22337,N_20534);
or U27022 (N_27022,N_22977,N_22134);
and U27023 (N_27023,N_21787,N_23502);
or U27024 (N_27024,N_23006,N_24745);
and U27025 (N_27025,N_22624,N_20661);
nor U27026 (N_27026,N_24044,N_20148);
nand U27027 (N_27027,N_22669,N_21357);
nand U27028 (N_27028,N_24793,N_20802);
nor U27029 (N_27029,N_24008,N_20982);
and U27030 (N_27030,N_22697,N_20268);
nor U27031 (N_27031,N_20658,N_21259);
and U27032 (N_27032,N_21831,N_23527);
or U27033 (N_27033,N_24041,N_23448);
or U27034 (N_27034,N_21227,N_23848);
nor U27035 (N_27035,N_24850,N_20311);
and U27036 (N_27036,N_20034,N_23292);
or U27037 (N_27037,N_23689,N_23861);
and U27038 (N_27038,N_22384,N_24127);
and U27039 (N_27039,N_24167,N_20757);
nand U27040 (N_27040,N_24413,N_21644);
nor U27041 (N_27041,N_20257,N_24498);
nand U27042 (N_27042,N_20841,N_21667);
xnor U27043 (N_27043,N_20869,N_21385);
nand U27044 (N_27044,N_23606,N_22210);
or U27045 (N_27045,N_22527,N_22811);
nor U27046 (N_27046,N_23196,N_20940);
nor U27047 (N_27047,N_22660,N_24778);
nand U27048 (N_27048,N_21906,N_20877);
nand U27049 (N_27049,N_22050,N_20553);
xor U27050 (N_27050,N_23922,N_20066);
nor U27051 (N_27051,N_21978,N_20419);
and U27052 (N_27052,N_21070,N_21344);
or U27053 (N_27053,N_24818,N_20814);
or U27054 (N_27054,N_24475,N_24250);
nand U27055 (N_27055,N_21883,N_24200);
nand U27056 (N_27056,N_24930,N_22001);
and U27057 (N_27057,N_21448,N_21696);
and U27058 (N_27058,N_23010,N_20161);
nand U27059 (N_27059,N_23835,N_21353);
nor U27060 (N_27060,N_22225,N_21687);
and U27061 (N_27061,N_22227,N_24663);
nor U27062 (N_27062,N_23045,N_23134);
and U27063 (N_27063,N_21588,N_20783);
and U27064 (N_27064,N_20337,N_21400);
and U27065 (N_27065,N_21517,N_24011);
and U27066 (N_27066,N_22973,N_24249);
nor U27067 (N_27067,N_20085,N_21368);
or U27068 (N_27068,N_24918,N_21556);
nor U27069 (N_27069,N_23351,N_22189);
nand U27070 (N_27070,N_22345,N_21539);
and U27071 (N_27071,N_22988,N_22271);
nor U27072 (N_27072,N_21840,N_22071);
and U27073 (N_27073,N_20144,N_22605);
or U27074 (N_27074,N_24114,N_23572);
nand U27075 (N_27075,N_21516,N_21413);
and U27076 (N_27076,N_20689,N_21629);
nand U27077 (N_27077,N_21078,N_20091);
nand U27078 (N_27078,N_22621,N_21874);
or U27079 (N_27079,N_24057,N_23821);
and U27080 (N_27080,N_23377,N_20829);
nor U27081 (N_27081,N_23808,N_21319);
and U27082 (N_27082,N_21965,N_23139);
nand U27083 (N_27083,N_21121,N_23162);
xnor U27084 (N_27084,N_22036,N_23086);
or U27085 (N_27085,N_20354,N_24949);
nand U27086 (N_27086,N_20826,N_22365);
xnor U27087 (N_27087,N_20300,N_20855);
nand U27088 (N_27088,N_20809,N_21392);
and U27089 (N_27089,N_20753,N_22960);
nand U27090 (N_27090,N_22661,N_20007);
nor U27091 (N_27091,N_20263,N_21105);
nor U27092 (N_27092,N_23986,N_20181);
nand U27093 (N_27093,N_22127,N_20761);
nand U27094 (N_27094,N_21096,N_24119);
nor U27095 (N_27095,N_20057,N_23510);
and U27096 (N_27096,N_20453,N_23945);
nor U27097 (N_27097,N_21201,N_23639);
xnor U27098 (N_27098,N_20597,N_21134);
and U27099 (N_27099,N_20222,N_22952);
nand U27100 (N_27100,N_22240,N_24217);
nor U27101 (N_27101,N_22539,N_23566);
nand U27102 (N_27102,N_20630,N_21551);
nand U27103 (N_27103,N_20316,N_24832);
nor U27104 (N_27104,N_23217,N_21534);
nand U27105 (N_27105,N_22804,N_23329);
nand U27106 (N_27106,N_21966,N_22808);
nand U27107 (N_27107,N_21920,N_24446);
nor U27108 (N_27108,N_24659,N_22570);
or U27109 (N_27109,N_20766,N_22662);
nand U27110 (N_27110,N_20202,N_21343);
and U27111 (N_27111,N_20755,N_24379);
nand U27112 (N_27112,N_22562,N_20050);
nand U27113 (N_27113,N_22686,N_23209);
and U27114 (N_27114,N_20154,N_24960);
nand U27115 (N_27115,N_22158,N_21285);
and U27116 (N_27116,N_24588,N_22689);
nor U27117 (N_27117,N_23007,N_20975);
or U27118 (N_27118,N_23908,N_22886);
and U27119 (N_27119,N_21150,N_20615);
nor U27120 (N_27120,N_21487,N_20054);
xnor U27121 (N_27121,N_23610,N_24809);
nor U27122 (N_27122,N_21850,N_20284);
nor U27123 (N_27123,N_22277,N_24092);
nor U27124 (N_27124,N_21880,N_22807);
and U27125 (N_27125,N_23915,N_21098);
nor U27126 (N_27126,N_21371,N_23775);
nand U27127 (N_27127,N_24341,N_21585);
and U27128 (N_27128,N_20294,N_21545);
or U27129 (N_27129,N_21555,N_22800);
or U27130 (N_27130,N_20775,N_21719);
nor U27131 (N_27131,N_24601,N_20804);
and U27132 (N_27132,N_24609,N_20721);
nand U27133 (N_27133,N_22677,N_22547);
nor U27134 (N_27134,N_21756,N_22427);
nor U27135 (N_27135,N_24414,N_21248);
nor U27136 (N_27136,N_21928,N_23355);
nand U27137 (N_27137,N_24245,N_20626);
or U27138 (N_27138,N_20430,N_22651);
and U27139 (N_27139,N_23665,N_22810);
and U27140 (N_27140,N_23366,N_24152);
and U27141 (N_27141,N_23298,N_22493);
and U27142 (N_27142,N_23678,N_20759);
xor U27143 (N_27143,N_20908,N_22462);
or U27144 (N_27144,N_24474,N_23804);
nand U27145 (N_27145,N_21115,N_24932);
nand U27146 (N_27146,N_22198,N_20341);
or U27147 (N_27147,N_22074,N_24043);
xor U27148 (N_27148,N_22913,N_22866);
nand U27149 (N_27149,N_22255,N_20651);
nor U27150 (N_27150,N_22418,N_20986);
nand U27151 (N_27151,N_23483,N_24388);
xnor U27152 (N_27152,N_22795,N_23919);
or U27153 (N_27153,N_24050,N_23869);
nand U27154 (N_27154,N_22380,N_23464);
or U27155 (N_27155,N_23307,N_21463);
and U27156 (N_27156,N_23357,N_22196);
nand U27157 (N_27157,N_21499,N_22779);
or U27158 (N_27158,N_21922,N_22261);
and U27159 (N_27159,N_21740,N_20929);
nor U27160 (N_27160,N_24240,N_20187);
and U27161 (N_27161,N_20273,N_22202);
nor U27162 (N_27162,N_20366,N_24404);
or U27163 (N_27163,N_20401,N_23582);
or U27164 (N_27164,N_22489,N_20404);
nand U27165 (N_27165,N_23051,N_23232);
and U27166 (N_27166,N_20000,N_23803);
nor U27167 (N_27167,N_24644,N_21907);
or U27168 (N_27168,N_24310,N_21583);
nand U27169 (N_27169,N_24915,N_24042);
and U27170 (N_27170,N_24891,N_20976);
nand U27171 (N_27171,N_22699,N_20998);
nand U27172 (N_27172,N_24081,N_20169);
nor U27173 (N_27173,N_22154,N_24387);
or U27174 (N_27174,N_23111,N_24680);
nor U27175 (N_27175,N_20782,N_24633);
and U27176 (N_27176,N_22595,N_23967);
nand U27177 (N_27177,N_23891,N_21209);
and U27178 (N_27178,N_20522,N_22221);
nor U27179 (N_27179,N_22220,N_24946);
or U27180 (N_27180,N_21396,N_21839);
nor U27181 (N_27181,N_20602,N_21877);
nor U27182 (N_27182,N_23581,N_22834);
nand U27183 (N_27183,N_24873,N_21665);
nor U27184 (N_27184,N_20745,N_24700);
nor U27185 (N_27185,N_22751,N_21449);
nor U27186 (N_27186,N_20447,N_24274);
nand U27187 (N_27187,N_20647,N_20487);
nand U27188 (N_27188,N_22907,N_20498);
and U27189 (N_27189,N_20089,N_24765);
nor U27190 (N_27190,N_22515,N_22408);
nand U27191 (N_27191,N_20997,N_23082);
and U27192 (N_27192,N_22827,N_21912);
nor U27193 (N_27193,N_20449,N_23756);
nor U27194 (N_27194,N_24756,N_20078);
and U27195 (N_27195,N_24987,N_22632);
nor U27196 (N_27196,N_24053,N_23547);
nor U27197 (N_27197,N_23988,N_22851);
or U27198 (N_27198,N_22860,N_24520);
nand U27199 (N_27199,N_22350,N_20360);
and U27200 (N_27200,N_21869,N_21859);
or U27201 (N_27201,N_23789,N_24418);
nand U27202 (N_27202,N_20789,N_23846);
and U27203 (N_27203,N_21387,N_24040);
nand U27204 (N_27204,N_22016,N_24939);
and U27205 (N_27205,N_21376,N_22057);
nor U27206 (N_27206,N_20340,N_20843);
nand U27207 (N_27207,N_21117,N_22525);
nand U27208 (N_27208,N_23309,N_21434);
nor U27209 (N_27209,N_24156,N_23325);
or U27210 (N_27210,N_20665,N_22638);
or U27211 (N_27211,N_23024,N_21625);
or U27212 (N_27212,N_23463,N_21261);
and U27213 (N_27213,N_23730,N_21136);
and U27214 (N_27214,N_21300,N_24281);
or U27215 (N_27215,N_24556,N_20137);
or U27216 (N_27216,N_20093,N_23950);
or U27217 (N_27217,N_22367,N_20055);
or U27218 (N_27218,N_20832,N_21058);
or U27219 (N_27219,N_24518,N_22979);
nor U27220 (N_27220,N_20012,N_20065);
xor U27221 (N_27221,N_23056,N_24261);
nand U27222 (N_27222,N_21481,N_20214);
or U27223 (N_27223,N_23303,N_22391);
nand U27224 (N_27224,N_22175,N_22692);
and U27225 (N_27225,N_20020,N_20373);
xor U27226 (N_27226,N_22487,N_20954);
nand U27227 (N_27227,N_23902,N_21825);
nor U27228 (N_27228,N_23033,N_23022);
nor U27229 (N_27229,N_20223,N_20387);
or U27230 (N_27230,N_21447,N_23636);
xor U27231 (N_27231,N_23965,N_24586);
or U27232 (N_27232,N_23983,N_21612);
and U27233 (N_27233,N_24628,N_23109);
or U27234 (N_27234,N_22161,N_21374);
or U27235 (N_27235,N_24242,N_20406);
nor U27236 (N_27236,N_22286,N_24158);
xnor U27237 (N_27237,N_20033,N_22420);
nand U27238 (N_27238,N_22131,N_21633);
nor U27239 (N_27239,N_20724,N_23014);
nor U27240 (N_27240,N_22246,N_24592);
or U27241 (N_27241,N_20864,N_20348);
nor U27242 (N_27242,N_24230,N_24559);
xnor U27243 (N_27243,N_20659,N_21747);
nor U27244 (N_27244,N_24270,N_24821);
or U27245 (N_27245,N_24205,N_21114);
nor U27246 (N_27246,N_23094,N_24630);
and U27247 (N_27247,N_20235,N_23136);
nand U27248 (N_27248,N_21223,N_24632);
nor U27249 (N_27249,N_20457,N_22985);
nor U27250 (N_27250,N_20562,N_23894);
nand U27251 (N_27251,N_20509,N_21712);
xor U27252 (N_27252,N_20853,N_21252);
and U27253 (N_27253,N_24329,N_22620);
nand U27254 (N_27254,N_22781,N_24533);
and U27255 (N_27255,N_20198,N_21913);
and U27256 (N_27256,N_23396,N_24186);
nor U27257 (N_27257,N_22889,N_21579);
or U27258 (N_27258,N_24571,N_24138);
nand U27259 (N_27259,N_23855,N_23687);
nor U27260 (N_27260,N_20796,N_24264);
or U27261 (N_27261,N_21389,N_24165);
nor U27262 (N_27262,N_23972,N_24608);
nand U27263 (N_27263,N_23208,N_21811);
xnor U27264 (N_27264,N_23063,N_22275);
and U27265 (N_27265,N_24375,N_22828);
or U27266 (N_27266,N_24029,N_24715);
nand U27267 (N_27267,N_24721,N_24219);
or U27268 (N_27268,N_23940,N_23585);
nand U27269 (N_27269,N_21601,N_23895);
nand U27270 (N_27270,N_24910,N_24675);
and U27271 (N_27271,N_22309,N_22244);
and U27272 (N_27272,N_20143,N_20983);
xor U27273 (N_27273,N_21272,N_24220);
nand U27274 (N_27274,N_21253,N_23982);
xor U27275 (N_27275,N_20208,N_24673);
nor U27276 (N_27276,N_23555,N_21862);
or U27277 (N_27277,N_21711,N_21010);
nor U27278 (N_27278,N_23412,N_20554);
or U27279 (N_27279,N_21118,N_24059);
or U27280 (N_27280,N_20865,N_20876);
xnor U27281 (N_27281,N_21302,N_20532);
and U27282 (N_27282,N_21924,N_24495);
nand U27283 (N_27283,N_20968,N_20673);
nand U27284 (N_27284,N_21412,N_24979);
or U27285 (N_27285,N_22445,N_22983);
and U27286 (N_27286,N_24722,N_22352);
or U27287 (N_27287,N_23723,N_21974);
or U27288 (N_27288,N_21164,N_23615);
or U27289 (N_27289,N_22159,N_20902);
or U27290 (N_27290,N_23191,N_24417);
or U27291 (N_27291,N_20548,N_22600);
nor U27292 (N_27292,N_23119,N_23805);
nand U27293 (N_27293,N_24993,N_23078);
xor U27294 (N_27294,N_20097,N_21668);
or U27295 (N_27295,N_22702,N_24259);
nor U27296 (N_27296,N_20462,N_22266);
and U27297 (N_27297,N_22406,N_24324);
nand U27298 (N_27298,N_21783,N_24162);
or U27299 (N_27299,N_20403,N_21679);
nand U27300 (N_27300,N_20884,N_24276);
nor U27301 (N_27301,N_21950,N_21384);
and U27302 (N_27302,N_21506,N_21704);
and U27303 (N_27303,N_23833,N_20664);
and U27304 (N_27304,N_20178,N_22925);
and U27305 (N_27305,N_20973,N_20999);
nor U27306 (N_27306,N_20592,N_21158);
xor U27307 (N_27307,N_22996,N_22732);
nand U27308 (N_27308,N_24515,N_23263);
nand U27309 (N_27309,N_24641,N_22612);
and U27310 (N_27310,N_20369,N_20195);
nor U27311 (N_27311,N_24197,N_24805);
nor U27312 (N_27312,N_21439,N_23860);
nor U27313 (N_27313,N_22905,N_23609);
or U27314 (N_27314,N_24614,N_24743);
and U27315 (N_27315,N_21079,N_22129);
nor U27316 (N_27316,N_23380,N_21986);
xnor U27317 (N_27317,N_23675,N_22566);
and U27318 (N_27318,N_23702,N_23211);
and U27319 (N_27319,N_24164,N_21845);
and U27320 (N_27320,N_22091,N_23561);
nor U27321 (N_27321,N_22455,N_24936);
nor U27322 (N_27322,N_21183,N_23233);
and U27323 (N_27323,N_21720,N_24706);
nor U27324 (N_27324,N_23699,N_23414);
or U27325 (N_27325,N_21304,N_21634);
nor U27326 (N_27326,N_20159,N_22453);
and U27327 (N_27327,N_23013,N_24431);
and U27328 (N_27328,N_21706,N_20734);
nand U27329 (N_27329,N_22226,N_23025);
nor U27330 (N_27330,N_22693,N_21414);
nor U27331 (N_27331,N_22639,N_22968);
nand U27332 (N_27332,N_21037,N_21202);
or U27333 (N_27333,N_24647,N_22411);
or U27334 (N_27334,N_22015,N_24409);
xnor U27335 (N_27335,N_22171,N_23809);
or U27336 (N_27336,N_24456,N_24492);
and U27337 (N_27337,N_23042,N_22583);
and U27338 (N_27338,N_24606,N_24191);
nand U27339 (N_27339,N_21792,N_20418);
nand U27340 (N_27340,N_21889,N_24851);
and U27341 (N_27341,N_20881,N_20892);
nor U27342 (N_27342,N_24508,N_21609);
xor U27343 (N_27343,N_23758,N_22980);
nand U27344 (N_27344,N_24583,N_22769);
and U27345 (N_27345,N_22156,N_24289);
nor U27346 (N_27346,N_21823,N_20177);
or U27347 (N_27347,N_20445,N_24740);
nor U27348 (N_27348,N_21422,N_24655);
nor U27349 (N_27349,N_20426,N_24997);
nand U27350 (N_27350,N_21762,N_24865);
or U27351 (N_27351,N_24791,N_21281);
nand U27352 (N_27352,N_22068,N_24640);
and U27353 (N_27353,N_24366,N_20516);
nand U27354 (N_27354,N_22217,N_20454);
and U27355 (N_27355,N_20692,N_21203);
nor U27356 (N_27356,N_22823,N_24768);
and U27357 (N_27357,N_21584,N_20646);
nor U27358 (N_27358,N_24776,N_21641);
and U27359 (N_27359,N_20236,N_23691);
or U27360 (N_27360,N_24947,N_24837);
or U27361 (N_27361,N_23570,N_24514);
nand U27362 (N_27362,N_21419,N_24378);
or U27363 (N_27363,N_22932,N_24895);
nand U27364 (N_27364,N_22774,N_20092);
nor U27365 (N_27365,N_20546,N_21995);
or U27366 (N_27366,N_24849,N_21894);
nor U27367 (N_27367,N_22152,N_23563);
nand U27368 (N_27368,N_21931,N_23468);
nand U27369 (N_27369,N_22744,N_20764);
xnor U27370 (N_27370,N_22123,N_21572);
and U27371 (N_27371,N_21664,N_22682);
and U27372 (N_27372,N_20246,N_23777);
nand U27373 (N_27373,N_24902,N_22957);
nor U27374 (N_27374,N_24061,N_20041);
nor U27375 (N_27375,N_21789,N_23324);
or U27376 (N_27376,N_21054,N_24868);
or U27377 (N_27377,N_23956,N_21510);
and U27378 (N_27378,N_20512,N_21871);
and U27379 (N_27379,N_20702,N_23096);
nor U27380 (N_27380,N_21273,N_24103);
xnor U27381 (N_27381,N_21035,N_21479);
and U27382 (N_27382,N_22874,N_21837);
nor U27383 (N_27383,N_24115,N_23553);
or U27384 (N_27384,N_23607,N_24080);
xnor U27385 (N_27385,N_21607,N_20163);
nand U27386 (N_27386,N_24635,N_21518);
nand U27387 (N_27387,N_23205,N_22546);
nand U27388 (N_27388,N_24852,N_22951);
or U27389 (N_27389,N_20781,N_20424);
nand U27390 (N_27390,N_23735,N_21558);
xor U27391 (N_27391,N_22483,N_20425);
nand U27392 (N_27392,N_23537,N_23416);
or U27393 (N_27393,N_20813,N_24585);
and U27394 (N_27394,N_21324,N_20045);
or U27395 (N_27395,N_24534,N_21700);
and U27396 (N_27396,N_20052,N_24555);
and U27397 (N_27397,N_22194,N_21784);
nand U27398 (N_27398,N_24658,N_20900);
or U27399 (N_27399,N_21363,N_20240);
xnor U27400 (N_27400,N_22315,N_21184);
and U27401 (N_27401,N_23823,N_24685);
nand U27402 (N_27402,N_22072,N_22020);
nor U27403 (N_27403,N_21122,N_21356);
or U27404 (N_27404,N_21716,N_22491);
or U27405 (N_27405,N_20838,N_20835);
nor U27406 (N_27406,N_22858,N_23896);
and U27407 (N_27407,N_20111,N_21046);
or U27408 (N_27408,N_23137,N_22000);
or U27409 (N_27409,N_23964,N_22415);
or U27410 (N_27410,N_24942,N_21836);
or U27411 (N_27411,N_20296,N_23496);
nor U27412 (N_27412,N_22892,N_23761);
or U27413 (N_27413,N_20605,N_23065);
nor U27414 (N_27414,N_21144,N_24123);
or U27415 (N_27415,N_20593,N_24253);
nand U27416 (N_27416,N_23097,N_24491);
nand U27417 (N_27417,N_20155,N_24542);
nor U27418 (N_27418,N_23052,N_24331);
nor U27419 (N_27419,N_24027,N_21685);
nor U27420 (N_27420,N_22592,N_20537);
or U27421 (N_27421,N_20017,N_23690);
nor U27422 (N_27422,N_20966,N_20818);
nor U27423 (N_27423,N_22135,N_22021);
nor U27424 (N_27424,N_23545,N_22274);
nor U27425 (N_27425,N_21346,N_24129);
nor U27426 (N_27426,N_21718,N_21917);
and U27427 (N_27427,N_23168,N_20179);
nor U27428 (N_27428,N_20743,N_24493);
or U27429 (N_27429,N_23375,N_22499);
or U27430 (N_27430,N_23517,N_23186);
nand U27431 (N_27431,N_23862,N_20937);
or U27432 (N_27432,N_24018,N_21288);
or U27433 (N_27433,N_23710,N_23551);
nand U27434 (N_27434,N_23847,N_21605);
and U27435 (N_27435,N_24610,N_22326);
nor U27436 (N_27436,N_24971,N_23912);
nand U27437 (N_27437,N_20286,N_20628);
or U27438 (N_27438,N_22854,N_24360);
or U27439 (N_27439,N_23713,N_20464);
and U27440 (N_27440,N_24333,N_24128);
nor U27441 (N_27441,N_21976,N_24626);
nor U27442 (N_27442,N_24783,N_20423);
nand U27443 (N_27443,N_22160,N_23444);
and U27444 (N_27444,N_24425,N_21157);
nand U27445 (N_27445,N_24549,N_23454);
nand U27446 (N_27446,N_23600,N_21576);
nand U27447 (N_27447,N_21143,N_22728);
nand U27448 (N_27448,N_20322,N_23348);
nor U27449 (N_27449,N_22410,N_24657);
nand U27450 (N_27450,N_22753,N_23258);
nand U27451 (N_27451,N_20226,N_22070);
and U27452 (N_27452,N_22183,N_22458);
nor U27453 (N_27453,N_21060,N_21210);
nand U27454 (N_27454,N_20248,N_21024);
nor U27455 (N_27455,N_22398,N_20506);
nor U27456 (N_27456,N_23185,N_22793);
nor U27457 (N_27457,N_21554,N_22419);
nor U27458 (N_27458,N_20014,N_21165);
or U27459 (N_27459,N_22471,N_20070);
xor U27460 (N_27460,N_20851,N_21072);
and U27461 (N_27461,N_21145,N_24239);
or U27462 (N_27462,N_23529,N_24988);
or U27463 (N_27463,N_20207,N_20149);
and U27464 (N_27464,N_20740,N_24973);
or U27465 (N_27465,N_24878,N_20086);
and U27466 (N_27466,N_21742,N_20635);
or U27467 (N_27467,N_20817,N_23650);
and U27468 (N_27468,N_24347,N_23559);
or U27469 (N_27469,N_22842,N_20409);
and U27470 (N_27470,N_22180,N_24154);
nor U27471 (N_27471,N_21829,N_21959);
nand U27472 (N_27472,N_21083,N_24451);
or U27473 (N_27473,N_24060,N_22619);
nand U27474 (N_27474,N_21048,N_20280);
nor U27475 (N_27475,N_22763,N_22289);
or U27476 (N_27476,N_21666,N_24813);
nor U27477 (N_27477,N_20846,N_20332);
and U27478 (N_27478,N_21800,N_22773);
xnor U27479 (N_27479,N_22470,N_20168);
and U27480 (N_27480,N_21345,N_23852);
or U27481 (N_27481,N_24406,N_23627);
xnor U27482 (N_27482,N_23286,N_20648);
or U27483 (N_27483,N_24698,N_23410);
xor U27484 (N_27484,N_23213,N_24480);
or U27485 (N_27485,N_22433,N_20455);
and U27486 (N_27486,N_22784,N_20933);
nor U27487 (N_27487,N_24996,N_24461);
and U27488 (N_27488,N_20823,N_23100);
or U27489 (N_27489,N_20132,N_20668);
and U27490 (N_27490,N_24339,N_22762);
or U27491 (N_27491,N_24986,N_23401);
or U27492 (N_27492,N_22943,N_23011);
or U27493 (N_27493,N_21139,N_23072);
or U27494 (N_27494,N_21065,N_20887);
and U27495 (N_27495,N_21895,N_21146);
nand U27496 (N_27496,N_24391,N_23419);
nor U27497 (N_27497,N_20282,N_22342);
nand U27498 (N_27498,N_21250,N_24098);
nand U27499 (N_27499,N_20882,N_21803);
or U27500 (N_27500,N_24784,N_22065);
nand U27501 (N_27501,N_23555,N_22502);
or U27502 (N_27502,N_22769,N_24136);
nor U27503 (N_27503,N_24811,N_23637);
nand U27504 (N_27504,N_23097,N_23783);
and U27505 (N_27505,N_21483,N_20039);
nand U27506 (N_27506,N_23394,N_21490);
or U27507 (N_27507,N_20818,N_23221);
nand U27508 (N_27508,N_22112,N_24821);
nor U27509 (N_27509,N_21240,N_20701);
and U27510 (N_27510,N_23009,N_22936);
or U27511 (N_27511,N_24590,N_23835);
nand U27512 (N_27512,N_22375,N_22859);
or U27513 (N_27513,N_20393,N_20349);
nand U27514 (N_27514,N_22446,N_24802);
xor U27515 (N_27515,N_20748,N_22357);
nor U27516 (N_27516,N_23353,N_24964);
nor U27517 (N_27517,N_22876,N_24543);
nor U27518 (N_27518,N_23608,N_23589);
xnor U27519 (N_27519,N_20176,N_21940);
nor U27520 (N_27520,N_22377,N_20362);
and U27521 (N_27521,N_21947,N_22146);
nor U27522 (N_27522,N_22115,N_24136);
xnor U27523 (N_27523,N_21818,N_20686);
and U27524 (N_27524,N_23537,N_22658);
or U27525 (N_27525,N_23835,N_23112);
xor U27526 (N_27526,N_23301,N_24824);
nand U27527 (N_27527,N_21613,N_24623);
nor U27528 (N_27528,N_20974,N_24989);
or U27529 (N_27529,N_23247,N_22252);
nand U27530 (N_27530,N_21439,N_22786);
nor U27531 (N_27531,N_23218,N_24463);
nand U27532 (N_27532,N_21286,N_22452);
and U27533 (N_27533,N_22612,N_24581);
nor U27534 (N_27534,N_20724,N_22072);
nand U27535 (N_27535,N_24542,N_21028);
nand U27536 (N_27536,N_24457,N_24015);
and U27537 (N_27537,N_24029,N_24082);
or U27538 (N_27538,N_23341,N_22573);
nor U27539 (N_27539,N_21948,N_24527);
and U27540 (N_27540,N_24118,N_20156);
nor U27541 (N_27541,N_22513,N_24077);
and U27542 (N_27542,N_22924,N_21400);
or U27543 (N_27543,N_24994,N_24087);
and U27544 (N_27544,N_24838,N_22238);
nand U27545 (N_27545,N_21630,N_22735);
nand U27546 (N_27546,N_22623,N_20317);
nand U27547 (N_27547,N_20562,N_22689);
nor U27548 (N_27548,N_20056,N_24625);
nand U27549 (N_27549,N_21370,N_22832);
and U27550 (N_27550,N_20309,N_24311);
and U27551 (N_27551,N_23174,N_23599);
nand U27552 (N_27552,N_21824,N_22640);
nor U27553 (N_27553,N_22445,N_23799);
and U27554 (N_27554,N_21739,N_21005);
nand U27555 (N_27555,N_22912,N_22198);
nand U27556 (N_27556,N_23968,N_23542);
and U27557 (N_27557,N_21928,N_24633);
and U27558 (N_27558,N_23439,N_22509);
nor U27559 (N_27559,N_21821,N_20790);
or U27560 (N_27560,N_21662,N_23814);
xor U27561 (N_27561,N_20586,N_23064);
xnor U27562 (N_27562,N_24121,N_22495);
nor U27563 (N_27563,N_24193,N_22399);
and U27564 (N_27564,N_21891,N_21886);
nand U27565 (N_27565,N_23321,N_21660);
or U27566 (N_27566,N_23724,N_20635);
or U27567 (N_27567,N_20756,N_20123);
and U27568 (N_27568,N_22014,N_22015);
nor U27569 (N_27569,N_21026,N_21888);
or U27570 (N_27570,N_20629,N_21160);
xnor U27571 (N_27571,N_20128,N_21445);
nor U27572 (N_27572,N_21316,N_20088);
or U27573 (N_27573,N_24904,N_20910);
nand U27574 (N_27574,N_21870,N_21242);
and U27575 (N_27575,N_23983,N_23838);
or U27576 (N_27576,N_24625,N_22197);
or U27577 (N_27577,N_24448,N_21259);
nand U27578 (N_27578,N_22895,N_24694);
and U27579 (N_27579,N_23367,N_23022);
nor U27580 (N_27580,N_20409,N_22407);
nor U27581 (N_27581,N_23287,N_23653);
nand U27582 (N_27582,N_24213,N_22865);
nor U27583 (N_27583,N_23941,N_22007);
nand U27584 (N_27584,N_22214,N_22814);
or U27585 (N_27585,N_23886,N_24770);
or U27586 (N_27586,N_22476,N_20054);
or U27587 (N_27587,N_20417,N_24013);
and U27588 (N_27588,N_24998,N_22498);
nor U27589 (N_27589,N_20994,N_22108);
nand U27590 (N_27590,N_20171,N_22063);
and U27591 (N_27591,N_21510,N_20973);
and U27592 (N_27592,N_24394,N_22825);
nand U27593 (N_27593,N_20986,N_22235);
xor U27594 (N_27594,N_24019,N_22149);
nor U27595 (N_27595,N_23655,N_20524);
nor U27596 (N_27596,N_22239,N_24204);
and U27597 (N_27597,N_24850,N_23316);
and U27598 (N_27598,N_24861,N_24101);
nand U27599 (N_27599,N_20633,N_20882);
and U27600 (N_27600,N_23543,N_21155);
and U27601 (N_27601,N_23657,N_21400);
or U27602 (N_27602,N_20700,N_23619);
or U27603 (N_27603,N_20391,N_23963);
and U27604 (N_27604,N_22416,N_21534);
and U27605 (N_27605,N_21228,N_22600);
nor U27606 (N_27606,N_21805,N_21656);
xor U27607 (N_27607,N_20893,N_20589);
and U27608 (N_27608,N_23291,N_23278);
nand U27609 (N_27609,N_20564,N_20313);
nand U27610 (N_27610,N_23616,N_24790);
and U27611 (N_27611,N_24235,N_24935);
or U27612 (N_27612,N_24133,N_23956);
xor U27613 (N_27613,N_24763,N_23669);
xnor U27614 (N_27614,N_23930,N_21592);
or U27615 (N_27615,N_21164,N_23347);
and U27616 (N_27616,N_21695,N_23350);
and U27617 (N_27617,N_21757,N_23792);
or U27618 (N_27618,N_20729,N_24024);
or U27619 (N_27619,N_24634,N_20123);
nor U27620 (N_27620,N_21210,N_24474);
nor U27621 (N_27621,N_23270,N_24469);
nor U27622 (N_27622,N_23680,N_24217);
nor U27623 (N_27623,N_23497,N_22446);
and U27624 (N_27624,N_21683,N_21651);
or U27625 (N_27625,N_24584,N_22607);
or U27626 (N_27626,N_22107,N_21075);
xnor U27627 (N_27627,N_21218,N_22352);
or U27628 (N_27628,N_23997,N_24628);
or U27629 (N_27629,N_24772,N_23813);
nor U27630 (N_27630,N_22089,N_20463);
or U27631 (N_27631,N_24591,N_21237);
nand U27632 (N_27632,N_22207,N_20863);
or U27633 (N_27633,N_20254,N_23829);
nand U27634 (N_27634,N_24794,N_20814);
or U27635 (N_27635,N_24722,N_24701);
nand U27636 (N_27636,N_22277,N_21547);
xor U27637 (N_27637,N_20403,N_23554);
nand U27638 (N_27638,N_22898,N_20347);
nor U27639 (N_27639,N_20188,N_23265);
xnor U27640 (N_27640,N_24132,N_24094);
nor U27641 (N_27641,N_24168,N_20638);
nand U27642 (N_27642,N_22231,N_21252);
and U27643 (N_27643,N_22836,N_21244);
or U27644 (N_27644,N_21163,N_21998);
and U27645 (N_27645,N_20280,N_24333);
nor U27646 (N_27646,N_22125,N_21353);
xor U27647 (N_27647,N_20337,N_20287);
nor U27648 (N_27648,N_22712,N_24633);
nor U27649 (N_27649,N_24283,N_22197);
nand U27650 (N_27650,N_20584,N_20940);
and U27651 (N_27651,N_24820,N_22492);
nand U27652 (N_27652,N_20552,N_22678);
nand U27653 (N_27653,N_21446,N_22582);
nor U27654 (N_27654,N_23208,N_21337);
nor U27655 (N_27655,N_21935,N_22917);
nor U27656 (N_27656,N_20659,N_20234);
and U27657 (N_27657,N_24545,N_20476);
nor U27658 (N_27658,N_24516,N_20424);
nor U27659 (N_27659,N_22458,N_23343);
and U27660 (N_27660,N_21009,N_24213);
nand U27661 (N_27661,N_24034,N_21502);
nand U27662 (N_27662,N_20244,N_22874);
xnor U27663 (N_27663,N_24678,N_20930);
or U27664 (N_27664,N_23469,N_24399);
nor U27665 (N_27665,N_21714,N_23232);
and U27666 (N_27666,N_24747,N_23553);
nand U27667 (N_27667,N_23907,N_22313);
nor U27668 (N_27668,N_24193,N_24182);
or U27669 (N_27669,N_20867,N_22697);
nor U27670 (N_27670,N_21449,N_23697);
nor U27671 (N_27671,N_20556,N_24395);
and U27672 (N_27672,N_20686,N_23170);
or U27673 (N_27673,N_20970,N_22212);
nand U27674 (N_27674,N_21918,N_22025);
nand U27675 (N_27675,N_21441,N_22974);
nor U27676 (N_27676,N_21319,N_22738);
nor U27677 (N_27677,N_24171,N_21060);
and U27678 (N_27678,N_24820,N_24386);
nor U27679 (N_27679,N_20577,N_24490);
nor U27680 (N_27680,N_21045,N_23048);
nand U27681 (N_27681,N_24371,N_21601);
nand U27682 (N_27682,N_24203,N_23958);
nor U27683 (N_27683,N_22823,N_24634);
nand U27684 (N_27684,N_23364,N_20314);
and U27685 (N_27685,N_20986,N_21403);
or U27686 (N_27686,N_24974,N_20422);
or U27687 (N_27687,N_22371,N_24824);
nand U27688 (N_27688,N_23826,N_23149);
or U27689 (N_27689,N_22338,N_22905);
nand U27690 (N_27690,N_20639,N_20828);
and U27691 (N_27691,N_22218,N_23682);
and U27692 (N_27692,N_22989,N_23008);
nand U27693 (N_27693,N_22565,N_22307);
nor U27694 (N_27694,N_22976,N_21046);
xor U27695 (N_27695,N_24689,N_24954);
nor U27696 (N_27696,N_22871,N_24059);
and U27697 (N_27697,N_24692,N_21967);
or U27698 (N_27698,N_23415,N_23968);
nor U27699 (N_27699,N_24053,N_22898);
or U27700 (N_27700,N_22752,N_22390);
nor U27701 (N_27701,N_24894,N_22036);
and U27702 (N_27702,N_21545,N_23234);
and U27703 (N_27703,N_23816,N_23621);
nand U27704 (N_27704,N_21108,N_21104);
nand U27705 (N_27705,N_22449,N_23928);
xnor U27706 (N_27706,N_20094,N_22311);
and U27707 (N_27707,N_24159,N_21625);
or U27708 (N_27708,N_20038,N_23879);
xnor U27709 (N_27709,N_22490,N_23706);
nor U27710 (N_27710,N_20989,N_20448);
nor U27711 (N_27711,N_22359,N_20872);
or U27712 (N_27712,N_24437,N_22531);
or U27713 (N_27713,N_24335,N_23311);
or U27714 (N_27714,N_21512,N_20974);
nor U27715 (N_27715,N_21079,N_23125);
nand U27716 (N_27716,N_23863,N_23224);
and U27717 (N_27717,N_20595,N_23747);
and U27718 (N_27718,N_20624,N_23781);
xnor U27719 (N_27719,N_20583,N_21036);
xnor U27720 (N_27720,N_22849,N_24955);
or U27721 (N_27721,N_22198,N_20416);
or U27722 (N_27722,N_23148,N_23198);
and U27723 (N_27723,N_21231,N_20064);
and U27724 (N_27724,N_20269,N_22780);
and U27725 (N_27725,N_24002,N_20006);
or U27726 (N_27726,N_24211,N_24282);
nand U27727 (N_27727,N_24374,N_24681);
or U27728 (N_27728,N_21934,N_21912);
nand U27729 (N_27729,N_20150,N_22754);
nand U27730 (N_27730,N_22750,N_24209);
or U27731 (N_27731,N_22422,N_24498);
or U27732 (N_27732,N_20680,N_23169);
nor U27733 (N_27733,N_21232,N_20052);
or U27734 (N_27734,N_21422,N_22759);
nor U27735 (N_27735,N_21604,N_20284);
and U27736 (N_27736,N_23061,N_20153);
or U27737 (N_27737,N_23011,N_24351);
nand U27738 (N_27738,N_21038,N_24183);
and U27739 (N_27739,N_23242,N_23878);
and U27740 (N_27740,N_24283,N_20626);
nand U27741 (N_27741,N_21393,N_22443);
nor U27742 (N_27742,N_21264,N_21151);
or U27743 (N_27743,N_21450,N_23924);
or U27744 (N_27744,N_23296,N_20577);
nand U27745 (N_27745,N_20184,N_20351);
nor U27746 (N_27746,N_21088,N_24776);
nand U27747 (N_27747,N_23231,N_23229);
nand U27748 (N_27748,N_23287,N_21059);
or U27749 (N_27749,N_23363,N_21447);
xnor U27750 (N_27750,N_23866,N_22699);
nor U27751 (N_27751,N_23109,N_24215);
or U27752 (N_27752,N_21466,N_24582);
or U27753 (N_27753,N_22945,N_22803);
or U27754 (N_27754,N_22612,N_21283);
and U27755 (N_27755,N_22244,N_24949);
nor U27756 (N_27756,N_20426,N_22345);
xor U27757 (N_27757,N_21768,N_22721);
or U27758 (N_27758,N_22961,N_24812);
nor U27759 (N_27759,N_21981,N_20451);
xor U27760 (N_27760,N_22895,N_22263);
nor U27761 (N_27761,N_21410,N_22387);
and U27762 (N_27762,N_21575,N_22220);
nand U27763 (N_27763,N_24939,N_22693);
and U27764 (N_27764,N_21274,N_21028);
nand U27765 (N_27765,N_24148,N_20337);
or U27766 (N_27766,N_22234,N_20149);
nor U27767 (N_27767,N_21726,N_23934);
nand U27768 (N_27768,N_20358,N_22010);
and U27769 (N_27769,N_23224,N_22604);
nor U27770 (N_27770,N_21294,N_23454);
nand U27771 (N_27771,N_23677,N_21217);
and U27772 (N_27772,N_23905,N_23293);
nor U27773 (N_27773,N_22205,N_23937);
nand U27774 (N_27774,N_22202,N_20515);
and U27775 (N_27775,N_20439,N_20798);
nor U27776 (N_27776,N_24564,N_23054);
nand U27777 (N_27777,N_24330,N_24868);
or U27778 (N_27778,N_22368,N_21017);
or U27779 (N_27779,N_24530,N_22713);
nor U27780 (N_27780,N_20986,N_22124);
nand U27781 (N_27781,N_24384,N_21362);
or U27782 (N_27782,N_24306,N_21287);
nor U27783 (N_27783,N_22229,N_24247);
and U27784 (N_27784,N_20155,N_21558);
nor U27785 (N_27785,N_21468,N_21842);
nor U27786 (N_27786,N_20700,N_23679);
or U27787 (N_27787,N_23080,N_22338);
nor U27788 (N_27788,N_21715,N_20905);
and U27789 (N_27789,N_23632,N_20843);
or U27790 (N_27790,N_21476,N_21938);
nand U27791 (N_27791,N_23670,N_24939);
nand U27792 (N_27792,N_22520,N_21495);
or U27793 (N_27793,N_20400,N_23129);
nor U27794 (N_27794,N_21884,N_20418);
xor U27795 (N_27795,N_24315,N_24063);
nor U27796 (N_27796,N_24767,N_24472);
nor U27797 (N_27797,N_20743,N_21563);
or U27798 (N_27798,N_22212,N_24182);
nor U27799 (N_27799,N_20471,N_20755);
nand U27800 (N_27800,N_24817,N_21389);
nor U27801 (N_27801,N_22182,N_22752);
and U27802 (N_27802,N_23714,N_24251);
or U27803 (N_27803,N_23066,N_20598);
nand U27804 (N_27804,N_24118,N_22001);
nand U27805 (N_27805,N_20211,N_22959);
or U27806 (N_27806,N_24452,N_21438);
nand U27807 (N_27807,N_23266,N_23574);
nand U27808 (N_27808,N_22422,N_22273);
or U27809 (N_27809,N_21380,N_21052);
and U27810 (N_27810,N_22612,N_22224);
or U27811 (N_27811,N_21205,N_23276);
and U27812 (N_27812,N_24393,N_24770);
nand U27813 (N_27813,N_20230,N_22852);
nand U27814 (N_27814,N_23394,N_21199);
nor U27815 (N_27815,N_23348,N_24954);
nor U27816 (N_27816,N_22294,N_23005);
nand U27817 (N_27817,N_22096,N_21413);
nor U27818 (N_27818,N_20615,N_21205);
and U27819 (N_27819,N_20612,N_21601);
or U27820 (N_27820,N_20825,N_21252);
and U27821 (N_27821,N_20342,N_23809);
nor U27822 (N_27822,N_22919,N_23644);
nor U27823 (N_27823,N_21763,N_22759);
nand U27824 (N_27824,N_20251,N_22098);
and U27825 (N_27825,N_23436,N_20355);
and U27826 (N_27826,N_24495,N_23655);
nor U27827 (N_27827,N_23658,N_20701);
and U27828 (N_27828,N_24935,N_24337);
and U27829 (N_27829,N_21630,N_21953);
or U27830 (N_27830,N_24991,N_21243);
xor U27831 (N_27831,N_24704,N_21939);
or U27832 (N_27832,N_22933,N_20103);
or U27833 (N_27833,N_24338,N_22005);
nor U27834 (N_27834,N_24175,N_23584);
or U27835 (N_27835,N_23731,N_24684);
xor U27836 (N_27836,N_24611,N_20800);
or U27837 (N_27837,N_22699,N_24848);
or U27838 (N_27838,N_20689,N_22080);
and U27839 (N_27839,N_20767,N_23920);
xnor U27840 (N_27840,N_21769,N_20978);
nor U27841 (N_27841,N_22192,N_24517);
nor U27842 (N_27842,N_23511,N_23339);
and U27843 (N_27843,N_20383,N_22612);
or U27844 (N_27844,N_21876,N_20389);
and U27845 (N_27845,N_21820,N_22619);
nor U27846 (N_27846,N_24508,N_23571);
nand U27847 (N_27847,N_24397,N_22005);
nor U27848 (N_27848,N_23623,N_24426);
nor U27849 (N_27849,N_20437,N_20171);
and U27850 (N_27850,N_22752,N_22725);
nor U27851 (N_27851,N_21815,N_23067);
xor U27852 (N_27852,N_21746,N_22644);
and U27853 (N_27853,N_24152,N_20450);
xnor U27854 (N_27854,N_20962,N_23424);
nand U27855 (N_27855,N_22169,N_23183);
nor U27856 (N_27856,N_24481,N_24757);
nand U27857 (N_27857,N_22796,N_21443);
nand U27858 (N_27858,N_20560,N_22172);
or U27859 (N_27859,N_24187,N_24103);
or U27860 (N_27860,N_23544,N_24203);
xnor U27861 (N_27861,N_24782,N_21704);
nand U27862 (N_27862,N_20037,N_23394);
and U27863 (N_27863,N_24434,N_22993);
and U27864 (N_27864,N_21084,N_23895);
or U27865 (N_27865,N_22525,N_22506);
nand U27866 (N_27866,N_23422,N_22146);
nand U27867 (N_27867,N_22701,N_20217);
or U27868 (N_27868,N_22492,N_23844);
nand U27869 (N_27869,N_20555,N_24783);
nor U27870 (N_27870,N_20859,N_24322);
or U27871 (N_27871,N_23064,N_23785);
nor U27872 (N_27872,N_22212,N_23957);
nand U27873 (N_27873,N_21542,N_23191);
nor U27874 (N_27874,N_22628,N_21122);
nor U27875 (N_27875,N_20987,N_23117);
and U27876 (N_27876,N_24717,N_22535);
nor U27877 (N_27877,N_24498,N_20792);
nor U27878 (N_27878,N_24026,N_23689);
xnor U27879 (N_27879,N_20262,N_21281);
nand U27880 (N_27880,N_22552,N_23075);
nand U27881 (N_27881,N_23484,N_20534);
xnor U27882 (N_27882,N_21880,N_22146);
and U27883 (N_27883,N_21615,N_23565);
nand U27884 (N_27884,N_22196,N_20174);
nand U27885 (N_27885,N_23478,N_21167);
nor U27886 (N_27886,N_20358,N_20377);
and U27887 (N_27887,N_21607,N_23508);
xor U27888 (N_27888,N_21348,N_23451);
nand U27889 (N_27889,N_21715,N_23055);
xor U27890 (N_27890,N_20248,N_23021);
or U27891 (N_27891,N_23050,N_24758);
nor U27892 (N_27892,N_22162,N_24276);
and U27893 (N_27893,N_20728,N_21548);
nand U27894 (N_27894,N_21531,N_23400);
and U27895 (N_27895,N_20802,N_22580);
and U27896 (N_27896,N_23225,N_21636);
or U27897 (N_27897,N_22393,N_24072);
nor U27898 (N_27898,N_23485,N_20066);
or U27899 (N_27899,N_23856,N_24563);
nand U27900 (N_27900,N_23746,N_20070);
and U27901 (N_27901,N_24993,N_22979);
or U27902 (N_27902,N_23735,N_22745);
nand U27903 (N_27903,N_24076,N_22284);
xor U27904 (N_27904,N_24336,N_20034);
nand U27905 (N_27905,N_21397,N_20800);
and U27906 (N_27906,N_21957,N_20298);
nand U27907 (N_27907,N_20963,N_22447);
or U27908 (N_27908,N_21053,N_20143);
xnor U27909 (N_27909,N_23353,N_22723);
nand U27910 (N_27910,N_20145,N_22291);
nor U27911 (N_27911,N_24723,N_20431);
and U27912 (N_27912,N_23955,N_24434);
and U27913 (N_27913,N_20119,N_21893);
and U27914 (N_27914,N_22404,N_21884);
nand U27915 (N_27915,N_24068,N_23430);
nand U27916 (N_27916,N_21317,N_23710);
nand U27917 (N_27917,N_22097,N_23356);
nor U27918 (N_27918,N_20448,N_21889);
and U27919 (N_27919,N_20745,N_23838);
or U27920 (N_27920,N_23984,N_20668);
or U27921 (N_27921,N_23846,N_24729);
or U27922 (N_27922,N_22938,N_20126);
or U27923 (N_27923,N_20086,N_20173);
nor U27924 (N_27924,N_21125,N_22633);
and U27925 (N_27925,N_23203,N_20695);
or U27926 (N_27926,N_23741,N_22808);
nand U27927 (N_27927,N_22415,N_23507);
and U27928 (N_27928,N_22128,N_20247);
or U27929 (N_27929,N_20937,N_21019);
or U27930 (N_27930,N_22334,N_20530);
nand U27931 (N_27931,N_21771,N_23469);
nand U27932 (N_27932,N_22565,N_20568);
nor U27933 (N_27933,N_23965,N_20116);
and U27934 (N_27934,N_22678,N_22776);
nor U27935 (N_27935,N_22509,N_24742);
xnor U27936 (N_27936,N_24424,N_23010);
or U27937 (N_27937,N_23839,N_24776);
nand U27938 (N_27938,N_22193,N_24963);
nand U27939 (N_27939,N_21404,N_24653);
and U27940 (N_27940,N_23867,N_20892);
or U27941 (N_27941,N_20585,N_24887);
xor U27942 (N_27942,N_21890,N_23419);
nor U27943 (N_27943,N_23161,N_21339);
nor U27944 (N_27944,N_20274,N_22356);
and U27945 (N_27945,N_23901,N_23407);
or U27946 (N_27946,N_23384,N_22977);
or U27947 (N_27947,N_20245,N_23222);
and U27948 (N_27948,N_20239,N_20673);
and U27949 (N_27949,N_20026,N_23024);
nor U27950 (N_27950,N_22635,N_24482);
nor U27951 (N_27951,N_24452,N_24653);
or U27952 (N_27952,N_20009,N_20132);
nand U27953 (N_27953,N_22272,N_20021);
nor U27954 (N_27954,N_20471,N_23271);
nand U27955 (N_27955,N_23396,N_24229);
nor U27956 (N_27956,N_24079,N_24180);
and U27957 (N_27957,N_23191,N_22249);
nand U27958 (N_27958,N_20778,N_24584);
and U27959 (N_27959,N_21720,N_20955);
nor U27960 (N_27960,N_20051,N_22322);
xor U27961 (N_27961,N_20962,N_23064);
or U27962 (N_27962,N_22151,N_20110);
xnor U27963 (N_27963,N_21089,N_24563);
or U27964 (N_27964,N_23047,N_20717);
nand U27965 (N_27965,N_23194,N_23846);
nor U27966 (N_27966,N_20130,N_24799);
or U27967 (N_27967,N_24933,N_22030);
nand U27968 (N_27968,N_20151,N_22516);
and U27969 (N_27969,N_20309,N_23133);
and U27970 (N_27970,N_21446,N_21501);
xnor U27971 (N_27971,N_21927,N_24110);
and U27972 (N_27972,N_23006,N_20587);
or U27973 (N_27973,N_21666,N_21307);
nor U27974 (N_27974,N_20451,N_21092);
nand U27975 (N_27975,N_23293,N_20962);
nor U27976 (N_27976,N_23501,N_20183);
nor U27977 (N_27977,N_24127,N_23416);
and U27978 (N_27978,N_24981,N_24098);
nor U27979 (N_27979,N_24883,N_21570);
and U27980 (N_27980,N_21775,N_24033);
and U27981 (N_27981,N_24800,N_24802);
or U27982 (N_27982,N_21318,N_24494);
and U27983 (N_27983,N_24506,N_21279);
nand U27984 (N_27984,N_21888,N_20866);
or U27985 (N_27985,N_24495,N_23127);
xnor U27986 (N_27986,N_24126,N_20989);
nand U27987 (N_27987,N_23860,N_23271);
or U27988 (N_27988,N_23648,N_24844);
and U27989 (N_27989,N_23781,N_20119);
nor U27990 (N_27990,N_21446,N_21368);
nor U27991 (N_27991,N_21559,N_20231);
nor U27992 (N_27992,N_24556,N_24822);
nand U27993 (N_27993,N_22156,N_20067);
xnor U27994 (N_27994,N_23419,N_23332);
or U27995 (N_27995,N_24108,N_22882);
nand U27996 (N_27996,N_21716,N_21170);
or U27997 (N_27997,N_21474,N_22438);
and U27998 (N_27998,N_24039,N_24819);
and U27999 (N_27999,N_22396,N_24469);
and U28000 (N_28000,N_23116,N_24641);
and U28001 (N_28001,N_21283,N_24727);
nor U28002 (N_28002,N_20892,N_20192);
nor U28003 (N_28003,N_20052,N_22711);
or U28004 (N_28004,N_20953,N_22063);
or U28005 (N_28005,N_20495,N_23956);
nand U28006 (N_28006,N_24064,N_23054);
or U28007 (N_28007,N_20755,N_23263);
or U28008 (N_28008,N_21316,N_22414);
or U28009 (N_28009,N_20787,N_22461);
nor U28010 (N_28010,N_22505,N_22330);
nand U28011 (N_28011,N_23445,N_20028);
or U28012 (N_28012,N_24442,N_23146);
nor U28013 (N_28013,N_21679,N_22470);
nor U28014 (N_28014,N_20025,N_23445);
and U28015 (N_28015,N_23474,N_24771);
nand U28016 (N_28016,N_24188,N_21876);
nand U28017 (N_28017,N_24661,N_21903);
nand U28018 (N_28018,N_22522,N_20474);
nor U28019 (N_28019,N_21501,N_20158);
or U28020 (N_28020,N_20070,N_24204);
nand U28021 (N_28021,N_23718,N_21486);
nand U28022 (N_28022,N_21428,N_24657);
or U28023 (N_28023,N_22054,N_23335);
nor U28024 (N_28024,N_23712,N_23701);
nand U28025 (N_28025,N_24541,N_22170);
xnor U28026 (N_28026,N_22332,N_22355);
nand U28027 (N_28027,N_20725,N_20543);
xor U28028 (N_28028,N_24722,N_23797);
nand U28029 (N_28029,N_20482,N_22953);
nor U28030 (N_28030,N_22387,N_21590);
or U28031 (N_28031,N_21486,N_21689);
or U28032 (N_28032,N_24847,N_24334);
xnor U28033 (N_28033,N_22547,N_24595);
and U28034 (N_28034,N_20087,N_21710);
or U28035 (N_28035,N_24969,N_20109);
nand U28036 (N_28036,N_21706,N_21779);
nand U28037 (N_28037,N_24348,N_23126);
or U28038 (N_28038,N_22327,N_22311);
or U28039 (N_28039,N_21129,N_20883);
or U28040 (N_28040,N_21855,N_24768);
nor U28041 (N_28041,N_20246,N_20214);
nand U28042 (N_28042,N_20377,N_23655);
nor U28043 (N_28043,N_22295,N_21455);
and U28044 (N_28044,N_24741,N_24484);
and U28045 (N_28045,N_23709,N_20565);
nand U28046 (N_28046,N_24908,N_21646);
nor U28047 (N_28047,N_20636,N_24684);
xor U28048 (N_28048,N_22432,N_22359);
nor U28049 (N_28049,N_24426,N_21580);
or U28050 (N_28050,N_20912,N_22737);
nor U28051 (N_28051,N_20096,N_22741);
nand U28052 (N_28052,N_23108,N_24040);
nand U28053 (N_28053,N_24252,N_23629);
xor U28054 (N_28054,N_24691,N_22459);
nor U28055 (N_28055,N_21375,N_22417);
nand U28056 (N_28056,N_22369,N_24291);
nor U28057 (N_28057,N_23312,N_24793);
and U28058 (N_28058,N_21526,N_20660);
nor U28059 (N_28059,N_24890,N_23094);
nor U28060 (N_28060,N_21436,N_23937);
and U28061 (N_28061,N_23250,N_24753);
nand U28062 (N_28062,N_23814,N_21441);
and U28063 (N_28063,N_20208,N_23704);
nand U28064 (N_28064,N_22652,N_23435);
or U28065 (N_28065,N_24395,N_20533);
and U28066 (N_28066,N_24211,N_20184);
nand U28067 (N_28067,N_21882,N_21356);
nand U28068 (N_28068,N_24661,N_22633);
nand U28069 (N_28069,N_20896,N_22998);
nor U28070 (N_28070,N_20418,N_22419);
nor U28071 (N_28071,N_24880,N_21193);
nand U28072 (N_28072,N_20550,N_21318);
nor U28073 (N_28073,N_20450,N_21996);
nand U28074 (N_28074,N_24716,N_20758);
or U28075 (N_28075,N_21305,N_23845);
xnor U28076 (N_28076,N_23099,N_20558);
nand U28077 (N_28077,N_22949,N_22477);
xnor U28078 (N_28078,N_24052,N_20902);
nor U28079 (N_28079,N_22008,N_21228);
and U28080 (N_28080,N_22356,N_20187);
or U28081 (N_28081,N_24347,N_20508);
and U28082 (N_28082,N_22333,N_22303);
nor U28083 (N_28083,N_24186,N_23456);
or U28084 (N_28084,N_21643,N_22073);
nand U28085 (N_28085,N_22682,N_20488);
or U28086 (N_28086,N_24080,N_23181);
nor U28087 (N_28087,N_22266,N_22501);
nand U28088 (N_28088,N_24811,N_22013);
xnor U28089 (N_28089,N_24012,N_23064);
and U28090 (N_28090,N_20026,N_21201);
xor U28091 (N_28091,N_21454,N_21122);
and U28092 (N_28092,N_21457,N_24391);
xor U28093 (N_28093,N_22395,N_24517);
and U28094 (N_28094,N_21456,N_21478);
nor U28095 (N_28095,N_23681,N_20387);
nor U28096 (N_28096,N_20328,N_24523);
or U28097 (N_28097,N_21855,N_24017);
xor U28098 (N_28098,N_23678,N_21737);
nor U28099 (N_28099,N_21179,N_20896);
and U28100 (N_28100,N_22839,N_23834);
xor U28101 (N_28101,N_21250,N_21365);
or U28102 (N_28102,N_23824,N_21094);
nor U28103 (N_28103,N_22619,N_21321);
nor U28104 (N_28104,N_20688,N_24025);
xnor U28105 (N_28105,N_22298,N_20566);
and U28106 (N_28106,N_21228,N_23570);
and U28107 (N_28107,N_21312,N_22752);
or U28108 (N_28108,N_24183,N_21958);
nor U28109 (N_28109,N_20982,N_22620);
or U28110 (N_28110,N_20372,N_20879);
and U28111 (N_28111,N_22002,N_23094);
and U28112 (N_28112,N_24968,N_22415);
nand U28113 (N_28113,N_24538,N_22095);
or U28114 (N_28114,N_23725,N_20924);
xor U28115 (N_28115,N_24985,N_23578);
nor U28116 (N_28116,N_21363,N_20182);
nor U28117 (N_28117,N_22308,N_24477);
and U28118 (N_28118,N_24694,N_24468);
nand U28119 (N_28119,N_20116,N_23666);
and U28120 (N_28120,N_20224,N_22517);
and U28121 (N_28121,N_21103,N_23228);
nand U28122 (N_28122,N_22354,N_21007);
or U28123 (N_28123,N_20632,N_20464);
or U28124 (N_28124,N_24720,N_21830);
and U28125 (N_28125,N_22402,N_20959);
and U28126 (N_28126,N_21687,N_24069);
and U28127 (N_28127,N_20630,N_24891);
nand U28128 (N_28128,N_24870,N_21790);
and U28129 (N_28129,N_21721,N_22199);
and U28130 (N_28130,N_23330,N_22347);
xor U28131 (N_28131,N_24212,N_20071);
xor U28132 (N_28132,N_22366,N_22332);
nand U28133 (N_28133,N_21516,N_20737);
nand U28134 (N_28134,N_21606,N_23044);
nand U28135 (N_28135,N_24134,N_20970);
nor U28136 (N_28136,N_21808,N_22879);
nand U28137 (N_28137,N_20297,N_20348);
nand U28138 (N_28138,N_22564,N_22092);
nor U28139 (N_28139,N_22022,N_23976);
nand U28140 (N_28140,N_21135,N_22439);
and U28141 (N_28141,N_23110,N_23221);
and U28142 (N_28142,N_24320,N_23705);
or U28143 (N_28143,N_24853,N_21966);
nand U28144 (N_28144,N_22157,N_21772);
nand U28145 (N_28145,N_21488,N_21186);
nor U28146 (N_28146,N_22474,N_21768);
xor U28147 (N_28147,N_21165,N_20194);
or U28148 (N_28148,N_21551,N_23917);
nand U28149 (N_28149,N_20522,N_20284);
or U28150 (N_28150,N_23928,N_23327);
nand U28151 (N_28151,N_20775,N_21886);
nand U28152 (N_28152,N_20931,N_23846);
xor U28153 (N_28153,N_23967,N_20930);
or U28154 (N_28154,N_20329,N_20110);
or U28155 (N_28155,N_24578,N_20587);
or U28156 (N_28156,N_20496,N_21625);
and U28157 (N_28157,N_21187,N_24479);
nand U28158 (N_28158,N_20279,N_20230);
or U28159 (N_28159,N_23179,N_24437);
nor U28160 (N_28160,N_20403,N_24843);
or U28161 (N_28161,N_21523,N_21054);
nand U28162 (N_28162,N_24841,N_22927);
nand U28163 (N_28163,N_20895,N_20703);
nand U28164 (N_28164,N_24915,N_20118);
or U28165 (N_28165,N_21138,N_23245);
or U28166 (N_28166,N_22191,N_20780);
xor U28167 (N_28167,N_22953,N_20319);
and U28168 (N_28168,N_20466,N_21844);
nand U28169 (N_28169,N_23894,N_24558);
nor U28170 (N_28170,N_24710,N_24421);
nor U28171 (N_28171,N_24503,N_20849);
or U28172 (N_28172,N_24308,N_23718);
and U28173 (N_28173,N_21375,N_21799);
and U28174 (N_28174,N_20560,N_22883);
nor U28175 (N_28175,N_21058,N_20812);
xor U28176 (N_28176,N_21091,N_22930);
and U28177 (N_28177,N_24342,N_20770);
nor U28178 (N_28178,N_22671,N_21130);
or U28179 (N_28179,N_24352,N_23870);
nand U28180 (N_28180,N_24657,N_22032);
and U28181 (N_28181,N_23456,N_23551);
xor U28182 (N_28182,N_22131,N_24488);
xor U28183 (N_28183,N_21724,N_20115);
nor U28184 (N_28184,N_22160,N_23719);
nor U28185 (N_28185,N_20626,N_22125);
nor U28186 (N_28186,N_20861,N_23203);
or U28187 (N_28187,N_23472,N_20432);
nor U28188 (N_28188,N_23206,N_22614);
xor U28189 (N_28189,N_24090,N_20316);
and U28190 (N_28190,N_21425,N_23402);
or U28191 (N_28191,N_23077,N_21301);
nand U28192 (N_28192,N_20953,N_21126);
or U28193 (N_28193,N_23000,N_24034);
and U28194 (N_28194,N_24176,N_22053);
nand U28195 (N_28195,N_20266,N_21129);
nand U28196 (N_28196,N_21945,N_21566);
nand U28197 (N_28197,N_22046,N_20978);
and U28198 (N_28198,N_22728,N_21788);
nand U28199 (N_28199,N_23285,N_22818);
and U28200 (N_28200,N_23919,N_23400);
or U28201 (N_28201,N_23239,N_20781);
and U28202 (N_28202,N_20555,N_20796);
nand U28203 (N_28203,N_23603,N_21661);
nand U28204 (N_28204,N_23961,N_24570);
and U28205 (N_28205,N_21792,N_22146);
xnor U28206 (N_28206,N_20355,N_24884);
nand U28207 (N_28207,N_21113,N_22552);
nand U28208 (N_28208,N_24779,N_22395);
or U28209 (N_28209,N_20181,N_23805);
nand U28210 (N_28210,N_20553,N_21542);
nor U28211 (N_28211,N_22116,N_20029);
and U28212 (N_28212,N_21665,N_24204);
and U28213 (N_28213,N_23175,N_24138);
or U28214 (N_28214,N_22018,N_22060);
and U28215 (N_28215,N_24280,N_21377);
and U28216 (N_28216,N_20502,N_21170);
nor U28217 (N_28217,N_21582,N_24882);
and U28218 (N_28218,N_21689,N_20193);
nand U28219 (N_28219,N_23787,N_24815);
nand U28220 (N_28220,N_22022,N_23051);
or U28221 (N_28221,N_21061,N_20790);
nand U28222 (N_28222,N_22563,N_24953);
or U28223 (N_28223,N_24416,N_23289);
nand U28224 (N_28224,N_24192,N_23008);
nand U28225 (N_28225,N_24249,N_23753);
and U28226 (N_28226,N_23494,N_24539);
or U28227 (N_28227,N_22310,N_24805);
nor U28228 (N_28228,N_20101,N_21058);
nor U28229 (N_28229,N_24640,N_22754);
and U28230 (N_28230,N_20025,N_23223);
nor U28231 (N_28231,N_22655,N_22344);
and U28232 (N_28232,N_22564,N_24221);
nor U28233 (N_28233,N_22634,N_21065);
nand U28234 (N_28234,N_21273,N_20780);
and U28235 (N_28235,N_21283,N_23350);
or U28236 (N_28236,N_20078,N_20666);
nor U28237 (N_28237,N_24434,N_21340);
nor U28238 (N_28238,N_24956,N_24853);
nor U28239 (N_28239,N_21243,N_22496);
nor U28240 (N_28240,N_23558,N_23384);
xor U28241 (N_28241,N_24836,N_20543);
nand U28242 (N_28242,N_20457,N_22938);
and U28243 (N_28243,N_22533,N_24076);
nand U28244 (N_28244,N_23818,N_21512);
xor U28245 (N_28245,N_22144,N_24971);
nor U28246 (N_28246,N_22634,N_20708);
nor U28247 (N_28247,N_20719,N_21215);
or U28248 (N_28248,N_21639,N_23878);
nand U28249 (N_28249,N_20486,N_22603);
xor U28250 (N_28250,N_22089,N_20713);
nor U28251 (N_28251,N_23499,N_22288);
xnor U28252 (N_28252,N_22114,N_22577);
or U28253 (N_28253,N_24425,N_23697);
or U28254 (N_28254,N_23323,N_24658);
nor U28255 (N_28255,N_24522,N_24365);
or U28256 (N_28256,N_21809,N_22534);
and U28257 (N_28257,N_20699,N_20703);
nor U28258 (N_28258,N_20880,N_22346);
or U28259 (N_28259,N_23027,N_24294);
or U28260 (N_28260,N_22679,N_22358);
nand U28261 (N_28261,N_23074,N_20360);
nor U28262 (N_28262,N_21145,N_23638);
or U28263 (N_28263,N_22139,N_24863);
nor U28264 (N_28264,N_23374,N_20182);
and U28265 (N_28265,N_22573,N_24186);
nor U28266 (N_28266,N_23146,N_23948);
or U28267 (N_28267,N_21455,N_23591);
nor U28268 (N_28268,N_20724,N_24989);
nand U28269 (N_28269,N_24148,N_24474);
nor U28270 (N_28270,N_22934,N_21079);
nor U28271 (N_28271,N_22489,N_21593);
nor U28272 (N_28272,N_20444,N_23234);
nand U28273 (N_28273,N_23720,N_20064);
or U28274 (N_28274,N_23891,N_20378);
or U28275 (N_28275,N_21838,N_23216);
nor U28276 (N_28276,N_20910,N_20333);
nor U28277 (N_28277,N_21158,N_24352);
xor U28278 (N_28278,N_20307,N_23669);
nor U28279 (N_28279,N_20492,N_21964);
nor U28280 (N_28280,N_22384,N_23256);
and U28281 (N_28281,N_20074,N_21265);
xor U28282 (N_28282,N_24369,N_21960);
and U28283 (N_28283,N_20923,N_22049);
and U28284 (N_28284,N_23478,N_23068);
or U28285 (N_28285,N_24215,N_24246);
nor U28286 (N_28286,N_20625,N_21829);
or U28287 (N_28287,N_20253,N_24584);
xor U28288 (N_28288,N_23919,N_22283);
nor U28289 (N_28289,N_23193,N_21926);
or U28290 (N_28290,N_24281,N_20551);
nand U28291 (N_28291,N_20226,N_20139);
nor U28292 (N_28292,N_22467,N_20698);
or U28293 (N_28293,N_23343,N_22228);
and U28294 (N_28294,N_24649,N_20208);
nor U28295 (N_28295,N_22806,N_24824);
or U28296 (N_28296,N_23180,N_21910);
nand U28297 (N_28297,N_24732,N_22019);
nor U28298 (N_28298,N_21872,N_21237);
nand U28299 (N_28299,N_24012,N_24882);
xnor U28300 (N_28300,N_22182,N_21016);
nor U28301 (N_28301,N_20484,N_23041);
nand U28302 (N_28302,N_23272,N_24117);
nand U28303 (N_28303,N_22873,N_20228);
nor U28304 (N_28304,N_21874,N_24754);
nand U28305 (N_28305,N_23270,N_20415);
xor U28306 (N_28306,N_24749,N_21086);
and U28307 (N_28307,N_24911,N_22456);
nor U28308 (N_28308,N_22639,N_23905);
or U28309 (N_28309,N_21967,N_22919);
and U28310 (N_28310,N_21779,N_22688);
or U28311 (N_28311,N_22199,N_24044);
nand U28312 (N_28312,N_21738,N_23764);
nor U28313 (N_28313,N_21321,N_24963);
and U28314 (N_28314,N_24335,N_23915);
or U28315 (N_28315,N_23424,N_22559);
nor U28316 (N_28316,N_21828,N_21164);
or U28317 (N_28317,N_22529,N_20325);
or U28318 (N_28318,N_22107,N_20004);
nand U28319 (N_28319,N_23434,N_21572);
and U28320 (N_28320,N_23888,N_21197);
xor U28321 (N_28321,N_21102,N_21186);
and U28322 (N_28322,N_20997,N_20216);
nor U28323 (N_28323,N_23874,N_22820);
or U28324 (N_28324,N_21920,N_24422);
nand U28325 (N_28325,N_23380,N_20503);
xor U28326 (N_28326,N_24379,N_22965);
nand U28327 (N_28327,N_22880,N_20088);
nor U28328 (N_28328,N_24508,N_24731);
or U28329 (N_28329,N_20246,N_22945);
nand U28330 (N_28330,N_24128,N_22765);
or U28331 (N_28331,N_20957,N_23192);
nand U28332 (N_28332,N_24742,N_23058);
or U28333 (N_28333,N_23034,N_21824);
and U28334 (N_28334,N_24298,N_21173);
nand U28335 (N_28335,N_21726,N_21252);
or U28336 (N_28336,N_22914,N_23695);
nor U28337 (N_28337,N_22774,N_24976);
nand U28338 (N_28338,N_23513,N_23618);
and U28339 (N_28339,N_22807,N_22504);
or U28340 (N_28340,N_23001,N_22990);
or U28341 (N_28341,N_21338,N_23894);
nand U28342 (N_28342,N_23328,N_22949);
nand U28343 (N_28343,N_21523,N_24913);
xor U28344 (N_28344,N_22131,N_21691);
xor U28345 (N_28345,N_22027,N_23439);
nor U28346 (N_28346,N_23167,N_20057);
nand U28347 (N_28347,N_22804,N_21556);
nand U28348 (N_28348,N_23064,N_24979);
nand U28349 (N_28349,N_20160,N_24854);
and U28350 (N_28350,N_20914,N_20023);
or U28351 (N_28351,N_21826,N_21583);
nor U28352 (N_28352,N_21702,N_23604);
nor U28353 (N_28353,N_20891,N_24352);
or U28354 (N_28354,N_21772,N_20137);
or U28355 (N_28355,N_21038,N_20180);
and U28356 (N_28356,N_21396,N_20263);
nor U28357 (N_28357,N_20365,N_22051);
nand U28358 (N_28358,N_22714,N_24028);
nand U28359 (N_28359,N_23131,N_20516);
nor U28360 (N_28360,N_24634,N_20681);
xnor U28361 (N_28361,N_24260,N_21526);
xnor U28362 (N_28362,N_23549,N_20043);
or U28363 (N_28363,N_20406,N_23294);
nor U28364 (N_28364,N_22964,N_21869);
xor U28365 (N_28365,N_21856,N_22885);
and U28366 (N_28366,N_22462,N_23258);
nor U28367 (N_28367,N_24932,N_24987);
nor U28368 (N_28368,N_21836,N_23387);
and U28369 (N_28369,N_22351,N_20643);
or U28370 (N_28370,N_22247,N_20452);
or U28371 (N_28371,N_22033,N_22258);
or U28372 (N_28372,N_21086,N_23393);
and U28373 (N_28373,N_20764,N_23246);
and U28374 (N_28374,N_21052,N_23099);
xnor U28375 (N_28375,N_20105,N_21290);
nand U28376 (N_28376,N_21085,N_22214);
or U28377 (N_28377,N_22247,N_22988);
or U28378 (N_28378,N_24870,N_22555);
or U28379 (N_28379,N_22112,N_21285);
nand U28380 (N_28380,N_20758,N_21604);
nand U28381 (N_28381,N_21068,N_23149);
nand U28382 (N_28382,N_23883,N_21753);
and U28383 (N_28383,N_20362,N_20146);
nand U28384 (N_28384,N_22072,N_23620);
nor U28385 (N_28385,N_21092,N_24290);
and U28386 (N_28386,N_20708,N_21376);
xor U28387 (N_28387,N_20043,N_20506);
and U28388 (N_28388,N_24378,N_21013);
nand U28389 (N_28389,N_21472,N_22336);
xor U28390 (N_28390,N_23778,N_20952);
and U28391 (N_28391,N_23022,N_22833);
nand U28392 (N_28392,N_24612,N_24233);
xor U28393 (N_28393,N_24516,N_23975);
or U28394 (N_28394,N_22954,N_24353);
nand U28395 (N_28395,N_24423,N_20105);
or U28396 (N_28396,N_24111,N_24691);
nor U28397 (N_28397,N_23469,N_24370);
nor U28398 (N_28398,N_20208,N_20470);
nand U28399 (N_28399,N_24678,N_20823);
and U28400 (N_28400,N_24943,N_22337);
nand U28401 (N_28401,N_21655,N_24896);
nand U28402 (N_28402,N_21038,N_21387);
nor U28403 (N_28403,N_21070,N_20258);
xnor U28404 (N_28404,N_22237,N_24007);
nor U28405 (N_28405,N_24248,N_23462);
or U28406 (N_28406,N_24738,N_23612);
xnor U28407 (N_28407,N_21005,N_21457);
or U28408 (N_28408,N_20725,N_23937);
nor U28409 (N_28409,N_23990,N_24024);
nor U28410 (N_28410,N_24846,N_23140);
nand U28411 (N_28411,N_21111,N_23804);
and U28412 (N_28412,N_23567,N_23417);
and U28413 (N_28413,N_21592,N_22738);
nand U28414 (N_28414,N_21400,N_22779);
xnor U28415 (N_28415,N_24919,N_21225);
or U28416 (N_28416,N_20059,N_24218);
nand U28417 (N_28417,N_21865,N_22146);
or U28418 (N_28418,N_20696,N_24419);
and U28419 (N_28419,N_24736,N_20788);
nand U28420 (N_28420,N_22485,N_22495);
nor U28421 (N_28421,N_24201,N_21503);
and U28422 (N_28422,N_24564,N_24041);
nand U28423 (N_28423,N_23459,N_22535);
nand U28424 (N_28424,N_23749,N_24782);
and U28425 (N_28425,N_24782,N_21539);
or U28426 (N_28426,N_23378,N_24394);
xnor U28427 (N_28427,N_24304,N_22377);
nand U28428 (N_28428,N_23725,N_23957);
and U28429 (N_28429,N_21034,N_23811);
nor U28430 (N_28430,N_21782,N_21978);
nor U28431 (N_28431,N_22848,N_23895);
or U28432 (N_28432,N_24583,N_21073);
nor U28433 (N_28433,N_20460,N_22662);
xor U28434 (N_28434,N_22062,N_24498);
and U28435 (N_28435,N_23895,N_23298);
nand U28436 (N_28436,N_23090,N_20254);
or U28437 (N_28437,N_23330,N_21577);
nand U28438 (N_28438,N_23002,N_23556);
nand U28439 (N_28439,N_23245,N_22050);
nor U28440 (N_28440,N_22206,N_20860);
nor U28441 (N_28441,N_20264,N_20686);
or U28442 (N_28442,N_23519,N_24911);
or U28443 (N_28443,N_21292,N_22843);
xnor U28444 (N_28444,N_20329,N_23845);
nand U28445 (N_28445,N_21685,N_20784);
and U28446 (N_28446,N_24669,N_22116);
and U28447 (N_28447,N_20487,N_20730);
xnor U28448 (N_28448,N_21402,N_22656);
nand U28449 (N_28449,N_23808,N_24167);
nand U28450 (N_28450,N_22375,N_23669);
nand U28451 (N_28451,N_22870,N_24757);
and U28452 (N_28452,N_21816,N_21691);
or U28453 (N_28453,N_21828,N_20952);
nor U28454 (N_28454,N_20370,N_24919);
nand U28455 (N_28455,N_21176,N_23462);
or U28456 (N_28456,N_20073,N_24339);
or U28457 (N_28457,N_20459,N_21024);
nor U28458 (N_28458,N_24944,N_22343);
nand U28459 (N_28459,N_24297,N_23982);
nor U28460 (N_28460,N_20438,N_22711);
nand U28461 (N_28461,N_20036,N_23623);
xnor U28462 (N_28462,N_21929,N_24265);
nor U28463 (N_28463,N_24190,N_24733);
or U28464 (N_28464,N_20732,N_22134);
or U28465 (N_28465,N_24005,N_21020);
nand U28466 (N_28466,N_23908,N_21882);
nor U28467 (N_28467,N_22120,N_23584);
nand U28468 (N_28468,N_24640,N_21982);
nor U28469 (N_28469,N_24286,N_21750);
nand U28470 (N_28470,N_23617,N_23925);
xor U28471 (N_28471,N_23412,N_23980);
nor U28472 (N_28472,N_20366,N_21754);
or U28473 (N_28473,N_21068,N_24375);
or U28474 (N_28474,N_23462,N_22763);
nor U28475 (N_28475,N_24526,N_24118);
nor U28476 (N_28476,N_22941,N_21998);
or U28477 (N_28477,N_22972,N_22199);
and U28478 (N_28478,N_21467,N_21235);
nor U28479 (N_28479,N_24768,N_23376);
nor U28480 (N_28480,N_24735,N_24418);
xnor U28481 (N_28481,N_21221,N_20000);
and U28482 (N_28482,N_21272,N_23240);
and U28483 (N_28483,N_23176,N_21241);
xnor U28484 (N_28484,N_21342,N_23303);
nand U28485 (N_28485,N_21558,N_21771);
or U28486 (N_28486,N_21601,N_22885);
and U28487 (N_28487,N_22846,N_23873);
or U28488 (N_28488,N_23909,N_23615);
nor U28489 (N_28489,N_23434,N_20346);
nor U28490 (N_28490,N_20648,N_21722);
nand U28491 (N_28491,N_23594,N_23563);
xor U28492 (N_28492,N_21934,N_22086);
or U28493 (N_28493,N_24804,N_20524);
or U28494 (N_28494,N_22107,N_21467);
xnor U28495 (N_28495,N_23013,N_24306);
nor U28496 (N_28496,N_20134,N_23364);
and U28497 (N_28497,N_23631,N_21688);
nor U28498 (N_28498,N_20586,N_20636);
nand U28499 (N_28499,N_20791,N_24028);
nor U28500 (N_28500,N_21957,N_21757);
nor U28501 (N_28501,N_20499,N_20401);
and U28502 (N_28502,N_24819,N_22173);
nor U28503 (N_28503,N_23957,N_23366);
or U28504 (N_28504,N_21733,N_24137);
and U28505 (N_28505,N_20155,N_22556);
or U28506 (N_28506,N_22692,N_24154);
xor U28507 (N_28507,N_21990,N_20468);
or U28508 (N_28508,N_23234,N_21587);
nor U28509 (N_28509,N_22238,N_20145);
or U28510 (N_28510,N_20286,N_20392);
nor U28511 (N_28511,N_24919,N_24253);
and U28512 (N_28512,N_23760,N_20318);
xnor U28513 (N_28513,N_24907,N_21108);
xor U28514 (N_28514,N_23818,N_22213);
or U28515 (N_28515,N_21984,N_23115);
xnor U28516 (N_28516,N_20067,N_23995);
and U28517 (N_28517,N_24388,N_21428);
nand U28518 (N_28518,N_20922,N_22694);
nand U28519 (N_28519,N_20841,N_24309);
or U28520 (N_28520,N_23278,N_23924);
and U28521 (N_28521,N_20621,N_21098);
or U28522 (N_28522,N_20838,N_20158);
and U28523 (N_28523,N_24463,N_21836);
or U28524 (N_28524,N_22069,N_22588);
xnor U28525 (N_28525,N_20892,N_20050);
nor U28526 (N_28526,N_22335,N_24914);
nor U28527 (N_28527,N_22723,N_21739);
nand U28528 (N_28528,N_20680,N_22337);
or U28529 (N_28529,N_21903,N_21124);
nor U28530 (N_28530,N_24383,N_22026);
or U28531 (N_28531,N_24453,N_23953);
nor U28532 (N_28532,N_20515,N_22976);
nand U28533 (N_28533,N_23404,N_24423);
and U28534 (N_28534,N_20890,N_24845);
nand U28535 (N_28535,N_24110,N_20936);
nand U28536 (N_28536,N_20614,N_24038);
or U28537 (N_28537,N_23996,N_23940);
nand U28538 (N_28538,N_23563,N_20994);
nand U28539 (N_28539,N_20931,N_20863);
or U28540 (N_28540,N_20676,N_21624);
or U28541 (N_28541,N_24383,N_22347);
nor U28542 (N_28542,N_24453,N_20314);
nand U28543 (N_28543,N_22744,N_20989);
nand U28544 (N_28544,N_22329,N_20877);
nor U28545 (N_28545,N_22153,N_24430);
and U28546 (N_28546,N_23476,N_20063);
or U28547 (N_28547,N_20378,N_21471);
or U28548 (N_28548,N_20162,N_22780);
or U28549 (N_28549,N_23705,N_22867);
nand U28550 (N_28550,N_21435,N_24736);
or U28551 (N_28551,N_22900,N_22523);
and U28552 (N_28552,N_23720,N_21090);
nand U28553 (N_28553,N_20400,N_24663);
nand U28554 (N_28554,N_24947,N_23924);
nand U28555 (N_28555,N_20020,N_24462);
nand U28556 (N_28556,N_21968,N_23202);
nor U28557 (N_28557,N_21050,N_20646);
nor U28558 (N_28558,N_21226,N_24558);
nor U28559 (N_28559,N_20842,N_21334);
nor U28560 (N_28560,N_20209,N_21001);
and U28561 (N_28561,N_24045,N_24088);
nor U28562 (N_28562,N_20080,N_23521);
or U28563 (N_28563,N_22050,N_23908);
and U28564 (N_28564,N_22375,N_21517);
and U28565 (N_28565,N_20032,N_24549);
or U28566 (N_28566,N_23891,N_22356);
nand U28567 (N_28567,N_20025,N_21273);
or U28568 (N_28568,N_23136,N_20485);
or U28569 (N_28569,N_24388,N_23886);
xor U28570 (N_28570,N_21572,N_21095);
nor U28571 (N_28571,N_21360,N_21425);
nor U28572 (N_28572,N_23501,N_21654);
or U28573 (N_28573,N_23311,N_22789);
nor U28574 (N_28574,N_22781,N_22958);
nor U28575 (N_28575,N_20095,N_21849);
and U28576 (N_28576,N_22417,N_23142);
xor U28577 (N_28577,N_22501,N_21815);
nand U28578 (N_28578,N_23671,N_24712);
or U28579 (N_28579,N_24745,N_20728);
nand U28580 (N_28580,N_20385,N_24990);
or U28581 (N_28581,N_21745,N_23174);
and U28582 (N_28582,N_24881,N_21746);
nor U28583 (N_28583,N_24151,N_22615);
nor U28584 (N_28584,N_22962,N_24961);
nand U28585 (N_28585,N_21401,N_20228);
xor U28586 (N_28586,N_23816,N_22317);
xnor U28587 (N_28587,N_20256,N_20316);
nor U28588 (N_28588,N_20595,N_24944);
nor U28589 (N_28589,N_24601,N_23234);
or U28590 (N_28590,N_24070,N_24637);
nand U28591 (N_28591,N_20594,N_20268);
and U28592 (N_28592,N_21889,N_24475);
or U28593 (N_28593,N_23702,N_20515);
xor U28594 (N_28594,N_22137,N_23344);
and U28595 (N_28595,N_24713,N_24289);
or U28596 (N_28596,N_24891,N_20408);
nor U28597 (N_28597,N_20460,N_24148);
nand U28598 (N_28598,N_20566,N_22911);
xnor U28599 (N_28599,N_21335,N_20203);
and U28600 (N_28600,N_20084,N_23207);
and U28601 (N_28601,N_20557,N_20445);
or U28602 (N_28602,N_22418,N_24967);
or U28603 (N_28603,N_22656,N_20667);
nand U28604 (N_28604,N_20329,N_24862);
or U28605 (N_28605,N_20986,N_21586);
nand U28606 (N_28606,N_21331,N_24079);
and U28607 (N_28607,N_21861,N_21289);
or U28608 (N_28608,N_22586,N_24729);
nand U28609 (N_28609,N_24169,N_20408);
nand U28610 (N_28610,N_21695,N_22858);
and U28611 (N_28611,N_23589,N_24970);
nor U28612 (N_28612,N_23058,N_20968);
or U28613 (N_28613,N_20788,N_21788);
and U28614 (N_28614,N_24811,N_22939);
nand U28615 (N_28615,N_24061,N_20748);
and U28616 (N_28616,N_21900,N_23543);
nor U28617 (N_28617,N_20170,N_21100);
or U28618 (N_28618,N_21224,N_22148);
and U28619 (N_28619,N_23075,N_24859);
and U28620 (N_28620,N_20251,N_24430);
and U28621 (N_28621,N_24018,N_22377);
nand U28622 (N_28622,N_22149,N_23930);
nand U28623 (N_28623,N_22580,N_24854);
nor U28624 (N_28624,N_24272,N_21206);
nand U28625 (N_28625,N_22287,N_21230);
and U28626 (N_28626,N_22443,N_22144);
and U28627 (N_28627,N_20614,N_23898);
nand U28628 (N_28628,N_22849,N_23608);
nor U28629 (N_28629,N_24381,N_22568);
nor U28630 (N_28630,N_21634,N_20005);
and U28631 (N_28631,N_20835,N_23791);
nand U28632 (N_28632,N_23871,N_20874);
xnor U28633 (N_28633,N_20698,N_24116);
nor U28634 (N_28634,N_20196,N_24572);
nand U28635 (N_28635,N_24041,N_20671);
xor U28636 (N_28636,N_22225,N_24365);
or U28637 (N_28637,N_24818,N_21268);
nand U28638 (N_28638,N_23919,N_20167);
nor U28639 (N_28639,N_22228,N_22060);
nand U28640 (N_28640,N_20608,N_21071);
nand U28641 (N_28641,N_24582,N_23936);
or U28642 (N_28642,N_21227,N_22285);
and U28643 (N_28643,N_24106,N_24400);
and U28644 (N_28644,N_23832,N_20565);
nand U28645 (N_28645,N_24370,N_20614);
nand U28646 (N_28646,N_21600,N_24887);
and U28647 (N_28647,N_20849,N_24606);
nand U28648 (N_28648,N_21622,N_24813);
xor U28649 (N_28649,N_21731,N_23570);
nor U28650 (N_28650,N_20669,N_23131);
nand U28651 (N_28651,N_22051,N_23745);
or U28652 (N_28652,N_20541,N_20818);
or U28653 (N_28653,N_23004,N_21935);
xor U28654 (N_28654,N_20580,N_22644);
or U28655 (N_28655,N_21806,N_24881);
xor U28656 (N_28656,N_22016,N_24824);
nor U28657 (N_28657,N_22108,N_24871);
or U28658 (N_28658,N_21378,N_22765);
or U28659 (N_28659,N_21533,N_20017);
nand U28660 (N_28660,N_24736,N_23768);
nor U28661 (N_28661,N_23291,N_20495);
nand U28662 (N_28662,N_20573,N_20047);
nand U28663 (N_28663,N_23438,N_23053);
nand U28664 (N_28664,N_22587,N_23851);
nand U28665 (N_28665,N_23032,N_23322);
nand U28666 (N_28666,N_22241,N_24905);
nor U28667 (N_28667,N_24239,N_22719);
nor U28668 (N_28668,N_24905,N_23425);
or U28669 (N_28669,N_20843,N_21705);
or U28670 (N_28670,N_22824,N_24694);
nor U28671 (N_28671,N_20876,N_22551);
or U28672 (N_28672,N_21485,N_24460);
nand U28673 (N_28673,N_21265,N_22853);
nor U28674 (N_28674,N_21624,N_23619);
nand U28675 (N_28675,N_21490,N_24693);
and U28676 (N_28676,N_24758,N_22825);
nand U28677 (N_28677,N_24574,N_21650);
nand U28678 (N_28678,N_21748,N_23827);
nor U28679 (N_28679,N_20447,N_23437);
or U28680 (N_28680,N_22657,N_21042);
nand U28681 (N_28681,N_24592,N_22236);
xnor U28682 (N_28682,N_21919,N_23715);
or U28683 (N_28683,N_22876,N_20404);
or U28684 (N_28684,N_23123,N_24430);
xor U28685 (N_28685,N_24952,N_20440);
nor U28686 (N_28686,N_23396,N_21251);
nor U28687 (N_28687,N_20381,N_20516);
nand U28688 (N_28688,N_23891,N_23374);
nor U28689 (N_28689,N_20904,N_24015);
nand U28690 (N_28690,N_20843,N_22896);
nor U28691 (N_28691,N_22203,N_21745);
or U28692 (N_28692,N_24894,N_22111);
xnor U28693 (N_28693,N_23551,N_22976);
nand U28694 (N_28694,N_22522,N_22146);
or U28695 (N_28695,N_24343,N_23421);
and U28696 (N_28696,N_23191,N_22668);
or U28697 (N_28697,N_23169,N_21739);
nor U28698 (N_28698,N_21284,N_20887);
nor U28699 (N_28699,N_21258,N_24504);
or U28700 (N_28700,N_24840,N_23303);
and U28701 (N_28701,N_23958,N_22862);
or U28702 (N_28702,N_23377,N_20238);
nand U28703 (N_28703,N_23766,N_22086);
and U28704 (N_28704,N_22758,N_23733);
and U28705 (N_28705,N_20191,N_22539);
nand U28706 (N_28706,N_23128,N_20636);
and U28707 (N_28707,N_21568,N_21992);
nand U28708 (N_28708,N_23812,N_20185);
nand U28709 (N_28709,N_20638,N_21444);
and U28710 (N_28710,N_22687,N_24126);
nand U28711 (N_28711,N_24755,N_24957);
nor U28712 (N_28712,N_21522,N_24779);
and U28713 (N_28713,N_24591,N_23212);
and U28714 (N_28714,N_24196,N_23411);
nor U28715 (N_28715,N_24898,N_21647);
or U28716 (N_28716,N_24158,N_23625);
or U28717 (N_28717,N_24278,N_23069);
or U28718 (N_28718,N_22870,N_22553);
and U28719 (N_28719,N_23918,N_22235);
or U28720 (N_28720,N_21106,N_20171);
or U28721 (N_28721,N_23981,N_22227);
xor U28722 (N_28722,N_21489,N_24908);
or U28723 (N_28723,N_22837,N_22817);
or U28724 (N_28724,N_20994,N_24726);
nand U28725 (N_28725,N_22942,N_22279);
nand U28726 (N_28726,N_23074,N_23150);
or U28727 (N_28727,N_20613,N_24506);
nand U28728 (N_28728,N_23607,N_20743);
nor U28729 (N_28729,N_20475,N_22003);
xnor U28730 (N_28730,N_23816,N_21405);
nand U28731 (N_28731,N_20123,N_21371);
nor U28732 (N_28732,N_21721,N_23442);
and U28733 (N_28733,N_23878,N_23580);
nand U28734 (N_28734,N_24543,N_23255);
nor U28735 (N_28735,N_21419,N_22705);
or U28736 (N_28736,N_20210,N_24930);
or U28737 (N_28737,N_22427,N_22767);
nor U28738 (N_28738,N_21080,N_22913);
nor U28739 (N_28739,N_24608,N_23701);
and U28740 (N_28740,N_22511,N_20085);
nand U28741 (N_28741,N_21922,N_20146);
nor U28742 (N_28742,N_24174,N_21169);
nor U28743 (N_28743,N_22733,N_22858);
or U28744 (N_28744,N_24100,N_20616);
nor U28745 (N_28745,N_21552,N_20362);
and U28746 (N_28746,N_21810,N_24860);
or U28747 (N_28747,N_22852,N_20283);
and U28748 (N_28748,N_22247,N_22901);
and U28749 (N_28749,N_22119,N_20754);
nor U28750 (N_28750,N_23271,N_22486);
or U28751 (N_28751,N_23950,N_23989);
nor U28752 (N_28752,N_20748,N_21124);
or U28753 (N_28753,N_23313,N_23834);
nor U28754 (N_28754,N_21773,N_20260);
and U28755 (N_28755,N_24189,N_24795);
nor U28756 (N_28756,N_20081,N_23791);
nor U28757 (N_28757,N_24990,N_23346);
xor U28758 (N_28758,N_22634,N_22955);
nor U28759 (N_28759,N_23426,N_22809);
and U28760 (N_28760,N_21413,N_24792);
nand U28761 (N_28761,N_24554,N_24507);
and U28762 (N_28762,N_21727,N_23864);
nand U28763 (N_28763,N_21170,N_22102);
xnor U28764 (N_28764,N_21952,N_23783);
or U28765 (N_28765,N_21274,N_20733);
nand U28766 (N_28766,N_24598,N_24343);
and U28767 (N_28767,N_20841,N_24562);
or U28768 (N_28768,N_24330,N_24858);
or U28769 (N_28769,N_22726,N_23269);
or U28770 (N_28770,N_20564,N_20456);
and U28771 (N_28771,N_24626,N_23916);
and U28772 (N_28772,N_22711,N_22051);
nand U28773 (N_28773,N_23456,N_23126);
or U28774 (N_28774,N_22656,N_20257);
nand U28775 (N_28775,N_21474,N_20980);
or U28776 (N_28776,N_20433,N_20842);
or U28777 (N_28777,N_22008,N_24536);
xor U28778 (N_28778,N_22797,N_24724);
nand U28779 (N_28779,N_21371,N_22869);
nand U28780 (N_28780,N_22982,N_21451);
and U28781 (N_28781,N_24305,N_20875);
and U28782 (N_28782,N_23962,N_24521);
or U28783 (N_28783,N_23125,N_24150);
nand U28784 (N_28784,N_23623,N_22191);
and U28785 (N_28785,N_22415,N_22192);
nor U28786 (N_28786,N_20000,N_21054);
nor U28787 (N_28787,N_20186,N_20987);
or U28788 (N_28788,N_22473,N_22384);
and U28789 (N_28789,N_24757,N_22915);
and U28790 (N_28790,N_23530,N_23059);
xnor U28791 (N_28791,N_21866,N_22846);
and U28792 (N_28792,N_21097,N_21756);
xnor U28793 (N_28793,N_22249,N_21563);
xnor U28794 (N_28794,N_21450,N_23582);
and U28795 (N_28795,N_23815,N_21590);
and U28796 (N_28796,N_24017,N_23735);
and U28797 (N_28797,N_24934,N_22750);
nor U28798 (N_28798,N_21666,N_20124);
or U28799 (N_28799,N_23335,N_20405);
and U28800 (N_28800,N_22079,N_20761);
nand U28801 (N_28801,N_20902,N_22022);
or U28802 (N_28802,N_24442,N_20297);
nand U28803 (N_28803,N_23475,N_23337);
xor U28804 (N_28804,N_20026,N_24105);
nor U28805 (N_28805,N_22239,N_22766);
or U28806 (N_28806,N_24877,N_22043);
or U28807 (N_28807,N_24433,N_23625);
nor U28808 (N_28808,N_24596,N_22816);
nor U28809 (N_28809,N_20510,N_22503);
xnor U28810 (N_28810,N_22233,N_20424);
or U28811 (N_28811,N_21839,N_21003);
xor U28812 (N_28812,N_23123,N_23489);
nand U28813 (N_28813,N_22326,N_24207);
nor U28814 (N_28814,N_20876,N_22758);
nand U28815 (N_28815,N_21722,N_24136);
or U28816 (N_28816,N_23133,N_20107);
or U28817 (N_28817,N_20520,N_22027);
nor U28818 (N_28818,N_21637,N_24314);
nand U28819 (N_28819,N_22307,N_24804);
and U28820 (N_28820,N_22063,N_24562);
nor U28821 (N_28821,N_20619,N_20013);
or U28822 (N_28822,N_24335,N_22458);
nor U28823 (N_28823,N_22541,N_20826);
and U28824 (N_28824,N_21479,N_20647);
or U28825 (N_28825,N_20590,N_22728);
nand U28826 (N_28826,N_24616,N_21162);
xor U28827 (N_28827,N_23843,N_20370);
nor U28828 (N_28828,N_22668,N_20031);
nand U28829 (N_28829,N_24661,N_23217);
and U28830 (N_28830,N_24398,N_20939);
or U28831 (N_28831,N_23653,N_24622);
or U28832 (N_28832,N_22839,N_23344);
nand U28833 (N_28833,N_23715,N_21362);
and U28834 (N_28834,N_23498,N_20977);
or U28835 (N_28835,N_21863,N_23196);
or U28836 (N_28836,N_20909,N_21187);
nor U28837 (N_28837,N_21853,N_20923);
xnor U28838 (N_28838,N_23345,N_24184);
or U28839 (N_28839,N_22832,N_21944);
nand U28840 (N_28840,N_24338,N_22685);
nor U28841 (N_28841,N_21404,N_24491);
or U28842 (N_28842,N_24117,N_22294);
or U28843 (N_28843,N_20340,N_24648);
or U28844 (N_28844,N_23193,N_20609);
nand U28845 (N_28845,N_23400,N_24284);
or U28846 (N_28846,N_21484,N_23112);
nand U28847 (N_28847,N_22550,N_22291);
nor U28848 (N_28848,N_23528,N_23040);
and U28849 (N_28849,N_23936,N_23673);
nand U28850 (N_28850,N_22008,N_21372);
or U28851 (N_28851,N_23505,N_23325);
nor U28852 (N_28852,N_20342,N_21529);
or U28853 (N_28853,N_24907,N_20774);
xnor U28854 (N_28854,N_20935,N_22601);
and U28855 (N_28855,N_24980,N_22538);
and U28856 (N_28856,N_24387,N_22030);
nor U28857 (N_28857,N_21852,N_24649);
and U28858 (N_28858,N_23568,N_23310);
nor U28859 (N_28859,N_21584,N_24805);
nand U28860 (N_28860,N_21944,N_23024);
nand U28861 (N_28861,N_21627,N_24730);
and U28862 (N_28862,N_24875,N_22437);
nand U28863 (N_28863,N_23727,N_22142);
nand U28864 (N_28864,N_24494,N_21632);
nand U28865 (N_28865,N_21752,N_24232);
nor U28866 (N_28866,N_20983,N_24917);
nand U28867 (N_28867,N_22218,N_24080);
nor U28868 (N_28868,N_24460,N_24209);
nor U28869 (N_28869,N_20082,N_22711);
or U28870 (N_28870,N_23465,N_24557);
xnor U28871 (N_28871,N_24850,N_20786);
and U28872 (N_28872,N_22849,N_20534);
xor U28873 (N_28873,N_24092,N_24838);
and U28874 (N_28874,N_21323,N_22732);
xor U28875 (N_28875,N_24705,N_20372);
xor U28876 (N_28876,N_22332,N_22789);
and U28877 (N_28877,N_24173,N_20378);
and U28878 (N_28878,N_20445,N_22951);
and U28879 (N_28879,N_20277,N_22841);
or U28880 (N_28880,N_24543,N_22664);
and U28881 (N_28881,N_21427,N_24240);
nand U28882 (N_28882,N_21304,N_23255);
or U28883 (N_28883,N_22515,N_24385);
or U28884 (N_28884,N_24302,N_24552);
or U28885 (N_28885,N_21125,N_24583);
and U28886 (N_28886,N_21223,N_21723);
and U28887 (N_28887,N_24440,N_24107);
or U28888 (N_28888,N_20107,N_22694);
nand U28889 (N_28889,N_23364,N_24867);
or U28890 (N_28890,N_22546,N_23460);
nor U28891 (N_28891,N_23506,N_23937);
nor U28892 (N_28892,N_20308,N_21090);
or U28893 (N_28893,N_23056,N_20543);
or U28894 (N_28894,N_22214,N_20813);
nand U28895 (N_28895,N_21485,N_24640);
nand U28896 (N_28896,N_24864,N_22613);
xor U28897 (N_28897,N_23793,N_21393);
or U28898 (N_28898,N_22034,N_20998);
or U28899 (N_28899,N_20323,N_24963);
nand U28900 (N_28900,N_20757,N_22612);
and U28901 (N_28901,N_24219,N_24964);
or U28902 (N_28902,N_23641,N_24993);
xor U28903 (N_28903,N_22406,N_24057);
xnor U28904 (N_28904,N_21120,N_23205);
or U28905 (N_28905,N_24686,N_23849);
and U28906 (N_28906,N_21303,N_23859);
xnor U28907 (N_28907,N_22189,N_20664);
nor U28908 (N_28908,N_21642,N_23401);
or U28909 (N_28909,N_23620,N_22916);
xor U28910 (N_28910,N_23559,N_20336);
nand U28911 (N_28911,N_22415,N_22508);
nand U28912 (N_28912,N_22988,N_20584);
or U28913 (N_28913,N_20825,N_20805);
and U28914 (N_28914,N_21251,N_24124);
and U28915 (N_28915,N_23027,N_23280);
nand U28916 (N_28916,N_22432,N_21293);
or U28917 (N_28917,N_21843,N_24711);
and U28918 (N_28918,N_22919,N_23907);
and U28919 (N_28919,N_21615,N_24082);
or U28920 (N_28920,N_20563,N_23443);
or U28921 (N_28921,N_21267,N_21971);
xor U28922 (N_28922,N_24433,N_23712);
and U28923 (N_28923,N_23251,N_24488);
and U28924 (N_28924,N_24877,N_21380);
xor U28925 (N_28925,N_22711,N_21320);
nand U28926 (N_28926,N_22552,N_23593);
nand U28927 (N_28927,N_24041,N_22066);
and U28928 (N_28928,N_20257,N_22001);
nand U28929 (N_28929,N_22405,N_20372);
nand U28930 (N_28930,N_20071,N_23173);
nor U28931 (N_28931,N_22316,N_22235);
nand U28932 (N_28932,N_21352,N_24185);
nor U28933 (N_28933,N_22716,N_21795);
and U28934 (N_28934,N_20146,N_24217);
and U28935 (N_28935,N_21835,N_22834);
xnor U28936 (N_28936,N_21160,N_20712);
or U28937 (N_28937,N_23689,N_24825);
xnor U28938 (N_28938,N_24917,N_21414);
or U28939 (N_28939,N_20624,N_23772);
nor U28940 (N_28940,N_20674,N_22122);
nand U28941 (N_28941,N_22242,N_23449);
or U28942 (N_28942,N_23121,N_21665);
nand U28943 (N_28943,N_20148,N_24193);
nor U28944 (N_28944,N_24615,N_23287);
nand U28945 (N_28945,N_22554,N_20293);
or U28946 (N_28946,N_21697,N_21616);
nor U28947 (N_28947,N_20229,N_24909);
xnor U28948 (N_28948,N_21196,N_23685);
nor U28949 (N_28949,N_21569,N_22868);
or U28950 (N_28950,N_20882,N_21632);
or U28951 (N_28951,N_21919,N_24796);
nand U28952 (N_28952,N_20237,N_21715);
nand U28953 (N_28953,N_22756,N_23395);
nor U28954 (N_28954,N_23342,N_21626);
nand U28955 (N_28955,N_22452,N_21358);
xnor U28956 (N_28956,N_21090,N_21460);
nor U28957 (N_28957,N_21938,N_24343);
nor U28958 (N_28958,N_20658,N_23234);
or U28959 (N_28959,N_21738,N_23505);
or U28960 (N_28960,N_21069,N_20070);
and U28961 (N_28961,N_23617,N_23411);
or U28962 (N_28962,N_23910,N_20543);
nor U28963 (N_28963,N_24900,N_23165);
or U28964 (N_28964,N_23316,N_22662);
and U28965 (N_28965,N_24615,N_23772);
xor U28966 (N_28966,N_21833,N_24661);
xnor U28967 (N_28967,N_24194,N_23412);
nand U28968 (N_28968,N_24751,N_24499);
nor U28969 (N_28969,N_23336,N_24594);
and U28970 (N_28970,N_22141,N_21732);
or U28971 (N_28971,N_20272,N_23080);
and U28972 (N_28972,N_20671,N_22631);
nor U28973 (N_28973,N_22077,N_22830);
or U28974 (N_28974,N_23962,N_23717);
nand U28975 (N_28975,N_22408,N_22848);
and U28976 (N_28976,N_20742,N_23848);
nor U28977 (N_28977,N_22014,N_21356);
nor U28978 (N_28978,N_23836,N_20442);
or U28979 (N_28979,N_23715,N_24441);
xor U28980 (N_28980,N_21105,N_21040);
nand U28981 (N_28981,N_20787,N_20413);
nor U28982 (N_28982,N_20196,N_22404);
nor U28983 (N_28983,N_21029,N_22637);
and U28984 (N_28984,N_20412,N_20063);
or U28985 (N_28985,N_20353,N_22629);
nand U28986 (N_28986,N_24731,N_21614);
and U28987 (N_28987,N_24618,N_24881);
and U28988 (N_28988,N_20368,N_24900);
nor U28989 (N_28989,N_21376,N_21065);
nor U28990 (N_28990,N_23307,N_22565);
nand U28991 (N_28991,N_21791,N_23502);
and U28992 (N_28992,N_24254,N_21607);
or U28993 (N_28993,N_21596,N_23582);
xnor U28994 (N_28994,N_21052,N_22226);
and U28995 (N_28995,N_21594,N_22492);
nand U28996 (N_28996,N_22304,N_23800);
nor U28997 (N_28997,N_20464,N_21387);
and U28998 (N_28998,N_22677,N_23134);
or U28999 (N_28999,N_23058,N_24973);
nand U29000 (N_29000,N_21006,N_20336);
or U29001 (N_29001,N_23479,N_20702);
and U29002 (N_29002,N_20622,N_22549);
and U29003 (N_29003,N_22614,N_22976);
and U29004 (N_29004,N_20631,N_24646);
or U29005 (N_29005,N_20506,N_21113);
or U29006 (N_29006,N_21887,N_22420);
xor U29007 (N_29007,N_21689,N_22997);
and U29008 (N_29008,N_23803,N_21371);
nand U29009 (N_29009,N_20778,N_20368);
or U29010 (N_29010,N_20281,N_24499);
or U29011 (N_29011,N_23087,N_21980);
nor U29012 (N_29012,N_23477,N_23123);
nor U29013 (N_29013,N_21350,N_20494);
or U29014 (N_29014,N_23322,N_21528);
or U29015 (N_29015,N_24037,N_23908);
or U29016 (N_29016,N_22586,N_21079);
and U29017 (N_29017,N_20455,N_20503);
nor U29018 (N_29018,N_22940,N_24814);
or U29019 (N_29019,N_20667,N_21010);
xnor U29020 (N_29020,N_23691,N_21904);
nor U29021 (N_29021,N_23329,N_23333);
nor U29022 (N_29022,N_20775,N_24372);
xnor U29023 (N_29023,N_21995,N_20619);
xnor U29024 (N_29024,N_24237,N_23034);
or U29025 (N_29025,N_24727,N_24332);
nand U29026 (N_29026,N_21163,N_22391);
and U29027 (N_29027,N_24331,N_20837);
nor U29028 (N_29028,N_23449,N_22442);
xnor U29029 (N_29029,N_24913,N_21916);
nor U29030 (N_29030,N_21722,N_20665);
nand U29031 (N_29031,N_20934,N_23673);
nor U29032 (N_29032,N_21661,N_21372);
or U29033 (N_29033,N_23154,N_20083);
nand U29034 (N_29034,N_21062,N_21203);
xnor U29035 (N_29035,N_23777,N_24618);
xnor U29036 (N_29036,N_21563,N_24002);
nor U29037 (N_29037,N_22788,N_20221);
nor U29038 (N_29038,N_22048,N_24842);
nand U29039 (N_29039,N_22859,N_24324);
nand U29040 (N_29040,N_20890,N_20018);
and U29041 (N_29041,N_21633,N_21388);
xor U29042 (N_29042,N_24321,N_24498);
or U29043 (N_29043,N_21603,N_20342);
nor U29044 (N_29044,N_20454,N_24708);
or U29045 (N_29045,N_22613,N_22417);
and U29046 (N_29046,N_22767,N_22291);
nor U29047 (N_29047,N_20600,N_21519);
nand U29048 (N_29048,N_23480,N_20729);
or U29049 (N_29049,N_21294,N_22133);
nor U29050 (N_29050,N_20344,N_23962);
nor U29051 (N_29051,N_21855,N_21581);
or U29052 (N_29052,N_24465,N_21359);
nor U29053 (N_29053,N_23252,N_23661);
and U29054 (N_29054,N_23627,N_23493);
nand U29055 (N_29055,N_20845,N_21070);
xnor U29056 (N_29056,N_20824,N_20854);
and U29057 (N_29057,N_23248,N_23672);
and U29058 (N_29058,N_21259,N_21537);
and U29059 (N_29059,N_21961,N_21300);
and U29060 (N_29060,N_23759,N_23520);
or U29061 (N_29061,N_20094,N_24852);
nor U29062 (N_29062,N_24232,N_23823);
or U29063 (N_29063,N_23836,N_21154);
nor U29064 (N_29064,N_24978,N_21073);
or U29065 (N_29065,N_23970,N_22781);
xnor U29066 (N_29066,N_20491,N_21353);
and U29067 (N_29067,N_21954,N_23548);
and U29068 (N_29068,N_21252,N_23596);
or U29069 (N_29069,N_24902,N_22875);
nand U29070 (N_29070,N_20968,N_24265);
nand U29071 (N_29071,N_24210,N_24902);
xor U29072 (N_29072,N_22288,N_20647);
nor U29073 (N_29073,N_20252,N_23164);
or U29074 (N_29074,N_23023,N_21975);
or U29075 (N_29075,N_20192,N_24191);
nand U29076 (N_29076,N_24532,N_22922);
nand U29077 (N_29077,N_21321,N_24936);
or U29078 (N_29078,N_23093,N_24309);
and U29079 (N_29079,N_21913,N_23897);
or U29080 (N_29080,N_20285,N_24428);
and U29081 (N_29081,N_21739,N_24574);
nor U29082 (N_29082,N_24099,N_22662);
nand U29083 (N_29083,N_21263,N_22976);
and U29084 (N_29084,N_21213,N_22741);
nand U29085 (N_29085,N_21647,N_20885);
and U29086 (N_29086,N_23177,N_23934);
and U29087 (N_29087,N_21886,N_23201);
xor U29088 (N_29088,N_22199,N_23444);
nor U29089 (N_29089,N_23130,N_20631);
or U29090 (N_29090,N_23485,N_23746);
and U29091 (N_29091,N_22883,N_21351);
and U29092 (N_29092,N_21616,N_20425);
xor U29093 (N_29093,N_20162,N_24865);
nor U29094 (N_29094,N_21315,N_21979);
xor U29095 (N_29095,N_20791,N_22925);
or U29096 (N_29096,N_23161,N_22074);
or U29097 (N_29097,N_23299,N_21335);
nand U29098 (N_29098,N_22061,N_22026);
or U29099 (N_29099,N_22798,N_21477);
nand U29100 (N_29100,N_24399,N_24181);
and U29101 (N_29101,N_21123,N_24657);
nor U29102 (N_29102,N_21896,N_24009);
or U29103 (N_29103,N_21115,N_20104);
and U29104 (N_29104,N_23183,N_20378);
nor U29105 (N_29105,N_20786,N_21479);
nand U29106 (N_29106,N_22622,N_20625);
and U29107 (N_29107,N_24645,N_23867);
nor U29108 (N_29108,N_23970,N_21829);
and U29109 (N_29109,N_24318,N_22090);
nor U29110 (N_29110,N_22022,N_20544);
and U29111 (N_29111,N_20489,N_21571);
nand U29112 (N_29112,N_21545,N_21160);
or U29113 (N_29113,N_20876,N_20274);
and U29114 (N_29114,N_22118,N_22754);
nor U29115 (N_29115,N_23700,N_22217);
nor U29116 (N_29116,N_21847,N_21838);
nand U29117 (N_29117,N_20683,N_24725);
nand U29118 (N_29118,N_23033,N_22979);
nand U29119 (N_29119,N_21626,N_24074);
and U29120 (N_29120,N_20685,N_24990);
xor U29121 (N_29121,N_23274,N_22989);
or U29122 (N_29122,N_23498,N_20457);
and U29123 (N_29123,N_20719,N_22202);
and U29124 (N_29124,N_22341,N_20828);
or U29125 (N_29125,N_24941,N_24418);
and U29126 (N_29126,N_20014,N_20269);
nand U29127 (N_29127,N_21348,N_23982);
or U29128 (N_29128,N_21981,N_22779);
nand U29129 (N_29129,N_21050,N_20689);
and U29130 (N_29130,N_20217,N_23905);
nand U29131 (N_29131,N_22127,N_22735);
nor U29132 (N_29132,N_20395,N_23708);
nor U29133 (N_29133,N_22586,N_21829);
nand U29134 (N_29134,N_21114,N_23540);
nor U29135 (N_29135,N_21404,N_20075);
and U29136 (N_29136,N_21360,N_21856);
nand U29137 (N_29137,N_24726,N_20080);
nand U29138 (N_29138,N_22811,N_22627);
or U29139 (N_29139,N_20279,N_20812);
nand U29140 (N_29140,N_24369,N_23073);
or U29141 (N_29141,N_20116,N_20825);
nand U29142 (N_29142,N_22426,N_22064);
and U29143 (N_29143,N_20440,N_23498);
or U29144 (N_29144,N_22249,N_20894);
nand U29145 (N_29145,N_23266,N_21363);
nor U29146 (N_29146,N_24201,N_20220);
nand U29147 (N_29147,N_24466,N_21814);
or U29148 (N_29148,N_22885,N_23213);
xnor U29149 (N_29149,N_20702,N_24347);
and U29150 (N_29150,N_23086,N_23175);
nor U29151 (N_29151,N_23013,N_20089);
nor U29152 (N_29152,N_21037,N_21793);
nor U29153 (N_29153,N_21849,N_21478);
nor U29154 (N_29154,N_21104,N_21532);
nand U29155 (N_29155,N_23028,N_24686);
or U29156 (N_29156,N_22958,N_20894);
nand U29157 (N_29157,N_21227,N_23109);
and U29158 (N_29158,N_24988,N_22492);
nor U29159 (N_29159,N_20294,N_20192);
nand U29160 (N_29160,N_23767,N_21117);
nand U29161 (N_29161,N_20827,N_22238);
nor U29162 (N_29162,N_21300,N_20266);
nor U29163 (N_29163,N_24426,N_24966);
or U29164 (N_29164,N_22873,N_23544);
and U29165 (N_29165,N_23149,N_24664);
nand U29166 (N_29166,N_20731,N_22889);
nand U29167 (N_29167,N_22685,N_23263);
nor U29168 (N_29168,N_20790,N_22918);
and U29169 (N_29169,N_20763,N_20741);
and U29170 (N_29170,N_24959,N_23308);
nor U29171 (N_29171,N_23110,N_23605);
nor U29172 (N_29172,N_23879,N_20528);
and U29173 (N_29173,N_21754,N_22597);
or U29174 (N_29174,N_20119,N_23142);
and U29175 (N_29175,N_24309,N_20890);
xnor U29176 (N_29176,N_20959,N_20411);
nor U29177 (N_29177,N_21181,N_22992);
or U29178 (N_29178,N_20633,N_22723);
nand U29179 (N_29179,N_20333,N_24676);
and U29180 (N_29180,N_21983,N_22075);
or U29181 (N_29181,N_23047,N_24885);
and U29182 (N_29182,N_24085,N_21581);
or U29183 (N_29183,N_22247,N_21972);
nor U29184 (N_29184,N_22085,N_23420);
nand U29185 (N_29185,N_22186,N_22224);
nand U29186 (N_29186,N_24126,N_21374);
or U29187 (N_29187,N_22879,N_22290);
nand U29188 (N_29188,N_20582,N_21995);
and U29189 (N_29189,N_20513,N_24901);
nand U29190 (N_29190,N_23294,N_24951);
or U29191 (N_29191,N_23075,N_21673);
xnor U29192 (N_29192,N_20396,N_21083);
and U29193 (N_29193,N_23531,N_21381);
and U29194 (N_29194,N_24337,N_24186);
nand U29195 (N_29195,N_20784,N_20550);
and U29196 (N_29196,N_24887,N_21155);
and U29197 (N_29197,N_21394,N_23693);
and U29198 (N_29198,N_22022,N_21805);
and U29199 (N_29199,N_24598,N_24433);
nor U29200 (N_29200,N_23794,N_21906);
nor U29201 (N_29201,N_21798,N_22969);
nand U29202 (N_29202,N_22741,N_24742);
nor U29203 (N_29203,N_24987,N_24753);
or U29204 (N_29204,N_24871,N_24608);
or U29205 (N_29205,N_24491,N_21257);
or U29206 (N_29206,N_22626,N_23556);
nand U29207 (N_29207,N_24258,N_23419);
or U29208 (N_29208,N_22841,N_21698);
nand U29209 (N_29209,N_22244,N_24928);
nand U29210 (N_29210,N_22732,N_21615);
nand U29211 (N_29211,N_23557,N_23870);
xnor U29212 (N_29212,N_20968,N_24794);
nor U29213 (N_29213,N_23038,N_21922);
and U29214 (N_29214,N_20078,N_24290);
or U29215 (N_29215,N_22806,N_23586);
and U29216 (N_29216,N_23807,N_21774);
or U29217 (N_29217,N_23992,N_20714);
and U29218 (N_29218,N_20136,N_22563);
or U29219 (N_29219,N_20801,N_20076);
and U29220 (N_29220,N_22299,N_22526);
nand U29221 (N_29221,N_21242,N_23702);
nor U29222 (N_29222,N_23200,N_22708);
xnor U29223 (N_29223,N_20738,N_23849);
nor U29224 (N_29224,N_20529,N_23202);
and U29225 (N_29225,N_24439,N_21247);
nor U29226 (N_29226,N_20716,N_22123);
nor U29227 (N_29227,N_21340,N_21190);
nand U29228 (N_29228,N_21746,N_23370);
nor U29229 (N_29229,N_21688,N_24276);
nor U29230 (N_29230,N_21733,N_21717);
nor U29231 (N_29231,N_24637,N_22137);
or U29232 (N_29232,N_22797,N_22100);
nand U29233 (N_29233,N_21186,N_21274);
nor U29234 (N_29234,N_23669,N_21615);
nand U29235 (N_29235,N_23547,N_24597);
nor U29236 (N_29236,N_21653,N_21867);
and U29237 (N_29237,N_24276,N_23940);
and U29238 (N_29238,N_20340,N_20919);
or U29239 (N_29239,N_24579,N_23222);
nand U29240 (N_29240,N_21509,N_23981);
nand U29241 (N_29241,N_23040,N_23084);
xor U29242 (N_29242,N_23585,N_21261);
or U29243 (N_29243,N_21969,N_24528);
and U29244 (N_29244,N_21658,N_21635);
nand U29245 (N_29245,N_22283,N_21194);
nand U29246 (N_29246,N_21862,N_22785);
nand U29247 (N_29247,N_20319,N_20264);
nand U29248 (N_29248,N_24095,N_24730);
or U29249 (N_29249,N_24751,N_20870);
or U29250 (N_29250,N_22859,N_22605);
nor U29251 (N_29251,N_24747,N_20861);
xnor U29252 (N_29252,N_20918,N_20936);
nor U29253 (N_29253,N_22650,N_22677);
nand U29254 (N_29254,N_24490,N_21359);
and U29255 (N_29255,N_23440,N_24503);
nand U29256 (N_29256,N_23692,N_20275);
nor U29257 (N_29257,N_21026,N_21919);
xor U29258 (N_29258,N_24767,N_23551);
nor U29259 (N_29259,N_20921,N_21591);
nand U29260 (N_29260,N_21272,N_21581);
nand U29261 (N_29261,N_21385,N_20415);
nand U29262 (N_29262,N_21321,N_23625);
nor U29263 (N_29263,N_23791,N_22567);
and U29264 (N_29264,N_20927,N_20009);
and U29265 (N_29265,N_20773,N_21868);
and U29266 (N_29266,N_22248,N_21804);
nand U29267 (N_29267,N_23477,N_22063);
xnor U29268 (N_29268,N_21481,N_24280);
nor U29269 (N_29269,N_22646,N_22699);
nand U29270 (N_29270,N_24071,N_24279);
xor U29271 (N_29271,N_24820,N_24647);
and U29272 (N_29272,N_20512,N_22831);
xnor U29273 (N_29273,N_24959,N_21535);
or U29274 (N_29274,N_23089,N_21321);
or U29275 (N_29275,N_23667,N_20614);
and U29276 (N_29276,N_24128,N_22929);
nand U29277 (N_29277,N_22971,N_20698);
or U29278 (N_29278,N_20074,N_23494);
nand U29279 (N_29279,N_24249,N_24725);
and U29280 (N_29280,N_20250,N_22038);
nand U29281 (N_29281,N_24222,N_20508);
and U29282 (N_29282,N_24469,N_20493);
nand U29283 (N_29283,N_20271,N_21438);
and U29284 (N_29284,N_20862,N_22991);
or U29285 (N_29285,N_23825,N_22862);
or U29286 (N_29286,N_22765,N_21886);
nor U29287 (N_29287,N_23938,N_23223);
or U29288 (N_29288,N_24311,N_23919);
or U29289 (N_29289,N_22851,N_24630);
and U29290 (N_29290,N_24141,N_21298);
xor U29291 (N_29291,N_24368,N_24610);
and U29292 (N_29292,N_24500,N_22299);
nand U29293 (N_29293,N_21424,N_22547);
nor U29294 (N_29294,N_20933,N_23011);
nor U29295 (N_29295,N_23972,N_24785);
xor U29296 (N_29296,N_20100,N_22336);
or U29297 (N_29297,N_23576,N_24255);
and U29298 (N_29298,N_23907,N_22705);
nor U29299 (N_29299,N_23212,N_23467);
or U29300 (N_29300,N_22448,N_24140);
nor U29301 (N_29301,N_21192,N_21330);
nor U29302 (N_29302,N_22503,N_20336);
nand U29303 (N_29303,N_22090,N_22879);
xor U29304 (N_29304,N_23439,N_21805);
xor U29305 (N_29305,N_20739,N_23152);
nand U29306 (N_29306,N_24023,N_23604);
and U29307 (N_29307,N_21609,N_20178);
and U29308 (N_29308,N_23630,N_20316);
and U29309 (N_29309,N_24375,N_21540);
xor U29310 (N_29310,N_21008,N_22157);
and U29311 (N_29311,N_24365,N_23161);
nand U29312 (N_29312,N_20812,N_24399);
or U29313 (N_29313,N_22024,N_20224);
nor U29314 (N_29314,N_20899,N_22343);
or U29315 (N_29315,N_21017,N_22560);
or U29316 (N_29316,N_22248,N_22318);
nor U29317 (N_29317,N_20076,N_20010);
nor U29318 (N_29318,N_20429,N_24422);
or U29319 (N_29319,N_21998,N_24312);
and U29320 (N_29320,N_24134,N_22392);
nand U29321 (N_29321,N_24443,N_24361);
or U29322 (N_29322,N_22038,N_21712);
xor U29323 (N_29323,N_22126,N_22231);
nand U29324 (N_29324,N_20178,N_22629);
or U29325 (N_29325,N_22515,N_22820);
or U29326 (N_29326,N_20014,N_21963);
nand U29327 (N_29327,N_20012,N_23744);
or U29328 (N_29328,N_20527,N_20880);
nor U29329 (N_29329,N_21387,N_24266);
or U29330 (N_29330,N_21726,N_24965);
nor U29331 (N_29331,N_20969,N_21875);
or U29332 (N_29332,N_22421,N_22074);
or U29333 (N_29333,N_24326,N_22499);
or U29334 (N_29334,N_22349,N_24073);
nor U29335 (N_29335,N_24926,N_23519);
nor U29336 (N_29336,N_21819,N_22180);
or U29337 (N_29337,N_21025,N_20050);
nor U29338 (N_29338,N_24179,N_23085);
or U29339 (N_29339,N_21828,N_21869);
nand U29340 (N_29340,N_20813,N_21310);
or U29341 (N_29341,N_23164,N_24907);
nor U29342 (N_29342,N_24577,N_21089);
nand U29343 (N_29343,N_20552,N_24454);
and U29344 (N_29344,N_23243,N_20311);
nor U29345 (N_29345,N_20642,N_21138);
nor U29346 (N_29346,N_21878,N_21542);
nor U29347 (N_29347,N_23420,N_20554);
or U29348 (N_29348,N_23583,N_24506);
xnor U29349 (N_29349,N_24955,N_24789);
nand U29350 (N_29350,N_23295,N_20603);
nand U29351 (N_29351,N_23316,N_22033);
and U29352 (N_29352,N_24540,N_22452);
xnor U29353 (N_29353,N_23938,N_23581);
nand U29354 (N_29354,N_22245,N_22892);
and U29355 (N_29355,N_20527,N_20623);
or U29356 (N_29356,N_23705,N_23977);
xnor U29357 (N_29357,N_20811,N_23849);
nand U29358 (N_29358,N_20210,N_21817);
and U29359 (N_29359,N_22001,N_23136);
or U29360 (N_29360,N_23021,N_24696);
and U29361 (N_29361,N_20134,N_22546);
and U29362 (N_29362,N_20060,N_21954);
nor U29363 (N_29363,N_21598,N_23281);
and U29364 (N_29364,N_20885,N_24727);
xnor U29365 (N_29365,N_21220,N_21050);
nor U29366 (N_29366,N_24723,N_23720);
nand U29367 (N_29367,N_22838,N_24048);
nor U29368 (N_29368,N_23994,N_23543);
and U29369 (N_29369,N_22009,N_21772);
nor U29370 (N_29370,N_24301,N_21710);
nor U29371 (N_29371,N_23283,N_21123);
xnor U29372 (N_29372,N_23718,N_23462);
or U29373 (N_29373,N_23149,N_21714);
and U29374 (N_29374,N_22836,N_22148);
nand U29375 (N_29375,N_22100,N_21558);
and U29376 (N_29376,N_24641,N_23925);
nand U29377 (N_29377,N_21583,N_23883);
or U29378 (N_29378,N_23200,N_23582);
or U29379 (N_29379,N_24030,N_20149);
and U29380 (N_29380,N_23846,N_23495);
nand U29381 (N_29381,N_23601,N_20941);
nor U29382 (N_29382,N_21900,N_22212);
nand U29383 (N_29383,N_23170,N_24119);
and U29384 (N_29384,N_22169,N_23049);
and U29385 (N_29385,N_23797,N_21530);
and U29386 (N_29386,N_20900,N_21976);
nand U29387 (N_29387,N_23698,N_22107);
or U29388 (N_29388,N_21846,N_24701);
or U29389 (N_29389,N_20173,N_23573);
or U29390 (N_29390,N_23322,N_23048);
or U29391 (N_29391,N_24894,N_20843);
nand U29392 (N_29392,N_21357,N_23112);
and U29393 (N_29393,N_21821,N_20265);
and U29394 (N_29394,N_20615,N_24390);
or U29395 (N_29395,N_20939,N_24456);
nor U29396 (N_29396,N_23795,N_21596);
nand U29397 (N_29397,N_22450,N_21062);
nor U29398 (N_29398,N_21106,N_24781);
or U29399 (N_29399,N_21012,N_21576);
nand U29400 (N_29400,N_23949,N_21075);
nor U29401 (N_29401,N_23913,N_22046);
or U29402 (N_29402,N_23684,N_21163);
nor U29403 (N_29403,N_21830,N_24277);
nand U29404 (N_29404,N_21240,N_21778);
nand U29405 (N_29405,N_21319,N_23807);
nor U29406 (N_29406,N_21155,N_22643);
xor U29407 (N_29407,N_22334,N_22843);
nor U29408 (N_29408,N_20399,N_21392);
or U29409 (N_29409,N_21755,N_20615);
nor U29410 (N_29410,N_22188,N_21964);
xnor U29411 (N_29411,N_21830,N_22197);
nor U29412 (N_29412,N_22059,N_21791);
xor U29413 (N_29413,N_23096,N_23409);
nand U29414 (N_29414,N_21782,N_22084);
nand U29415 (N_29415,N_23550,N_22498);
nor U29416 (N_29416,N_20778,N_21227);
xnor U29417 (N_29417,N_21751,N_22200);
nand U29418 (N_29418,N_22863,N_20974);
nor U29419 (N_29419,N_21048,N_21931);
nor U29420 (N_29420,N_24088,N_24087);
or U29421 (N_29421,N_23924,N_20982);
xnor U29422 (N_29422,N_22260,N_20073);
nand U29423 (N_29423,N_23144,N_23322);
or U29424 (N_29424,N_20793,N_22561);
nor U29425 (N_29425,N_20766,N_21918);
and U29426 (N_29426,N_22796,N_24644);
and U29427 (N_29427,N_22023,N_21423);
nand U29428 (N_29428,N_24311,N_24259);
or U29429 (N_29429,N_20439,N_22790);
nor U29430 (N_29430,N_22592,N_24175);
or U29431 (N_29431,N_20194,N_20604);
and U29432 (N_29432,N_20604,N_22498);
nand U29433 (N_29433,N_21376,N_23887);
xnor U29434 (N_29434,N_23152,N_21960);
or U29435 (N_29435,N_20137,N_21848);
and U29436 (N_29436,N_20763,N_24931);
or U29437 (N_29437,N_22403,N_21225);
or U29438 (N_29438,N_22899,N_20744);
xor U29439 (N_29439,N_22040,N_23630);
and U29440 (N_29440,N_20197,N_24071);
xnor U29441 (N_29441,N_23667,N_23754);
nor U29442 (N_29442,N_21926,N_22879);
nand U29443 (N_29443,N_22360,N_22623);
nor U29444 (N_29444,N_22398,N_23055);
or U29445 (N_29445,N_23334,N_23222);
nor U29446 (N_29446,N_24483,N_20668);
xor U29447 (N_29447,N_23994,N_21431);
nor U29448 (N_29448,N_20884,N_22953);
and U29449 (N_29449,N_24820,N_24261);
and U29450 (N_29450,N_22772,N_23313);
nand U29451 (N_29451,N_21834,N_23597);
nand U29452 (N_29452,N_23329,N_22034);
and U29453 (N_29453,N_24157,N_22965);
and U29454 (N_29454,N_23560,N_21532);
or U29455 (N_29455,N_20190,N_21064);
and U29456 (N_29456,N_23895,N_21699);
nand U29457 (N_29457,N_24661,N_22468);
xor U29458 (N_29458,N_20768,N_22164);
and U29459 (N_29459,N_22773,N_22436);
or U29460 (N_29460,N_23950,N_21651);
and U29461 (N_29461,N_20677,N_21120);
and U29462 (N_29462,N_21222,N_24834);
or U29463 (N_29463,N_22590,N_24843);
nand U29464 (N_29464,N_24266,N_21629);
or U29465 (N_29465,N_20898,N_24408);
nor U29466 (N_29466,N_22515,N_22375);
nor U29467 (N_29467,N_21427,N_23110);
and U29468 (N_29468,N_23462,N_22632);
nand U29469 (N_29469,N_20852,N_21925);
xor U29470 (N_29470,N_21286,N_21659);
and U29471 (N_29471,N_21819,N_21446);
or U29472 (N_29472,N_23163,N_22854);
or U29473 (N_29473,N_22498,N_21694);
nand U29474 (N_29474,N_23590,N_21069);
nand U29475 (N_29475,N_20292,N_23559);
nand U29476 (N_29476,N_24779,N_23215);
nand U29477 (N_29477,N_22629,N_20102);
and U29478 (N_29478,N_22677,N_24079);
or U29479 (N_29479,N_24796,N_22358);
or U29480 (N_29480,N_21695,N_22644);
xor U29481 (N_29481,N_20642,N_23692);
or U29482 (N_29482,N_23076,N_23381);
and U29483 (N_29483,N_23429,N_23112);
nand U29484 (N_29484,N_20261,N_24684);
nand U29485 (N_29485,N_21971,N_20186);
nor U29486 (N_29486,N_22956,N_24177);
nand U29487 (N_29487,N_22109,N_22174);
or U29488 (N_29488,N_20295,N_22588);
and U29489 (N_29489,N_21598,N_20898);
nor U29490 (N_29490,N_20727,N_20449);
nor U29491 (N_29491,N_22515,N_22009);
and U29492 (N_29492,N_23096,N_21269);
or U29493 (N_29493,N_20328,N_22534);
nor U29494 (N_29494,N_20641,N_23658);
or U29495 (N_29495,N_24977,N_21321);
and U29496 (N_29496,N_24951,N_24677);
and U29497 (N_29497,N_23281,N_23388);
or U29498 (N_29498,N_22946,N_24856);
nor U29499 (N_29499,N_23817,N_21441);
and U29500 (N_29500,N_24473,N_22195);
or U29501 (N_29501,N_22413,N_21051);
nor U29502 (N_29502,N_22263,N_20453);
or U29503 (N_29503,N_23483,N_23165);
nor U29504 (N_29504,N_22810,N_20650);
nand U29505 (N_29505,N_22687,N_20053);
or U29506 (N_29506,N_23378,N_20440);
nand U29507 (N_29507,N_22952,N_20854);
nand U29508 (N_29508,N_20557,N_23599);
nor U29509 (N_29509,N_21721,N_21098);
nand U29510 (N_29510,N_21446,N_20185);
nand U29511 (N_29511,N_21073,N_22754);
and U29512 (N_29512,N_22043,N_24316);
or U29513 (N_29513,N_23103,N_22229);
xor U29514 (N_29514,N_20136,N_23857);
and U29515 (N_29515,N_21274,N_21445);
nor U29516 (N_29516,N_21403,N_20840);
nor U29517 (N_29517,N_22724,N_20495);
nand U29518 (N_29518,N_21280,N_22789);
and U29519 (N_29519,N_21069,N_20330);
and U29520 (N_29520,N_24927,N_24219);
or U29521 (N_29521,N_24075,N_21160);
nor U29522 (N_29522,N_23535,N_20985);
or U29523 (N_29523,N_24615,N_22787);
and U29524 (N_29524,N_20184,N_23518);
or U29525 (N_29525,N_22233,N_20102);
and U29526 (N_29526,N_23312,N_24752);
xnor U29527 (N_29527,N_22622,N_20621);
nand U29528 (N_29528,N_23968,N_24943);
xor U29529 (N_29529,N_21033,N_21197);
nand U29530 (N_29530,N_23757,N_21567);
nand U29531 (N_29531,N_21137,N_20841);
xor U29532 (N_29532,N_21840,N_20303);
and U29533 (N_29533,N_21386,N_20273);
and U29534 (N_29534,N_23078,N_23830);
nand U29535 (N_29535,N_23297,N_24607);
and U29536 (N_29536,N_24046,N_21607);
nor U29537 (N_29537,N_23436,N_22349);
nor U29538 (N_29538,N_22199,N_21720);
xor U29539 (N_29539,N_20200,N_23564);
and U29540 (N_29540,N_20302,N_24279);
nand U29541 (N_29541,N_21377,N_22681);
or U29542 (N_29542,N_21973,N_23404);
nand U29543 (N_29543,N_23468,N_20852);
xnor U29544 (N_29544,N_22705,N_23183);
nor U29545 (N_29545,N_24097,N_21615);
and U29546 (N_29546,N_21449,N_24770);
xnor U29547 (N_29547,N_20414,N_20679);
xnor U29548 (N_29548,N_23800,N_21348);
nand U29549 (N_29549,N_24382,N_23438);
or U29550 (N_29550,N_21553,N_21607);
or U29551 (N_29551,N_21490,N_23114);
and U29552 (N_29552,N_20501,N_22910);
nand U29553 (N_29553,N_24020,N_23209);
and U29554 (N_29554,N_22308,N_20243);
nor U29555 (N_29555,N_22595,N_20146);
and U29556 (N_29556,N_21763,N_22267);
or U29557 (N_29557,N_21542,N_24386);
nand U29558 (N_29558,N_21751,N_23368);
and U29559 (N_29559,N_24096,N_23064);
nor U29560 (N_29560,N_20726,N_21578);
xor U29561 (N_29561,N_22210,N_22853);
xor U29562 (N_29562,N_20850,N_24505);
nor U29563 (N_29563,N_23257,N_21974);
nand U29564 (N_29564,N_24119,N_21594);
and U29565 (N_29565,N_21971,N_20986);
and U29566 (N_29566,N_23856,N_23220);
and U29567 (N_29567,N_23184,N_21208);
or U29568 (N_29568,N_23683,N_22018);
and U29569 (N_29569,N_21145,N_20396);
nand U29570 (N_29570,N_21717,N_24771);
nor U29571 (N_29571,N_21529,N_22550);
nand U29572 (N_29572,N_22304,N_21876);
and U29573 (N_29573,N_23531,N_21866);
nand U29574 (N_29574,N_24973,N_23987);
or U29575 (N_29575,N_24267,N_20643);
nand U29576 (N_29576,N_23664,N_23784);
nand U29577 (N_29577,N_21591,N_20740);
and U29578 (N_29578,N_24970,N_20770);
nor U29579 (N_29579,N_21976,N_20837);
xnor U29580 (N_29580,N_23476,N_23083);
or U29581 (N_29581,N_20004,N_21871);
nor U29582 (N_29582,N_23033,N_24006);
or U29583 (N_29583,N_21270,N_21706);
or U29584 (N_29584,N_20985,N_21924);
nor U29585 (N_29585,N_22276,N_20508);
and U29586 (N_29586,N_24216,N_24460);
or U29587 (N_29587,N_20836,N_21583);
xor U29588 (N_29588,N_22880,N_20374);
and U29589 (N_29589,N_22608,N_23049);
nand U29590 (N_29590,N_24651,N_24032);
nand U29591 (N_29591,N_23947,N_23198);
and U29592 (N_29592,N_23619,N_23687);
and U29593 (N_29593,N_24559,N_20365);
nor U29594 (N_29594,N_21641,N_23036);
nor U29595 (N_29595,N_23625,N_20610);
nand U29596 (N_29596,N_24671,N_22874);
and U29597 (N_29597,N_21796,N_23337);
and U29598 (N_29598,N_20781,N_20939);
or U29599 (N_29599,N_24267,N_24750);
and U29600 (N_29600,N_20042,N_24288);
nand U29601 (N_29601,N_23723,N_22852);
nor U29602 (N_29602,N_22448,N_22795);
nor U29603 (N_29603,N_23221,N_20398);
and U29604 (N_29604,N_23048,N_24676);
nand U29605 (N_29605,N_21269,N_21970);
nand U29606 (N_29606,N_23346,N_20840);
nand U29607 (N_29607,N_22545,N_22640);
xor U29608 (N_29608,N_22318,N_23198);
xor U29609 (N_29609,N_23450,N_23081);
nor U29610 (N_29610,N_24463,N_22382);
xor U29611 (N_29611,N_22922,N_24957);
and U29612 (N_29612,N_24053,N_21336);
nor U29613 (N_29613,N_22317,N_23469);
nor U29614 (N_29614,N_22934,N_20256);
or U29615 (N_29615,N_24211,N_20021);
nand U29616 (N_29616,N_23374,N_21120);
xor U29617 (N_29617,N_21978,N_24361);
xnor U29618 (N_29618,N_20898,N_20340);
or U29619 (N_29619,N_21032,N_20627);
xor U29620 (N_29620,N_22057,N_23573);
xor U29621 (N_29621,N_20888,N_24613);
nand U29622 (N_29622,N_22217,N_22121);
nor U29623 (N_29623,N_20223,N_21537);
and U29624 (N_29624,N_20199,N_21723);
and U29625 (N_29625,N_20508,N_23451);
and U29626 (N_29626,N_23861,N_24626);
nor U29627 (N_29627,N_20103,N_21537);
nand U29628 (N_29628,N_24430,N_21645);
and U29629 (N_29629,N_20960,N_20966);
nand U29630 (N_29630,N_21939,N_22321);
and U29631 (N_29631,N_23992,N_23555);
and U29632 (N_29632,N_22043,N_23035);
nor U29633 (N_29633,N_20835,N_24047);
and U29634 (N_29634,N_20611,N_22509);
nor U29635 (N_29635,N_20812,N_24648);
nand U29636 (N_29636,N_21671,N_23591);
nor U29637 (N_29637,N_22464,N_21180);
or U29638 (N_29638,N_23575,N_20822);
nor U29639 (N_29639,N_22605,N_22920);
nor U29640 (N_29640,N_22515,N_20783);
and U29641 (N_29641,N_22302,N_21939);
nor U29642 (N_29642,N_21886,N_23792);
and U29643 (N_29643,N_21161,N_23681);
nand U29644 (N_29644,N_24435,N_23990);
or U29645 (N_29645,N_24838,N_21507);
or U29646 (N_29646,N_20298,N_24295);
and U29647 (N_29647,N_23754,N_24591);
xnor U29648 (N_29648,N_20397,N_20598);
or U29649 (N_29649,N_20013,N_22262);
nand U29650 (N_29650,N_23883,N_24841);
xnor U29651 (N_29651,N_20554,N_21082);
xor U29652 (N_29652,N_23343,N_20028);
nand U29653 (N_29653,N_23697,N_21991);
nand U29654 (N_29654,N_20662,N_23621);
nor U29655 (N_29655,N_20846,N_21982);
nand U29656 (N_29656,N_24858,N_21050);
nor U29657 (N_29657,N_24781,N_20177);
nor U29658 (N_29658,N_21430,N_22577);
nor U29659 (N_29659,N_21119,N_24811);
nand U29660 (N_29660,N_24733,N_23549);
or U29661 (N_29661,N_23035,N_21529);
nor U29662 (N_29662,N_22935,N_24675);
or U29663 (N_29663,N_20340,N_21127);
nor U29664 (N_29664,N_23423,N_23700);
nand U29665 (N_29665,N_20181,N_20648);
or U29666 (N_29666,N_22662,N_21260);
nor U29667 (N_29667,N_24941,N_23634);
and U29668 (N_29668,N_24079,N_23711);
nand U29669 (N_29669,N_20919,N_20208);
xnor U29670 (N_29670,N_21637,N_23820);
nor U29671 (N_29671,N_20489,N_22219);
and U29672 (N_29672,N_24157,N_21952);
xnor U29673 (N_29673,N_20414,N_24030);
nand U29674 (N_29674,N_23385,N_22937);
and U29675 (N_29675,N_24625,N_22990);
and U29676 (N_29676,N_24541,N_24946);
and U29677 (N_29677,N_24512,N_24563);
or U29678 (N_29678,N_23061,N_20652);
or U29679 (N_29679,N_20857,N_22506);
and U29680 (N_29680,N_23697,N_21711);
nor U29681 (N_29681,N_23588,N_24724);
or U29682 (N_29682,N_20374,N_23254);
or U29683 (N_29683,N_24016,N_23901);
nor U29684 (N_29684,N_24988,N_22016);
and U29685 (N_29685,N_24014,N_24536);
and U29686 (N_29686,N_23156,N_21779);
nand U29687 (N_29687,N_23529,N_20238);
nor U29688 (N_29688,N_24545,N_20094);
or U29689 (N_29689,N_20789,N_20830);
nand U29690 (N_29690,N_21718,N_24539);
nand U29691 (N_29691,N_22179,N_22564);
and U29692 (N_29692,N_22611,N_20956);
xnor U29693 (N_29693,N_20605,N_24107);
nand U29694 (N_29694,N_21799,N_24399);
or U29695 (N_29695,N_22950,N_21987);
xnor U29696 (N_29696,N_23238,N_22972);
nand U29697 (N_29697,N_22489,N_21992);
or U29698 (N_29698,N_21093,N_24111);
nor U29699 (N_29699,N_23690,N_22135);
nand U29700 (N_29700,N_22431,N_21686);
nand U29701 (N_29701,N_21915,N_24318);
nand U29702 (N_29702,N_21057,N_24932);
nand U29703 (N_29703,N_22198,N_23470);
nand U29704 (N_29704,N_23985,N_22544);
and U29705 (N_29705,N_20897,N_22517);
nor U29706 (N_29706,N_21559,N_22754);
xnor U29707 (N_29707,N_20792,N_21656);
or U29708 (N_29708,N_24210,N_23147);
nand U29709 (N_29709,N_23193,N_21409);
nor U29710 (N_29710,N_21918,N_23714);
or U29711 (N_29711,N_21332,N_22829);
nand U29712 (N_29712,N_22871,N_23715);
nand U29713 (N_29713,N_20716,N_22003);
nand U29714 (N_29714,N_21852,N_23884);
and U29715 (N_29715,N_22308,N_22902);
nand U29716 (N_29716,N_21140,N_21157);
and U29717 (N_29717,N_21397,N_20627);
and U29718 (N_29718,N_23248,N_21339);
xor U29719 (N_29719,N_24441,N_21629);
nor U29720 (N_29720,N_20483,N_21286);
nor U29721 (N_29721,N_24024,N_23546);
nand U29722 (N_29722,N_24642,N_20230);
or U29723 (N_29723,N_21269,N_23795);
or U29724 (N_29724,N_21425,N_22359);
and U29725 (N_29725,N_20726,N_22129);
xor U29726 (N_29726,N_23593,N_21157);
nand U29727 (N_29727,N_22652,N_23985);
nor U29728 (N_29728,N_22605,N_20389);
xor U29729 (N_29729,N_24400,N_23972);
and U29730 (N_29730,N_23239,N_22719);
or U29731 (N_29731,N_21483,N_22937);
nand U29732 (N_29732,N_22118,N_23449);
xnor U29733 (N_29733,N_24485,N_20588);
and U29734 (N_29734,N_20301,N_22169);
xnor U29735 (N_29735,N_22909,N_21302);
and U29736 (N_29736,N_24993,N_20107);
nor U29737 (N_29737,N_22203,N_21975);
xor U29738 (N_29738,N_22998,N_20324);
and U29739 (N_29739,N_21278,N_23843);
nor U29740 (N_29740,N_22977,N_21297);
or U29741 (N_29741,N_20300,N_22119);
nand U29742 (N_29742,N_20938,N_23381);
and U29743 (N_29743,N_21189,N_24182);
nand U29744 (N_29744,N_24356,N_24607);
or U29745 (N_29745,N_24571,N_22047);
nor U29746 (N_29746,N_20132,N_21470);
nor U29747 (N_29747,N_23049,N_24027);
xor U29748 (N_29748,N_21997,N_22979);
nor U29749 (N_29749,N_23490,N_24479);
nor U29750 (N_29750,N_24844,N_21158);
nand U29751 (N_29751,N_21226,N_24033);
and U29752 (N_29752,N_22656,N_21472);
nor U29753 (N_29753,N_24503,N_23792);
nor U29754 (N_29754,N_24012,N_24769);
nand U29755 (N_29755,N_21732,N_21272);
and U29756 (N_29756,N_21347,N_24120);
and U29757 (N_29757,N_21986,N_20706);
and U29758 (N_29758,N_23871,N_22882);
and U29759 (N_29759,N_20072,N_21646);
and U29760 (N_29760,N_22670,N_20187);
xor U29761 (N_29761,N_23133,N_21643);
nand U29762 (N_29762,N_23088,N_22127);
and U29763 (N_29763,N_21273,N_21791);
or U29764 (N_29764,N_21926,N_22800);
or U29765 (N_29765,N_24786,N_22773);
nand U29766 (N_29766,N_22449,N_23907);
nand U29767 (N_29767,N_21749,N_24533);
and U29768 (N_29768,N_24782,N_20421);
nor U29769 (N_29769,N_20894,N_21537);
nand U29770 (N_29770,N_23255,N_24911);
and U29771 (N_29771,N_20421,N_21366);
nor U29772 (N_29772,N_24433,N_24278);
xor U29773 (N_29773,N_22213,N_22415);
or U29774 (N_29774,N_20047,N_24265);
nand U29775 (N_29775,N_23197,N_23121);
or U29776 (N_29776,N_24850,N_21494);
or U29777 (N_29777,N_20356,N_20491);
nand U29778 (N_29778,N_22652,N_24026);
and U29779 (N_29779,N_22921,N_20397);
and U29780 (N_29780,N_21218,N_20705);
and U29781 (N_29781,N_23597,N_21667);
and U29782 (N_29782,N_20254,N_21885);
or U29783 (N_29783,N_21395,N_24278);
nor U29784 (N_29784,N_22616,N_20310);
or U29785 (N_29785,N_21510,N_22152);
nand U29786 (N_29786,N_22846,N_22616);
nand U29787 (N_29787,N_23165,N_24983);
and U29788 (N_29788,N_20448,N_22816);
and U29789 (N_29789,N_21951,N_22370);
or U29790 (N_29790,N_22679,N_22560);
or U29791 (N_29791,N_23924,N_21682);
and U29792 (N_29792,N_24404,N_21781);
and U29793 (N_29793,N_20977,N_20780);
or U29794 (N_29794,N_24706,N_20250);
or U29795 (N_29795,N_23592,N_24314);
or U29796 (N_29796,N_24966,N_21120);
nand U29797 (N_29797,N_21209,N_23299);
xor U29798 (N_29798,N_22070,N_23777);
xor U29799 (N_29799,N_24940,N_21365);
xnor U29800 (N_29800,N_21900,N_23992);
nand U29801 (N_29801,N_22192,N_24461);
nor U29802 (N_29802,N_24154,N_20754);
nor U29803 (N_29803,N_21507,N_24149);
xor U29804 (N_29804,N_23485,N_20401);
or U29805 (N_29805,N_21960,N_21567);
and U29806 (N_29806,N_24143,N_23130);
or U29807 (N_29807,N_20929,N_20046);
nor U29808 (N_29808,N_24990,N_21705);
nand U29809 (N_29809,N_20398,N_24344);
and U29810 (N_29810,N_21959,N_23920);
nand U29811 (N_29811,N_23504,N_24472);
nor U29812 (N_29812,N_21317,N_22068);
nand U29813 (N_29813,N_23389,N_23086);
nor U29814 (N_29814,N_23254,N_20562);
nand U29815 (N_29815,N_21048,N_22702);
nand U29816 (N_29816,N_24252,N_23981);
nand U29817 (N_29817,N_22563,N_22480);
xor U29818 (N_29818,N_24906,N_21459);
or U29819 (N_29819,N_24851,N_21965);
nor U29820 (N_29820,N_21100,N_21651);
nand U29821 (N_29821,N_21518,N_22735);
nand U29822 (N_29822,N_20059,N_21870);
and U29823 (N_29823,N_20883,N_20740);
nor U29824 (N_29824,N_21384,N_23919);
nor U29825 (N_29825,N_22917,N_21071);
or U29826 (N_29826,N_23182,N_24296);
nor U29827 (N_29827,N_22402,N_20292);
nor U29828 (N_29828,N_21376,N_21145);
xor U29829 (N_29829,N_23881,N_21111);
xnor U29830 (N_29830,N_23893,N_20004);
nor U29831 (N_29831,N_23215,N_24925);
and U29832 (N_29832,N_22371,N_20640);
and U29833 (N_29833,N_22991,N_20604);
nand U29834 (N_29834,N_24839,N_21650);
or U29835 (N_29835,N_24359,N_23954);
and U29836 (N_29836,N_24694,N_22146);
nand U29837 (N_29837,N_20835,N_24633);
nand U29838 (N_29838,N_20455,N_23970);
nand U29839 (N_29839,N_23566,N_24781);
or U29840 (N_29840,N_24969,N_20817);
or U29841 (N_29841,N_21377,N_23579);
nand U29842 (N_29842,N_22509,N_24321);
and U29843 (N_29843,N_23208,N_21017);
nor U29844 (N_29844,N_20285,N_22954);
nor U29845 (N_29845,N_23188,N_20106);
xnor U29846 (N_29846,N_21318,N_23315);
nor U29847 (N_29847,N_22256,N_24564);
or U29848 (N_29848,N_22521,N_24858);
nor U29849 (N_29849,N_22155,N_21876);
nand U29850 (N_29850,N_20238,N_23803);
nand U29851 (N_29851,N_20556,N_23733);
and U29852 (N_29852,N_21578,N_23980);
or U29853 (N_29853,N_23717,N_22219);
nor U29854 (N_29854,N_23537,N_23740);
or U29855 (N_29855,N_21911,N_23215);
nand U29856 (N_29856,N_20753,N_22173);
nand U29857 (N_29857,N_22197,N_23732);
nor U29858 (N_29858,N_20386,N_21057);
or U29859 (N_29859,N_23465,N_24935);
and U29860 (N_29860,N_23286,N_23582);
nand U29861 (N_29861,N_21531,N_24793);
xor U29862 (N_29862,N_24559,N_22553);
nand U29863 (N_29863,N_22092,N_21332);
nor U29864 (N_29864,N_24920,N_23408);
nor U29865 (N_29865,N_23388,N_23254);
nand U29866 (N_29866,N_21489,N_20679);
or U29867 (N_29867,N_21603,N_22045);
xor U29868 (N_29868,N_20943,N_20997);
nor U29869 (N_29869,N_23576,N_20975);
nor U29870 (N_29870,N_22525,N_24979);
and U29871 (N_29871,N_24239,N_24202);
nor U29872 (N_29872,N_24813,N_22942);
and U29873 (N_29873,N_24092,N_22897);
nor U29874 (N_29874,N_20063,N_22446);
or U29875 (N_29875,N_22218,N_22792);
and U29876 (N_29876,N_22282,N_20731);
nand U29877 (N_29877,N_24536,N_24192);
nand U29878 (N_29878,N_24900,N_21858);
and U29879 (N_29879,N_24591,N_24122);
nor U29880 (N_29880,N_24590,N_22013);
nand U29881 (N_29881,N_23584,N_20565);
or U29882 (N_29882,N_20633,N_23348);
or U29883 (N_29883,N_20517,N_24359);
nor U29884 (N_29884,N_23180,N_21892);
xor U29885 (N_29885,N_21891,N_21977);
and U29886 (N_29886,N_23314,N_23445);
nor U29887 (N_29887,N_21662,N_22677);
or U29888 (N_29888,N_23226,N_23608);
and U29889 (N_29889,N_20262,N_20106);
nand U29890 (N_29890,N_24080,N_24792);
and U29891 (N_29891,N_23017,N_24082);
nor U29892 (N_29892,N_24341,N_24978);
nand U29893 (N_29893,N_22020,N_23215);
nor U29894 (N_29894,N_21469,N_20087);
nand U29895 (N_29895,N_23617,N_21185);
and U29896 (N_29896,N_21978,N_21839);
or U29897 (N_29897,N_22253,N_24818);
xnor U29898 (N_29898,N_20054,N_21678);
or U29899 (N_29899,N_23442,N_23075);
nor U29900 (N_29900,N_22769,N_22776);
nor U29901 (N_29901,N_24026,N_24092);
and U29902 (N_29902,N_22081,N_22512);
nand U29903 (N_29903,N_22753,N_24984);
nand U29904 (N_29904,N_23402,N_22398);
nand U29905 (N_29905,N_24596,N_23107);
xnor U29906 (N_29906,N_20920,N_21121);
nand U29907 (N_29907,N_20823,N_24566);
and U29908 (N_29908,N_23378,N_20628);
nand U29909 (N_29909,N_24049,N_21279);
nand U29910 (N_29910,N_20826,N_23976);
and U29911 (N_29911,N_20942,N_20898);
nor U29912 (N_29912,N_23438,N_20678);
nor U29913 (N_29913,N_22017,N_23667);
xnor U29914 (N_29914,N_23655,N_22360);
and U29915 (N_29915,N_20103,N_22803);
nor U29916 (N_29916,N_20118,N_24977);
nand U29917 (N_29917,N_24928,N_20666);
and U29918 (N_29918,N_24379,N_21694);
nand U29919 (N_29919,N_22188,N_21229);
nand U29920 (N_29920,N_20523,N_24905);
nand U29921 (N_29921,N_22813,N_20570);
or U29922 (N_29922,N_21304,N_23744);
nor U29923 (N_29923,N_22098,N_24952);
nor U29924 (N_29924,N_20027,N_23793);
nor U29925 (N_29925,N_21240,N_20775);
or U29926 (N_29926,N_24411,N_22565);
xnor U29927 (N_29927,N_21719,N_24630);
nand U29928 (N_29928,N_22300,N_22298);
or U29929 (N_29929,N_22222,N_22289);
and U29930 (N_29930,N_20829,N_23760);
nor U29931 (N_29931,N_22803,N_21625);
nand U29932 (N_29932,N_20163,N_24197);
nor U29933 (N_29933,N_20887,N_24051);
nor U29934 (N_29934,N_23871,N_24016);
or U29935 (N_29935,N_23450,N_24183);
and U29936 (N_29936,N_21865,N_24059);
nand U29937 (N_29937,N_24317,N_21390);
nand U29938 (N_29938,N_20674,N_22084);
and U29939 (N_29939,N_20212,N_24780);
nor U29940 (N_29940,N_21655,N_20930);
or U29941 (N_29941,N_20930,N_23061);
xor U29942 (N_29942,N_22465,N_20365);
nor U29943 (N_29943,N_23005,N_21559);
xor U29944 (N_29944,N_24118,N_21777);
and U29945 (N_29945,N_24689,N_24924);
and U29946 (N_29946,N_22045,N_20386);
nand U29947 (N_29947,N_20087,N_21971);
xor U29948 (N_29948,N_24460,N_22504);
nor U29949 (N_29949,N_23844,N_20158);
nand U29950 (N_29950,N_24256,N_23037);
nand U29951 (N_29951,N_21664,N_22483);
nor U29952 (N_29952,N_21033,N_20811);
nand U29953 (N_29953,N_20032,N_24658);
nand U29954 (N_29954,N_24212,N_22303);
nor U29955 (N_29955,N_23766,N_24264);
xnor U29956 (N_29956,N_22941,N_22556);
or U29957 (N_29957,N_23482,N_24402);
or U29958 (N_29958,N_20437,N_24061);
and U29959 (N_29959,N_20130,N_21204);
nor U29960 (N_29960,N_24411,N_24030);
xor U29961 (N_29961,N_20350,N_24358);
xor U29962 (N_29962,N_21947,N_21711);
nand U29963 (N_29963,N_24873,N_22573);
xnor U29964 (N_29964,N_21407,N_20393);
nand U29965 (N_29965,N_21404,N_23505);
or U29966 (N_29966,N_20703,N_22867);
and U29967 (N_29967,N_24032,N_20312);
nand U29968 (N_29968,N_22497,N_22390);
nand U29969 (N_29969,N_20165,N_20101);
or U29970 (N_29970,N_24726,N_22826);
nor U29971 (N_29971,N_22641,N_20390);
nor U29972 (N_29972,N_24124,N_23955);
or U29973 (N_29973,N_20762,N_21637);
or U29974 (N_29974,N_23333,N_22105);
and U29975 (N_29975,N_21312,N_21146);
or U29976 (N_29976,N_20619,N_22887);
nand U29977 (N_29977,N_22236,N_23619);
or U29978 (N_29978,N_23814,N_22099);
nor U29979 (N_29979,N_21475,N_22713);
nand U29980 (N_29980,N_24250,N_21675);
nand U29981 (N_29981,N_21714,N_20415);
nor U29982 (N_29982,N_24690,N_22144);
nor U29983 (N_29983,N_20013,N_21038);
nor U29984 (N_29984,N_22289,N_20157);
and U29985 (N_29985,N_22649,N_21919);
nand U29986 (N_29986,N_21214,N_20672);
and U29987 (N_29987,N_20852,N_23324);
nand U29988 (N_29988,N_21840,N_21276);
or U29989 (N_29989,N_20731,N_21225);
and U29990 (N_29990,N_20785,N_21108);
and U29991 (N_29991,N_23842,N_22187);
or U29992 (N_29992,N_20722,N_22896);
or U29993 (N_29993,N_23231,N_21622);
and U29994 (N_29994,N_20141,N_22374);
nand U29995 (N_29995,N_22741,N_21381);
nor U29996 (N_29996,N_21051,N_23997);
nand U29997 (N_29997,N_23537,N_24613);
nand U29998 (N_29998,N_23462,N_24349);
nor U29999 (N_29999,N_23427,N_20006);
nor UO_0 (O_0,N_27977,N_26177);
xor UO_1 (O_1,N_27802,N_25549);
nor UO_2 (O_2,N_25772,N_26323);
and UO_3 (O_3,N_29675,N_25458);
nor UO_4 (O_4,N_28568,N_29665);
nor UO_5 (O_5,N_28877,N_29033);
nand UO_6 (O_6,N_25661,N_25156);
or UO_7 (O_7,N_27450,N_25228);
nor UO_8 (O_8,N_28050,N_26231);
nor UO_9 (O_9,N_25226,N_26201);
nand UO_10 (O_10,N_29276,N_29397);
and UO_11 (O_11,N_27241,N_25183);
and UO_12 (O_12,N_27925,N_29588);
xor UO_13 (O_13,N_26998,N_26984);
nand UO_14 (O_14,N_27082,N_26339);
and UO_15 (O_15,N_27867,N_26937);
or UO_16 (O_16,N_25330,N_29892);
and UO_17 (O_17,N_28858,N_27668);
nor UO_18 (O_18,N_26544,N_27787);
nor UO_19 (O_19,N_26977,N_28509);
and UO_20 (O_20,N_28150,N_28441);
or UO_21 (O_21,N_28940,N_25711);
or UO_22 (O_22,N_28166,N_26550);
and UO_23 (O_23,N_28604,N_29332);
or UO_24 (O_24,N_26356,N_27100);
nand UO_25 (O_25,N_26746,N_28643);
nand UO_26 (O_26,N_25396,N_25860);
nand UO_27 (O_27,N_29346,N_26238);
nor UO_28 (O_28,N_26508,N_26331);
xor UO_29 (O_29,N_27114,N_26052);
nor UO_30 (O_30,N_28693,N_27215);
nor UO_31 (O_31,N_29520,N_27859);
nor UO_32 (O_32,N_25512,N_29654);
and UO_33 (O_33,N_28437,N_26855);
and UO_34 (O_34,N_25022,N_27547);
or UO_35 (O_35,N_27843,N_28861);
or UO_36 (O_36,N_25197,N_28577);
xor UO_37 (O_37,N_28987,N_27799);
or UO_38 (O_38,N_25361,N_25247);
nor UO_39 (O_39,N_28903,N_29202);
or UO_40 (O_40,N_28692,N_28424);
nor UO_41 (O_41,N_25749,N_26887);
or UO_42 (O_42,N_25457,N_26686);
or UO_43 (O_43,N_28070,N_25249);
nand UO_44 (O_44,N_28589,N_28325);
xnor UO_45 (O_45,N_26466,N_29615);
or UO_46 (O_46,N_28075,N_29471);
nor UO_47 (O_47,N_26532,N_28175);
and UO_48 (O_48,N_29339,N_28979);
xor UO_49 (O_49,N_28576,N_28765);
or UO_50 (O_50,N_29240,N_26140);
or UO_51 (O_51,N_27755,N_27663);
nor UO_52 (O_52,N_28550,N_28746);
nor UO_53 (O_53,N_26512,N_26056);
and UO_54 (O_54,N_25400,N_25444);
or UO_55 (O_55,N_28905,N_25878);
or UO_56 (O_56,N_27421,N_25121);
or UO_57 (O_57,N_27360,N_27273);
nor UO_58 (O_58,N_27600,N_29645);
nand UO_59 (O_59,N_25912,N_25826);
nor UO_60 (O_60,N_29028,N_26458);
nand UO_61 (O_61,N_25532,N_28885);
nand UO_62 (O_62,N_29526,N_29481);
nand UO_63 (O_63,N_27329,N_25871);
nor UO_64 (O_64,N_28217,N_26216);
nor UO_65 (O_65,N_28446,N_28431);
and UO_66 (O_66,N_28822,N_27839);
or UO_67 (O_67,N_28695,N_29600);
or UO_68 (O_68,N_28279,N_28481);
and UO_69 (O_69,N_28892,N_26452);
nor UO_70 (O_70,N_28219,N_25016);
and UO_71 (O_71,N_29705,N_29174);
and UO_72 (O_72,N_25962,N_28821);
nand UO_73 (O_73,N_28596,N_29924);
and UO_74 (O_74,N_29823,N_27151);
and UO_75 (O_75,N_29528,N_28878);
or UO_76 (O_76,N_25271,N_29025);
or UO_77 (O_77,N_26509,N_29385);
and UO_78 (O_78,N_29484,N_26061);
nand UO_79 (O_79,N_26946,N_29296);
and UO_80 (O_80,N_29795,N_25803);
nand UO_81 (O_81,N_29487,N_29170);
nor UO_82 (O_82,N_25092,N_28447);
and UO_83 (O_83,N_25304,N_28908);
and UO_84 (O_84,N_28356,N_25779);
or UO_85 (O_85,N_29144,N_28241);
nor UO_86 (O_86,N_27800,N_27063);
nor UO_87 (O_87,N_29218,N_27637);
or UO_88 (O_88,N_28027,N_25148);
and UO_89 (O_89,N_27850,N_25339);
nor UO_90 (O_90,N_25392,N_28571);
nor UO_91 (O_91,N_25657,N_29749);
and UO_92 (O_92,N_29546,N_29418);
or UO_93 (O_93,N_25964,N_26552);
nor UO_94 (O_94,N_25069,N_25072);
xnor UO_95 (O_95,N_27549,N_28803);
nor UO_96 (O_96,N_29522,N_27861);
or UO_97 (O_97,N_26758,N_27906);
nor UO_98 (O_98,N_28439,N_26963);
nor UO_99 (O_99,N_27455,N_27030);
nor UO_100 (O_100,N_26801,N_29466);
nor UO_101 (O_101,N_25329,N_25869);
and UO_102 (O_102,N_28257,N_29623);
or UO_103 (O_103,N_29779,N_27775);
or UO_104 (O_104,N_29716,N_29669);
nand UO_105 (O_105,N_27411,N_26065);
or UO_106 (O_106,N_28713,N_29848);
nor UO_107 (O_107,N_25623,N_29959);
nor UO_108 (O_108,N_29052,N_28873);
and UO_109 (O_109,N_27310,N_29162);
and UO_110 (O_110,N_26173,N_25681);
nand UO_111 (O_111,N_28687,N_25793);
and UO_112 (O_112,N_25483,N_28683);
nor UO_113 (O_113,N_26921,N_26266);
and UO_114 (O_114,N_28379,N_29245);
nor UO_115 (O_115,N_27276,N_28637);
and UO_116 (O_116,N_25331,N_28718);
and UO_117 (O_117,N_25647,N_27871);
nand UO_118 (O_118,N_25917,N_27390);
xor UO_119 (O_119,N_28579,N_26793);
nand UO_120 (O_120,N_28993,N_26881);
nor UO_121 (O_121,N_27845,N_25105);
and UO_122 (O_122,N_29045,N_26500);
or UO_123 (O_123,N_28240,N_28463);
xnor UO_124 (O_124,N_27333,N_25041);
or UO_125 (O_125,N_29209,N_27192);
and UO_126 (O_126,N_25527,N_27161);
nand UO_127 (O_127,N_25059,N_27443);
xnor UO_128 (O_128,N_28763,N_25068);
nor UO_129 (O_129,N_26308,N_26971);
nor UO_130 (O_130,N_26545,N_26955);
or UO_131 (O_131,N_27228,N_29474);
or UO_132 (O_132,N_25785,N_25787);
and UO_133 (O_133,N_28267,N_28278);
nor UO_134 (O_134,N_26272,N_26920);
nand UO_135 (O_135,N_26611,N_25642);
or UO_136 (O_136,N_25874,N_29506);
and UO_137 (O_137,N_27482,N_25216);
nor UO_138 (O_138,N_29225,N_29902);
nand UO_139 (O_139,N_29783,N_26625);
nor UO_140 (O_140,N_27902,N_25238);
nand UO_141 (O_141,N_26197,N_27499);
and UO_142 (O_142,N_27579,N_25309);
nor UO_143 (O_143,N_29662,N_26541);
nor UO_144 (O_144,N_25096,N_26012);
nand UO_145 (O_145,N_28244,N_25859);
or UO_146 (O_146,N_27693,N_29246);
nand UO_147 (O_147,N_27036,N_27319);
or UO_148 (O_148,N_28332,N_25705);
or UO_149 (O_149,N_26415,N_25628);
nor UO_150 (O_150,N_25524,N_27983);
nor UO_151 (O_151,N_28101,N_27020);
nor UO_152 (O_152,N_26904,N_29476);
xnor UO_153 (O_153,N_27269,N_29255);
and UO_154 (O_154,N_26363,N_29835);
nor UO_155 (O_155,N_26291,N_29119);
and UO_156 (O_156,N_25316,N_27229);
xnor UO_157 (O_157,N_26181,N_28696);
or UO_158 (O_158,N_25338,N_25544);
or UO_159 (O_159,N_29023,N_28002);
and UO_160 (O_160,N_26134,N_28033);
nand UO_161 (O_161,N_26411,N_28706);
nor UO_162 (O_162,N_25990,N_29248);
nor UO_163 (O_163,N_29929,N_26326);
and UO_164 (O_164,N_25486,N_29403);
nor UO_165 (O_165,N_28078,N_27572);
and UO_166 (O_166,N_27400,N_27289);
nand UO_167 (O_167,N_25560,N_27836);
nor UO_168 (O_168,N_27467,N_25935);
nand UO_169 (O_169,N_28962,N_26546);
or UO_170 (O_170,N_27338,N_29816);
or UO_171 (O_171,N_28677,N_28483);
nor UO_172 (O_172,N_25499,N_29211);
nand UO_173 (O_173,N_26093,N_27658);
nor UO_174 (O_174,N_28256,N_27890);
nor UO_175 (O_175,N_26751,N_27986);
nor UO_176 (O_176,N_27051,N_25149);
xnor UO_177 (O_177,N_26547,N_26410);
and UO_178 (O_178,N_29518,N_26351);
or UO_179 (O_179,N_27331,N_29353);
and UO_180 (O_180,N_25938,N_25175);
xor UO_181 (O_181,N_25176,N_26076);
nand UO_182 (O_182,N_27284,N_26613);
and UO_183 (O_183,N_25649,N_25612);
and UO_184 (O_184,N_25144,N_25375);
or UO_185 (O_185,N_29782,N_29989);
and UO_186 (O_186,N_27440,N_27089);
nand UO_187 (O_187,N_26381,N_29789);
nor UO_188 (O_188,N_25876,N_27560);
and UO_189 (O_189,N_25502,N_26107);
xnor UO_190 (O_190,N_26264,N_29495);
and UO_191 (O_191,N_25492,N_25154);
nand UO_192 (O_192,N_27138,N_28128);
nor UO_193 (O_193,N_28270,N_27757);
and UO_194 (O_194,N_27248,N_28700);
xor UO_195 (O_195,N_26837,N_26092);
nor UO_196 (O_196,N_27199,N_27277);
nand UO_197 (O_197,N_26344,N_26641);
nand UO_198 (O_198,N_28805,N_29190);
nand UO_199 (O_199,N_25360,N_27334);
nor UO_200 (O_200,N_28773,N_27261);
nor UO_201 (O_201,N_26262,N_28585);
nor UO_202 (O_202,N_27785,N_29389);
nand UO_203 (O_203,N_29679,N_29786);
or UO_204 (O_204,N_26191,N_29291);
or UO_205 (O_205,N_28393,N_29047);
nor UO_206 (O_206,N_25881,N_25870);
and UO_207 (O_207,N_26587,N_29521);
xor UO_208 (O_208,N_25212,N_27777);
and UO_209 (O_209,N_29633,N_29777);
nor UO_210 (O_210,N_26401,N_26103);
or UO_211 (O_211,N_29696,N_26205);
and UO_212 (O_212,N_29371,N_26814);
or UO_213 (O_213,N_25719,N_28848);
nor UO_214 (O_214,N_28381,N_29009);
nand UO_215 (O_215,N_29960,N_27381);
nand UO_216 (O_216,N_26919,N_29290);
nand UO_217 (O_217,N_25841,N_26354);
or UO_218 (O_218,N_27472,N_26617);
nor UO_219 (O_219,N_27872,N_29204);
nand UO_220 (O_220,N_27827,N_29269);
nand UO_221 (O_221,N_29860,N_25231);
nand UO_222 (O_222,N_27251,N_27096);
and UO_223 (O_223,N_26529,N_28627);
nand UO_224 (O_224,N_26962,N_27741);
nor UO_225 (O_225,N_27570,N_25384);
or UO_226 (O_226,N_29392,N_28732);
nand UO_227 (O_227,N_25958,N_25007);
nand UO_228 (O_228,N_28062,N_27683);
and UO_229 (O_229,N_27092,N_27893);
nand UO_230 (O_230,N_25614,N_26969);
nand UO_231 (O_231,N_25203,N_26757);
nor UO_232 (O_232,N_28768,N_27997);
nand UO_233 (O_233,N_27501,N_27109);
or UO_234 (O_234,N_25752,N_27529);
or UO_235 (O_235,N_26894,N_25426);
nand UO_236 (O_236,N_27474,N_27217);
xor UO_237 (O_237,N_27681,N_26108);
nand UO_238 (O_238,N_29948,N_26008);
or UO_239 (O_239,N_26554,N_25145);
nand UO_240 (O_240,N_25159,N_25662);
nand UO_241 (O_241,N_28015,N_29056);
nand UO_242 (O_242,N_29272,N_26853);
or UO_243 (O_243,N_26035,N_29844);
and UO_244 (O_244,N_26324,N_29559);
and UO_245 (O_245,N_26465,N_29817);
xor UO_246 (O_246,N_28544,N_28348);
nand UO_247 (O_247,N_25459,N_29130);
nand UO_248 (O_248,N_28512,N_27825);
nor UO_249 (O_249,N_28127,N_26408);
nor UO_250 (O_250,N_26114,N_28974);
xor UO_251 (O_251,N_25721,N_28239);
nand UO_252 (O_252,N_29871,N_26852);
and UO_253 (O_253,N_28941,N_25116);
and UO_254 (O_254,N_29672,N_26959);
or UO_255 (O_255,N_26276,N_29415);
or UO_256 (O_256,N_25823,N_27520);
nand UO_257 (O_257,N_27690,N_28832);
and UO_258 (O_258,N_25606,N_28880);
nand UO_259 (O_259,N_26553,N_25673);
or UO_260 (O_260,N_28083,N_29193);
nor UO_261 (O_261,N_28841,N_28835);
nand UO_262 (O_262,N_26772,N_29124);
and UO_263 (O_263,N_28375,N_28022);
and UO_264 (O_264,N_25018,N_27582);
nor UO_265 (O_265,N_27098,N_27924);
or UO_266 (O_266,N_28798,N_25748);
or UO_267 (O_267,N_25056,N_27704);
xnor UO_268 (O_268,N_26933,N_27708);
and UO_269 (O_269,N_29996,N_26283);
or UO_270 (O_270,N_25890,N_28281);
or UO_271 (O_271,N_28008,N_28206);
nand UO_272 (O_272,N_26599,N_26212);
and UO_273 (O_273,N_28222,N_28890);
nand UO_274 (O_274,N_28158,N_29912);
or UO_275 (O_275,N_27946,N_27569);
nor UO_276 (O_276,N_26528,N_28052);
nor UO_277 (O_277,N_27300,N_27599);
and UO_278 (O_278,N_27208,N_25202);
nand UO_279 (O_279,N_26188,N_27728);
xor UO_280 (O_280,N_25344,N_28567);
nor UO_281 (O_281,N_28864,N_26676);
and UO_282 (O_282,N_27196,N_26637);
nand UO_283 (O_283,N_29102,N_27876);
nand UO_284 (O_284,N_26213,N_27999);
nand UO_285 (O_285,N_28546,N_25346);
nor UO_286 (O_286,N_27971,N_29992);
nand UO_287 (O_287,N_27789,N_27259);
nand UO_288 (O_288,N_29165,N_25843);
and UO_289 (O_289,N_27067,N_25218);
nand UO_290 (O_290,N_25872,N_25633);
or UO_291 (O_291,N_28777,N_27088);
and UO_292 (O_292,N_27714,N_28020);
and UO_293 (O_293,N_28421,N_29208);
xor UO_294 (O_294,N_28262,N_25577);
nand UO_295 (O_295,N_28895,N_27072);
and UO_296 (O_296,N_27466,N_28642);
or UO_297 (O_297,N_26876,N_25213);
or UO_298 (O_298,N_28436,N_26386);
xor UO_299 (O_299,N_27631,N_25842);
nor UO_300 (O_300,N_29440,N_27901);
nand UO_301 (O_301,N_28871,N_29096);
and UO_302 (O_302,N_29723,N_26385);
and UO_303 (O_303,N_27065,N_27015);
xnor UO_304 (O_304,N_25828,N_28775);
xor UO_305 (O_305,N_27973,N_25634);
nor UO_306 (O_306,N_28112,N_29910);
and UO_307 (O_307,N_27780,N_25619);
or UO_308 (O_308,N_25794,N_29406);
nor UO_309 (O_309,N_29821,N_29523);
or UO_310 (O_310,N_26388,N_28337);
or UO_311 (O_311,N_25750,N_25366);
and UO_312 (O_312,N_27561,N_28238);
or UO_313 (O_313,N_26961,N_29216);
or UO_314 (O_314,N_28742,N_29350);
nand UO_315 (O_315,N_29529,N_27522);
nor UO_316 (O_316,N_26217,N_25497);
or UO_317 (O_317,N_29465,N_29838);
and UO_318 (O_318,N_27214,N_27689);
and UO_319 (O_319,N_27152,N_29362);
and UO_320 (O_320,N_29906,N_27527);
nand UO_321 (O_321,N_29320,N_29067);
nor UO_322 (O_322,N_26384,N_28183);
and UO_323 (O_323,N_29981,N_25783);
or UO_324 (O_324,N_29062,N_29808);
or UO_325 (O_325,N_27605,N_26902);
nand UO_326 (O_326,N_26690,N_25674);
nand UO_327 (O_327,N_27166,N_26194);
nor UO_328 (O_328,N_29311,N_28413);
and UO_329 (O_329,N_29220,N_29555);
and UO_330 (O_330,N_25235,N_29812);
and UO_331 (O_331,N_25579,N_28235);
or UO_332 (O_332,N_27727,N_26062);
and UO_333 (O_333,N_26475,N_28074);
and UO_334 (O_334,N_29066,N_26234);
nor UO_335 (O_335,N_25519,N_26708);
nor UO_336 (O_336,N_29088,N_26517);
xor UO_337 (O_337,N_27242,N_26137);
nand UO_338 (O_338,N_25971,N_28939);
nor UO_339 (O_339,N_28556,N_29420);
xor UO_340 (O_340,N_29525,N_29046);
nor UO_341 (O_341,N_26631,N_29562);
nor UO_342 (O_342,N_25908,N_26460);
nand UO_343 (O_343,N_28931,N_27090);
nor UO_344 (O_344,N_27804,N_26441);
and UO_345 (O_345,N_27205,N_25731);
or UO_346 (O_346,N_26536,N_29718);
nor UO_347 (O_347,N_29927,N_26737);
or UO_348 (O_348,N_25933,N_26704);
nand UO_349 (O_349,N_25911,N_25185);
xnor UO_350 (O_350,N_25272,N_26871);
and UO_351 (O_351,N_28610,N_26476);
nor UO_352 (O_352,N_28527,N_29772);
nor UO_353 (O_353,N_29370,N_26168);
nor UO_354 (O_354,N_25780,N_27703);
or UO_355 (O_355,N_29937,N_26828);
nand UO_356 (O_356,N_28747,N_26202);
or UO_357 (O_357,N_29122,N_29087);
nor UO_358 (O_358,N_29863,N_28387);
nor UO_359 (O_359,N_28738,N_27254);
and UO_360 (O_360,N_28559,N_28759);
and UO_361 (O_361,N_28060,N_26586);
or UO_362 (O_362,N_26808,N_29444);
and UO_363 (O_363,N_28723,N_29509);
nand UO_364 (O_364,N_28419,N_27954);
and UO_365 (O_365,N_29507,N_26718);
nand UO_366 (O_366,N_27771,N_27190);
and UO_367 (O_367,N_29148,N_26319);
nand UO_368 (O_368,N_29452,N_25740);
nor UO_369 (O_369,N_27723,N_27788);
nor UO_370 (O_370,N_28384,N_26387);
nand UO_371 (O_371,N_28784,N_29285);
xnor UO_372 (O_372,N_25540,N_26899);
nand UO_373 (O_373,N_29135,N_27340);
and UO_374 (O_374,N_28819,N_28520);
or UO_375 (O_375,N_26754,N_25369);
and UO_376 (O_376,N_25941,N_27385);
nor UO_377 (O_377,N_29818,N_26342);
nor UO_378 (O_378,N_26159,N_27460);
nand UO_379 (O_379,N_28095,N_26600);
and UO_380 (O_380,N_26169,N_27327);
and UO_381 (O_381,N_26488,N_29417);
and UO_382 (O_382,N_27431,N_29651);
nor UO_383 (O_383,N_25528,N_25024);
nor UO_384 (O_384,N_29702,N_28160);
nand UO_385 (O_385,N_28553,N_28164);
nand UO_386 (O_386,N_28981,N_26986);
nand UO_387 (O_387,N_27833,N_28162);
nand UO_388 (O_388,N_26446,N_26095);
or UO_389 (O_389,N_26932,N_25677);
and UO_390 (O_390,N_25776,N_29595);
or UO_391 (O_391,N_29974,N_29439);
and UO_392 (O_392,N_27136,N_26633);
or UO_393 (O_393,N_28657,N_25124);
xor UO_394 (O_394,N_29176,N_25298);
nor UO_395 (O_395,N_25952,N_28492);
nor UO_396 (O_396,N_29990,N_28552);
and UO_397 (O_397,N_25363,N_29897);
or UO_398 (O_398,N_29915,N_29003);
and UO_399 (O_399,N_25452,N_25863);
nor UO_400 (O_400,N_29398,N_27315);
or UO_401 (O_401,N_29940,N_28029);
nor UO_402 (O_402,N_25365,N_29508);
xor UO_403 (O_403,N_28521,N_29970);
and UO_404 (O_404,N_28678,N_27210);
nand UO_405 (O_405,N_29012,N_27206);
or UO_406 (O_406,N_25586,N_25289);
and UO_407 (O_407,N_29911,N_29407);
nand UO_408 (O_408,N_28490,N_27252);
or UO_409 (O_409,N_26778,N_27688);
and UO_410 (O_410,N_27456,N_25136);
nand UO_411 (O_411,N_27618,N_28331);
or UO_412 (O_412,N_27058,N_28109);
nand UO_413 (O_413,N_29748,N_29853);
nor UO_414 (O_414,N_26254,N_27651);
and UO_415 (O_415,N_29053,N_27480);
nand UO_416 (O_416,N_27953,N_27243);
nor UO_417 (O_417,N_27744,N_29472);
or UO_418 (O_418,N_28006,N_25376);
nor UO_419 (O_419,N_27677,N_28064);
nand UO_420 (O_420,N_28839,N_26243);
xnor UO_421 (O_421,N_28644,N_27620);
and UO_422 (O_422,N_26333,N_27669);
and UO_423 (O_423,N_26560,N_26141);
nor UO_424 (O_424,N_28757,N_28287);
and UO_425 (O_425,N_29198,N_26214);
and UO_426 (O_426,N_27674,N_26653);
or UO_427 (O_427,N_28350,N_27162);
xor UO_428 (O_428,N_29329,N_29873);
and UO_429 (O_429,N_25478,N_28992);
and UO_430 (O_430,N_28796,N_29249);
nor UO_431 (O_431,N_29570,N_26789);
nand UO_432 (O_432,N_29118,N_27519);
and UO_433 (O_433,N_27389,N_27892);
nor UO_434 (O_434,N_28724,N_27235);
and UO_435 (O_435,N_29334,N_29963);
nor UO_436 (O_436,N_26530,N_27323);
and UO_437 (O_437,N_27075,N_27678);
and UO_438 (O_438,N_26094,N_27132);
and UO_439 (O_439,N_29792,N_26121);
nor UO_440 (O_440,N_28364,N_29950);
nor UO_441 (O_441,N_26588,N_29068);
and UO_442 (O_442,N_25034,N_27120);
and UO_443 (O_443,N_27649,N_28476);
xnor UO_444 (O_444,N_26736,N_28828);
or UO_445 (O_445,N_25222,N_26534);
and UO_446 (O_446,N_28690,N_29813);
or UO_447 (O_447,N_25617,N_25132);
xor UO_448 (O_448,N_26563,N_25118);
nor UO_449 (O_449,N_26997,N_27006);
or UO_450 (O_450,N_27819,N_28333);
xnor UO_451 (O_451,N_29297,N_29113);
nand UO_452 (O_452,N_27970,N_28352);
and UO_453 (O_453,N_29707,N_26002);
nor UO_454 (O_454,N_27324,N_29323);
nand UO_455 (O_455,N_27609,N_29836);
nand UO_456 (O_456,N_29300,N_28850);
and UO_457 (O_457,N_28883,N_26082);
or UO_458 (O_458,N_28725,N_27991);
nor UO_459 (O_459,N_27332,N_29676);
nor UO_460 (O_460,N_29728,N_25195);
and UO_461 (O_461,N_27477,N_29458);
or UO_462 (O_462,N_28231,N_29447);
nand UO_463 (O_463,N_26485,N_27398);
or UO_464 (O_464,N_27023,N_28748);
nor UO_465 (O_465,N_29120,N_27057);
or UO_466 (O_466,N_25137,N_27308);
or UO_467 (O_467,N_28028,N_26765);
and UO_468 (O_468,N_27919,N_28435);
and UO_469 (O_469,N_28602,N_26505);
nor UO_470 (O_470,N_28651,N_25265);
xnor UO_471 (O_471,N_28174,N_28087);
nand UO_472 (O_472,N_25561,N_25811);
and UO_473 (O_473,N_27271,N_27626);
nor UO_474 (O_474,N_25322,N_27039);
and UO_475 (O_475,N_29738,N_27948);
and UO_476 (O_476,N_29237,N_29629);
and UO_477 (O_477,N_27375,N_29899);
or UO_478 (O_478,N_27179,N_27950);
and UO_479 (O_479,N_28252,N_29223);
nand UO_480 (O_480,N_27724,N_25857);
and UO_481 (O_481,N_26489,N_25485);
nor UO_482 (O_482,N_28912,N_28360);
nor UO_483 (O_483,N_26750,N_26972);
xor UO_484 (O_484,N_27025,N_25021);
and UO_485 (O_485,N_29464,N_25209);
nand UO_486 (O_486,N_27347,N_28462);
and UO_487 (O_487,N_28597,N_25758);
and UO_488 (O_488,N_27290,N_28261);
and UO_489 (O_489,N_29031,N_27134);
and UO_490 (O_490,N_26005,N_28135);
nor UO_491 (O_491,N_26773,N_27733);
and UO_492 (O_492,N_26826,N_25390);
and UO_493 (O_493,N_28915,N_25281);
and UO_494 (O_494,N_27258,N_26183);
and UO_495 (O_495,N_25670,N_28729);
nand UO_496 (O_496,N_26368,N_28433);
nand UO_497 (O_497,N_29172,N_26392);
and UO_498 (O_498,N_27664,N_27142);
or UO_499 (O_499,N_25201,N_25127);
nand UO_500 (O_500,N_25208,N_26184);
nand UO_501 (O_501,N_25080,N_26526);
and UO_502 (O_502,N_26727,N_29184);
and UO_503 (O_503,N_25777,N_28283);
nor UO_504 (O_504,N_29513,N_28632);
or UO_505 (O_505,N_26261,N_26644);
and UO_506 (O_506,N_25425,N_26629);
or UO_507 (O_507,N_25953,N_27070);
nand UO_508 (O_508,N_27917,N_28391);
and UO_509 (O_509,N_29188,N_27961);
or UO_510 (O_510,N_29746,N_29405);
xor UO_511 (O_511,N_26379,N_29644);
nor UO_512 (O_512,N_25389,N_27805);
and UO_513 (O_513,N_28203,N_29598);
and UO_514 (O_514,N_28118,N_28380);
nor UO_515 (O_515,N_29427,N_25162);
xor UO_516 (O_516,N_25755,N_27557);
nand UO_517 (O_517,N_26456,N_29424);
xnor UO_518 (O_518,N_28976,N_27884);
and UO_519 (O_519,N_29335,N_28788);
nand UO_520 (O_520,N_26666,N_29874);
or UO_521 (O_521,N_26311,N_26843);
or UO_522 (O_522,N_25342,N_27439);
nor UO_523 (O_523,N_25773,N_25654);
nand UO_524 (O_524,N_28804,N_26229);
xnor UO_525 (O_525,N_28025,N_29628);
nand UO_526 (O_526,N_25481,N_29008);
nand UO_527 (O_527,N_29081,N_28534);
nor UO_528 (O_528,N_27750,N_26480);
and UO_529 (O_529,N_28192,N_27987);
or UO_530 (O_530,N_26287,N_25261);
and UO_531 (O_531,N_27128,N_26285);
nor UO_532 (O_532,N_28163,N_25802);
nor UO_533 (O_533,N_29826,N_28921);
or UO_534 (O_534,N_25253,N_28415);
nand UO_535 (O_535,N_29150,N_25172);
nand UO_536 (O_536,N_25009,N_25393);
or UO_537 (O_537,N_28361,N_26559);
nand UO_538 (O_538,N_28731,N_26719);
nand UO_539 (O_539,N_27099,N_29374);
or UO_540 (O_540,N_27445,N_25480);
or UO_541 (O_541,N_27103,N_29064);
and UO_542 (O_542,N_28698,N_27594);
and UO_543 (O_543,N_27113,N_26090);
and UO_544 (O_544,N_27470,N_25055);
nand UO_545 (O_545,N_28897,N_26252);
and UO_546 (O_546,N_26706,N_29268);
or UO_547 (O_547,N_27007,N_26548);
nor UO_548 (O_548,N_26848,N_29670);
and UO_549 (O_549,N_27153,N_27856);
and UO_550 (O_550,N_29463,N_27189);
or UO_551 (O_551,N_29267,N_26551);
or UO_552 (O_552,N_26200,N_28849);
nor UO_553 (O_553,N_27763,N_25276);
xnor UO_554 (O_554,N_29129,N_29326);
xor UO_555 (O_555,N_25621,N_25967);
nor UO_556 (O_556,N_25925,N_27191);
nor UO_557 (O_557,N_29467,N_25367);
nor UO_558 (O_558,N_29071,N_27428);
and UO_559 (O_559,N_26148,N_25408);
or UO_560 (O_560,N_29757,N_26888);
nor UO_561 (O_561,N_27635,N_27083);
or UO_562 (O_562,N_27469,N_27168);
or UO_563 (O_563,N_25134,N_28619);
and UO_564 (O_564,N_25013,N_25582);
and UO_565 (O_565,N_25296,N_27822);
and UO_566 (O_566,N_29040,N_29827);
and UO_567 (O_567,N_26729,N_25804);
and UO_568 (O_568,N_25545,N_27364);
nor UO_569 (O_569,N_27040,N_29840);
nand UO_570 (O_570,N_29342,N_25251);
nand UO_571 (O_571,N_25275,N_29044);
nor UO_572 (O_572,N_25926,N_26377);
nand UO_573 (O_573,N_25340,N_29308);
xnor UO_574 (O_574,N_26976,N_26027);
nor UO_575 (O_575,N_26598,N_26928);
or UO_576 (O_576,N_27653,N_29214);
and UO_577 (O_577,N_27234,N_29995);
or UO_578 (O_578,N_27048,N_27359);
nor UO_579 (O_579,N_25094,N_29709);
and UO_580 (O_580,N_26618,N_26979);
nor UO_581 (O_581,N_29128,N_26503);
nor UO_582 (O_582,N_28321,N_25567);
nor UO_583 (O_583,N_28980,N_26926);
and UO_584 (O_584,N_29341,N_28376);
xnor UO_585 (O_585,N_28782,N_27004);
or UO_586 (O_586,N_28667,N_29425);
nand UO_587 (O_587,N_28829,N_25191);
or UO_588 (O_588,N_28530,N_27821);
nand UO_589 (O_589,N_28755,N_29791);
and UO_590 (O_590,N_25525,N_27309);
or UO_591 (O_591,N_26756,N_29236);
and UO_592 (O_592,N_27401,N_29475);
nor UO_593 (O_593,N_26775,N_26863);
nand UO_594 (O_594,N_29413,N_27768);
or UO_595 (O_595,N_27812,N_26841);
nor UO_596 (O_596,N_29136,N_27233);
or UO_597 (O_597,N_25113,N_27506);
nor UO_598 (O_598,N_28031,N_29433);
nor UO_599 (O_599,N_28478,N_27033);
and UO_600 (O_600,N_25844,N_26178);
xor UO_601 (O_601,N_27602,N_29759);
and UO_602 (O_602,N_25301,N_25484);
or UO_603 (O_603,N_28058,N_28504);
or UO_604 (O_604,N_25865,N_29361);
and UO_605 (O_605,N_26113,N_25495);
and UO_606 (O_606,N_25587,N_28336);
and UO_607 (O_607,N_26337,N_25703);
xor UO_608 (O_608,N_26382,N_29183);
nor UO_609 (O_609,N_26336,N_29489);
nor UO_610 (O_610,N_25608,N_27931);
nor UO_611 (O_611,N_25259,N_27274);
or UO_612 (O_612,N_27554,N_29093);
or UO_613 (O_613,N_27280,N_25627);
and UO_614 (O_614,N_29256,N_25746);
or UO_615 (O_615,N_27478,N_29271);
nand UO_616 (O_616,N_28392,N_27598);
xor UO_617 (O_617,N_29318,N_28685);
nand UO_618 (O_618,N_28089,N_25693);
nand UO_619 (O_619,N_29175,N_25968);
or UO_620 (O_620,N_25576,N_25814);
xor UO_621 (O_621,N_25308,N_29804);
and UO_622 (O_622,N_27513,N_27776);
and UO_623 (O_623,N_26893,N_29185);
nor UO_624 (O_624,N_27388,N_25796);
or UO_625 (O_625,N_28195,N_25727);
nand UO_626 (O_626,N_28558,N_27177);
and UO_627 (O_627,N_25115,N_26985);
and UO_628 (O_628,N_26230,N_29007);
nand UO_629 (O_629,N_29253,N_29577);
nor UO_630 (O_630,N_29745,N_28679);
nor UO_631 (O_631,N_27049,N_26910);
or UO_632 (O_632,N_27815,N_26739);
nor UO_633 (O_633,N_25819,N_26543);
and UO_634 (O_634,N_29719,N_25089);
nand UO_635 (O_635,N_25321,N_25707);
nand UO_636 (O_636,N_25541,N_27348);
xor UO_637 (O_637,N_28416,N_26603);
xor UO_638 (O_638,N_28872,N_28898);
nand UO_639 (O_639,N_26978,N_28013);
nand UO_640 (O_640,N_29658,N_26301);
nand UO_641 (O_641,N_27278,N_28856);
nor UO_642 (O_642,N_29714,N_28769);
nor UO_643 (O_643,N_26567,N_26353);
nand UO_644 (O_644,N_27646,N_28229);
or UO_645 (O_645,N_27444,N_25725);
and UO_646 (O_646,N_26792,N_27245);
and UO_647 (O_647,N_29002,N_27641);
xnor UO_648 (O_648,N_28182,N_28484);
and UO_649 (O_649,N_28019,N_27968);
nand UO_650 (O_650,N_26759,N_28290);
and UO_651 (O_651,N_26809,N_28622);
nand UO_652 (O_652,N_25460,N_29163);
xnor UO_653 (O_653,N_25146,N_25875);
nand UO_654 (O_654,N_25897,N_29480);
nor UO_655 (O_655,N_27005,N_25759);
and UO_656 (O_656,N_26610,N_25575);
or UO_657 (O_657,N_25883,N_28491);
nor UO_658 (O_658,N_28096,N_25867);
or UO_659 (O_659,N_28794,N_28102);
or UO_660 (O_660,N_29961,N_28432);
or UO_661 (O_661,N_28857,N_27201);
nand UO_662 (O_662,N_28586,N_26112);
and UO_663 (O_663,N_28053,N_27370);
and UO_664 (O_664,N_25572,N_26156);
nand UO_665 (O_665,N_26846,N_27122);
and UO_666 (O_666,N_26996,N_25382);
and UO_667 (O_667,N_25315,N_27496);
nand UO_668 (O_668,N_29074,N_27667);
and UO_669 (O_669,N_26215,N_28090);
xnor UO_670 (O_670,N_29152,N_28345);
nand UO_671 (O_671,N_25445,N_29139);
nor UO_672 (O_672,N_26072,N_28314);
nor UO_673 (O_673,N_29345,N_25450);
and UO_674 (O_674,N_26627,N_25078);
nor UO_675 (O_675,N_28477,N_28296);
nand UO_676 (O_676,N_29829,N_27671);
nand UO_677 (O_677,N_29095,N_26364);
nor UO_678 (O_678,N_29436,N_26555);
nor UO_679 (O_679,N_26332,N_25433);
nor UO_680 (O_680,N_26590,N_28684);
or UO_681 (O_681,N_25760,N_29455);
nor UO_682 (O_682,N_29978,N_28218);
and UO_683 (O_683,N_25464,N_28396);
nand UO_684 (O_684,N_28499,N_25120);
nor UO_685 (O_685,N_26391,N_28480);
or UO_686 (O_686,N_27864,N_26882);
nand UO_687 (O_687,N_28220,N_26300);
or UO_688 (O_688,N_26835,N_28474);
nand UO_689 (O_689,N_26664,N_28515);
nor UO_690 (O_690,N_28951,N_29862);
and UO_691 (O_691,N_25409,N_26009);
xnor UO_692 (O_692,N_25358,N_29275);
nand UO_693 (O_693,N_29098,N_27294);
nand UO_694 (O_694,N_28444,N_28430);
and UO_695 (O_695,N_26046,N_25913);
nand UO_696 (O_696,N_25631,N_25822);
nand UO_697 (O_697,N_25932,N_26218);
and UO_698 (O_698,N_26747,N_28273);
and UO_699 (O_699,N_25928,N_25676);
nand UO_700 (O_700,N_29377,N_27905);
nand UO_701 (O_701,N_28372,N_29312);
nor UO_702 (O_702,N_29490,N_26688);
nand UO_703 (O_703,N_25651,N_25836);
and UO_704 (O_704,N_26802,N_29886);
nor UO_705 (O_705,N_27770,N_26060);
and UO_706 (O_706,N_25355,N_25036);
nand UO_707 (O_707,N_27022,N_27110);
and UO_708 (O_708,N_28578,N_27003);
nand UO_709 (O_709,N_29428,N_26699);
xor UO_710 (O_710,N_25632,N_25002);
nor UO_711 (O_711,N_26248,N_25026);
nor UO_712 (O_712,N_28378,N_28461);
or UO_713 (O_713,N_26934,N_29182);
or UO_714 (O_714,N_26794,N_29945);
or UO_715 (O_715,N_27402,N_28170);
nor UO_716 (O_716,N_27781,N_27630);
nor UO_717 (O_717,N_26717,N_29197);
nor UO_718 (O_718,N_29164,N_26891);
and UO_719 (O_719,N_25751,N_29514);
nor UO_720 (O_720,N_29438,N_28442);
nand UO_721 (O_721,N_28402,N_27998);
xnor UO_722 (O_722,N_25683,N_29222);
nor UO_723 (O_723,N_27739,N_26044);
nor UO_724 (O_724,N_25372,N_28831);
nand UO_725 (O_725,N_25155,N_28038);
nand UO_726 (O_726,N_29479,N_25742);
xor UO_727 (O_727,N_26063,N_26649);
and UO_728 (O_728,N_26373,N_27223);
and UO_729 (O_729,N_29360,N_27372);
nor UO_730 (O_730,N_29712,N_28404);
xor UO_731 (O_731,N_25050,N_27197);
nand UO_732 (O_732,N_28704,N_27988);
and UO_733 (O_733,N_27652,N_28525);
nand UO_734 (O_734,N_29556,N_28092);
and UO_735 (O_735,N_26620,N_28913);
nand UO_736 (O_736,N_27124,N_26069);
nand UO_737 (O_737,N_25548,N_27073);
or UO_738 (O_738,N_28147,N_28072);
and UO_739 (O_739,N_26579,N_28370);
nand UO_740 (O_740,N_29865,N_25454);
nand UO_741 (O_741,N_29322,N_25550);
xnor UO_742 (O_742,N_28582,N_29295);
nor UO_743 (O_743,N_25000,N_26347);
nor UO_744 (O_744,N_28168,N_26105);
and UO_745 (O_745,N_25030,N_25093);
nand UO_746 (O_746,N_25989,N_26568);
or UO_747 (O_747,N_27357,N_25001);
and UO_748 (O_748,N_28117,N_26165);
and UO_749 (O_749,N_27369,N_29277);
nor UO_750 (O_750,N_28427,N_26036);
or UO_751 (O_751,N_27155,N_25701);
nand UO_752 (O_752,N_28973,N_27544);
nor UO_753 (O_753,N_27820,N_29338);
nand UO_754 (O_754,N_25515,N_28843);
and UO_755 (O_755,N_28004,N_27001);
nand UO_756 (O_756,N_29212,N_27851);
nor UO_757 (O_757,N_25687,N_28590);
nand UO_758 (O_758,N_27227,N_29020);
nor UO_759 (O_759,N_27147,N_27555);
nor UO_760 (O_760,N_25558,N_28854);
and UO_761 (O_761,N_28855,N_28612);
or UO_762 (O_762,N_27221,N_27160);
and UO_763 (O_763,N_26806,N_27404);
nor UO_764 (O_764,N_26619,N_25268);
or UO_765 (O_765,N_28084,N_28984);
and UO_766 (O_766,N_27042,N_28395);
or UO_767 (O_767,N_26862,N_28711);
nand UO_768 (O_768,N_28989,N_25774);
nand UO_769 (O_769,N_28816,N_25141);
or UO_770 (O_770,N_28201,N_26658);
and UO_771 (O_771,N_27721,N_25111);
nor UO_772 (O_772,N_25595,N_26507);
nor UO_773 (O_773,N_26409,N_26164);
or UO_774 (O_774,N_28744,N_25158);
nand UO_775 (O_775,N_27533,N_26827);
nand UO_776 (O_776,N_26031,N_28324);
nor UO_777 (O_777,N_26463,N_27880);
nand UO_778 (O_778,N_28752,N_28010);
nand UO_779 (O_779,N_27434,N_25232);
or UO_780 (O_780,N_25607,N_27575);
nand UO_781 (O_781,N_27659,N_25234);
nor UO_782 (O_782,N_28297,N_26683);
or UO_783 (O_783,N_27226,N_27525);
nand UO_784 (O_784,N_27841,N_25482);
or UO_785 (O_785,N_27350,N_26030);
and UO_786 (O_786,N_25109,N_25534);
or UO_787 (O_787,N_25747,N_25994);
and UO_788 (O_788,N_29107,N_28440);
nor UO_789 (O_789,N_28793,N_29073);
or UO_790 (O_790,N_27935,N_29419);
nand UO_791 (O_791,N_29279,N_28634);
or UO_792 (O_792,N_25142,N_29706);
nand UO_793 (O_793,N_29624,N_26461);
and UO_794 (O_794,N_25206,N_28100);
or UO_795 (O_795,N_26493,N_26694);
nor UO_796 (O_796,N_29593,N_28294);
and UO_797 (O_797,N_29657,N_25604);
or UO_798 (O_798,N_26224,N_29121);
and UO_799 (O_799,N_25286,N_28714);
nand UO_800 (O_800,N_29396,N_28024);
and UO_801 (O_801,N_25960,N_27000);
xor UO_802 (O_802,N_26174,N_27380);
or UO_803 (O_803,N_26078,N_25194);
nor UO_804 (O_804,N_26582,N_25992);
or UO_805 (O_805,N_26692,N_28786);
or UO_806 (O_806,N_25104,N_29394);
nor UO_807 (O_807,N_29578,N_27219);
or UO_808 (O_808,N_28464,N_25493);
nor UO_809 (O_809,N_26761,N_28814);
nor UO_810 (O_810,N_29281,N_26523);
and UO_811 (O_811,N_25061,N_29072);
nor UO_812 (O_812,N_28251,N_25487);
and UO_813 (O_813,N_27891,N_29699);
and UO_814 (O_814,N_25214,N_29896);
nor UO_815 (O_815,N_27863,N_29179);
or UO_816 (O_816,N_28733,N_26481);
nand UO_817 (O_817,N_27339,N_28561);
nand UO_818 (O_818,N_28658,N_28954);
and UO_819 (O_819,N_25110,N_25679);
nand UO_820 (O_820,N_27459,N_29355);
and UO_821 (O_821,N_26790,N_25991);
nor UO_822 (O_822,N_25060,N_29411);
or UO_823 (O_823,N_26484,N_25349);
and UO_824 (O_824,N_26538,N_27542);
xor UO_825 (O_825,N_27321,N_28626);
and UO_826 (O_826,N_28566,N_27170);
and UO_827 (O_827,N_25704,N_28669);
or UO_828 (O_828,N_25999,N_26908);
xnor UO_829 (O_829,N_27979,N_29574);
nor UO_830 (O_830,N_28236,N_25738);
nor UO_831 (O_831,N_27037,N_26042);
and UO_832 (O_832,N_26885,N_26677);
nor UO_833 (O_833,N_26235,N_29687);
or UO_834 (O_834,N_25570,N_26371);
nor UO_835 (O_835,N_29969,N_25220);
or UO_836 (O_836,N_26204,N_27796);
nand UO_837 (O_837,N_28093,N_29549);
nand UO_838 (O_838,N_29869,N_27383);
nand UO_839 (O_839,N_26219,N_25861);
and UO_840 (O_840,N_25432,N_27912);
xnor UO_841 (O_841,N_29258,N_28263);
or UO_842 (O_842,N_25592,N_26923);
or UO_843 (O_843,N_28507,N_26524);
and UO_844 (O_844,N_28286,N_29830);
nand UO_845 (O_845,N_28303,N_28488);
nand UO_846 (O_846,N_25691,N_26085);
and UO_847 (O_847,N_27080,N_25161);
or UO_848 (O_848,N_29536,N_27951);
nor UO_849 (O_849,N_28401,N_27650);
or UO_850 (O_850,N_27665,N_25398);
nand UO_851 (O_851,N_29976,N_26715);
nand UO_852 (O_852,N_28343,N_27580);
nand UO_853 (O_853,N_25423,N_29443);
nor UO_854 (O_854,N_29317,N_27848);
nand UO_855 (O_855,N_27611,N_27517);
and UO_856 (O_856,N_29333,N_28918);
xor UO_857 (O_857,N_28063,N_25192);
nand UO_858 (O_858,N_27510,N_27387);
xor UO_859 (O_859,N_29516,N_29743);
nor UO_860 (O_860,N_27975,N_28129);
nor UO_861 (O_861,N_29936,N_29918);
nor UO_862 (O_862,N_28105,N_25629);
nor UO_863 (O_863,N_28307,N_27373);
nor UO_864 (O_864,N_25456,N_25943);
nor UO_865 (O_865,N_29468,N_27268);
nand UO_866 (O_866,N_28264,N_25291);
xor UO_867 (O_867,N_28495,N_25734);
or UO_868 (O_868,N_29085,N_29469);
xnor UO_869 (O_869,N_26854,N_25402);
nor UO_870 (O_870,N_29701,N_27511);
nor UO_871 (O_871,N_27314,N_28383);
nor UO_872 (O_872,N_29319,N_27608);
or UO_873 (O_873,N_26850,N_27766);
and UO_874 (O_874,N_27053,N_27509);
xor UO_875 (O_875,N_26817,N_27002);
and UO_876 (O_876,N_28448,N_28340);
or UO_877 (O_877,N_26818,N_29254);
nand UO_878 (O_878,N_28928,N_26020);
nand UO_879 (O_879,N_27619,N_25672);
and UO_880 (O_880,N_26004,N_27032);
nor UO_881 (O_881,N_25494,N_29390);
and UO_882 (O_882,N_27376,N_25507);
or UO_883 (O_883,N_25496,N_28648);
or UO_884 (O_884,N_26345,N_26158);
and UO_885 (O_885,N_26665,N_29832);
and UO_886 (O_886,N_26075,N_29643);
nand UO_887 (O_887,N_27115,N_29939);
and UO_888 (O_888,N_26839,N_29357);
or UO_889 (O_889,N_29270,N_28409);
nor UO_890 (O_890,N_29524,N_27516);
nand UO_891 (O_891,N_25590,N_25431);
nor UO_892 (O_892,N_28670,N_29441);
or UO_893 (O_893,N_25082,N_28097);
or UO_894 (O_894,N_27409,N_26457);
nor UO_895 (O_895,N_26430,N_25948);
nor UO_896 (O_896,N_27897,N_29767);
nand UO_897 (O_897,N_25103,N_27071);
or UO_898 (O_898,N_29566,N_29854);
nor UO_899 (O_899,N_25979,N_29932);
nand UO_900 (O_900,N_26019,N_25079);
or UO_901 (O_901,N_26010,N_26520);
nand UO_902 (O_902,N_26874,N_28455);
nand UO_903 (O_903,N_25603,N_28210);
or UO_904 (O_904,N_27297,N_26397);
or UO_905 (O_905,N_29903,N_25053);
and UO_906 (O_906,N_29530,N_28945);
and UO_907 (O_907,N_27043,N_29841);
and UO_908 (O_908,N_28139,N_28212);
nand UO_909 (O_909,N_26434,N_28518);
nor UO_910 (O_910,N_29586,N_25531);
and UO_911 (O_911,N_29365,N_25479);
nor UO_912 (O_912,N_27077,N_27495);
nand UO_913 (O_913,N_29614,N_29953);
nor UO_914 (O_914,N_29001,N_29755);
or UO_915 (O_915,N_26896,N_29126);
and UO_916 (O_916,N_28457,N_28914);
nor UO_917 (O_917,N_27250,N_27587);
nand UO_918 (O_918,N_29855,N_27807);
or UO_919 (O_919,N_26459,N_25065);
or UO_920 (O_920,N_25901,N_26098);
nor UO_921 (O_921,N_26310,N_29395);
xnor UO_922 (O_922,N_29875,N_28737);
xor UO_923 (O_923,N_27823,N_29082);
or UO_924 (O_924,N_27922,N_26478);
nor UO_925 (O_925,N_28902,N_25624);
xor UO_926 (O_926,N_28815,N_26557);
nand UO_927 (O_927,N_26661,N_25099);
nand UO_928 (O_928,N_26437,N_29880);
nor UO_929 (O_929,N_27305,N_27272);
nand UO_930 (O_930,N_27105,N_29647);
nand UO_931 (O_931,N_27942,N_25035);
nor UO_932 (O_932,N_26510,N_29132);
nor UO_933 (O_933,N_28144,N_26299);
nor UO_934 (O_934,N_28120,N_28119);
nand UO_935 (O_935,N_25813,N_26483);
nor UO_936 (O_936,N_28452,N_26126);
and UO_937 (O_937,N_25660,N_28807);
and UO_938 (O_938,N_28132,N_26130);
and UO_939 (O_939,N_27596,N_26689);
nand UO_940 (O_940,N_29678,N_27169);
or UO_941 (O_941,N_28970,N_25466);
nand UO_942 (O_942,N_26284,N_29999);
or UO_943 (O_943,N_26865,N_29266);
or UO_944 (O_944,N_27644,N_28403);
nand UO_945 (O_945,N_27437,N_29201);
and UO_946 (O_946,N_29703,N_26348);
nor UO_947 (O_947,N_26147,N_27623);
or UO_948 (O_948,N_25569,N_25838);
nand UO_949 (O_949,N_29029,N_29226);
nor UO_950 (O_950,N_27521,N_25373);
nor UO_951 (O_951,N_28126,N_27782);
nand UO_952 (O_952,N_25410,N_29315);
nor UO_953 (O_953,N_25529,N_27028);
or UO_954 (O_954,N_29347,N_29449);
and UO_955 (O_955,N_26742,N_28344);
nand UO_956 (O_956,N_29569,N_27875);
and UO_957 (O_957,N_26470,N_25038);
or UO_958 (O_958,N_27713,N_28284);
and UO_959 (O_959,N_27737,N_27414);
or UO_960 (O_960,N_26245,N_25307);
and UO_961 (O_961,N_26957,N_26605);
or UO_962 (O_962,N_25045,N_25424);
nor UO_963 (O_963,N_27616,N_28197);
nand UO_964 (O_964,N_29192,N_25039);
or UO_965 (O_965,N_29596,N_26438);
and UO_966 (O_966,N_29510,N_27927);
and UO_967 (O_967,N_26506,N_28812);
and UO_968 (O_968,N_25107,N_26767);
nor UO_969 (O_969,N_29650,N_26413);
xor UO_970 (O_970,N_27920,N_25864);
and UO_971 (O_971,N_26535,N_27415);
or UO_972 (O_972,N_29579,N_28767);
nor UO_973 (O_973,N_28365,N_26592);
nor UO_974 (O_974,N_27452,N_29885);
nand UO_975 (O_975,N_26680,N_27353);
or UO_976 (O_976,N_28354,N_26516);
and UO_977 (O_977,N_29196,N_25343);
xnor UO_978 (O_978,N_25171,N_27625);
and UO_979 (O_979,N_25547,N_28479);
nand UO_980 (O_980,N_25380,N_29343);
nand UO_981 (O_981,N_27107,N_29942);
or UO_982 (O_982,N_27397,N_29760);
and UO_983 (O_983,N_29026,N_29916);
or UO_984 (O_984,N_29620,N_29878);
or UO_985 (O_985,N_26125,N_25697);
and UO_986 (O_986,N_27831,N_25313);
nor UO_987 (O_987,N_26258,N_29887);
and UO_988 (O_988,N_28082,N_26735);
and UO_989 (O_989,N_26732,N_27087);
or UO_990 (O_990,N_27574,N_25788);
and UO_991 (O_991,N_25014,N_26395);
or UO_992 (O_992,N_29247,N_28863);
or UO_993 (O_993,N_25896,N_27676);
or UO_994 (O_994,N_27774,N_26810);
nand UO_995 (O_995,N_25332,N_29187);
or UO_996 (O_996,N_28847,N_26856);
or UO_997 (O_997,N_25187,N_25437);
or UO_998 (O_998,N_29773,N_28347);
or UO_999 (O_999,N_25824,N_28572);
nor UO_1000 (O_1000,N_25260,N_26054);
nor UO_1001 (O_1001,N_26487,N_27438);
and UO_1002 (O_1002,N_25557,N_27972);
and UO_1003 (O_1003,N_29260,N_27150);
nor UO_1004 (O_1004,N_28785,N_26947);
nand UO_1005 (O_1005,N_27532,N_25555);
and UO_1006 (O_1006,N_27211,N_28057);
and UO_1007 (O_1007,N_29558,N_26674);
nor UO_1008 (O_1008,N_27500,N_29146);
or UO_1009 (O_1009,N_26738,N_25306);
nand UO_1010 (O_1010,N_26829,N_28875);
xnor UO_1011 (O_1011,N_28400,N_26981);
nor UO_1012 (O_1012,N_26634,N_28694);
or UO_1013 (O_1013,N_28486,N_25598);
nand UO_1014 (O_1014,N_28656,N_26872);
or UO_1015 (O_1015,N_29985,N_25599);
nand UO_1016 (O_1016,N_25791,N_25983);
or UO_1017 (O_1017,N_28911,N_25978);
nor UO_1018 (O_1018,N_28285,N_28631);
nand UO_1019 (O_1019,N_26622,N_25385);
or UO_1020 (O_1020,N_26943,N_25613);
nand UO_1021 (O_1021,N_29625,N_28137);
and UO_1022 (O_1022,N_28428,N_25939);
or UO_1023 (O_1023,N_26712,N_28584);
or UO_1024 (O_1024,N_26203,N_27747);
and UO_1025 (O_1025,N_29800,N_29605);
nand UO_1026 (O_1026,N_25513,N_29519);
or UO_1027 (O_1027,N_26417,N_27903);
and UO_1028 (O_1028,N_25091,N_27066);
or UO_1029 (O_1029,N_27108,N_27673);
or UO_1030 (O_1030,N_26949,N_25616);
nand UO_1031 (O_1031,N_27335,N_25653);
nand UO_1032 (O_1032,N_26341,N_25381);
nand UO_1033 (O_1033,N_29076,N_25877);
xor UO_1034 (O_1034,N_26028,N_26753);
nand UO_1035 (O_1035,N_27955,N_28406);
xor UO_1036 (O_1036,N_28676,N_26256);
and UO_1037 (O_1037,N_26905,N_29765);
or UO_1038 (O_1038,N_25327,N_27240);
nand UO_1039 (O_1039,N_29230,N_25981);
or UO_1040 (O_1040,N_26436,N_27786);
and UO_1041 (O_1041,N_26994,N_25729);
nor UO_1042 (O_1042,N_29901,N_27965);
nor UO_1043 (O_1043,N_25448,N_26074);
nor UO_1044 (O_1044,N_25334,N_29962);
xnor UO_1045 (O_1045,N_29561,N_26740);
nor UO_1046 (O_1046,N_26328,N_26733);
nor UO_1047 (O_1047,N_28649,N_28820);
or UO_1048 (O_1048,N_28169,N_29584);
nor UO_1049 (O_1049,N_26447,N_25593);
and UO_1050 (O_1050,N_29781,N_29344);
nand UO_1051 (O_1051,N_27427,N_25368);
and UO_1052 (O_1052,N_29664,N_28313);
xnor UO_1053 (O_1053,N_28537,N_29221);
nor UO_1054 (O_1054,N_29191,N_26650);
or UO_1055 (O_1055,N_28107,N_28852);
xnor UO_1056 (O_1056,N_26741,N_29741);
and UO_1057 (O_1057,N_26681,N_26182);
or UO_1058 (O_1058,N_25957,N_26847);
nand UO_1059 (O_1059,N_25644,N_26187);
or UO_1060 (O_1060,N_26857,N_28997);
nor UO_1061 (O_1061,N_29366,N_25084);
or UO_1062 (O_1062,N_25976,N_25010);
and UO_1063 (O_1063,N_25403,N_29935);
nor UO_1064 (O_1064,N_28538,N_28888);
or UO_1065 (O_1065,N_29442,N_25128);
and UO_1066 (O_1066,N_29400,N_26651);
nor UO_1067 (O_1067,N_26129,N_29720);
and UO_1068 (O_1068,N_27990,N_25954);
or UO_1069 (O_1069,N_29432,N_25521);
xor UO_1070 (O_1070,N_25766,N_29951);
or UO_1071 (O_1071,N_27291,N_26119);
and UO_1072 (O_1072,N_27283,N_28358);
xnor UO_1073 (O_1073,N_25108,N_26499);
and UO_1074 (O_1074,N_29534,N_29055);
nand UO_1075 (O_1075,N_27200,N_26170);
or UO_1076 (O_1076,N_29806,N_27325);
or UO_1077 (O_1077,N_26734,N_29601);
or UO_1078 (O_1078,N_28373,N_28374);
xnor UO_1079 (O_1079,N_29861,N_26455);
nor UO_1080 (O_1080,N_26672,N_29682);
nand UO_1081 (O_1081,N_29607,N_28454);
nand UO_1082 (O_1082,N_27287,N_26760);
nor UO_1083 (O_1083,N_27175,N_28712);
nand UO_1084 (O_1084,N_26951,N_27194);
and UO_1085 (O_1085,N_25717,N_25475);
or UO_1086 (O_1086,N_28338,N_26440);
or UO_1087 (O_1087,N_25645,N_27638);
nor UO_1088 (O_1088,N_27494,N_28870);
nand UO_1089 (O_1089,N_28280,N_27230);
nand UO_1090 (O_1090,N_29540,N_28003);
nor UO_1091 (O_1091,N_29648,N_26246);
xnor UO_1092 (O_1092,N_29302,N_26771);
nor UO_1093 (O_1093,N_25638,N_27418);
nand UO_1094 (O_1094,N_25211,N_26233);
nand UO_1095 (O_1095,N_28429,N_29717);
or UO_1096 (O_1096,N_27546,N_27502);
or UO_1097 (O_1097,N_25429,N_28045);
or UO_1098 (O_1098,N_27485,N_26823);
nand UO_1099 (O_1099,N_28772,N_29734);
nand UO_1100 (O_1100,N_29108,N_27817);
or UO_1101 (O_1101,N_25337,N_28616);
or UO_1102 (O_1102,N_27512,N_29282);
and UO_1103 (O_1103,N_25414,N_28716);
nand UO_1104 (O_1104,N_28629,N_27934);
and UO_1105 (O_1105,N_26185,N_29688);
and UO_1106 (O_1106,N_25922,N_28526);
nor UO_1107 (O_1107,N_28535,N_29758);
and UO_1108 (O_1108,N_29234,N_28389);
nand UO_1109 (O_1109,N_26128,N_27426);
nand UO_1110 (O_1110,N_25310,N_25317);
nand UO_1111 (O_1111,N_29372,N_26025);
nand UO_1112 (O_1112,N_25919,N_26050);
and UO_1113 (O_1113,N_27722,N_29117);
nor UO_1114 (O_1114,N_25893,N_27534);
or UO_1115 (O_1115,N_26176,N_25708);
and UO_1116 (O_1116,N_29938,N_26366);
xnor UO_1117 (O_1117,N_26669,N_26525);
nor UO_1118 (O_1118,N_27111,N_25739);
or UO_1119 (O_1119,N_25044,N_25415);
nand UO_1120 (O_1120,N_25537,N_25659);
or UO_1121 (O_1121,N_29434,N_27129);
and UO_1122 (O_1122,N_28603,N_27222);
and UO_1123 (O_1123,N_27783,N_25641);
and UO_1124 (O_1124,N_25439,N_28202);
nor UO_1125 (O_1125,N_29511,N_28673);
or UO_1126 (O_1126,N_29224,N_29497);
or UO_1127 (O_1127,N_27603,N_27076);
and UO_1128 (O_1128,N_27275,N_26198);
and UO_1129 (O_1129,N_27978,N_25354);
nor UO_1130 (O_1130,N_27016,N_27127);
xnor UO_1131 (O_1131,N_25236,N_28564);
or UO_1132 (O_1132,N_25884,N_29049);
and UO_1133 (O_1133,N_27832,N_29725);
nor UO_1134 (O_1134,N_29550,N_25090);
or UO_1135 (O_1135,N_29695,N_29097);
and UO_1136 (O_1136,N_27895,N_27266);
xor UO_1137 (O_1137,N_28007,N_27068);
xor UO_1138 (O_1138,N_27959,N_28869);
nor UO_1139 (O_1139,N_27209,N_27430);
nor UO_1140 (O_1140,N_25806,N_26355);
or UO_1141 (O_1141,N_26196,N_28124);
or UO_1142 (O_1142,N_27330,N_27497);
nand UO_1143 (O_1143,N_25086,N_29048);
and UO_1144 (O_1144,N_26084,N_26662);
nor UO_1145 (O_1145,N_27492,N_25946);
or UO_1146 (O_1146,N_28560,N_26313);
or UO_1147 (O_1147,N_29721,N_26192);
and UO_1148 (O_1148,N_26043,N_28496);
or UO_1149 (O_1149,N_29078,N_27910);
and UO_1150 (O_1150,N_28026,N_26866);
nand UO_1151 (O_1151,N_25965,N_28860);
or UO_1152 (O_1152,N_27700,N_26766);
and UO_1153 (O_1153,N_29606,N_26964);
or UO_1154 (O_1154,N_28274,N_25583);
or UO_1155 (O_1155,N_28959,N_26967);
nand UO_1156 (O_1156,N_28734,N_27969);
and UO_1157 (O_1157,N_25551,N_27336);
nor UO_1158 (O_1158,N_27589,N_27503);
and UO_1159 (O_1159,N_29454,N_29386);
nand UO_1160 (O_1160,N_25886,N_29778);
nand UO_1161 (O_1161,N_28275,N_29106);
nand UO_1162 (O_1162,N_29019,N_27628);
or UO_1163 (O_1163,N_26150,N_26001);
xnor UO_1164 (O_1164,N_26724,N_26428);
and UO_1165 (O_1165,N_25862,N_29968);
nor UO_1166 (O_1166,N_28149,N_27801);
nor UO_1167 (O_1167,N_27119,N_27701);
xor UO_1168 (O_1168,N_25357,N_28116);
nand UO_1169 (O_1169,N_29014,N_27285);
and UO_1170 (O_1170,N_29373,N_29766);
nor UO_1171 (O_1171,N_27866,N_25419);
and UO_1172 (O_1172,N_26469,N_29314);
or UO_1173 (O_1173,N_27236,N_25610);
nor UO_1174 (O_1174,N_25809,N_27454);
xnor UO_1175 (O_1175,N_27882,N_27146);
xor UO_1176 (O_1176,N_27311,N_28211);
nand UO_1177 (O_1177,N_27433,N_25723);
nand UO_1178 (O_1178,N_28023,N_27773);
nand UO_1179 (O_1179,N_26492,N_25769);
or UO_1180 (O_1180,N_29866,N_28771);
and UO_1181 (O_1181,N_28056,N_28929);
or UO_1182 (O_1182,N_29697,N_28080);
and UO_1183 (O_1183,N_29611,N_27116);
nor UO_1184 (O_1184,N_26917,N_27476);
or UO_1185 (O_1185,N_25879,N_29898);
and UO_1186 (O_1186,N_26709,N_28171);
and UO_1187 (O_1187,N_25678,N_27174);
and UO_1188 (O_1188,N_26306,N_28562);
nand UO_1189 (O_1189,N_29203,N_28000);
nand UO_1190 (O_1190,N_26412,N_26330);
or UO_1191 (O_1191,N_27416,N_28722);
and UO_1192 (O_1192,N_26038,N_28155);
xor UO_1193 (O_1193,N_26021,N_28845);
nor UO_1194 (O_1194,N_28245,N_26645);
or UO_1195 (O_1195,N_26824,N_27125);
and UO_1196 (O_1196,N_25637,N_28764);
nand UO_1197 (O_1197,N_25100,N_29330);
or UO_1198 (O_1198,N_27064,N_27907);
or UO_1199 (O_1199,N_25266,N_25909);
or UO_1200 (O_1200,N_25371,N_27255);
or UO_1201 (O_1201,N_25955,N_29043);
or UO_1202 (O_1202,N_28647,N_29305);
nand UO_1203 (O_1203,N_25284,N_26260);
and UO_1204 (O_1204,N_25771,N_25052);
xnor UO_1205 (O_1205,N_26189,N_27424);
or UO_1206 (O_1206,N_27758,N_28386);
nand UO_1207 (O_1207,N_25488,N_26807);
and UO_1208 (O_1208,N_25139,N_26684);
nand UO_1209 (O_1209,N_25903,N_26297);
nor UO_1210 (O_1210,N_28048,N_29798);
nor UO_1211 (O_1211,N_29635,N_28573);
xor UO_1212 (O_1212,N_28140,N_27026);
xor UO_1213 (O_1213,N_28181,N_27699);
xnor UO_1214 (O_1214,N_27790,N_26104);
and UO_1215 (O_1215,N_26825,N_26573);
xor UO_1216 (O_1216,N_25173,N_26369);
nor UO_1217 (O_1217,N_27928,N_25898);
and UO_1218 (O_1218,N_28234,N_29833);
nor UO_1219 (O_1219,N_27041,N_26722);
or UO_1220 (O_1220,N_26639,N_25710);
nor UO_1221 (O_1221,N_29831,N_26193);
xnor UO_1222 (O_1222,N_26179,N_26139);
nand UO_1223 (O_1223,N_29889,N_26350);
nand UO_1224 (O_1224,N_29847,N_26255);
or UO_1225 (O_1225,N_26956,N_26429);
nand UO_1226 (O_1226,N_26540,N_26058);
and UO_1227 (O_1227,N_29104,N_27578);
nand UO_1228 (O_1228,N_29036,N_26720);
nor UO_1229 (O_1229,N_25795,N_28988);
nor UO_1230 (O_1230,N_26175,N_28443);
and UO_1231 (O_1231,N_29594,N_25181);
nor UO_1232 (O_1232,N_28186,N_25868);
or UO_1233 (O_1233,N_27767,N_27538);
and UO_1234 (O_1234,N_25636,N_26303);
nor UO_1235 (O_1235,N_27738,N_28660);
or UO_1236 (O_1236,N_26340,N_25279);
or UO_1237 (O_1237,N_27745,N_25921);
nand UO_1238 (O_1238,N_27185,N_26697);
and UO_1239 (O_1239,N_25510,N_28399);
and UO_1240 (O_1240,N_28214,N_28661);
nand UO_1241 (O_1241,N_29895,N_26991);
nand UO_1242 (O_1242,N_27568,N_25163);
nor UO_1243 (O_1243,N_26549,N_28138);
nor UO_1244 (O_1244,N_26786,N_26378);
or UO_1245 (O_1245,N_26199,N_25386);
or UO_1246 (O_1246,N_28532,N_29070);
nand UO_1247 (O_1247,N_25379,N_26640);
or UO_1248 (O_1248,N_29842,N_25461);
and UO_1249 (O_1249,N_28368,N_25668);
and UO_1250 (O_1250,N_25498,N_26298);
or UO_1251 (O_1251,N_27803,N_26628);
and UO_1252 (O_1252,N_25596,N_29378);
xnor UO_1253 (O_1253,N_25230,N_27140);
nand UO_1254 (O_1254,N_28232,N_27670);
nor UO_1255 (O_1255,N_26155,N_26897);
nor UO_1256 (O_1256,N_28246,N_25553);
and UO_1257 (O_1257,N_25730,N_25906);
and UO_1258 (O_1258,N_29292,N_26419);
nand UO_1259 (O_1259,N_27909,N_27858);
nor UO_1260 (O_1260,N_27712,N_25589);
nand UO_1261 (O_1261,N_25169,N_25387);
nand UO_1262 (O_1262,N_25427,N_28639);
or UO_1263 (O_1263,N_27994,N_29685);
nand UO_1264 (O_1264,N_27944,N_26504);
or UO_1265 (O_1265,N_29502,N_29387);
nand UO_1266 (O_1266,N_26832,N_25501);
nand UO_1267 (O_1267,N_27396,N_26089);
nand UO_1268 (O_1268,N_28276,N_29796);
and UO_1269 (O_1269,N_25578,N_28887);
or UO_1270 (O_1270,N_26990,N_26396);
xnor UO_1271 (O_1271,N_27855,N_26585);
nor UO_1272 (O_1272,N_27034,N_29259);
nand UO_1273 (O_1273,N_28408,N_28468);
nor UO_1274 (O_1274,N_25075,N_26779);
nor UO_1275 (O_1275,N_29492,N_28565);
nor UO_1276 (O_1276,N_29732,N_27943);
and UO_1277 (O_1277,N_27887,N_26003);
and UO_1278 (O_1278,N_27661,N_29327);
and UO_1279 (O_1279,N_26247,N_27881);
or UO_1280 (O_1280,N_29864,N_25336);
or UO_1281 (O_1281,N_27698,N_25293);
nand UO_1282 (O_1282,N_25825,N_25067);
and UO_1283 (O_1283,N_26821,N_25058);
xor UO_1284 (O_1284,N_29944,N_25753);
nor UO_1285 (O_1285,N_27995,N_26811);
and UO_1286 (O_1286,N_26791,N_29157);
and UO_1287 (O_1287,N_28802,N_27564);
and UO_1288 (O_1288,N_28282,N_29331);
nor UO_1289 (O_1289,N_29543,N_28489);
and UO_1290 (O_1290,N_28874,N_28310);
xor UO_1291 (O_1291,N_25151,N_27195);
and UO_1292 (O_1292,N_25963,N_28065);
and UO_1293 (O_1293,N_25383,N_26707);
nand UO_1294 (O_1294,N_25422,N_28740);
xor UO_1295 (O_1295,N_29363,N_28018);
or UO_1296 (O_1296,N_26296,N_29393);
nor UO_1297 (O_1297,N_25264,N_26531);
or UO_1298 (O_1298,N_27980,N_29822);
nand UO_1299 (O_1299,N_27292,N_28743);
nand UO_1300 (O_1300,N_29639,N_28316);
nor UO_1301 (O_1301,N_25449,N_25207);
nor UO_1302 (O_1302,N_28943,N_25352);
nand UO_1303 (O_1303,N_26982,N_28739);
and UO_1304 (O_1304,N_28011,N_29824);
nor UO_1305 (O_1305,N_27488,N_25564);
xnor UO_1306 (O_1306,N_27017,N_27610);
or UO_1307 (O_1307,N_25051,N_29751);
and UO_1308 (O_1308,N_29736,N_28681);
and UO_1309 (O_1309,N_26879,N_29060);
and UO_1310 (O_1310,N_29498,N_29689);
nor UO_1311 (O_1311,N_26049,N_25474);
nand UO_1312 (O_1312,N_28306,N_27778);
nor UO_1313 (O_1313,N_28776,N_29079);
or UO_1314 (O_1314,N_28193,N_29065);
or UO_1315 (O_1315,N_28249,N_25421);
nor UO_1316 (O_1316,N_27813,N_27834);
nand UO_1317 (O_1317,N_28191,N_28593);
nor UO_1318 (O_1318,N_28756,N_26011);
nor UO_1319 (O_1319,N_29774,N_29352);
and UO_1320 (O_1320,N_25326,N_27490);
and UO_1321 (O_1321,N_29988,N_25848);
nor UO_1322 (O_1322,N_27760,N_25846);
and UO_1323 (O_1323,N_27084,N_29354);
or UO_1324 (O_1324,N_29160,N_28787);
or UO_1325 (O_1325,N_26501,N_27585);
or UO_1326 (O_1326,N_28592,N_26322);
nand UO_1327 (O_1327,N_27371,N_29110);
nand UO_1328 (O_1328,N_28216,N_29904);
or UO_1329 (O_1329,N_25818,N_26952);
and UO_1330 (O_1330,N_28867,N_28068);
and UO_1331 (O_1331,N_26834,N_27936);
xnor UO_1332 (O_1332,N_28668,N_25325);
or UO_1333 (O_1333,N_29219,N_27597);
nand UO_1334 (O_1334,N_28836,N_28641);
xnor UO_1335 (O_1335,N_27312,N_29456);
and UO_1336 (O_1336,N_25914,N_26120);
and UO_1337 (O_1337,N_25311,N_27345);
nand UO_1338 (O_1338,N_25193,N_29849);
and UO_1339 (O_1339,N_28611,N_25015);
and UO_1340 (O_1340,N_25436,N_27860);
or UO_1341 (O_1341,N_26693,N_25102);
nor UO_1342 (O_1342,N_28620,N_29964);
or UO_1343 (O_1343,N_27463,N_28924);
nor UO_1344 (O_1344,N_27246,N_27491);
nand UO_1345 (O_1345,N_28051,N_25737);
nor UO_1346 (O_1346,N_26014,N_28645);
xor UO_1347 (O_1347,N_28506,N_26685);
nand UO_1348 (O_1348,N_29535,N_26195);
xor UO_1349 (O_1349,N_26404,N_28630);
and UO_1350 (O_1350,N_29058,N_26884);
nand UO_1351 (O_1351,N_26271,N_25600);
and UO_1352 (O_1352,N_25714,N_25123);
nor UO_1353 (O_1353,N_29039,N_26309);
xnor UO_1354 (O_1354,N_29883,N_26941);
nor UO_1355 (O_1355,N_27857,N_25522);
nor UO_1356 (O_1356,N_29100,N_29986);
or UO_1357 (O_1357,N_29294,N_26358);
xor UO_1358 (O_1358,N_26110,N_27008);
and UO_1359 (O_1359,N_25258,N_26352);
and UO_1360 (O_1360,N_25198,N_26604);
xnor UO_1361 (O_1361,N_26157,N_27216);
xnor UO_1362 (O_1362,N_25130,N_29993);
nor UO_1363 (O_1363,N_28594,N_28328);
or UO_1364 (O_1364,N_28172,N_25170);
and UO_1365 (O_1365,N_27213,N_27835);
and UO_1366 (O_1366,N_29410,N_28106);
and UO_1367 (O_1367,N_29634,N_25057);
and UO_1368 (O_1368,N_25428,N_27394);
nor UO_1369 (O_1369,N_25188,N_29488);
nand UO_1370 (O_1370,N_28157,N_28749);
nand UO_1371 (O_1371,N_27846,N_26439);
nor UO_1372 (O_1372,N_27095,N_29724);
nor UO_1373 (O_1373,N_28255,N_27420);
xnor UO_1374 (O_1374,N_27352,N_28304);
and UO_1375 (O_1375,N_26575,N_27182);
and UO_1376 (O_1376,N_27453,N_29461);
and UO_1377 (O_1377,N_26402,N_28199);
and UO_1378 (O_1378,N_27933,N_26875);
nand UO_1379 (O_1379,N_29301,N_25807);
xor UO_1380 (O_1380,N_28405,N_27102);
nor UO_1381 (O_1381,N_25973,N_25031);
nor UO_1382 (O_1382,N_26359,N_29437);
nand UO_1383 (O_1383,N_26418,N_26936);
nand UO_1384 (O_1384,N_27682,N_29810);
nor UO_1385 (O_1385,N_25011,N_25319);
nand UO_1386 (O_1386,N_28319,N_25131);
nand UO_1387 (O_1387,N_28549,N_26039);
or UO_1388 (O_1388,N_28986,N_26584);
nor UO_1389 (O_1389,N_25936,N_25506);
nor UO_1390 (O_1390,N_27952,N_28152);
and UO_1391 (O_1391,N_29512,N_25520);
nand UO_1392 (O_1392,N_27736,N_28809);
or UO_1393 (O_1393,N_26770,N_26675);
nand UO_1394 (O_1394,N_25243,N_25199);
or UO_1395 (O_1395,N_26820,N_28952);
or UO_1396 (O_1396,N_29257,N_27915);
and UO_1397 (O_1397,N_25277,N_29802);
or UO_1398 (O_1398,N_29138,N_26236);
nand UO_1399 (O_1399,N_26973,N_29955);
and UO_1400 (O_1400,N_29094,N_25239);
nand UO_1401 (O_1401,N_26696,N_27031);
nand UO_1402 (O_1402,N_29137,N_28173);
and UO_1403 (O_1403,N_29206,N_27441);
and UO_1404 (O_1404,N_28035,N_25465);
nand UO_1405 (O_1405,N_25434,N_29153);
and UO_1406 (O_1406,N_27985,N_26153);
nand UO_1407 (O_1407,N_25996,N_25451);
nand UO_1408 (O_1408,N_27508,N_29722);
or UO_1409 (O_1409,N_27811,N_25784);
or UO_1410 (O_1410,N_29032,N_27344);
xnor UO_1411 (O_1411,N_25215,N_29542);
nand UO_1412 (O_1412,N_27393,N_28213);
or UO_1413 (O_1413,N_25287,N_28961);
xnor UO_1414 (O_1414,N_27377,N_28503);
nor UO_1415 (O_1415,N_28851,N_27945);
and UO_1416 (O_1416,N_26748,N_27286);
xor UO_1417 (O_1417,N_27157,N_25391);
or UO_1418 (O_1418,N_29531,N_25097);
nor UO_1419 (O_1419,N_29575,N_25591);
or UO_1420 (O_1420,N_27949,N_27976);
nand UO_1421 (O_1421,N_26115,N_27826);
nor UO_1422 (O_1422,N_27967,N_25147);
nand UO_1423 (O_1423,N_29762,N_27588);
or UO_1424 (O_1424,N_25318,N_28607);
xor UO_1425 (O_1425,N_25927,N_27982);
nor UO_1426 (O_1426,N_29814,N_27551);
nor UO_1427 (O_1427,N_27869,N_27993);
nand UO_1428 (O_1428,N_28956,N_27224);
nor UO_1429 (O_1429,N_28165,N_26721);
nor UO_1430 (O_1430,N_26451,N_29470);
or UO_1431 (O_1431,N_26636,N_28014);
nor UO_1432 (O_1432,N_26077,N_27029);
and UO_1433 (O_1433,N_27672,N_25643);
and UO_1434 (O_1434,N_28896,N_25395);
or UO_1435 (O_1435,N_29328,N_26916);
xnor UO_1436 (O_1436,N_26670,N_25972);
nor UO_1437 (O_1437,N_28300,N_25987);
nor UO_1438 (O_1438,N_27592,N_26263);
or UO_1439 (O_1439,N_28547,N_27849);
nor UO_1440 (O_1440,N_27366,N_26127);
nor UO_1441 (O_1441,N_26400,N_28932);
or UO_1442 (O_1442,N_25356,N_29656);
nor UO_1443 (O_1443,N_28985,N_28420);
nand UO_1444 (O_1444,N_25126,N_28909);
nand UO_1445 (O_1445,N_26781,N_26975);
and UO_1446 (O_1446,N_28697,N_26307);
nor UO_1447 (O_1447,N_28482,N_29666);
nand UO_1448 (O_1448,N_26925,N_29416);
or UO_1449 (O_1449,N_28581,N_27762);
and UO_1450 (O_1450,N_29947,N_27941);
nand UO_1451 (O_1451,N_26314,N_27992);
nor UO_1452 (O_1452,N_25378,N_29694);
xor UO_1453 (O_1453,N_26878,N_25401);
or UO_1454 (O_1454,N_26626,N_29763);
and UO_1455 (O_1455,N_29668,N_29116);
and UO_1456 (O_1456,N_27794,N_26454);
or UO_1457 (O_1457,N_25761,N_25902);
or UO_1458 (O_1458,N_25574,N_29627);
nand UO_1459 (O_1459,N_26211,N_28254);
and UO_1460 (O_1460,N_26679,N_26278);
nand UO_1461 (O_1461,N_26097,N_29952);
or UO_1462 (O_1462,N_27791,N_25974);
xor UO_1463 (O_1463,N_28609,N_28818);
nand UO_1464 (O_1464,N_27247,N_26898);
or UO_1465 (O_1465,N_28780,N_27711);
nor UO_1466 (O_1466,N_27926,N_28680);
or UO_1467 (O_1467,N_28806,N_28103);
nor UO_1468 (O_1468,N_27218,N_25895);
or UO_1469 (O_1469,N_28036,N_27244);
nor UO_1470 (O_1470,N_29867,N_29537);
nor UO_1471 (O_1471,N_25837,N_26420);
nor UO_1472 (O_1472,N_26521,N_25233);
nand UO_1473 (O_1473,N_28094,N_26468);
nor UO_1474 (O_1474,N_25833,N_25975);
or UO_1475 (O_1475,N_29446,N_28500);
nand UO_1476 (O_1476,N_25270,N_26873);
or UO_1477 (O_1477,N_26944,N_28289);
nand UO_1478 (O_1478,N_27705,N_26574);
nand UO_1479 (O_1479,N_27358,N_26698);
nand UO_1480 (O_1480,N_28686,N_27612);
nor UO_1481 (O_1481,N_25350,N_27237);
nor UO_1482 (O_1482,N_28039,N_29457);
and UO_1483 (O_1483,N_29532,N_29933);
nand UO_1484 (O_1484,N_26380,N_29691);
and UO_1485 (O_1485,N_28366,N_29274);
nand UO_1486 (O_1486,N_27391,N_26007);
nor UO_1487 (O_1487,N_28493,N_26691);
and UO_1488 (O_1488,N_28601,N_27874);
nand UO_1489 (O_1489,N_28617,N_29042);
nor UO_1490 (O_1490,N_29637,N_25542);
and UO_1491 (O_1491,N_27989,N_25916);
or UO_1492 (O_1492,N_27996,N_28750);
nor UO_1493 (O_1493,N_28972,N_26394);
nand UO_1494 (O_1494,N_26160,N_27615);
nor UO_1495 (O_1495,N_26225,N_26744);
and UO_1496 (O_1496,N_26022,N_25947);
nor UO_1497 (O_1497,N_27622,N_26274);
and UO_1498 (O_1498,N_27320,N_25762);
nor UO_1499 (O_1499,N_26913,N_27716);
nor UO_1500 (O_1500,N_28327,N_29553);
nand UO_1501 (O_1501,N_27956,N_25473);
xnor UO_1502 (O_1502,N_29740,N_26989);
nand UO_1503 (O_1503,N_26869,N_26830);
or UO_1504 (O_1504,N_29402,N_25070);
or UO_1505 (O_1505,N_27764,N_25210);
nor UO_1506 (O_1506,N_29674,N_26730);
xnor UO_1507 (O_1507,N_27830,N_29894);
nor UO_1508 (O_1508,N_29228,N_26895);
or UO_1509 (O_1509,N_26678,N_27295);
and UO_1510 (O_1510,N_25852,N_25278);
and UO_1511 (O_1511,N_28946,N_25244);
nor UO_1512 (O_1512,N_29358,N_26892);
nor UO_1513 (O_1513,N_26859,N_27326);
or UO_1514 (O_1514,N_29430,N_26797);
xor UO_1515 (O_1515,N_29972,N_26606);
nor UO_1516 (O_1516,N_28242,N_29105);
nand UO_1517 (O_1517,N_26784,N_26886);
or UO_1518 (O_1518,N_26318,N_28907);
xnor UO_1519 (O_1519,N_27581,N_29092);
nor UO_1520 (O_1520,N_27484,N_29580);
or UO_1521 (O_1521,N_25019,N_29631);
and UO_1522 (O_1522,N_28043,N_28761);
and UO_1523 (O_1523,N_27349,N_25255);
nor UO_1524 (O_1524,N_27725,N_27937);
and UO_1525 (O_1525,N_25669,N_27754);
nor UO_1526 (O_1526,N_26860,N_29030);
and UO_1527 (O_1527,N_27518,N_28085);
or UO_1528 (O_1528,N_29551,N_26305);
xnor UO_1529 (O_1529,N_29680,N_25345);
or UO_1530 (O_1530,N_28005,N_28691);
or UO_1531 (O_1531,N_28042,N_28999);
or UO_1532 (O_1532,N_29077,N_26833);
nor UO_1533 (O_1533,N_26527,N_28311);
or UO_1534 (O_1534,N_27593,N_27966);
nor UO_1535 (O_1535,N_26111,N_25546);
or UO_1536 (O_1536,N_26755,N_26083);
nor UO_1537 (O_1537,N_28960,N_26840);
xnor UO_1538 (O_1538,N_26295,N_29931);
and UO_1539 (O_1539,N_25299,N_28055);
or UO_1540 (O_1540,N_29504,N_26533);
and UO_1541 (O_1541,N_28037,N_26812);
or UO_1542 (O_1542,N_26621,N_26900);
nand UO_1543 (O_1543,N_27647,N_29309);
nor UO_1544 (O_1544,N_26251,N_28827);
nand UO_1545 (O_1545,N_27838,N_27749);
nor UO_1546 (O_1546,N_25858,N_27918);
and UO_1547 (O_1547,N_28423,N_26302);
or UO_1548 (O_1548,N_25997,N_26958);
nand UO_1549 (O_1549,N_25062,N_27021);
and UO_1550 (O_1550,N_29287,N_28682);
and UO_1551 (O_1551,N_26206,N_28188);
and UO_1552 (O_1552,N_25119,N_28813);
nand UO_1553 (O_1553,N_25227,N_26542);
nand UO_1554 (O_1554,N_27685,N_29617);
xnor UO_1555 (O_1555,N_27591,N_27408);
xor UO_1556 (O_1556,N_29010,N_27365);
and UO_1557 (O_1557,N_26474,N_26671);
nor UO_1558 (O_1558,N_29984,N_29391);
and UO_1559 (O_1559,N_26655,N_25798);
or UO_1560 (O_1560,N_27666,N_29189);
xnor UO_1561 (O_1561,N_29870,N_26966);
xnor UO_1562 (O_1562,N_26647,N_26635);
or UO_1563 (O_1563,N_27583,N_26450);
or UO_1564 (O_1564,N_25394,N_29784);
or UO_1565 (O_1565,N_25982,N_29429);
or UO_1566 (O_1566,N_28533,N_27614);
or UO_1567 (O_1567,N_26100,N_27317);
or UO_1568 (O_1568,N_29379,N_27198);
and UO_1569 (O_1569,N_27094,N_25267);
nand UO_1570 (O_1570,N_29602,N_26315);
nor UO_1571 (O_1571,N_25112,N_27019);
and UO_1572 (O_1572,N_25671,N_26522);
or UO_1573 (O_1573,N_29917,N_29893);
nand UO_1574 (O_1574,N_26491,N_29618);
or UO_1575 (O_1575,N_27981,N_26449);
or UO_1576 (O_1576,N_28511,N_28473);
or UO_1577 (O_1577,N_25122,N_29215);
or UO_1578 (O_1578,N_28377,N_27837);
or UO_1579 (O_1579,N_25320,N_25880);
or UO_1580 (O_1580,N_25028,N_28487);
nand UO_1581 (O_1581,N_26144,N_25718);
or UO_1582 (O_1582,N_28357,N_26286);
or UO_1583 (O_1583,N_29243,N_25970);
and UO_1584 (O_1584,N_27231,N_27898);
xnor UO_1585 (O_1585,N_26240,N_29375);
nand UO_1586 (O_1586,N_26519,N_27710);
nor UO_1587 (O_1587,N_26210,N_29803);
and UO_1588 (O_1588,N_28247,N_27958);
or UO_1589 (O_1589,N_27074,N_29155);
nor UO_1590 (O_1590,N_25046,N_25959);
nor UO_1591 (O_1591,N_29473,N_26851);
xor UO_1592 (O_1592,N_28925,N_28638);
nor UO_1593 (O_1593,N_28762,N_29501);
or UO_1594 (O_1594,N_28899,N_27914);
and UO_1595 (O_1595,N_25348,N_26228);
xnor UO_1596 (O_1596,N_29756,N_27963);
or UO_1597 (O_1597,N_26769,N_25285);
xnor UO_1598 (O_1598,N_25969,N_28079);
and UO_1599 (O_1599,N_26593,N_27106);
and UO_1600 (O_1600,N_27403,N_26495);
nor UO_1601 (O_1601,N_25765,N_28398);
nor UO_1602 (O_1602,N_25568,N_26844);
nand UO_1603 (O_1603,N_28949,N_27795);
nand UO_1604 (O_1604,N_25735,N_28919);
nand UO_1605 (O_1605,N_27085,N_25040);
and UO_1606 (O_1606,N_27584,N_29582);
or UO_1607 (O_1607,N_25489,N_28177);
or UO_1608 (O_1608,N_26638,N_28702);
nand UO_1609 (O_1609,N_25305,N_25114);
and UO_1610 (O_1610,N_28098,N_29143);
nor UO_1611 (O_1611,N_25552,N_28528);
and UO_1612 (O_1612,N_28146,N_29851);
nand UO_1613 (O_1613,N_29655,N_26016);
or UO_1614 (O_1614,N_29273,N_29213);
nor UO_1615 (O_1615,N_26883,N_27586);
nor UO_1616 (O_1616,N_28808,N_25889);
or UO_1617 (O_1617,N_25282,N_25625);
and UO_1618 (O_1618,N_26088,N_25966);
nor UO_1619 (O_1619,N_28032,N_25174);
nor UO_1620 (O_1620,N_28151,N_25566);
nand UO_1621 (O_1621,N_27806,N_28134);
or UO_1622 (O_1622,N_26646,N_28497);
and UO_1623 (O_1623,N_28133,N_27279);
nand UO_1624 (O_1624,N_29195,N_25328);
or UO_1625 (O_1625,N_27984,N_27662);
nand UO_1626 (O_1626,N_27097,N_28073);
nand UO_1627 (O_1627,N_26924,N_29819);
nor UO_1628 (O_1628,N_25832,N_28969);
and UO_1629 (O_1629,N_29289,N_26053);
nand UO_1630 (O_1630,N_26787,N_29780);
nand UO_1631 (O_1631,N_25648,N_26257);
and UO_1632 (O_1632,N_29013,N_27079);
nor UO_1633 (O_1633,N_25827,N_27865);
or UO_1634 (O_1634,N_27044,N_26393);
nor UO_1635 (O_1635,N_26066,N_29922);
and UO_1636 (O_1636,N_27238,N_29888);
xnor UO_1637 (O_1637,N_25150,N_27239);
or UO_1638 (O_1638,N_29920,N_28789);
nor UO_1639 (O_1639,N_25143,N_28459);
nand UO_1640 (O_1640,N_25706,N_29926);
xor UO_1641 (O_1641,N_26513,N_26131);
or UO_1642 (O_1642,N_27553,N_29154);
nand UO_1643 (O_1643,N_25744,N_26242);
nor UO_1644 (O_1644,N_25797,N_25585);
nor UO_1645 (O_1645,N_27842,N_26051);
nand UO_1646 (O_1646,N_29876,N_27743);
or UO_1647 (O_1647,N_29149,N_29921);
and UO_1648 (O_1648,N_25469,N_29399);
xnor UO_1649 (O_1649,N_25290,N_28472);
and UO_1650 (O_1650,N_29690,N_27657);
nor UO_1651 (O_1651,N_28720,N_29286);
nand UO_1652 (O_1652,N_27883,N_29348);
or UO_1653 (O_1653,N_28580,N_28388);
and UO_1654 (O_1654,N_26317,N_29973);
nor UO_1655 (O_1655,N_29038,N_26133);
nor UO_1656 (O_1656,N_27731,N_28471);
nand UO_1657 (O_1657,N_27011,N_27567);
and UO_1658 (O_1658,N_25012,N_26868);
and UO_1659 (O_1659,N_28179,N_29587);
and UO_1660 (O_1660,N_27604,N_25685);
nor UO_1661 (O_1661,N_27069,N_27473);
nand UO_1662 (O_1662,N_26906,N_26612);
nand UO_1663 (O_1663,N_26652,N_29698);
or UO_1664 (O_1664,N_25135,N_29057);
nor UO_1665 (O_1665,N_25063,N_26032);
nor UO_1666 (O_1666,N_26490,N_28689);
nand UO_1667 (O_1667,N_26086,N_29284);
xor UO_1668 (O_1668,N_25359,N_29022);
and UO_1669 (O_1669,N_25288,N_26427);
and UO_1670 (O_1670,N_26803,N_26580);
xor UO_1671 (O_1671,N_26080,N_25666);
nor UO_1672 (O_1672,N_29381,N_26338);
nor UO_1673 (O_1673,N_25417,N_25891);
and UO_1674 (O_1674,N_27639,N_27792);
xor UO_1675 (O_1675,N_26782,N_28417);
and UO_1676 (O_1676,N_29140,N_25817);
or UO_1677 (O_1677,N_28800,N_26591);
nor UO_1678 (O_1678,N_28995,N_29050);
and UO_1679 (O_1679,N_29868,N_28570);
nor UO_1680 (O_1680,N_27173,N_26798);
and UO_1681 (O_1681,N_29217,N_25930);
and UO_1682 (O_1682,N_27640,N_26569);
nor UO_1683 (O_1683,N_26146,N_26407);
nor UO_1684 (O_1684,N_25745,N_26166);
nand UO_1685 (O_1685,N_26034,N_29941);
nand UO_1686 (O_1686,N_28614,N_26571);
xnor UO_1687 (O_1687,N_29737,N_29293);
and UO_1688 (O_1688,N_28975,N_27253);
or UO_1689 (O_1689,N_27093,N_27121);
nor UO_1690 (O_1690,N_29401,N_25597);
and UO_1691 (O_1691,N_26728,N_27889);
nand UO_1692 (O_1692,N_25280,N_26795);
nor UO_1693 (O_1693,N_26055,N_28367);
nand UO_1694 (O_1694,N_28190,N_28122);
or UO_1695 (O_1695,N_25377,N_28557);
nor UO_1696 (O_1696,N_28049,N_27818);
or UO_1697 (O_1697,N_28510,N_28299);
and UO_1698 (O_1698,N_27707,N_25412);
and UO_1699 (O_1699,N_27054,N_29404);
or UO_1700 (O_1700,N_25129,N_28688);
nand UO_1701 (O_1701,N_25471,N_27422);
nor UO_1702 (O_1702,N_26227,N_29568);
nor UO_1703 (O_1703,N_28834,N_25246);
and UO_1704 (O_1704,N_26163,N_26601);
nand UO_1705 (O_1705,N_27465,N_28650);
or UO_1706 (O_1706,N_29304,N_28382);
or UO_1707 (O_1707,N_29683,N_27493);
nor UO_1708 (O_1708,N_26607,N_27078);
nor UO_1709 (O_1709,N_26374,N_28224);
or UO_1710 (O_1710,N_26244,N_25699);
nand UO_1711 (O_1711,N_26432,N_25323);
and UO_1712 (O_1712,N_29086,N_28523);
and UO_1713 (O_1713,N_29884,N_29557);
xor UO_1714 (O_1714,N_26124,N_26424);
nor UO_1715 (O_1715,N_27351,N_26648);
or UO_1716 (O_1716,N_27930,N_25950);
and UO_1717 (O_1717,N_29199,N_28531);
nand UO_1718 (O_1718,N_29839,N_27695);
nand UO_1719 (O_1719,N_28542,N_25855);
or UO_1720 (O_1720,N_27052,N_28978);
or UO_1721 (O_1721,N_29034,N_27765);
xor UO_1722 (O_1722,N_26816,N_27854);
xor UO_1723 (O_1723,N_29011,N_27164);
nand UO_1724 (O_1724,N_29367,N_28334);
nand UO_1725 (O_1725,N_25164,N_27548);
and UO_1726 (O_1726,N_25088,N_26293);
or UO_1727 (O_1727,N_27188,N_26335);
nand UO_1728 (O_1728,N_27304,N_25646);
or UO_1729 (O_1729,N_28625,N_25333);
or UO_1730 (O_1730,N_25420,N_29729);
nand UO_1731 (O_1731,N_29041,N_26578);
nand UO_1732 (O_1732,N_27537,N_27172);
nand UO_1733 (O_1733,N_25834,N_27756);
nor UO_1734 (O_1734,N_26289,N_25688);
nand UO_1735 (O_1735,N_26774,N_27392);
or UO_1736 (O_1736,N_27627,N_29147);
and UO_1737 (O_1737,N_28541,N_26938);
nand UO_1738 (O_1738,N_27536,N_25689);
nor UO_1739 (O_1739,N_28243,N_27363);
nor UO_1740 (O_1740,N_26383,N_29583);
or UO_1741 (O_1741,N_25083,N_27793);
nand UO_1742 (O_1742,N_29303,N_27911);
nor UO_1743 (O_1743,N_28253,N_27617);
nand UO_1744 (O_1744,N_26842,N_25977);
or UO_1745 (O_1745,N_25764,N_29982);
and UO_1746 (O_1746,N_28230,N_28485);
and UO_1747 (O_1747,N_25961,N_25724);
nor UO_1748 (O_1748,N_29265,N_27888);
nor UO_1749 (O_1749,N_26327,N_26282);
nor UO_1750 (O_1750,N_29949,N_26716);
and UO_1751 (O_1751,N_25508,N_27706);
nor UO_1752 (O_1752,N_27293,N_29200);
or UO_1753 (O_1753,N_25500,N_25894);
nand UO_1754 (O_1754,N_28894,N_25594);
and UO_1755 (O_1755,N_28884,N_27316);
or UO_1756 (O_1756,N_29630,N_26453);
and UO_1757 (O_1757,N_29837,N_28906);
nor UO_1758 (O_1758,N_26597,N_28494);
and UO_1759 (O_1759,N_25845,N_29590);
or UO_1760 (O_1760,N_27691,N_27515);
nor UO_1761 (O_1761,N_29114,N_26907);
and UO_1762 (O_1762,N_27462,N_25074);
or UO_1763 (O_1763,N_28543,N_29503);
nand UO_1764 (O_1764,N_29412,N_28529);
or UO_1765 (O_1765,N_25728,N_27413);
or UO_1766 (O_1766,N_25698,N_25463);
nand UO_1767 (O_1767,N_29946,N_26288);
or UO_1768 (O_1768,N_28965,N_29288);
nand UO_1769 (O_1769,N_28671,N_26253);
and UO_1770 (O_1770,N_27797,N_28599);
nand UO_1771 (O_1771,N_25252,N_28108);
or UO_1772 (O_1772,N_25274,N_25554);
nand UO_1773 (O_1773,N_26361,N_26570);
and UO_1774 (O_1774,N_28305,N_29261);
or UO_1775 (O_1775,N_29384,N_26710);
nand UO_1776 (O_1776,N_29649,N_25509);
and UO_1777 (O_1777,N_27232,N_29517);
and UO_1778 (O_1778,N_27530,N_28208);
nor UO_1779 (O_1779,N_27171,N_27921);
nand UO_1780 (O_1780,N_27613,N_29306);
nand UO_1781 (O_1781,N_29477,N_27483);
and UO_1782 (O_1782,N_27808,N_27940);
and UO_1783 (O_1783,N_29435,N_29547);
and UO_1784 (O_1784,N_29843,N_29900);
or UO_1785 (O_1785,N_29186,N_26357);
or UO_1786 (O_1786,N_25165,N_28044);
nand UO_1787 (O_1787,N_27648,N_26576);
and UO_1788 (O_1788,N_25756,N_26539);
and UO_1789 (O_1789,N_25399,N_28810);
nand UO_1790 (O_1790,N_29925,N_27303);
nor UO_1791 (O_1791,N_28817,N_27425);
and UO_1792 (O_1792,N_29801,N_29636);
or UO_1793 (O_1793,N_28942,N_29731);
or UO_1794 (O_1794,N_29744,N_28335);
and UO_1795 (O_1795,N_26186,N_27590);
xor UO_1796 (O_1796,N_28407,N_29325);
and UO_1797 (O_1797,N_25684,N_25757);
or UO_1798 (O_1798,N_25799,N_29907);
or UO_1799 (O_1799,N_27307,N_26081);
and UO_1800 (O_1800,N_27908,N_29560);
or UO_1801 (O_1801,N_27601,N_29646);
nand UO_1802 (O_1802,N_25937,N_29109);
and UO_1803 (O_1803,N_27322,N_27081);
xor UO_1804 (O_1804,N_26583,N_25462);
nand UO_1805 (O_1805,N_25517,N_28886);
and UO_1806 (O_1806,N_28958,N_25351);
nor UO_1807 (O_1807,N_29307,N_27313);
nor UO_1808 (O_1808,N_28200,N_27154);
nand UO_1809 (O_1809,N_27894,N_27257);
nor UO_1810 (O_1810,N_26162,N_26304);
nor UO_1811 (O_1811,N_28633,N_29805);
or UO_1812 (O_1812,N_29608,N_26657);
or UO_1813 (O_1813,N_25047,N_29422);
nand UO_1814 (O_1814,N_28901,N_26477);
and UO_1815 (O_1815,N_28318,N_29178);
nor UO_1816 (O_1816,N_27489,N_29708);
xnor UO_1817 (O_1817,N_26334,N_27436);
nand UO_1818 (O_1818,N_28266,N_29035);
nor UO_1819 (O_1819,N_25256,N_27539);
nor UO_1820 (O_1820,N_26067,N_27405);
or UO_1821 (O_1821,N_28889,N_28021);
and UO_1822 (O_1822,N_27145,N_29145);
xor UO_1823 (O_1823,N_29975,N_29591);
or UO_1824 (O_1824,N_26616,N_27471);
or UO_1825 (O_1825,N_28783,N_26780);
nor UO_1826 (O_1826,N_28076,N_26399);
nand UO_1827 (O_1827,N_26889,N_28675);
and UO_1828 (O_1828,N_28111,N_25829);
nand UO_1829 (O_1829,N_27281,N_26018);
and UO_1830 (O_1830,N_28936,N_26346);
or UO_1831 (O_1831,N_27435,N_29450);
nand UO_1832 (O_1832,N_27126,N_25900);
or UO_1833 (O_1833,N_27187,N_25476);
or UO_1834 (O_1834,N_29017,N_29141);
nand UO_1835 (O_1835,N_29882,N_25781);
nand UO_1836 (O_1836,N_26930,N_29499);
or UO_1837 (O_1837,N_25283,N_28450);
xnor UO_1838 (O_1838,N_26745,N_27163);
xor UO_1839 (O_1839,N_27526,N_28588);
xor UO_1840 (O_1840,N_27885,N_27726);
xor UO_1841 (O_1841,N_29091,N_26047);
nor UO_1842 (O_1842,N_25805,N_26482);
nor UO_1843 (O_1843,N_27135,N_27654);
nand UO_1844 (O_1844,N_27342,N_29845);
xor UO_1845 (O_1845,N_27810,N_29021);
nor UO_1846 (O_1846,N_26723,N_28067);
and UO_1847 (O_1847,N_28727,N_25225);
and UO_1848 (O_1848,N_29239,N_27130);
or UO_1849 (O_1849,N_25998,N_25993);
nand UO_1850 (O_1850,N_28719,N_28145);
nor UO_1851 (O_1851,N_26223,N_29764);
nor UO_1852 (O_1852,N_25071,N_26608);
nor UO_1853 (O_1853,N_27686,N_29478);
or UO_1854 (O_1854,N_25470,N_29486);
nor UO_1855 (O_1855,N_27709,N_26023);
and UO_1856 (O_1856,N_25048,N_26725);
and UO_1857 (O_1857,N_26776,N_25254);
and UO_1858 (O_1858,N_29084,N_28508);
xor UO_1859 (O_1859,N_25851,N_26912);
or UO_1860 (O_1860,N_26365,N_25882);
or UO_1861 (O_1861,N_28228,N_26059);
and UO_1862 (O_1862,N_25003,N_29811);
nor UO_1863 (O_1863,N_29571,N_25023);
nor UO_1864 (O_1864,N_29262,N_26462);
nand UO_1865 (O_1865,N_25179,N_25622);
and UO_1866 (O_1866,N_28795,N_28130);
or UO_1867 (O_1867,N_27060,N_28933);
or UO_1868 (O_1868,N_26701,N_28826);
nand UO_1869 (O_1869,N_28269,N_28059);
and UO_1870 (O_1870,N_28205,N_27718);
or UO_1871 (O_1871,N_25931,N_27541);
nor UO_1872 (O_1872,N_25133,N_27528);
and UO_1873 (O_1873,N_29264,N_29573);
nand UO_1874 (O_1874,N_26656,N_26045);
or UO_1875 (O_1875,N_29788,N_29089);
and UO_1876 (O_1876,N_26190,N_27355);
and UO_1877 (O_1877,N_27056,N_29527);
or UO_1878 (O_1878,N_27595,N_28811);
xnor UO_1879 (O_1879,N_26909,N_26562);
and UO_1880 (O_1880,N_29890,N_27562);
nor UO_1881 (O_1881,N_26813,N_25543);
nor UO_1882 (O_1882,N_28674,N_29790);
nand UO_1883 (O_1883,N_27423,N_26017);
or UO_1884 (O_1884,N_27301,N_29576);
and UO_1885 (O_1885,N_28944,N_26015);
and UO_1886 (O_1886,N_27507,N_28475);
and UO_1887 (O_1887,N_26149,N_26558);
or UO_1888 (O_1888,N_26057,N_28665);
or UO_1889 (O_1889,N_26208,N_28555);
or UO_1890 (O_1890,N_29980,N_25229);
or UO_1891 (O_1891,N_26079,N_28426);
nand UO_1892 (O_1892,N_25407,N_28323);
or UO_1893 (O_1893,N_28221,N_27059);
nor UO_1894 (O_1894,N_25032,N_27629);
or UO_1895 (O_1895,N_25477,N_28469);
or UO_1896 (O_1896,N_26423,N_28646);
or UO_1897 (O_1897,N_25153,N_29027);
nor UO_1898 (O_1898,N_26360,N_26362);
or UO_1899 (O_1899,N_27204,N_27270);
nand UO_1900 (O_1900,N_29710,N_28536);
nand UO_1901 (O_1901,N_29943,N_25800);
xnor UO_1902 (O_1902,N_25167,N_29622);
nand UO_1903 (O_1903,N_27143,N_27543);
or UO_1904 (O_1904,N_28292,N_28844);
and UO_1905 (O_1905,N_29991,N_29711);
xnor UO_1906 (O_1906,N_28227,N_29671);
xnor UO_1907 (O_1907,N_29733,N_28445);
or UO_1908 (O_1908,N_26241,N_27900);
and UO_1909 (O_1909,N_28369,N_28414);
and UO_1910 (O_1910,N_28624,N_25314);
xnor UO_1911 (O_1911,N_25085,N_27202);
nand UO_1912 (O_1912,N_25217,N_27050);
or UO_1913 (O_1913,N_27407,N_26497);
nand UO_1914 (O_1914,N_27014,N_28948);
and UO_1915 (O_1915,N_27550,N_25665);
or UO_1916 (O_1916,N_28185,N_28293);
nor UO_1917 (O_1917,N_28209,N_28699);
nand UO_1918 (O_1918,N_26290,N_26743);
and UO_1919 (O_1919,N_29846,N_28866);
or UO_1920 (O_1920,N_27288,N_27361);
or UO_1921 (O_1921,N_25043,N_25341);
nand UO_1922 (O_1922,N_27735,N_28539);
or UO_1923 (O_1923,N_25081,N_25168);
nand UO_1924 (O_1924,N_25741,N_28233);
nand UO_1925 (O_1925,N_27559,N_26777);
nand UO_1926 (O_1926,N_25984,N_27449);
nor UO_1927 (O_1927,N_27468,N_25262);
xor UO_1928 (O_1928,N_29340,N_28994);
xor UO_1929 (O_1929,N_26435,N_28204);
nor UO_1930 (O_1930,N_27487,N_27367);
nor UO_1931 (O_1931,N_28554,N_27225);
nand UO_1932 (O_1932,N_26663,N_29194);
nor UO_1933 (O_1933,N_29872,N_29787);
and UO_1934 (O_1934,N_25455,N_26101);
nor UO_1935 (O_1935,N_26992,N_27734);
nor UO_1936 (O_1936,N_28329,N_28223);
nor UO_1937 (O_1937,N_25899,N_29101);
or UO_1938 (O_1938,N_26726,N_27117);
nand UO_1939 (O_1939,N_26096,N_28778);
or UO_1940 (O_1940,N_27149,N_27702);
or UO_1941 (O_1941,N_25033,N_27742);
nor UO_1942 (O_1942,N_25910,N_29103);
and UO_1943 (O_1943,N_25505,N_28456);
nor UO_1944 (O_1944,N_28618,N_26764);
or UO_1945 (O_1945,N_28957,N_28876);
nor UO_1946 (O_1946,N_25397,N_29538);
and UO_1947 (O_1947,N_28927,N_28326);
nor UO_1948 (O_1948,N_25854,N_25905);
nor UO_1949 (O_1949,N_28838,N_28466);
or UO_1950 (O_1950,N_27913,N_26269);
nand UO_1951 (O_1951,N_29123,N_25655);
nand UO_1952 (O_1952,N_27545,N_29565);
and UO_1953 (O_1953,N_28330,N_27624);
nor UO_1954 (O_1954,N_25620,N_29852);
nor UO_1955 (O_1955,N_26267,N_28271);
xor UO_1956 (O_1956,N_27879,N_27263);
nor UO_1957 (O_1957,N_25416,N_26935);
or UO_1958 (O_1958,N_29156,N_28353);
nor UO_1959 (O_1959,N_26659,N_27923);
or UO_1960 (O_1960,N_26954,N_29059);
nor UO_1961 (O_1961,N_29173,N_28054);
nor UO_1962 (O_1962,N_27656,N_26804);
or UO_1963 (O_1963,N_28088,N_27899);
nor UO_1964 (O_1964,N_27027,N_28001);
nor UO_1965 (O_1965,N_25140,N_26965);
nand UO_1966 (O_1966,N_28309,N_25686);
and UO_1967 (O_1967,N_27761,N_28655);
and UO_1968 (O_1968,N_26564,N_29987);
nor UO_1969 (O_1969,N_26068,N_25292);
and UO_1970 (O_1970,N_27186,N_27938);
nand UO_1971 (O_1971,N_27607,N_25920);
nand UO_1972 (O_1972,N_26180,N_26403);
and UO_1973 (O_1973,N_28363,N_28104);
xor UO_1974 (O_1974,N_28709,N_27045);
nand UO_1975 (O_1975,N_25518,N_26502);
nand UO_1976 (O_1976,N_29966,N_26464);
nor UO_1977 (O_1977,N_28194,N_28277);
nand UO_1978 (O_1978,N_29640,N_28636);
and UO_1979 (O_1979,N_26805,N_29914);
or UO_1980 (O_1980,N_27844,N_29612);
nor UO_1981 (O_1981,N_25716,N_25312);
nand UO_1982 (O_1982,N_27137,N_29638);
or UO_1983 (O_1983,N_26414,N_27262);
nor UO_1984 (O_1984,N_28799,N_27645);
nand UO_1985 (O_1985,N_29581,N_28298);
nor UO_1986 (O_1986,N_28751,N_27504);
and UO_1987 (O_1987,N_26714,N_29770);
nor UO_1988 (O_1988,N_25087,N_29998);
and UO_1989 (O_1989,N_27302,N_29616);
and UO_1990 (O_1990,N_29169,N_28953);
nor UO_1991 (O_1991,N_29544,N_26070);
nor UO_1992 (O_1992,N_26431,N_27730);
and UO_1993 (O_1993,N_27180,N_26275);
or UO_1994 (O_1994,N_28041,N_25160);
nor UO_1995 (O_1995,N_27896,N_25609);
and UO_1996 (O_1996,N_26122,N_27753);
nand UO_1997 (O_1997,N_27853,N_28613);
nand UO_1998 (O_1998,N_29967,N_29351);
nor UO_1999 (O_1999,N_29080,N_25101);
and UO_2000 (O_2000,N_27840,N_25353);
nor UO_2001 (O_2001,N_28312,N_28148);
and UO_2002 (O_2002,N_25347,N_29610);
nand UO_2003 (O_2003,N_26442,N_25664);
or UO_2004 (O_2004,N_26731,N_26642);
or UO_2005 (O_2005,N_28342,N_26006);
nand UO_2006 (O_2006,N_27809,N_27178);
xnor UO_2007 (O_2007,N_28143,N_28666);
nand UO_2008 (O_2008,N_29663,N_25887);
xor UO_2009 (O_2009,N_25778,N_25581);
and UO_2010 (O_2010,N_27886,N_29336);
and UO_2011 (O_2011,N_25364,N_25098);
nand UO_2012 (O_2012,N_28879,N_25934);
nor UO_2013 (O_2013,N_26953,N_27535);
xnor UO_2014 (O_2014,N_25297,N_25413);
xnor UO_2015 (O_2015,N_28563,N_26577);
nand UO_2016 (O_2016,N_29977,N_27362);
nor UO_2017 (O_2017,N_28654,N_25945);
or UO_2018 (O_2018,N_25995,N_26565);
and UO_2019 (O_2019,N_26537,N_28237);
or UO_2020 (O_2020,N_26864,N_26145);
nand UO_2021 (O_2021,N_25467,N_27565);
nor UO_2022 (O_2022,N_29280,N_29515);
or UO_2023 (O_2023,N_26161,N_29850);
and UO_2024 (O_2024,N_29750,N_29621);
nor UO_2025 (O_2025,N_25435,N_28114);
or UO_2026 (O_2026,N_29054,N_26425);
xor UO_2027 (O_2027,N_29451,N_28792);
nor UO_2028 (O_2028,N_28315,N_29905);
and UO_2029 (O_2029,N_25257,N_26695);
and UO_2030 (O_2030,N_25269,N_26349);
nor UO_2031 (O_2031,N_27419,N_25680);
nor UO_2032 (O_2032,N_26980,N_27346);
nand UO_2033 (O_2033,N_29283,N_29131);
nor UO_2034 (O_2034,N_26630,N_28167);
or UO_2035 (O_2035,N_25029,N_28672);
nand UO_2036 (O_2036,N_26901,N_25985);
nand UO_2037 (O_2037,N_29928,N_26643);
nand UO_2038 (O_2038,N_27112,N_26220);
nand UO_2039 (O_2039,N_26615,N_26890);
nand UO_2040 (O_2040,N_29181,N_26700);
or UO_2041 (O_2041,N_25588,N_25694);
or UO_2042 (O_2042,N_25618,N_28833);
and UO_2043 (O_2043,N_29768,N_27540);
and UO_2044 (O_2044,N_28653,N_29024);
nand UO_2045 (O_2045,N_26443,N_29409);
or UO_2046 (O_2046,N_26796,N_29408);
or UO_2047 (O_2047,N_29310,N_29426);
or UO_2048 (O_2048,N_29075,N_26433);
nor UO_2049 (O_2049,N_27183,N_27748);
xor UO_2050 (O_2050,N_27772,N_28605);
and UO_2051 (O_2051,N_26632,N_26151);
nand UO_2052 (O_2052,N_25709,N_27451);
or UO_2053 (O_2053,N_25904,N_26970);
nand UO_2054 (O_2054,N_27552,N_28930);
or UO_2055 (O_2055,N_29491,N_25005);
and UO_2056 (O_2056,N_28904,N_29693);
nand UO_2057 (O_2057,N_27687,N_25535);
and UO_2058 (O_2058,N_28250,N_26518);
or UO_2059 (O_2059,N_29459,N_26940);
or UO_2060 (O_2060,N_26033,N_25241);
or UO_2061 (O_2061,N_29983,N_25696);
nor UO_2062 (O_2062,N_25248,N_27798);
or UO_2063 (O_2063,N_27481,N_25626);
or UO_2064 (O_2064,N_29061,N_27265);
and UO_2065 (O_2065,N_26654,N_26405);
nor UO_2066 (O_2066,N_27939,N_25563);
nor UO_2067 (O_2067,N_29250,N_28825);
xor UO_2068 (O_2068,N_28640,N_28937);
nor UO_2069 (O_2069,N_28066,N_29099);
or UO_2070 (O_2070,N_27118,N_26609);
nand UO_2071 (O_2071,N_28598,N_28362);
nor UO_2072 (O_2072,N_29445,N_29500);
and UO_2073 (O_2073,N_26822,N_27406);
or UO_2074 (O_2074,N_29592,N_25580);
nor UO_2075 (O_2075,N_29423,N_25853);
and UO_2076 (O_2076,N_29752,N_26498);
nand UO_2077 (O_2077,N_29585,N_25986);
or UO_2078 (O_2078,N_29383,N_25106);
xnor UO_2079 (O_2079,N_26232,N_25713);
nor UO_2080 (O_2080,N_25849,N_29232);
or UO_2081 (O_2081,N_28868,N_29652);
or UO_2082 (O_2082,N_27013,N_28659);
and UO_2083 (O_2083,N_27862,N_29496);
nand UO_2084 (O_2084,N_25712,N_25443);
nand UO_2085 (O_2085,N_28470,N_26783);
nor UO_2086 (O_2086,N_27012,N_27498);
or UO_2087 (O_2087,N_25767,N_25808);
and UO_2088 (O_2088,N_29482,N_28412);
xnor UO_2089 (O_2089,N_25856,N_25006);
nor UO_2090 (O_2090,N_26117,N_26515);
or UO_2091 (O_2091,N_29913,N_25601);
or UO_2092 (O_2092,N_26614,N_26048);
nand UO_2093 (O_2093,N_25504,N_29667);
xor UO_2094 (O_2094,N_29747,N_29016);
or UO_2095 (O_2095,N_28351,N_25690);
xnor UO_2096 (O_2096,N_29954,N_25559);
and UO_2097 (O_2097,N_25152,N_25536);
or UO_2098 (O_2098,N_27675,N_26870);
nand UO_2099 (O_2099,N_27715,N_25816);
xnor UO_2100 (O_2100,N_28040,N_25565);
nand UO_2101 (O_2101,N_27264,N_29539);
nand UO_2102 (O_2102,N_29660,N_28837);
nand UO_2103 (O_2103,N_26999,N_26799);
nor UO_2104 (O_2104,N_27563,N_29965);
nor UO_2105 (O_2105,N_29730,N_29069);
nor UO_2106 (O_2106,N_29684,N_29554);
and UO_2107 (O_2107,N_29244,N_28569);
and UO_2108 (O_2108,N_26277,N_26836);
nand UO_2109 (O_2109,N_28652,N_26000);
or UO_2110 (O_2110,N_29453,N_26911);
nor UO_2111 (O_2111,N_25754,N_29589);
or UO_2112 (O_2112,N_27212,N_28971);
and UO_2113 (O_2113,N_25770,N_26914);
nand UO_2114 (O_2114,N_27356,N_26762);
xor UO_2115 (O_2115,N_27386,N_26942);
and UO_2116 (O_2116,N_26858,N_28758);
nor UO_2117 (O_2117,N_29229,N_28113);
nand UO_2118 (O_2118,N_28663,N_28991);
xnor UO_2119 (O_2119,N_26594,N_26370);
nand UO_2120 (O_2120,N_27249,N_28161);
or UO_2121 (O_2121,N_26668,N_28916);
or UO_2122 (O_2122,N_25446,N_25219);
or UO_2123 (O_2123,N_28259,N_29563);
or UO_2124 (O_2124,N_25182,N_25924);
nand UO_2125 (O_2125,N_29958,N_27193);
nor UO_2126 (O_2126,N_25468,N_28853);
or UO_2127 (O_2127,N_25866,N_26172);
nand UO_2128 (O_2128,N_26270,N_27184);
nand UO_2129 (O_2129,N_28540,N_26596);
nor UO_2130 (O_2130,N_28086,N_27123);
nand UO_2131 (O_2131,N_25720,N_29177);
or UO_2132 (O_2132,N_28882,N_25242);
or UO_2133 (O_2133,N_26703,N_25362);
nand UO_2134 (O_2134,N_27181,N_28159);
nor UO_2135 (O_2135,N_28583,N_25956);
nor UO_2136 (O_2136,N_27684,N_28968);
nor UO_2137 (O_2137,N_28824,N_29754);
or UO_2138 (O_2138,N_26071,N_27606);
xor UO_2139 (O_2139,N_28187,N_27632);
or UO_2140 (O_2140,N_28524,N_29686);
or UO_2141 (O_2141,N_25847,N_29715);
nor UO_2142 (O_2142,N_26073,N_28301);
and UO_2143 (O_2143,N_28397,N_28030);
nor UO_2144 (O_2144,N_25605,N_28766);
nand UO_2145 (O_2145,N_28248,N_29299);
and UO_2146 (O_2146,N_25004,N_29207);
or UO_2147 (O_2147,N_27642,N_27828);
nand UO_2148 (O_2148,N_27847,N_25951);
and UO_2149 (O_2149,N_25411,N_25533);
and UO_2150 (O_2150,N_26116,N_26209);
and UO_2151 (O_2151,N_29642,N_25907);
nor UO_2152 (O_2152,N_28545,N_25812);
nor UO_2153 (O_2153,N_27904,N_25138);
nor UO_2154 (O_2154,N_29807,N_28302);
or UO_2155 (O_2155,N_28575,N_29090);
nand UO_2156 (O_2156,N_26167,N_29704);
or UO_2157 (O_2157,N_27256,N_25491);
or UO_2158 (O_2158,N_28308,N_26572);
nand UO_2159 (O_2159,N_28983,N_28355);
and UO_2160 (O_2160,N_28121,N_26329);
nand UO_2161 (O_2161,N_27964,N_25640);
and UO_2162 (O_2162,N_27732,N_28621);
nor UO_2163 (O_2163,N_28735,N_28272);
nand UO_2164 (O_2164,N_29771,N_28268);
xnor UO_2165 (O_2165,N_29431,N_25695);
and UO_2166 (O_2166,N_29180,N_29115);
nor UO_2167 (O_2167,N_25370,N_26800);
and UO_2168 (O_2168,N_26687,N_29263);
or UO_2169 (O_2169,N_26064,N_27720);
or UO_2170 (O_2170,N_29713,N_28458);
nand UO_2171 (O_2171,N_26421,N_27852);
nand UO_2172 (O_2172,N_27633,N_25702);
nor UO_2173 (O_2173,N_29112,N_28034);
or UO_2174 (O_2174,N_25516,N_29799);
or UO_2175 (O_2175,N_28754,N_27457);
or UO_2176 (O_2176,N_26325,N_27410);
xnor UO_2177 (O_2177,N_28938,N_26763);
xor UO_2178 (O_2178,N_28394,N_27328);
nand UO_2179 (O_2179,N_26931,N_29613);
nand UO_2180 (O_2180,N_26673,N_27870);
or UO_2181 (O_2181,N_27573,N_29238);
nor UO_2182 (O_2182,N_29739,N_28514);
nor UO_2183 (O_2183,N_28099,N_27479);
or UO_2184 (O_2184,N_28934,N_25885);
nor UO_2185 (O_2185,N_25453,N_26948);
nor UO_2186 (O_2186,N_28215,N_27877);
and UO_2187 (O_2187,N_29834,N_29742);
or UO_2188 (O_2188,N_26995,N_26486);
nand UO_2189 (O_2189,N_28587,N_25775);
xor UO_2190 (O_2190,N_26867,N_28859);
nand UO_2191 (O_2191,N_28016,N_28966);
or UO_2192 (O_2192,N_26472,N_25667);
and UO_2193 (O_2193,N_29632,N_26993);
and UO_2194 (O_2194,N_27694,N_25820);
or UO_2195 (O_2195,N_29934,N_29956);
and UO_2196 (O_2196,N_25611,N_26785);
nand UO_2197 (O_2197,N_29168,N_26426);
nor UO_2198 (O_2198,N_26445,N_28341);
nand UO_2199 (O_2199,N_29483,N_26903);
xnor UO_2200 (O_2200,N_28196,N_25658);
nand UO_2201 (O_2201,N_28069,N_29368);
nor UO_2202 (O_2202,N_27829,N_29659);
nand UO_2203 (O_2203,N_28505,N_29700);
nor UO_2204 (O_2204,N_26496,N_25630);
or UO_2205 (O_2205,N_25184,N_29380);
nand UO_2206 (O_2206,N_28922,N_25573);
xnor UO_2207 (O_2207,N_28453,N_25440);
nand UO_2208 (O_2208,N_25786,N_28339);
nor UO_2209 (O_2209,N_25263,N_27558);
nand UO_2210 (O_2210,N_28781,N_26918);
or UO_2211 (O_2211,N_28574,N_28046);
or UO_2212 (O_2212,N_29448,N_26660);
xnor UO_2213 (O_2213,N_27091,N_29908);
or UO_2214 (O_2214,N_26013,N_26280);
or UO_2215 (O_2215,N_29382,N_27566);
or UO_2216 (O_2216,N_29877,N_29161);
or UO_2217 (O_2217,N_29567,N_26988);
and UO_2218 (O_2218,N_25066,N_28501);
and UO_2219 (O_2219,N_27207,N_27009);
or UO_2220 (O_2220,N_26222,N_29159);
xnor UO_2221 (O_2221,N_25388,N_26511);
nand UO_2222 (O_2222,N_25789,N_29858);
xnor UO_2223 (O_2223,N_27692,N_25189);
nand UO_2224 (O_2224,N_26123,N_28225);
nand UO_2225 (O_2225,N_27719,N_27318);
and UO_2226 (O_2226,N_29133,N_26406);
or UO_2227 (O_2227,N_26259,N_25178);
nand UO_2228 (O_2228,N_26915,N_25204);
nand UO_2229 (O_2229,N_25821,N_28955);
nor UO_2230 (O_2230,N_27974,N_27298);
and UO_2231 (O_2231,N_28422,N_26711);
nand UO_2232 (O_2232,N_25405,N_25221);
and UO_2233 (O_2233,N_27384,N_29252);
and UO_2234 (O_2234,N_27104,N_29572);
xor UO_2235 (O_2235,N_26398,N_29857);
nor UO_2236 (O_2236,N_28178,N_29994);
nor UO_2237 (O_2237,N_25523,N_29337);
or UO_2238 (O_2238,N_26788,N_25008);
nand UO_2239 (O_2239,N_26702,N_25743);
or UO_2240 (O_2240,N_25447,N_29797);
xor UO_2241 (O_2241,N_25733,N_28465);
nand UO_2242 (O_2242,N_28434,N_28498);
nand UO_2243 (O_2243,N_28628,N_29820);
nor UO_2244 (O_2244,N_28136,N_27141);
nand UO_2245 (O_2245,N_26316,N_29604);
xnor UO_2246 (O_2246,N_28707,N_28317);
nand UO_2247 (O_2247,N_25768,N_29037);
nor UO_2248 (O_2248,N_28522,N_28842);
nand UO_2249 (O_2249,N_28154,N_28061);
nand UO_2250 (O_2250,N_28893,N_27267);
and UO_2251 (O_2251,N_28730,N_27636);
and UO_2252 (O_2252,N_27571,N_27378);
nor UO_2253 (O_2253,N_28123,N_26040);
and UO_2254 (O_2254,N_25054,N_25839);
xnor UO_2255 (O_2255,N_29597,N_26749);
nor UO_2256 (O_2256,N_25438,N_26221);
xnor UO_2257 (O_2257,N_27957,N_26037);
xor UO_2258 (O_2258,N_29142,N_26312);
nor UO_2259 (O_2259,N_28865,N_28184);
and UO_2260 (O_2260,N_27524,N_27144);
nor UO_2261 (O_2261,N_28801,N_29278);
and UO_2262 (O_2262,N_27696,N_29909);
and UO_2263 (O_2263,N_29825,N_26561);
and UO_2264 (O_2264,N_28153,N_25526);
or UO_2265 (O_2265,N_27929,N_28411);
nor UO_2266 (O_2266,N_29661,N_28790);
and UO_2267 (O_2267,N_28715,N_27475);
and UO_2268 (O_2268,N_26250,N_25020);
nor UO_2269 (O_2269,N_28964,N_27282);
nor UO_2270 (O_2270,N_25830,N_28982);
and UO_2271 (O_2271,N_29125,N_29815);
nand UO_2272 (O_2272,N_27047,N_27621);
or UO_2273 (O_2273,N_29879,N_28741);
nor UO_2274 (O_2274,N_27873,N_26581);
nand UO_2275 (O_2275,N_25562,N_27399);
or UO_2276 (O_2276,N_26623,N_28320);
xor UO_2277 (O_2277,N_28009,N_26026);
xnor UO_2278 (O_2278,N_29541,N_27679);
or UO_2279 (O_2279,N_28830,N_25530);
and UO_2280 (O_2280,N_28349,N_26880);
nor UO_2281 (O_2281,N_26479,N_25511);
nand UO_2282 (O_2282,N_29919,N_28606);
or UO_2283 (O_2283,N_27159,N_27643);
nand UO_2284 (O_2284,N_28207,N_27417);
and UO_2285 (O_2285,N_27024,N_26102);
nor UO_2286 (O_2286,N_26091,N_26514);
and UO_2287 (O_2287,N_26422,N_27176);
nor UO_2288 (O_2288,N_28967,N_29359);
and UO_2289 (O_2289,N_28840,N_26226);
nand UO_2290 (O_2290,N_29793,N_29493);
nand UO_2291 (O_2291,N_25615,N_29251);
and UO_2292 (O_2292,N_27751,N_27055);
nand UO_2293 (O_2293,N_28923,N_26960);
xor UO_2294 (O_2294,N_28728,N_25736);
xnor UO_2295 (O_2295,N_28770,N_27814);
or UO_2296 (O_2296,N_25404,N_28926);
nand UO_2297 (O_2297,N_26595,N_26143);
and UO_2298 (O_2298,N_27523,N_28595);
nor UO_2299 (O_2299,N_25025,N_25892);
nand UO_2300 (O_2300,N_27461,N_28451);
nor UO_2301 (O_2301,N_28947,N_28862);
or UO_2302 (O_2302,N_26849,N_28891);
or UO_2303 (O_2303,N_27779,N_27447);
or UO_2304 (O_2304,N_28047,N_29785);
nor UO_2305 (O_2305,N_26376,N_29388);
nor UO_2306 (O_2306,N_26268,N_26768);
nand UO_2307 (O_2307,N_29462,N_25037);
nand UO_2308 (O_2308,N_25177,N_29015);
nand UO_2309 (O_2309,N_26471,N_26968);
xor UO_2310 (O_2310,N_27412,N_26249);
nand UO_2311 (O_2311,N_26118,N_26927);
nor UO_2312 (O_2312,N_28779,N_28823);
or UO_2313 (O_2313,N_29018,N_25835);
or UO_2314 (O_2314,N_29000,N_28963);
nand UO_2315 (O_2315,N_29673,N_29564);
nand UO_2316 (O_2316,N_28176,N_28920);
nor UO_2317 (O_2317,N_27947,N_26448);
or UO_2318 (O_2318,N_28156,N_25682);
or UO_2319 (O_2319,N_29313,N_28760);
nand UO_2320 (O_2320,N_29603,N_28438);
xnor UO_2321 (O_2321,N_27868,N_28662);
and UO_2322 (O_2322,N_26372,N_29083);
nor UO_2323 (O_2323,N_25556,N_27932);
nor UO_2324 (O_2324,N_26987,N_29210);
or UO_2325 (O_2325,N_26142,N_25196);
nor UO_2326 (O_2326,N_25652,N_29321);
or UO_2327 (O_2327,N_29231,N_27148);
and UO_2328 (O_2328,N_29923,N_26473);
nor UO_2329 (O_2329,N_25294,N_28551);
or UO_2330 (O_2330,N_25503,N_27260);
nand UO_2331 (O_2331,N_29809,N_25374);
and UO_2332 (O_2332,N_28091,N_25815);
or UO_2333 (O_2333,N_25077,N_26494);
nor UO_2334 (O_2334,N_25790,N_25406);
or UO_2335 (O_2335,N_25980,N_26321);
nor UO_2336 (O_2336,N_26132,N_26024);
and UO_2337 (O_2337,N_26152,N_28467);
nand UO_2338 (O_2338,N_27505,N_26861);
nor UO_2339 (O_2339,N_28189,N_29233);
xnor UO_2340 (O_2340,N_26041,N_27299);
and UO_2341 (O_2341,N_27046,N_29324);
or UO_2342 (O_2342,N_25186,N_25430);
and UO_2343 (O_2343,N_29735,N_26171);
and UO_2344 (O_2344,N_28996,N_25095);
xnor UO_2345 (O_2345,N_27634,N_29227);
or UO_2346 (O_2346,N_25303,N_28615);
and UO_2347 (O_2347,N_29891,N_25732);
or UO_2348 (O_2348,N_28726,N_25639);
nand UO_2349 (O_2349,N_27577,N_27306);
nor UO_2350 (O_2350,N_27395,N_29369);
and UO_2351 (O_2351,N_25888,N_29828);
or UO_2352 (O_2352,N_27916,N_28291);
xnor UO_2353 (O_2353,N_25801,N_28071);
nand UO_2354 (O_2354,N_29349,N_29609);
and UO_2355 (O_2355,N_29421,N_27960);
nor UO_2356 (O_2356,N_29681,N_25571);
and UO_2357 (O_2357,N_28260,N_27759);
or UO_2358 (O_2358,N_25675,N_28701);
xnor UO_2359 (O_2359,N_28449,N_27018);
nand UO_2360 (O_2360,N_27086,N_25650);
nand UO_2361 (O_2361,N_28141,N_29599);
or UO_2362 (O_2362,N_25918,N_27038);
nand UO_2363 (O_2363,N_26320,N_28077);
nor UO_2364 (O_2364,N_25635,N_25205);
nand UO_2365 (O_2365,N_26831,N_26929);
or UO_2366 (O_2366,N_28346,N_29794);
xnor UO_2367 (O_2367,N_27816,N_25027);
xor UO_2368 (O_2368,N_25988,N_29505);
nand UO_2369 (O_2369,N_29414,N_28519);
nand UO_2370 (O_2370,N_27655,N_26705);
or UO_2371 (O_2371,N_26265,N_28703);
or UO_2372 (O_2372,N_26029,N_28460);
nor UO_2373 (O_2373,N_28710,N_27139);
nand UO_2374 (O_2374,N_29494,N_27382);
and UO_2375 (O_2375,N_25076,N_29241);
nor UO_2376 (O_2376,N_27343,N_28410);
nand UO_2377 (O_2377,N_27458,N_28385);
nor UO_2378 (O_2378,N_27341,N_29364);
or UO_2379 (O_2379,N_28705,N_25442);
nor UO_2380 (O_2380,N_26239,N_28774);
nand UO_2381 (O_2381,N_27442,N_27368);
nor UO_2382 (O_2382,N_25017,N_27062);
nand UO_2383 (O_2383,N_25240,N_28265);
and UO_2384 (O_2384,N_28322,N_28591);
nor UO_2385 (O_2385,N_28371,N_28635);
nor UO_2386 (O_2386,N_28115,N_29677);
and UO_2387 (O_2387,N_26109,N_25166);
or UO_2388 (O_2388,N_27878,N_26389);
or UO_2389 (O_2389,N_25763,N_29166);
nand UO_2390 (O_2390,N_27167,N_29753);
nand UO_2391 (O_2391,N_26950,N_28295);
nand UO_2392 (O_2392,N_28736,N_25873);
nor UO_2393 (O_2393,N_29376,N_25324);
xor UO_2394 (O_2394,N_28359,N_27962);
nor UO_2395 (O_2395,N_25792,N_28017);
nand UO_2396 (O_2396,N_26682,N_25117);
nand UO_2397 (O_2397,N_25180,N_25940);
and UO_2398 (O_2398,N_29727,N_28288);
or UO_2399 (O_2399,N_26752,N_27156);
nand UO_2400 (O_2400,N_29726,N_28502);
nand UO_2401 (O_2401,N_27131,N_27374);
nor UO_2402 (O_2402,N_27576,N_27784);
nor UO_2403 (O_2403,N_29460,N_27660);
and UO_2404 (O_2404,N_29205,N_28753);
nand UO_2405 (O_2405,N_29997,N_26939);
or UO_2406 (O_2406,N_26877,N_26945);
nor UO_2407 (O_2407,N_25831,N_29134);
and UO_2408 (O_2408,N_26845,N_25584);
and UO_2409 (O_2409,N_29626,N_26556);
nor UO_2410 (O_2410,N_28081,N_28623);
or UO_2411 (O_2411,N_29127,N_25237);
or UO_2412 (O_2412,N_26922,N_29641);
nand UO_2413 (O_2413,N_28797,N_29856);
and UO_2414 (O_2414,N_26106,N_27061);
xor UO_2415 (O_2415,N_27680,N_27717);
nand UO_2416 (O_2416,N_26983,N_28881);
nor UO_2417 (O_2417,N_29356,N_28721);
nor UO_2418 (O_2418,N_25064,N_29761);
nor UO_2419 (O_2419,N_27010,N_28791);
and UO_2420 (O_2420,N_29151,N_28012);
nand UO_2421 (O_2421,N_29485,N_29235);
or UO_2422 (O_2422,N_26367,N_27158);
nor UO_2423 (O_2423,N_25942,N_28910);
or UO_2424 (O_2424,N_27556,N_29769);
nor UO_2425 (O_2425,N_25949,N_27035);
nand UO_2426 (O_2426,N_26087,N_28180);
or UO_2427 (O_2427,N_25073,N_27133);
nor UO_2428 (O_2428,N_28513,N_27432);
or UO_2429 (O_2429,N_27165,N_25944);
and UO_2430 (O_2430,N_29063,N_29051);
and UO_2431 (O_2431,N_28125,N_26838);
or UO_2432 (O_2432,N_28935,N_25663);
nor UO_2433 (O_2433,N_27697,N_26467);
nand UO_2434 (O_2434,N_29111,N_29004);
or UO_2435 (O_2435,N_29242,N_27429);
xor UO_2436 (O_2436,N_28745,N_26624);
or UO_2437 (O_2437,N_25490,N_25157);
nor UO_2438 (O_2438,N_25200,N_26136);
nor UO_2439 (O_2439,N_29979,N_29171);
xnor UO_2440 (O_2440,N_26099,N_26602);
nand UO_2441 (O_2441,N_25441,N_25125);
or UO_2442 (O_2442,N_27486,N_27824);
nor UO_2443 (O_2443,N_29005,N_26815);
nor UO_2444 (O_2444,N_27514,N_28258);
nand UO_2445 (O_2445,N_29776,N_27464);
xnor UO_2446 (O_2446,N_26273,N_25602);
nor UO_2447 (O_2447,N_27446,N_25250);
nor UO_2448 (O_2448,N_27740,N_25539);
and UO_2449 (O_2449,N_27337,N_25923);
or UO_2450 (O_2450,N_28708,N_26207);
nor UO_2451 (O_2451,N_26279,N_29957);
or UO_2452 (O_2452,N_29859,N_28418);
and UO_2453 (O_2453,N_28917,N_29692);
nand UO_2454 (O_2454,N_29653,N_25656);
or UO_2455 (O_2455,N_25850,N_26343);
nand UO_2456 (O_2456,N_29167,N_28608);
nor UO_2457 (O_2457,N_27729,N_29006);
nand UO_2458 (O_2458,N_26713,N_28846);
and UO_2459 (O_2459,N_25245,N_28198);
xor UO_2460 (O_2460,N_25726,N_29298);
or UO_2461 (O_2461,N_27752,N_25514);
nor UO_2462 (O_2462,N_25049,N_26135);
xnor UO_2463 (O_2463,N_28900,N_26294);
nand UO_2464 (O_2464,N_25223,N_26589);
nor UO_2465 (O_2465,N_25295,N_25042);
nor UO_2466 (O_2466,N_28131,N_26138);
and UO_2467 (O_2467,N_28950,N_27448);
nand UO_2468 (O_2468,N_25190,N_26974);
or UO_2469 (O_2469,N_26375,N_27354);
nor UO_2470 (O_2470,N_26237,N_25472);
nor UO_2471 (O_2471,N_25538,N_25224);
xor UO_2472 (O_2472,N_29619,N_27379);
or UO_2473 (O_2473,N_25418,N_28548);
or UO_2474 (O_2474,N_26667,N_27769);
and UO_2475 (O_2475,N_28600,N_29552);
nand UO_2476 (O_2476,N_29930,N_25840);
or UO_2477 (O_2477,N_28664,N_29533);
nor UO_2478 (O_2478,N_28390,N_26444);
or UO_2479 (O_2479,N_28226,N_26566);
or UO_2480 (O_2480,N_29881,N_28998);
and UO_2481 (O_2481,N_25273,N_25335);
or UO_2482 (O_2482,N_29548,N_26416);
xor UO_2483 (O_2483,N_28717,N_25700);
or UO_2484 (O_2484,N_29316,N_28110);
and UO_2485 (O_2485,N_27746,N_28990);
nor UO_2486 (O_2486,N_29775,N_25692);
nor UO_2487 (O_2487,N_28977,N_29545);
nand UO_2488 (O_2488,N_28142,N_25782);
nand UO_2489 (O_2489,N_25300,N_25810);
nand UO_2490 (O_2490,N_27531,N_27203);
xnor UO_2491 (O_2491,N_25715,N_25929);
and UO_2492 (O_2492,N_27101,N_25915);
or UO_2493 (O_2493,N_27296,N_29971);
nor UO_2494 (O_2494,N_28517,N_29158);
nor UO_2495 (O_2495,N_28516,N_27220);
nand UO_2496 (O_2496,N_26390,N_25302);
nand UO_2497 (O_2497,N_28425,N_26819);
and UO_2498 (O_2498,N_26154,N_25722);
nand UO_2499 (O_2499,N_26292,N_26281);
or UO_2500 (O_2500,N_29176,N_27357);
nor UO_2501 (O_2501,N_27913,N_26320);
or UO_2502 (O_2502,N_26944,N_28384);
or UO_2503 (O_2503,N_28190,N_27426);
nor UO_2504 (O_2504,N_26243,N_25122);
and UO_2505 (O_2505,N_29075,N_26382);
and UO_2506 (O_2506,N_27498,N_27391);
nor UO_2507 (O_2507,N_25525,N_26633);
xnor UO_2508 (O_2508,N_26635,N_28164);
or UO_2509 (O_2509,N_29608,N_25723);
xor UO_2510 (O_2510,N_25457,N_27651);
and UO_2511 (O_2511,N_25421,N_26460);
or UO_2512 (O_2512,N_28136,N_28842);
and UO_2513 (O_2513,N_29069,N_28533);
xnor UO_2514 (O_2514,N_26713,N_28808);
nand UO_2515 (O_2515,N_27448,N_28071);
or UO_2516 (O_2516,N_26642,N_27396);
nand UO_2517 (O_2517,N_29928,N_29419);
nor UO_2518 (O_2518,N_29672,N_27892);
xnor UO_2519 (O_2519,N_25548,N_29669);
or UO_2520 (O_2520,N_25262,N_26988);
nor UO_2521 (O_2521,N_25466,N_26621);
nand UO_2522 (O_2522,N_27652,N_25774);
or UO_2523 (O_2523,N_26967,N_25583);
or UO_2524 (O_2524,N_25291,N_26063);
or UO_2525 (O_2525,N_29441,N_29642);
nor UO_2526 (O_2526,N_27993,N_28511);
or UO_2527 (O_2527,N_26520,N_25629);
or UO_2528 (O_2528,N_27813,N_26096);
or UO_2529 (O_2529,N_29162,N_26334);
nand UO_2530 (O_2530,N_27690,N_26917);
and UO_2531 (O_2531,N_27958,N_29619);
and UO_2532 (O_2532,N_28663,N_26856);
nand UO_2533 (O_2533,N_26037,N_28321);
or UO_2534 (O_2534,N_26432,N_28180);
nor UO_2535 (O_2535,N_26203,N_26427);
or UO_2536 (O_2536,N_25025,N_29240);
and UO_2537 (O_2537,N_26713,N_29116);
nand UO_2538 (O_2538,N_29892,N_29142);
nand UO_2539 (O_2539,N_26042,N_29330);
nor UO_2540 (O_2540,N_26654,N_25922);
and UO_2541 (O_2541,N_26714,N_27414);
and UO_2542 (O_2542,N_27615,N_28760);
nor UO_2543 (O_2543,N_27248,N_27808);
nand UO_2544 (O_2544,N_26354,N_28432);
nor UO_2545 (O_2545,N_29087,N_29820);
nand UO_2546 (O_2546,N_29993,N_28677);
nand UO_2547 (O_2547,N_29188,N_28909);
or UO_2548 (O_2548,N_26047,N_25704);
or UO_2549 (O_2549,N_28077,N_26151);
xor UO_2550 (O_2550,N_27009,N_25156);
nor UO_2551 (O_2551,N_28671,N_26546);
or UO_2552 (O_2552,N_25098,N_29822);
and UO_2553 (O_2553,N_28039,N_25429);
nand UO_2554 (O_2554,N_26748,N_29142);
nand UO_2555 (O_2555,N_26503,N_28621);
nand UO_2556 (O_2556,N_27970,N_27247);
or UO_2557 (O_2557,N_28228,N_25793);
or UO_2558 (O_2558,N_26624,N_26821);
nor UO_2559 (O_2559,N_26660,N_28558);
nand UO_2560 (O_2560,N_25497,N_29237);
and UO_2561 (O_2561,N_28642,N_28212);
nor UO_2562 (O_2562,N_27333,N_28987);
nand UO_2563 (O_2563,N_28209,N_27725);
or UO_2564 (O_2564,N_27718,N_28297);
xor UO_2565 (O_2565,N_28992,N_28747);
or UO_2566 (O_2566,N_25078,N_27507);
nand UO_2567 (O_2567,N_26089,N_25456);
xnor UO_2568 (O_2568,N_26449,N_26325);
nand UO_2569 (O_2569,N_26275,N_29189);
or UO_2570 (O_2570,N_25741,N_27785);
nor UO_2571 (O_2571,N_27308,N_29976);
nand UO_2572 (O_2572,N_26796,N_28842);
nand UO_2573 (O_2573,N_27929,N_27379);
or UO_2574 (O_2574,N_29574,N_25413);
or UO_2575 (O_2575,N_25173,N_29329);
nor UO_2576 (O_2576,N_28759,N_29567);
nand UO_2577 (O_2577,N_25762,N_26769);
or UO_2578 (O_2578,N_27993,N_26499);
nand UO_2579 (O_2579,N_26029,N_28591);
and UO_2580 (O_2580,N_28603,N_27479);
and UO_2581 (O_2581,N_28944,N_28276);
nor UO_2582 (O_2582,N_28777,N_28457);
nand UO_2583 (O_2583,N_25656,N_29492);
nor UO_2584 (O_2584,N_29212,N_26596);
and UO_2585 (O_2585,N_26206,N_29103);
nand UO_2586 (O_2586,N_27253,N_25598);
or UO_2587 (O_2587,N_25556,N_26567);
nor UO_2588 (O_2588,N_26843,N_29493);
or UO_2589 (O_2589,N_28674,N_29112);
and UO_2590 (O_2590,N_27850,N_29810);
nand UO_2591 (O_2591,N_27683,N_26966);
nor UO_2592 (O_2592,N_29303,N_28574);
nand UO_2593 (O_2593,N_26483,N_25779);
nand UO_2594 (O_2594,N_27514,N_28328);
xor UO_2595 (O_2595,N_29523,N_29446);
nor UO_2596 (O_2596,N_28551,N_27205);
xor UO_2597 (O_2597,N_28658,N_29172);
nor UO_2598 (O_2598,N_25553,N_26033);
and UO_2599 (O_2599,N_25251,N_25774);
or UO_2600 (O_2600,N_25568,N_28028);
nor UO_2601 (O_2601,N_25774,N_26819);
and UO_2602 (O_2602,N_27303,N_29842);
nor UO_2603 (O_2603,N_27095,N_27699);
and UO_2604 (O_2604,N_27081,N_25614);
and UO_2605 (O_2605,N_25085,N_27211);
and UO_2606 (O_2606,N_28812,N_28604);
or UO_2607 (O_2607,N_25185,N_28253);
nor UO_2608 (O_2608,N_25393,N_27473);
nor UO_2609 (O_2609,N_27942,N_26389);
nor UO_2610 (O_2610,N_27439,N_29014);
and UO_2611 (O_2611,N_28944,N_29914);
and UO_2612 (O_2612,N_27674,N_28393);
nor UO_2613 (O_2613,N_28508,N_29304);
nor UO_2614 (O_2614,N_25649,N_29665);
nand UO_2615 (O_2615,N_29698,N_26918);
nand UO_2616 (O_2616,N_26046,N_25746);
nor UO_2617 (O_2617,N_28001,N_28712);
nand UO_2618 (O_2618,N_27658,N_29815);
nor UO_2619 (O_2619,N_28687,N_27745);
xnor UO_2620 (O_2620,N_27511,N_25655);
nand UO_2621 (O_2621,N_25317,N_28084);
xor UO_2622 (O_2622,N_27276,N_27158);
nor UO_2623 (O_2623,N_27228,N_25017);
xnor UO_2624 (O_2624,N_27960,N_29906);
xnor UO_2625 (O_2625,N_25877,N_28583);
or UO_2626 (O_2626,N_26949,N_27368);
xor UO_2627 (O_2627,N_28106,N_29797);
xor UO_2628 (O_2628,N_28858,N_26363);
nand UO_2629 (O_2629,N_29425,N_26213);
and UO_2630 (O_2630,N_26430,N_29426);
or UO_2631 (O_2631,N_29614,N_29214);
and UO_2632 (O_2632,N_26183,N_28366);
nor UO_2633 (O_2633,N_27552,N_26985);
nand UO_2634 (O_2634,N_28520,N_26353);
xor UO_2635 (O_2635,N_29461,N_28250);
and UO_2636 (O_2636,N_25078,N_25268);
or UO_2637 (O_2637,N_28469,N_26108);
or UO_2638 (O_2638,N_25155,N_27467);
nand UO_2639 (O_2639,N_25689,N_28681);
nor UO_2640 (O_2640,N_26605,N_28547);
xnor UO_2641 (O_2641,N_26390,N_28277);
nor UO_2642 (O_2642,N_29892,N_29572);
and UO_2643 (O_2643,N_28371,N_28763);
nand UO_2644 (O_2644,N_29851,N_26627);
nor UO_2645 (O_2645,N_27712,N_25796);
xnor UO_2646 (O_2646,N_29188,N_27663);
and UO_2647 (O_2647,N_26268,N_29164);
or UO_2648 (O_2648,N_26126,N_25377);
nor UO_2649 (O_2649,N_29504,N_26630);
and UO_2650 (O_2650,N_25836,N_27855);
xor UO_2651 (O_2651,N_25612,N_26444);
nand UO_2652 (O_2652,N_29475,N_25246);
and UO_2653 (O_2653,N_28814,N_28411);
or UO_2654 (O_2654,N_25056,N_28239);
and UO_2655 (O_2655,N_26333,N_27934);
nand UO_2656 (O_2656,N_29670,N_29354);
nor UO_2657 (O_2657,N_25049,N_28865);
and UO_2658 (O_2658,N_28514,N_28843);
or UO_2659 (O_2659,N_28805,N_29951);
nor UO_2660 (O_2660,N_28116,N_26556);
xor UO_2661 (O_2661,N_25538,N_29549);
or UO_2662 (O_2662,N_29300,N_25978);
or UO_2663 (O_2663,N_26928,N_26178);
nor UO_2664 (O_2664,N_26558,N_29965);
and UO_2665 (O_2665,N_25674,N_28720);
and UO_2666 (O_2666,N_25756,N_29340);
nand UO_2667 (O_2667,N_25371,N_28712);
nor UO_2668 (O_2668,N_29192,N_29489);
or UO_2669 (O_2669,N_27032,N_27096);
nand UO_2670 (O_2670,N_29541,N_27975);
nor UO_2671 (O_2671,N_28994,N_29093);
or UO_2672 (O_2672,N_27617,N_26104);
nand UO_2673 (O_2673,N_28340,N_26131);
nand UO_2674 (O_2674,N_29499,N_29479);
or UO_2675 (O_2675,N_28430,N_28985);
or UO_2676 (O_2676,N_28689,N_29914);
nor UO_2677 (O_2677,N_26984,N_25247);
nand UO_2678 (O_2678,N_29946,N_27500);
nand UO_2679 (O_2679,N_28351,N_28690);
and UO_2680 (O_2680,N_28258,N_28540);
or UO_2681 (O_2681,N_29960,N_25095);
or UO_2682 (O_2682,N_27513,N_27548);
nor UO_2683 (O_2683,N_28318,N_29893);
nor UO_2684 (O_2684,N_27211,N_28788);
nor UO_2685 (O_2685,N_29564,N_26462);
or UO_2686 (O_2686,N_25609,N_28505);
xnor UO_2687 (O_2687,N_28314,N_29619);
nand UO_2688 (O_2688,N_26586,N_28972);
nand UO_2689 (O_2689,N_27159,N_27794);
and UO_2690 (O_2690,N_27513,N_26870);
or UO_2691 (O_2691,N_29671,N_29355);
nand UO_2692 (O_2692,N_27911,N_27286);
or UO_2693 (O_2693,N_25055,N_28826);
or UO_2694 (O_2694,N_27102,N_27082);
nor UO_2695 (O_2695,N_28492,N_29229);
nor UO_2696 (O_2696,N_29442,N_25466);
and UO_2697 (O_2697,N_25537,N_25078);
and UO_2698 (O_2698,N_27261,N_28097);
nand UO_2699 (O_2699,N_27038,N_29611);
or UO_2700 (O_2700,N_25232,N_27390);
nand UO_2701 (O_2701,N_29789,N_28632);
and UO_2702 (O_2702,N_25003,N_28624);
or UO_2703 (O_2703,N_26251,N_25649);
or UO_2704 (O_2704,N_27555,N_26615);
nor UO_2705 (O_2705,N_26514,N_29471);
and UO_2706 (O_2706,N_29007,N_25783);
nor UO_2707 (O_2707,N_25631,N_25470);
xnor UO_2708 (O_2708,N_29319,N_28217);
and UO_2709 (O_2709,N_28022,N_28267);
or UO_2710 (O_2710,N_26909,N_25404);
xnor UO_2711 (O_2711,N_29302,N_28090);
or UO_2712 (O_2712,N_26124,N_29552);
xor UO_2713 (O_2713,N_28919,N_26688);
nand UO_2714 (O_2714,N_28507,N_28620);
nand UO_2715 (O_2715,N_25415,N_27567);
nand UO_2716 (O_2716,N_27767,N_29339);
or UO_2717 (O_2717,N_25877,N_28541);
nor UO_2718 (O_2718,N_27131,N_29062);
or UO_2719 (O_2719,N_27492,N_29842);
or UO_2720 (O_2720,N_26848,N_25701);
nor UO_2721 (O_2721,N_25016,N_25401);
and UO_2722 (O_2722,N_29920,N_27207);
and UO_2723 (O_2723,N_28860,N_25422);
or UO_2724 (O_2724,N_28583,N_27966);
or UO_2725 (O_2725,N_29918,N_28252);
xor UO_2726 (O_2726,N_26347,N_27172);
nand UO_2727 (O_2727,N_28319,N_27018);
xnor UO_2728 (O_2728,N_27581,N_28119);
xnor UO_2729 (O_2729,N_28002,N_27429);
nor UO_2730 (O_2730,N_25637,N_27954);
nand UO_2731 (O_2731,N_26475,N_26332);
and UO_2732 (O_2732,N_25474,N_29301);
nor UO_2733 (O_2733,N_25047,N_29499);
or UO_2734 (O_2734,N_27875,N_26494);
nor UO_2735 (O_2735,N_29998,N_25175);
or UO_2736 (O_2736,N_26723,N_27255);
nand UO_2737 (O_2737,N_25286,N_29609);
nand UO_2738 (O_2738,N_28063,N_27885);
or UO_2739 (O_2739,N_25573,N_28250);
or UO_2740 (O_2740,N_26479,N_28863);
or UO_2741 (O_2741,N_26662,N_29036);
and UO_2742 (O_2742,N_28728,N_25244);
and UO_2743 (O_2743,N_28940,N_26167);
and UO_2744 (O_2744,N_28128,N_27189);
nand UO_2745 (O_2745,N_26247,N_27991);
xnor UO_2746 (O_2746,N_29348,N_25660);
nor UO_2747 (O_2747,N_27031,N_25807);
nor UO_2748 (O_2748,N_28443,N_29071);
or UO_2749 (O_2749,N_25766,N_25780);
xor UO_2750 (O_2750,N_26480,N_28023);
or UO_2751 (O_2751,N_26325,N_27352);
and UO_2752 (O_2752,N_28585,N_26096);
and UO_2753 (O_2753,N_28598,N_25144);
nand UO_2754 (O_2754,N_28525,N_26379);
nor UO_2755 (O_2755,N_28636,N_29680);
nand UO_2756 (O_2756,N_27573,N_25721);
nor UO_2757 (O_2757,N_25904,N_26404);
or UO_2758 (O_2758,N_28303,N_28546);
and UO_2759 (O_2759,N_29853,N_28906);
nand UO_2760 (O_2760,N_27910,N_28801);
xnor UO_2761 (O_2761,N_28480,N_26242);
nor UO_2762 (O_2762,N_28254,N_26161);
and UO_2763 (O_2763,N_26886,N_26750);
and UO_2764 (O_2764,N_25686,N_27694);
or UO_2765 (O_2765,N_27586,N_25824);
and UO_2766 (O_2766,N_25496,N_29852);
and UO_2767 (O_2767,N_25217,N_27798);
xnor UO_2768 (O_2768,N_27536,N_28035);
nor UO_2769 (O_2769,N_25428,N_29016);
or UO_2770 (O_2770,N_25325,N_27893);
and UO_2771 (O_2771,N_26779,N_29554);
and UO_2772 (O_2772,N_26805,N_27460);
xor UO_2773 (O_2773,N_25596,N_26465);
nand UO_2774 (O_2774,N_26255,N_28096);
nor UO_2775 (O_2775,N_28239,N_26665);
nor UO_2776 (O_2776,N_28966,N_26141);
or UO_2777 (O_2777,N_26805,N_26079);
nand UO_2778 (O_2778,N_26170,N_26558);
and UO_2779 (O_2779,N_26438,N_25052);
nor UO_2780 (O_2780,N_29634,N_29163);
nand UO_2781 (O_2781,N_26159,N_27084);
nor UO_2782 (O_2782,N_29900,N_26083);
nand UO_2783 (O_2783,N_26291,N_29529);
xnor UO_2784 (O_2784,N_27409,N_26206);
and UO_2785 (O_2785,N_26750,N_29726);
xor UO_2786 (O_2786,N_28294,N_28340);
and UO_2787 (O_2787,N_28879,N_27775);
and UO_2788 (O_2788,N_28781,N_27655);
or UO_2789 (O_2789,N_29108,N_26225);
nand UO_2790 (O_2790,N_25647,N_25058);
and UO_2791 (O_2791,N_28842,N_25596);
and UO_2792 (O_2792,N_29544,N_25751);
nor UO_2793 (O_2793,N_27676,N_28275);
nand UO_2794 (O_2794,N_28149,N_29394);
nor UO_2795 (O_2795,N_25550,N_27179);
and UO_2796 (O_2796,N_26050,N_29286);
xnor UO_2797 (O_2797,N_28870,N_25942);
nand UO_2798 (O_2798,N_29423,N_28919);
nand UO_2799 (O_2799,N_26783,N_28322);
xor UO_2800 (O_2800,N_29667,N_29452);
nor UO_2801 (O_2801,N_28346,N_26310);
and UO_2802 (O_2802,N_29131,N_28041);
or UO_2803 (O_2803,N_28930,N_28167);
xnor UO_2804 (O_2804,N_28909,N_26233);
nand UO_2805 (O_2805,N_29832,N_26480);
nand UO_2806 (O_2806,N_26699,N_25545);
nor UO_2807 (O_2807,N_26048,N_28019);
nand UO_2808 (O_2808,N_29061,N_29514);
nand UO_2809 (O_2809,N_27037,N_27543);
and UO_2810 (O_2810,N_29711,N_26344);
nor UO_2811 (O_2811,N_29446,N_28245);
and UO_2812 (O_2812,N_27788,N_29156);
and UO_2813 (O_2813,N_28684,N_29775);
nand UO_2814 (O_2814,N_27047,N_28477);
nor UO_2815 (O_2815,N_27264,N_28549);
or UO_2816 (O_2816,N_26585,N_29237);
and UO_2817 (O_2817,N_29473,N_29163);
nand UO_2818 (O_2818,N_27919,N_29406);
and UO_2819 (O_2819,N_28572,N_25965);
or UO_2820 (O_2820,N_25124,N_25120);
and UO_2821 (O_2821,N_27356,N_28659);
or UO_2822 (O_2822,N_29063,N_27410);
or UO_2823 (O_2823,N_28179,N_28952);
or UO_2824 (O_2824,N_27918,N_27993);
nand UO_2825 (O_2825,N_25876,N_26690);
and UO_2826 (O_2826,N_26005,N_25497);
and UO_2827 (O_2827,N_28258,N_28025);
nand UO_2828 (O_2828,N_28572,N_27037);
nor UO_2829 (O_2829,N_26444,N_28566);
nor UO_2830 (O_2830,N_27321,N_28402);
and UO_2831 (O_2831,N_28329,N_26922);
nand UO_2832 (O_2832,N_26972,N_26799);
and UO_2833 (O_2833,N_29394,N_25976);
or UO_2834 (O_2834,N_27323,N_26600);
nor UO_2835 (O_2835,N_28972,N_25578);
or UO_2836 (O_2836,N_25771,N_29050);
and UO_2837 (O_2837,N_25244,N_27449);
nor UO_2838 (O_2838,N_25926,N_26577);
and UO_2839 (O_2839,N_25751,N_28213);
or UO_2840 (O_2840,N_27247,N_27007);
and UO_2841 (O_2841,N_28325,N_25820);
xnor UO_2842 (O_2842,N_26086,N_25416);
nor UO_2843 (O_2843,N_25154,N_26998);
and UO_2844 (O_2844,N_28365,N_28402);
nand UO_2845 (O_2845,N_26309,N_25869);
nand UO_2846 (O_2846,N_25759,N_26423);
nand UO_2847 (O_2847,N_26269,N_27953);
or UO_2848 (O_2848,N_28423,N_25730);
nor UO_2849 (O_2849,N_28133,N_25078);
and UO_2850 (O_2850,N_28056,N_25600);
nand UO_2851 (O_2851,N_25058,N_29244);
or UO_2852 (O_2852,N_28887,N_29214);
nand UO_2853 (O_2853,N_28421,N_27724);
and UO_2854 (O_2854,N_25005,N_28518);
or UO_2855 (O_2855,N_28499,N_26472);
and UO_2856 (O_2856,N_29242,N_27131);
or UO_2857 (O_2857,N_29304,N_29200);
nand UO_2858 (O_2858,N_27706,N_26377);
or UO_2859 (O_2859,N_28251,N_26816);
nor UO_2860 (O_2860,N_29232,N_26676);
xnor UO_2861 (O_2861,N_26494,N_25858);
nor UO_2862 (O_2862,N_28148,N_27328);
nand UO_2863 (O_2863,N_25889,N_29504);
or UO_2864 (O_2864,N_25696,N_25255);
and UO_2865 (O_2865,N_29750,N_28374);
nand UO_2866 (O_2866,N_29420,N_28981);
or UO_2867 (O_2867,N_29866,N_29089);
nor UO_2868 (O_2868,N_28232,N_27813);
nor UO_2869 (O_2869,N_26730,N_26251);
nand UO_2870 (O_2870,N_27155,N_28675);
xnor UO_2871 (O_2871,N_25626,N_27523);
xnor UO_2872 (O_2872,N_29745,N_26784);
and UO_2873 (O_2873,N_26771,N_26617);
nor UO_2874 (O_2874,N_27784,N_28769);
or UO_2875 (O_2875,N_28408,N_28254);
nand UO_2876 (O_2876,N_25835,N_25808);
or UO_2877 (O_2877,N_29168,N_28024);
and UO_2878 (O_2878,N_25204,N_29710);
or UO_2879 (O_2879,N_27376,N_28998);
nand UO_2880 (O_2880,N_27778,N_27206);
nor UO_2881 (O_2881,N_29876,N_26038);
nor UO_2882 (O_2882,N_25798,N_27412);
and UO_2883 (O_2883,N_25201,N_29940);
xor UO_2884 (O_2884,N_27741,N_25607);
nor UO_2885 (O_2885,N_26891,N_28589);
nor UO_2886 (O_2886,N_25156,N_29666);
and UO_2887 (O_2887,N_25038,N_25711);
and UO_2888 (O_2888,N_25556,N_28579);
and UO_2889 (O_2889,N_29793,N_27515);
nand UO_2890 (O_2890,N_26624,N_25504);
nand UO_2891 (O_2891,N_28854,N_28824);
xnor UO_2892 (O_2892,N_29662,N_28532);
and UO_2893 (O_2893,N_26560,N_26017);
xnor UO_2894 (O_2894,N_26524,N_26976);
and UO_2895 (O_2895,N_27027,N_29631);
nor UO_2896 (O_2896,N_28832,N_27581);
nor UO_2897 (O_2897,N_29015,N_25463);
xor UO_2898 (O_2898,N_25716,N_29166);
xnor UO_2899 (O_2899,N_25936,N_29649);
or UO_2900 (O_2900,N_25243,N_29780);
xor UO_2901 (O_2901,N_28375,N_25212);
or UO_2902 (O_2902,N_27207,N_25788);
and UO_2903 (O_2903,N_25549,N_25236);
or UO_2904 (O_2904,N_29022,N_29696);
and UO_2905 (O_2905,N_29000,N_26187);
nor UO_2906 (O_2906,N_26329,N_29364);
nor UO_2907 (O_2907,N_27205,N_25783);
or UO_2908 (O_2908,N_25856,N_29859);
nor UO_2909 (O_2909,N_29170,N_25512);
or UO_2910 (O_2910,N_28386,N_27403);
nand UO_2911 (O_2911,N_26995,N_27451);
nor UO_2912 (O_2912,N_26930,N_27037);
or UO_2913 (O_2913,N_28226,N_28171);
or UO_2914 (O_2914,N_28831,N_28989);
or UO_2915 (O_2915,N_29871,N_26607);
and UO_2916 (O_2916,N_26385,N_28608);
nor UO_2917 (O_2917,N_28886,N_26664);
or UO_2918 (O_2918,N_25149,N_25955);
nor UO_2919 (O_2919,N_25461,N_25106);
or UO_2920 (O_2920,N_28610,N_28051);
or UO_2921 (O_2921,N_28073,N_28016);
nand UO_2922 (O_2922,N_27202,N_27165);
or UO_2923 (O_2923,N_29916,N_28534);
xnor UO_2924 (O_2924,N_28668,N_27471);
nor UO_2925 (O_2925,N_28046,N_25649);
nor UO_2926 (O_2926,N_25617,N_29343);
nor UO_2927 (O_2927,N_26617,N_27097);
nor UO_2928 (O_2928,N_29651,N_27936);
xnor UO_2929 (O_2929,N_26977,N_25100);
nand UO_2930 (O_2930,N_25662,N_27932);
nand UO_2931 (O_2931,N_27222,N_25785);
and UO_2932 (O_2932,N_28639,N_29633);
or UO_2933 (O_2933,N_25928,N_27283);
nor UO_2934 (O_2934,N_29701,N_29741);
nor UO_2935 (O_2935,N_29543,N_26759);
xnor UO_2936 (O_2936,N_28920,N_28522);
or UO_2937 (O_2937,N_29967,N_25152);
nand UO_2938 (O_2938,N_28917,N_26782);
xnor UO_2939 (O_2939,N_25473,N_29990);
xor UO_2940 (O_2940,N_29960,N_25251);
and UO_2941 (O_2941,N_27519,N_29214);
or UO_2942 (O_2942,N_29274,N_25581);
xor UO_2943 (O_2943,N_29981,N_29487);
nand UO_2944 (O_2944,N_29735,N_28560);
nand UO_2945 (O_2945,N_25850,N_25716);
nand UO_2946 (O_2946,N_27010,N_26947);
nand UO_2947 (O_2947,N_29653,N_25503);
nand UO_2948 (O_2948,N_27315,N_28166);
and UO_2949 (O_2949,N_27124,N_27833);
or UO_2950 (O_2950,N_26670,N_29773);
and UO_2951 (O_2951,N_29422,N_29502);
or UO_2952 (O_2952,N_25135,N_26291);
or UO_2953 (O_2953,N_28392,N_29807);
xnor UO_2954 (O_2954,N_28895,N_29984);
or UO_2955 (O_2955,N_29211,N_25134);
nand UO_2956 (O_2956,N_29780,N_27517);
xnor UO_2957 (O_2957,N_25873,N_27195);
or UO_2958 (O_2958,N_28619,N_26902);
xor UO_2959 (O_2959,N_25440,N_27194);
and UO_2960 (O_2960,N_29189,N_29409);
and UO_2961 (O_2961,N_25635,N_27290);
xnor UO_2962 (O_2962,N_25899,N_25829);
and UO_2963 (O_2963,N_29531,N_28651);
nand UO_2964 (O_2964,N_26697,N_29321);
nand UO_2965 (O_2965,N_27587,N_28649);
xnor UO_2966 (O_2966,N_28905,N_25744);
nor UO_2967 (O_2967,N_26498,N_26605);
nand UO_2968 (O_2968,N_27889,N_27763);
and UO_2969 (O_2969,N_28711,N_27328);
nand UO_2970 (O_2970,N_28284,N_25878);
or UO_2971 (O_2971,N_25900,N_29584);
or UO_2972 (O_2972,N_25260,N_26281);
xnor UO_2973 (O_2973,N_27152,N_28557);
nand UO_2974 (O_2974,N_26820,N_26800);
and UO_2975 (O_2975,N_29134,N_28900);
nand UO_2976 (O_2976,N_27894,N_25877);
nand UO_2977 (O_2977,N_28355,N_26254);
nor UO_2978 (O_2978,N_25664,N_25451);
nor UO_2979 (O_2979,N_25420,N_29837);
and UO_2980 (O_2980,N_27148,N_29402);
nor UO_2981 (O_2981,N_27745,N_29941);
nand UO_2982 (O_2982,N_28936,N_28812);
or UO_2983 (O_2983,N_25366,N_26887);
nand UO_2984 (O_2984,N_28384,N_27529);
and UO_2985 (O_2985,N_28090,N_27987);
nand UO_2986 (O_2986,N_29174,N_25761);
and UO_2987 (O_2987,N_26603,N_26904);
nand UO_2988 (O_2988,N_28192,N_26370);
nand UO_2989 (O_2989,N_28222,N_25447);
nor UO_2990 (O_2990,N_27742,N_25603);
nand UO_2991 (O_2991,N_28773,N_27967);
and UO_2992 (O_2992,N_28332,N_28883);
or UO_2993 (O_2993,N_28184,N_29923);
or UO_2994 (O_2994,N_25787,N_29526);
nand UO_2995 (O_2995,N_26992,N_28607);
nand UO_2996 (O_2996,N_26773,N_25744);
and UO_2997 (O_2997,N_25228,N_25061);
nand UO_2998 (O_2998,N_26091,N_27300);
or UO_2999 (O_2999,N_27006,N_29002);
nor UO_3000 (O_3000,N_29089,N_26242);
xor UO_3001 (O_3001,N_28285,N_25967);
xor UO_3002 (O_3002,N_29802,N_28583);
and UO_3003 (O_3003,N_27658,N_26913);
nand UO_3004 (O_3004,N_28869,N_29913);
and UO_3005 (O_3005,N_25053,N_28888);
nor UO_3006 (O_3006,N_26491,N_27396);
nand UO_3007 (O_3007,N_29297,N_26568);
nand UO_3008 (O_3008,N_27710,N_28766);
nand UO_3009 (O_3009,N_25314,N_25403);
nor UO_3010 (O_3010,N_29773,N_26809);
xor UO_3011 (O_3011,N_29022,N_28325);
nor UO_3012 (O_3012,N_28119,N_27638);
nand UO_3013 (O_3013,N_25366,N_25467);
and UO_3014 (O_3014,N_25229,N_28031);
or UO_3015 (O_3015,N_29320,N_27851);
nand UO_3016 (O_3016,N_27453,N_25026);
nand UO_3017 (O_3017,N_29041,N_25787);
and UO_3018 (O_3018,N_25588,N_28393);
xnor UO_3019 (O_3019,N_29229,N_26611);
or UO_3020 (O_3020,N_29743,N_27497);
and UO_3021 (O_3021,N_28435,N_27747);
and UO_3022 (O_3022,N_25570,N_28110);
or UO_3023 (O_3023,N_26435,N_29805);
and UO_3024 (O_3024,N_26858,N_26910);
nor UO_3025 (O_3025,N_28094,N_28095);
nand UO_3026 (O_3026,N_25975,N_27363);
or UO_3027 (O_3027,N_25985,N_26003);
xor UO_3028 (O_3028,N_25336,N_27883);
nor UO_3029 (O_3029,N_28496,N_25978);
xnor UO_3030 (O_3030,N_29473,N_26267);
nand UO_3031 (O_3031,N_28095,N_25234);
and UO_3032 (O_3032,N_29969,N_29456);
nor UO_3033 (O_3033,N_26581,N_27051);
xnor UO_3034 (O_3034,N_29601,N_29992);
nand UO_3035 (O_3035,N_27825,N_29299);
or UO_3036 (O_3036,N_29655,N_27429);
nor UO_3037 (O_3037,N_28540,N_26658);
xor UO_3038 (O_3038,N_27372,N_28010);
or UO_3039 (O_3039,N_25792,N_29691);
xor UO_3040 (O_3040,N_27309,N_25334);
and UO_3041 (O_3041,N_29684,N_27017);
and UO_3042 (O_3042,N_25871,N_26534);
xor UO_3043 (O_3043,N_27258,N_29210);
nor UO_3044 (O_3044,N_29223,N_26565);
nor UO_3045 (O_3045,N_28774,N_25701);
nand UO_3046 (O_3046,N_29912,N_28784);
nand UO_3047 (O_3047,N_28377,N_26029);
nand UO_3048 (O_3048,N_28088,N_25365);
and UO_3049 (O_3049,N_26996,N_25718);
xnor UO_3050 (O_3050,N_27439,N_27152);
or UO_3051 (O_3051,N_29747,N_25189);
or UO_3052 (O_3052,N_25493,N_25255);
xnor UO_3053 (O_3053,N_28724,N_25780);
and UO_3054 (O_3054,N_28327,N_28041);
nor UO_3055 (O_3055,N_26075,N_29234);
nand UO_3056 (O_3056,N_29185,N_27649);
xor UO_3057 (O_3057,N_25785,N_27340);
xor UO_3058 (O_3058,N_25935,N_28489);
nor UO_3059 (O_3059,N_28593,N_25348);
nor UO_3060 (O_3060,N_29553,N_29801);
and UO_3061 (O_3061,N_25937,N_26311);
xor UO_3062 (O_3062,N_25483,N_28884);
nand UO_3063 (O_3063,N_29490,N_28007);
nand UO_3064 (O_3064,N_27531,N_27036);
or UO_3065 (O_3065,N_28612,N_28169);
or UO_3066 (O_3066,N_29457,N_26675);
or UO_3067 (O_3067,N_27703,N_27633);
nor UO_3068 (O_3068,N_26325,N_29925);
nand UO_3069 (O_3069,N_25788,N_25540);
and UO_3070 (O_3070,N_25412,N_27783);
nor UO_3071 (O_3071,N_28545,N_26587);
xnor UO_3072 (O_3072,N_26195,N_28913);
or UO_3073 (O_3073,N_26902,N_29785);
nand UO_3074 (O_3074,N_27843,N_27182);
and UO_3075 (O_3075,N_26480,N_28638);
nor UO_3076 (O_3076,N_27877,N_26996);
nor UO_3077 (O_3077,N_26142,N_26963);
nand UO_3078 (O_3078,N_29829,N_27655);
nor UO_3079 (O_3079,N_27723,N_29355);
nand UO_3080 (O_3080,N_28483,N_29986);
and UO_3081 (O_3081,N_27191,N_29227);
xor UO_3082 (O_3082,N_27556,N_27778);
nand UO_3083 (O_3083,N_25081,N_29939);
and UO_3084 (O_3084,N_28748,N_25686);
nand UO_3085 (O_3085,N_28172,N_25325);
xor UO_3086 (O_3086,N_28958,N_25280);
nand UO_3087 (O_3087,N_26474,N_29574);
nand UO_3088 (O_3088,N_28137,N_25638);
or UO_3089 (O_3089,N_29812,N_26334);
nor UO_3090 (O_3090,N_27406,N_29613);
or UO_3091 (O_3091,N_26686,N_28456);
nand UO_3092 (O_3092,N_25225,N_26534);
and UO_3093 (O_3093,N_26495,N_26530);
or UO_3094 (O_3094,N_26315,N_29789);
nand UO_3095 (O_3095,N_29617,N_25329);
nand UO_3096 (O_3096,N_29430,N_28297);
nand UO_3097 (O_3097,N_28219,N_29180);
nand UO_3098 (O_3098,N_28258,N_29571);
and UO_3099 (O_3099,N_28412,N_28552);
nor UO_3100 (O_3100,N_27218,N_29459);
and UO_3101 (O_3101,N_26958,N_29726);
and UO_3102 (O_3102,N_29791,N_25329);
xor UO_3103 (O_3103,N_27868,N_27919);
or UO_3104 (O_3104,N_27379,N_28643);
nand UO_3105 (O_3105,N_25256,N_26068);
nor UO_3106 (O_3106,N_28969,N_27193);
and UO_3107 (O_3107,N_27621,N_26105);
or UO_3108 (O_3108,N_25432,N_26881);
xor UO_3109 (O_3109,N_25407,N_28221);
nor UO_3110 (O_3110,N_29190,N_26480);
and UO_3111 (O_3111,N_26477,N_27595);
and UO_3112 (O_3112,N_28466,N_29335);
xnor UO_3113 (O_3113,N_28654,N_28239);
or UO_3114 (O_3114,N_28407,N_29744);
or UO_3115 (O_3115,N_29132,N_25163);
nor UO_3116 (O_3116,N_25856,N_26254);
nor UO_3117 (O_3117,N_26569,N_28630);
xnor UO_3118 (O_3118,N_28905,N_26446);
or UO_3119 (O_3119,N_26877,N_29884);
and UO_3120 (O_3120,N_28214,N_28910);
or UO_3121 (O_3121,N_29003,N_27711);
nor UO_3122 (O_3122,N_27698,N_26104);
xnor UO_3123 (O_3123,N_25661,N_29052);
nand UO_3124 (O_3124,N_26032,N_27860);
or UO_3125 (O_3125,N_29948,N_25215);
and UO_3126 (O_3126,N_25323,N_25007);
xnor UO_3127 (O_3127,N_25291,N_28510);
nand UO_3128 (O_3128,N_27515,N_29506);
and UO_3129 (O_3129,N_27295,N_26238);
nor UO_3130 (O_3130,N_27204,N_29092);
and UO_3131 (O_3131,N_25778,N_26422);
and UO_3132 (O_3132,N_28231,N_27404);
nand UO_3133 (O_3133,N_25772,N_28461);
or UO_3134 (O_3134,N_29767,N_28726);
and UO_3135 (O_3135,N_28549,N_28233);
or UO_3136 (O_3136,N_28019,N_27814);
nor UO_3137 (O_3137,N_27600,N_28121);
nor UO_3138 (O_3138,N_28586,N_29577);
and UO_3139 (O_3139,N_26016,N_26778);
nor UO_3140 (O_3140,N_26958,N_28947);
or UO_3141 (O_3141,N_27831,N_25679);
and UO_3142 (O_3142,N_29168,N_28866);
xor UO_3143 (O_3143,N_28186,N_26649);
and UO_3144 (O_3144,N_29308,N_27371);
or UO_3145 (O_3145,N_25194,N_25542);
or UO_3146 (O_3146,N_28194,N_25006);
or UO_3147 (O_3147,N_27901,N_26073);
and UO_3148 (O_3148,N_28201,N_27293);
xnor UO_3149 (O_3149,N_28410,N_29592);
nand UO_3150 (O_3150,N_29203,N_28918);
nand UO_3151 (O_3151,N_29403,N_25606);
nor UO_3152 (O_3152,N_27595,N_27856);
nand UO_3153 (O_3153,N_29858,N_28230);
and UO_3154 (O_3154,N_26508,N_29827);
and UO_3155 (O_3155,N_27899,N_26680);
or UO_3156 (O_3156,N_29095,N_26873);
xor UO_3157 (O_3157,N_25152,N_26194);
xnor UO_3158 (O_3158,N_28782,N_29263);
nor UO_3159 (O_3159,N_25730,N_29585);
and UO_3160 (O_3160,N_26411,N_26383);
or UO_3161 (O_3161,N_28881,N_27250);
and UO_3162 (O_3162,N_25065,N_25567);
nor UO_3163 (O_3163,N_27923,N_29892);
or UO_3164 (O_3164,N_26685,N_25915);
nand UO_3165 (O_3165,N_28377,N_27656);
or UO_3166 (O_3166,N_26456,N_25562);
or UO_3167 (O_3167,N_28383,N_27064);
nor UO_3168 (O_3168,N_25804,N_26625);
nand UO_3169 (O_3169,N_27488,N_29177);
or UO_3170 (O_3170,N_28654,N_28263);
nor UO_3171 (O_3171,N_28532,N_28367);
and UO_3172 (O_3172,N_25905,N_27939);
nand UO_3173 (O_3173,N_27873,N_29461);
or UO_3174 (O_3174,N_29705,N_29772);
nand UO_3175 (O_3175,N_25524,N_25970);
nor UO_3176 (O_3176,N_25058,N_25075);
or UO_3177 (O_3177,N_26840,N_26038);
nor UO_3178 (O_3178,N_27476,N_28801);
or UO_3179 (O_3179,N_26914,N_29057);
and UO_3180 (O_3180,N_28391,N_25557);
or UO_3181 (O_3181,N_28849,N_26729);
or UO_3182 (O_3182,N_27353,N_28628);
nand UO_3183 (O_3183,N_27360,N_27973);
and UO_3184 (O_3184,N_28590,N_26316);
or UO_3185 (O_3185,N_27216,N_27957);
or UO_3186 (O_3186,N_26205,N_28313);
or UO_3187 (O_3187,N_28217,N_29628);
or UO_3188 (O_3188,N_25503,N_29228);
nand UO_3189 (O_3189,N_29622,N_26771);
nor UO_3190 (O_3190,N_27658,N_25442);
or UO_3191 (O_3191,N_28639,N_27509);
nor UO_3192 (O_3192,N_26582,N_27905);
xnor UO_3193 (O_3193,N_27641,N_26677);
and UO_3194 (O_3194,N_27545,N_25106);
nor UO_3195 (O_3195,N_26339,N_27274);
or UO_3196 (O_3196,N_25928,N_27436);
or UO_3197 (O_3197,N_29392,N_28030);
or UO_3198 (O_3198,N_27464,N_27399);
nor UO_3199 (O_3199,N_26407,N_27702);
and UO_3200 (O_3200,N_28134,N_28210);
nand UO_3201 (O_3201,N_28862,N_28919);
xnor UO_3202 (O_3202,N_28692,N_26806);
nand UO_3203 (O_3203,N_25574,N_28718);
nor UO_3204 (O_3204,N_29612,N_25532);
or UO_3205 (O_3205,N_26410,N_28406);
nor UO_3206 (O_3206,N_25650,N_26714);
and UO_3207 (O_3207,N_29941,N_25379);
nand UO_3208 (O_3208,N_26863,N_27936);
and UO_3209 (O_3209,N_28735,N_27561);
nor UO_3210 (O_3210,N_28485,N_26463);
and UO_3211 (O_3211,N_27601,N_29991);
or UO_3212 (O_3212,N_27100,N_29258);
nand UO_3213 (O_3213,N_27622,N_25565);
nand UO_3214 (O_3214,N_25523,N_29869);
nor UO_3215 (O_3215,N_25444,N_29790);
nor UO_3216 (O_3216,N_25037,N_27556);
xnor UO_3217 (O_3217,N_29516,N_27956);
nor UO_3218 (O_3218,N_27098,N_27496);
nor UO_3219 (O_3219,N_25363,N_27110);
and UO_3220 (O_3220,N_27208,N_29230);
nor UO_3221 (O_3221,N_27024,N_27865);
and UO_3222 (O_3222,N_29499,N_25754);
nor UO_3223 (O_3223,N_28936,N_28823);
or UO_3224 (O_3224,N_25978,N_28814);
or UO_3225 (O_3225,N_28081,N_25268);
and UO_3226 (O_3226,N_27591,N_25583);
xor UO_3227 (O_3227,N_28496,N_26648);
or UO_3228 (O_3228,N_27993,N_26154);
or UO_3229 (O_3229,N_28799,N_27750);
or UO_3230 (O_3230,N_28080,N_27863);
or UO_3231 (O_3231,N_26898,N_29587);
xor UO_3232 (O_3232,N_25995,N_29978);
nand UO_3233 (O_3233,N_29540,N_28784);
or UO_3234 (O_3234,N_25023,N_29913);
and UO_3235 (O_3235,N_27476,N_26042);
or UO_3236 (O_3236,N_28446,N_25284);
or UO_3237 (O_3237,N_26579,N_27137);
xor UO_3238 (O_3238,N_26632,N_26178);
nor UO_3239 (O_3239,N_27871,N_28288);
nand UO_3240 (O_3240,N_25991,N_29124);
and UO_3241 (O_3241,N_26034,N_26514);
nor UO_3242 (O_3242,N_25239,N_28691);
nor UO_3243 (O_3243,N_26285,N_26449);
nor UO_3244 (O_3244,N_27965,N_25059);
or UO_3245 (O_3245,N_25957,N_29800);
nor UO_3246 (O_3246,N_26814,N_29494);
nand UO_3247 (O_3247,N_26235,N_26010);
nand UO_3248 (O_3248,N_26278,N_27441);
nor UO_3249 (O_3249,N_25873,N_29968);
and UO_3250 (O_3250,N_25882,N_29997);
or UO_3251 (O_3251,N_27747,N_28357);
or UO_3252 (O_3252,N_26645,N_25042);
nor UO_3253 (O_3253,N_29010,N_28440);
xor UO_3254 (O_3254,N_28126,N_28474);
nor UO_3255 (O_3255,N_27417,N_29603);
nand UO_3256 (O_3256,N_27812,N_27108);
nand UO_3257 (O_3257,N_28367,N_27373);
nor UO_3258 (O_3258,N_25969,N_27637);
nand UO_3259 (O_3259,N_26882,N_25234);
nor UO_3260 (O_3260,N_27224,N_27118);
nor UO_3261 (O_3261,N_25956,N_27019);
nand UO_3262 (O_3262,N_26642,N_27456);
nand UO_3263 (O_3263,N_28035,N_28379);
or UO_3264 (O_3264,N_27951,N_28274);
or UO_3265 (O_3265,N_26302,N_26351);
nor UO_3266 (O_3266,N_25148,N_28932);
nor UO_3267 (O_3267,N_27881,N_28039);
nor UO_3268 (O_3268,N_27079,N_28225);
or UO_3269 (O_3269,N_28583,N_28407);
and UO_3270 (O_3270,N_27604,N_28380);
and UO_3271 (O_3271,N_28877,N_28127);
and UO_3272 (O_3272,N_26948,N_26405);
and UO_3273 (O_3273,N_29134,N_27415);
and UO_3274 (O_3274,N_29512,N_27181);
xor UO_3275 (O_3275,N_25304,N_29615);
and UO_3276 (O_3276,N_25155,N_27212);
nand UO_3277 (O_3277,N_25250,N_29320);
nor UO_3278 (O_3278,N_26642,N_29707);
and UO_3279 (O_3279,N_29615,N_29301);
nand UO_3280 (O_3280,N_29384,N_28543);
nand UO_3281 (O_3281,N_29216,N_27360);
nand UO_3282 (O_3282,N_29470,N_26129);
nand UO_3283 (O_3283,N_27690,N_28195);
nand UO_3284 (O_3284,N_28876,N_25285);
or UO_3285 (O_3285,N_27219,N_29325);
and UO_3286 (O_3286,N_26933,N_28695);
or UO_3287 (O_3287,N_26242,N_29455);
nand UO_3288 (O_3288,N_26442,N_26180);
xnor UO_3289 (O_3289,N_28650,N_25602);
nand UO_3290 (O_3290,N_26563,N_25612);
and UO_3291 (O_3291,N_29035,N_26092);
nand UO_3292 (O_3292,N_27553,N_29570);
or UO_3293 (O_3293,N_27991,N_25155);
and UO_3294 (O_3294,N_28613,N_29819);
nor UO_3295 (O_3295,N_27519,N_25670);
xor UO_3296 (O_3296,N_25056,N_26192);
and UO_3297 (O_3297,N_25518,N_25522);
xnor UO_3298 (O_3298,N_25480,N_29127);
or UO_3299 (O_3299,N_26274,N_29889);
nand UO_3300 (O_3300,N_25128,N_29675);
or UO_3301 (O_3301,N_26112,N_25053);
nor UO_3302 (O_3302,N_29775,N_29708);
or UO_3303 (O_3303,N_28014,N_25468);
xnor UO_3304 (O_3304,N_25094,N_26487);
nand UO_3305 (O_3305,N_28145,N_29802);
or UO_3306 (O_3306,N_29233,N_26581);
xnor UO_3307 (O_3307,N_28750,N_28655);
nor UO_3308 (O_3308,N_26544,N_29279);
and UO_3309 (O_3309,N_26895,N_25644);
or UO_3310 (O_3310,N_25423,N_27264);
nor UO_3311 (O_3311,N_29573,N_29800);
nand UO_3312 (O_3312,N_26528,N_29892);
nor UO_3313 (O_3313,N_28749,N_28484);
and UO_3314 (O_3314,N_27341,N_27529);
nand UO_3315 (O_3315,N_27033,N_27373);
and UO_3316 (O_3316,N_25576,N_29007);
nand UO_3317 (O_3317,N_28073,N_28877);
or UO_3318 (O_3318,N_28685,N_25676);
nor UO_3319 (O_3319,N_29667,N_27085);
or UO_3320 (O_3320,N_27464,N_28513);
nor UO_3321 (O_3321,N_28301,N_28755);
or UO_3322 (O_3322,N_25985,N_26239);
nor UO_3323 (O_3323,N_26554,N_26523);
or UO_3324 (O_3324,N_27189,N_27105);
or UO_3325 (O_3325,N_28539,N_29589);
and UO_3326 (O_3326,N_26985,N_27803);
nor UO_3327 (O_3327,N_28400,N_25213);
nand UO_3328 (O_3328,N_26494,N_29957);
or UO_3329 (O_3329,N_29233,N_29196);
and UO_3330 (O_3330,N_28516,N_25144);
nor UO_3331 (O_3331,N_28847,N_29096);
or UO_3332 (O_3332,N_27321,N_25690);
nand UO_3333 (O_3333,N_26361,N_27962);
xor UO_3334 (O_3334,N_28784,N_25040);
and UO_3335 (O_3335,N_27759,N_25830);
nand UO_3336 (O_3336,N_25769,N_26370);
nand UO_3337 (O_3337,N_26048,N_29800);
or UO_3338 (O_3338,N_25095,N_29003);
nand UO_3339 (O_3339,N_25829,N_25696);
and UO_3340 (O_3340,N_27263,N_28899);
and UO_3341 (O_3341,N_28916,N_28626);
and UO_3342 (O_3342,N_27869,N_26002);
nor UO_3343 (O_3343,N_29426,N_28042);
nor UO_3344 (O_3344,N_26804,N_26990);
nand UO_3345 (O_3345,N_27219,N_26860);
or UO_3346 (O_3346,N_29436,N_26557);
nand UO_3347 (O_3347,N_28669,N_29273);
xnor UO_3348 (O_3348,N_28356,N_25342);
and UO_3349 (O_3349,N_25383,N_29625);
xnor UO_3350 (O_3350,N_28448,N_26412);
nor UO_3351 (O_3351,N_27837,N_29396);
and UO_3352 (O_3352,N_25163,N_26578);
nand UO_3353 (O_3353,N_27054,N_25662);
or UO_3354 (O_3354,N_28200,N_28275);
nor UO_3355 (O_3355,N_28556,N_29649);
or UO_3356 (O_3356,N_26107,N_28935);
nand UO_3357 (O_3357,N_26871,N_25945);
and UO_3358 (O_3358,N_29287,N_25310);
or UO_3359 (O_3359,N_27950,N_26427);
xnor UO_3360 (O_3360,N_28317,N_25394);
or UO_3361 (O_3361,N_28144,N_25935);
or UO_3362 (O_3362,N_29042,N_29179);
nand UO_3363 (O_3363,N_25529,N_27708);
nand UO_3364 (O_3364,N_25505,N_26767);
nor UO_3365 (O_3365,N_25141,N_25830);
and UO_3366 (O_3366,N_28285,N_27712);
xor UO_3367 (O_3367,N_26345,N_26397);
and UO_3368 (O_3368,N_25859,N_28780);
or UO_3369 (O_3369,N_26523,N_29402);
and UO_3370 (O_3370,N_25611,N_27560);
nand UO_3371 (O_3371,N_25466,N_25027);
xor UO_3372 (O_3372,N_25794,N_28198);
nand UO_3373 (O_3373,N_25533,N_29327);
nor UO_3374 (O_3374,N_26014,N_28623);
nand UO_3375 (O_3375,N_28565,N_29661);
xor UO_3376 (O_3376,N_27371,N_28540);
and UO_3377 (O_3377,N_26197,N_28184);
nor UO_3378 (O_3378,N_27534,N_28289);
nand UO_3379 (O_3379,N_29932,N_26716);
nand UO_3380 (O_3380,N_27780,N_28043);
xor UO_3381 (O_3381,N_26210,N_27288);
or UO_3382 (O_3382,N_29891,N_29717);
and UO_3383 (O_3383,N_27827,N_25571);
nand UO_3384 (O_3384,N_25485,N_25615);
and UO_3385 (O_3385,N_25682,N_25902);
nand UO_3386 (O_3386,N_27046,N_26232);
and UO_3387 (O_3387,N_29155,N_29058);
or UO_3388 (O_3388,N_25648,N_27899);
nand UO_3389 (O_3389,N_27743,N_29746);
and UO_3390 (O_3390,N_26511,N_28407);
or UO_3391 (O_3391,N_27304,N_28179);
or UO_3392 (O_3392,N_27827,N_27599);
or UO_3393 (O_3393,N_29025,N_29086);
nor UO_3394 (O_3394,N_25845,N_28558);
and UO_3395 (O_3395,N_29786,N_29242);
nor UO_3396 (O_3396,N_27188,N_29508);
xnor UO_3397 (O_3397,N_25061,N_28727);
or UO_3398 (O_3398,N_25591,N_28598);
or UO_3399 (O_3399,N_27913,N_25106);
nand UO_3400 (O_3400,N_27775,N_28062);
nand UO_3401 (O_3401,N_27046,N_25747);
nor UO_3402 (O_3402,N_28938,N_28495);
and UO_3403 (O_3403,N_27779,N_26233);
and UO_3404 (O_3404,N_25834,N_27724);
nand UO_3405 (O_3405,N_25210,N_25604);
nor UO_3406 (O_3406,N_29322,N_25251);
nor UO_3407 (O_3407,N_29037,N_28041);
nand UO_3408 (O_3408,N_26898,N_28072);
nand UO_3409 (O_3409,N_29107,N_25571);
nand UO_3410 (O_3410,N_27060,N_27753);
nor UO_3411 (O_3411,N_29312,N_29189);
nor UO_3412 (O_3412,N_28299,N_26880);
nor UO_3413 (O_3413,N_26043,N_29377);
or UO_3414 (O_3414,N_28583,N_25634);
nand UO_3415 (O_3415,N_27566,N_27487);
nand UO_3416 (O_3416,N_25502,N_26515);
nor UO_3417 (O_3417,N_25749,N_27082);
nand UO_3418 (O_3418,N_25855,N_29471);
or UO_3419 (O_3419,N_27007,N_26688);
or UO_3420 (O_3420,N_26014,N_26537);
and UO_3421 (O_3421,N_28229,N_26120);
and UO_3422 (O_3422,N_29608,N_27621);
nand UO_3423 (O_3423,N_25274,N_26653);
nand UO_3424 (O_3424,N_28796,N_25029);
or UO_3425 (O_3425,N_26531,N_28297);
and UO_3426 (O_3426,N_27014,N_29477);
and UO_3427 (O_3427,N_26057,N_27699);
xor UO_3428 (O_3428,N_25155,N_27759);
nand UO_3429 (O_3429,N_29634,N_27718);
or UO_3430 (O_3430,N_25054,N_25593);
and UO_3431 (O_3431,N_25776,N_29041);
or UO_3432 (O_3432,N_29323,N_26390);
nor UO_3433 (O_3433,N_26215,N_26224);
nand UO_3434 (O_3434,N_29507,N_29680);
nor UO_3435 (O_3435,N_26321,N_26176);
and UO_3436 (O_3436,N_28680,N_27458);
and UO_3437 (O_3437,N_27843,N_29451);
nand UO_3438 (O_3438,N_29064,N_27797);
nor UO_3439 (O_3439,N_27159,N_26231);
and UO_3440 (O_3440,N_26567,N_29231);
and UO_3441 (O_3441,N_29245,N_29175);
xor UO_3442 (O_3442,N_29836,N_29524);
or UO_3443 (O_3443,N_25209,N_29685);
nand UO_3444 (O_3444,N_27044,N_25030);
and UO_3445 (O_3445,N_25947,N_28245);
or UO_3446 (O_3446,N_27336,N_26744);
nand UO_3447 (O_3447,N_27517,N_28125);
xor UO_3448 (O_3448,N_29509,N_27856);
and UO_3449 (O_3449,N_26661,N_26356);
nand UO_3450 (O_3450,N_25262,N_28629);
and UO_3451 (O_3451,N_26921,N_28361);
or UO_3452 (O_3452,N_25985,N_26668);
or UO_3453 (O_3453,N_28890,N_27065);
nand UO_3454 (O_3454,N_28625,N_28992);
nor UO_3455 (O_3455,N_27828,N_27212);
and UO_3456 (O_3456,N_29802,N_28556);
nor UO_3457 (O_3457,N_25892,N_27220);
nand UO_3458 (O_3458,N_28001,N_29011);
nor UO_3459 (O_3459,N_27020,N_27715);
and UO_3460 (O_3460,N_28752,N_27229);
nor UO_3461 (O_3461,N_27138,N_25348);
xnor UO_3462 (O_3462,N_28586,N_29930);
xnor UO_3463 (O_3463,N_26253,N_29528);
or UO_3464 (O_3464,N_25729,N_28545);
or UO_3465 (O_3465,N_27864,N_28739);
nand UO_3466 (O_3466,N_25948,N_29839);
or UO_3467 (O_3467,N_28036,N_25722);
xnor UO_3468 (O_3468,N_29872,N_25476);
and UO_3469 (O_3469,N_27893,N_26662);
xor UO_3470 (O_3470,N_25734,N_29924);
and UO_3471 (O_3471,N_25713,N_27756);
or UO_3472 (O_3472,N_28489,N_28052);
or UO_3473 (O_3473,N_27093,N_29834);
or UO_3474 (O_3474,N_26332,N_29737);
or UO_3475 (O_3475,N_29109,N_27791);
nand UO_3476 (O_3476,N_27265,N_25738);
xnor UO_3477 (O_3477,N_26992,N_25783);
or UO_3478 (O_3478,N_26983,N_26566);
nand UO_3479 (O_3479,N_29651,N_27347);
or UO_3480 (O_3480,N_29263,N_29102);
and UO_3481 (O_3481,N_26684,N_27408);
xnor UO_3482 (O_3482,N_27287,N_29694);
nor UO_3483 (O_3483,N_29461,N_25396);
nand UO_3484 (O_3484,N_28732,N_29322);
xor UO_3485 (O_3485,N_25758,N_26706);
and UO_3486 (O_3486,N_27183,N_25350);
nor UO_3487 (O_3487,N_26347,N_25934);
xnor UO_3488 (O_3488,N_27329,N_28330);
nand UO_3489 (O_3489,N_27635,N_27410);
nand UO_3490 (O_3490,N_29490,N_27710);
or UO_3491 (O_3491,N_26440,N_26710);
and UO_3492 (O_3492,N_29265,N_27138);
nand UO_3493 (O_3493,N_28521,N_28281);
or UO_3494 (O_3494,N_25885,N_27316);
and UO_3495 (O_3495,N_26601,N_25854);
nor UO_3496 (O_3496,N_25083,N_26564);
and UO_3497 (O_3497,N_29260,N_28595);
nand UO_3498 (O_3498,N_28306,N_27970);
and UO_3499 (O_3499,N_26110,N_25865);
endmodule