module basic_5000_50000_5000_50_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xor U0 (N_0,In_3761,In_4575);
and U1 (N_1,In_4454,In_3271);
nor U2 (N_2,In_2897,In_282);
or U3 (N_3,In_4466,In_627);
and U4 (N_4,In_345,In_4422);
and U5 (N_5,In_301,In_2507);
or U6 (N_6,In_3145,In_4498);
xnor U7 (N_7,In_3028,In_1767);
xor U8 (N_8,In_2950,In_239);
or U9 (N_9,In_2488,In_4407);
xnor U10 (N_10,In_1691,In_506);
nor U11 (N_11,In_3735,In_143);
or U12 (N_12,In_288,In_626);
nand U13 (N_13,In_3019,In_2016);
and U14 (N_14,In_2241,In_2988);
or U15 (N_15,In_2165,In_4260);
xnor U16 (N_16,In_3723,In_218);
xnor U17 (N_17,In_231,In_4935);
nand U18 (N_18,In_3798,In_1915);
nor U19 (N_19,In_3232,In_4238);
or U20 (N_20,In_144,In_2482);
and U21 (N_21,In_50,In_4144);
and U22 (N_22,In_4763,In_1633);
nor U23 (N_23,In_4428,In_1173);
nand U24 (N_24,In_4630,In_1384);
nor U25 (N_25,In_4767,In_2112);
and U26 (N_26,In_1496,In_1155);
nor U27 (N_27,In_2145,In_949);
and U28 (N_28,In_286,In_3379);
xor U29 (N_29,In_1279,In_3186);
xnor U30 (N_30,In_584,In_362);
and U31 (N_31,In_4294,In_2375);
and U32 (N_32,In_4887,In_1082);
xor U33 (N_33,In_188,In_68);
or U34 (N_34,In_78,In_3704);
nor U35 (N_35,In_443,In_3925);
or U36 (N_36,In_4692,In_2152);
or U37 (N_37,In_1324,In_258);
or U38 (N_38,In_3225,In_1490);
xnor U39 (N_39,In_4863,In_2104);
nand U40 (N_40,In_3133,In_354);
nor U41 (N_41,In_3577,In_94);
or U42 (N_42,In_3080,In_4636);
nand U43 (N_43,In_4751,In_547);
or U44 (N_44,In_2775,In_1945);
xor U45 (N_45,In_3468,In_2329);
nand U46 (N_46,In_2652,In_2749);
xnor U47 (N_47,In_369,In_487);
nor U48 (N_48,In_3156,In_930);
xor U49 (N_49,In_1164,In_3500);
or U50 (N_50,In_3491,In_564);
nand U51 (N_51,In_2952,In_1076);
and U52 (N_52,In_2810,In_3516);
and U53 (N_53,In_4180,In_2416);
xor U54 (N_54,In_1649,In_2940);
or U55 (N_55,In_174,In_1162);
nor U56 (N_56,In_3119,In_3948);
xnor U57 (N_57,In_338,In_330);
nor U58 (N_58,In_464,In_3520);
nor U59 (N_59,In_2039,In_2703);
nor U60 (N_60,In_482,In_1905);
nand U61 (N_61,In_79,In_2843);
xor U62 (N_62,In_944,In_2074);
and U63 (N_63,In_2984,In_2334);
or U64 (N_64,In_2317,In_2849);
nor U65 (N_65,In_3327,In_1329);
xnor U66 (N_66,In_2006,In_510);
xor U67 (N_67,In_1723,In_1015);
and U68 (N_68,In_2777,In_1798);
nor U69 (N_69,In_3878,In_4765);
or U70 (N_70,In_2421,In_1434);
nor U71 (N_71,In_348,In_3780);
nor U72 (N_72,In_3239,In_1535);
nand U73 (N_73,In_3994,In_4477);
and U74 (N_74,In_3876,In_334);
nand U75 (N_75,In_2427,In_3698);
nor U76 (N_76,In_4043,In_4006);
xnor U77 (N_77,In_844,In_204);
nor U78 (N_78,In_1614,In_3078);
nand U79 (N_79,In_1152,In_4328);
and U80 (N_80,In_977,In_2218);
and U81 (N_81,In_1834,In_3634);
and U82 (N_82,In_3788,In_2604);
xor U83 (N_83,In_3482,In_817);
and U84 (N_84,In_420,In_419);
or U85 (N_85,In_4307,In_1621);
nor U86 (N_86,In_4452,In_4184);
nand U87 (N_87,In_3715,In_3640);
nand U88 (N_88,In_4233,In_724);
nand U89 (N_89,In_417,In_3218);
nor U90 (N_90,In_2522,In_1780);
nand U91 (N_91,In_4173,In_4136);
nand U92 (N_92,In_4662,In_404);
xnor U93 (N_93,In_2598,In_2282);
and U94 (N_94,In_167,In_1119);
and U95 (N_95,In_579,In_4270);
and U96 (N_96,In_3966,In_2455);
nand U97 (N_97,In_1656,In_3845);
xnor U98 (N_98,In_447,In_4571);
nor U99 (N_99,In_4993,In_3662);
and U100 (N_100,In_901,In_4083);
xor U101 (N_101,In_1703,In_851);
nand U102 (N_102,In_4595,In_3782);
or U103 (N_103,In_4803,In_3466);
nand U104 (N_104,In_1244,In_1438);
nor U105 (N_105,In_349,In_3487);
or U106 (N_106,In_3739,In_480);
and U107 (N_107,In_2127,In_3787);
xor U108 (N_108,In_1852,In_2811);
nand U109 (N_109,In_2666,In_2237);
xor U110 (N_110,In_1335,In_1377);
nor U111 (N_111,In_4387,In_4500);
and U112 (N_112,In_4483,In_612);
xor U113 (N_113,In_2322,In_767);
and U114 (N_114,In_4783,In_545);
and U115 (N_115,In_2069,In_1681);
xnor U116 (N_116,In_849,In_2757);
nor U117 (N_117,In_1031,In_4673);
and U118 (N_118,In_792,In_1089);
and U119 (N_119,In_1085,In_2226);
nor U120 (N_120,In_1894,In_4316);
nand U121 (N_121,In_4378,In_1188);
nor U122 (N_122,In_3840,In_3934);
nor U123 (N_123,In_2702,In_858);
nor U124 (N_124,In_1243,In_717);
and U125 (N_125,In_4102,In_3674);
xnor U126 (N_126,In_4178,In_505);
or U127 (N_127,In_4790,In_3969);
or U128 (N_128,In_3774,In_4310);
nand U129 (N_129,In_3033,In_4964);
and U130 (N_130,In_1371,In_1499);
xnor U131 (N_131,In_1247,In_964);
xnor U132 (N_132,In_4738,In_2187);
nand U133 (N_133,In_4653,In_2568);
nor U134 (N_134,In_1799,In_3884);
and U135 (N_135,In_4998,In_2013);
and U136 (N_136,In_4977,In_3248);
nor U137 (N_137,In_1385,In_769);
nand U138 (N_138,In_3441,In_1998);
and U139 (N_139,In_3766,In_2788);
nor U140 (N_140,In_3978,In_2414);
and U141 (N_141,In_3067,In_2677);
xor U142 (N_142,In_2361,In_2883);
and U143 (N_143,In_1380,In_500);
and U144 (N_144,In_3973,In_4137);
and U145 (N_145,In_1558,In_1120);
xor U146 (N_146,In_164,In_4440);
or U147 (N_147,In_2668,In_1070);
or U148 (N_148,In_4099,In_192);
or U149 (N_149,In_2139,In_3373);
nor U150 (N_150,In_789,In_1319);
nand U151 (N_151,In_2186,In_4481);
and U152 (N_152,In_316,In_3307);
and U153 (N_153,In_4832,In_3877);
nand U154 (N_154,In_179,In_1849);
nand U155 (N_155,In_4755,In_3712);
xor U156 (N_156,In_1716,In_3034);
nand U157 (N_157,In_3895,In_557);
nor U158 (N_158,In_4325,In_1645);
xor U159 (N_159,In_3786,In_2303);
xor U160 (N_160,In_4097,In_4888);
nand U161 (N_161,In_115,In_3283);
xnor U162 (N_162,In_958,In_2767);
and U163 (N_163,In_1174,In_3660);
or U164 (N_164,In_721,In_4731);
nand U165 (N_165,In_581,In_2559);
nor U166 (N_166,In_2182,In_3542);
xnor U167 (N_167,In_1124,In_642);
xor U168 (N_168,In_693,In_2873);
nor U169 (N_169,In_1638,In_153);
nor U170 (N_170,In_2937,In_4112);
nor U171 (N_171,In_712,In_4346);
or U172 (N_172,In_60,In_3191);
nor U173 (N_173,In_1725,In_2624);
xnor U174 (N_174,In_3536,In_1757);
nand U175 (N_175,In_4701,In_1447);
nor U176 (N_176,In_4411,In_2132);
xnor U177 (N_177,In_2599,In_2618);
nor U178 (N_178,In_4643,In_4134);
or U179 (N_179,In_2826,In_967);
nor U180 (N_180,In_4757,In_791);
nor U181 (N_181,In_2501,In_868);
nor U182 (N_182,In_3850,In_3518);
and U183 (N_183,In_1215,In_559);
xor U184 (N_184,In_1333,In_714);
nor U185 (N_185,In_732,In_2257);
and U186 (N_186,In_1880,In_507);
nor U187 (N_187,In_3820,In_4080);
and U188 (N_188,In_3639,In_1121);
or U189 (N_189,In_4107,In_1273);
nand U190 (N_190,In_3515,In_1451);
and U191 (N_191,In_3110,In_4929);
or U192 (N_192,In_1442,In_2617);
nor U193 (N_193,In_1940,In_27);
xor U194 (N_194,In_3250,In_2866);
and U195 (N_195,In_4904,In_3154);
or U196 (N_196,In_3641,In_2217);
xnor U197 (N_197,In_3773,In_3809);
or U198 (N_198,In_1557,In_2480);
or U199 (N_199,In_854,In_1906);
and U200 (N_200,In_1183,In_249);
or U201 (N_201,In_574,In_2856);
and U202 (N_202,In_3830,In_3419);
nor U203 (N_203,In_555,In_2449);
nand U204 (N_204,In_1724,In_4305);
or U205 (N_205,In_1840,In_3407);
nand U206 (N_206,In_2960,In_4192);
nand U207 (N_207,In_253,In_2298);
nor U208 (N_208,In_2300,In_3429);
nor U209 (N_209,In_4526,In_4988);
or U210 (N_210,In_1635,In_2909);
and U211 (N_211,In_1470,In_965);
or U212 (N_212,In_2281,In_1437);
and U213 (N_213,In_536,In_3962);
nand U214 (N_214,In_313,In_202);
or U215 (N_215,In_4577,In_790);
xnor U216 (N_216,In_698,In_892);
nor U217 (N_217,In_1398,In_4649);
or U218 (N_218,In_535,In_3880);
nor U219 (N_219,In_670,In_3294);
and U220 (N_220,In_2641,In_3);
xor U221 (N_221,In_1025,In_2922);
or U222 (N_222,In_77,In_490);
or U223 (N_223,In_808,In_4179);
and U224 (N_224,In_908,In_4009);
and U225 (N_225,In_3908,In_3696);
and U226 (N_226,In_4811,In_2662);
and U227 (N_227,In_414,In_839);
nand U228 (N_228,In_1202,In_758);
nand U229 (N_229,In_2235,In_1521);
and U230 (N_230,In_1257,In_2957);
xnor U231 (N_231,In_4172,In_2294);
xor U232 (N_232,In_128,In_2423);
nor U233 (N_233,In_307,In_2064);
or U234 (N_234,In_4810,In_1396);
nor U235 (N_235,In_4063,In_669);
xor U236 (N_236,In_678,In_4947);
or U237 (N_237,In_934,In_2289);
nand U238 (N_238,In_2879,In_3164);
nor U239 (N_239,In_4700,In_227);
or U240 (N_240,In_3134,In_2080);
xnor U241 (N_241,In_3977,In_895);
nor U242 (N_242,In_4956,In_1465);
and U243 (N_243,In_277,In_652);
nand U244 (N_244,In_3550,In_2975);
or U245 (N_245,In_3082,In_914);
nor U246 (N_246,In_3216,In_69);
or U247 (N_247,In_1797,In_4282);
nor U248 (N_248,In_435,In_2025);
nand U249 (N_249,In_2902,In_2590);
and U250 (N_250,In_3902,In_707);
xor U251 (N_251,In_3143,In_1440);
nand U252 (N_252,In_1886,In_3358);
nor U253 (N_253,In_2209,In_2660);
or U254 (N_254,In_3335,In_1560);
xnor U255 (N_255,In_3437,In_4594);
nor U256 (N_256,In_951,In_4259);
and U257 (N_257,In_2711,In_3063);
and U258 (N_258,In_2242,In_328);
xnor U259 (N_259,In_828,In_666);
and U260 (N_260,In_1844,In_4502);
xor U261 (N_261,In_2718,In_4196);
nand U262 (N_262,In_1843,In_755);
xnor U263 (N_263,In_4779,In_2676);
or U264 (N_264,In_1373,In_3293);
nor U265 (N_265,In_1190,In_3776);
or U266 (N_266,In_2981,In_1900);
or U267 (N_267,In_690,In_2266);
and U268 (N_268,In_1974,In_2318);
nand U269 (N_269,In_677,In_3184);
and U270 (N_270,In_2272,In_4072);
nand U271 (N_271,In_592,In_120);
and U272 (N_272,In_2963,In_2787);
nor U273 (N_273,In_3302,In_2830);
or U274 (N_274,In_2397,In_1837);
xnor U275 (N_275,In_1893,In_830);
xnor U276 (N_276,In_3514,In_3657);
or U277 (N_277,In_1730,In_3747);
nor U278 (N_278,In_2188,In_4671);
xor U279 (N_279,In_1430,In_2792);
or U280 (N_280,In_3593,In_961);
and U281 (N_281,In_2386,In_1310);
and U282 (N_282,In_4531,In_1232);
nand U283 (N_283,In_4312,In_4185);
or U284 (N_284,In_2932,In_4802);
or U285 (N_285,In_3201,In_2908);
or U286 (N_286,In_3177,In_2531);
xnor U287 (N_287,In_1779,In_3541);
and U288 (N_288,In_1203,In_2847);
or U289 (N_289,In_803,In_1925);
and U290 (N_290,In_2486,In_4710);
or U291 (N_291,In_2601,In_2752);
and U292 (N_292,In_516,In_4908);
and U293 (N_293,In_3044,In_2889);
xor U294 (N_294,In_3277,In_2556);
xor U295 (N_295,In_124,In_4482);
nand U296 (N_296,In_1048,In_1166);
xnor U297 (N_297,In_4835,In_1315);
and U298 (N_298,In_2672,In_1588);
and U299 (N_299,In_3924,In_4774);
nor U300 (N_300,In_1427,In_3269);
and U301 (N_301,In_2831,In_1805);
and U302 (N_302,In_4031,In_3226);
nor U303 (N_303,In_1801,In_4916);
xnor U304 (N_304,In_1765,In_1472);
xnor U305 (N_305,In_2939,In_1127);
nor U306 (N_306,In_236,In_3176);
or U307 (N_307,In_4961,In_2644);
or U308 (N_308,In_2762,In_4223);
or U309 (N_309,In_3118,In_2686);
xnor U310 (N_310,In_180,In_1771);
nor U311 (N_311,In_3822,In_1734);
xor U312 (N_312,In_4773,In_2555);
xnor U313 (N_313,In_3719,In_826);
or U314 (N_314,In_2532,In_1710);
and U315 (N_315,In_996,In_1585);
and U316 (N_316,In_880,In_4759);
and U317 (N_317,In_216,In_1059);
nor U318 (N_318,In_2934,In_4979);
or U319 (N_319,In_1911,In_4749);
or U320 (N_320,In_2948,In_387);
xnor U321 (N_321,In_2185,In_3434);
xor U322 (N_322,In_1566,In_210);
nand U323 (N_323,In_3794,In_322);
nand U324 (N_324,In_3728,In_4403);
nand U325 (N_325,In_881,In_566);
or U326 (N_326,In_2207,In_3693);
or U327 (N_327,In_4532,In_1822);
and U328 (N_328,In_2580,In_1807);
nand U329 (N_329,In_1748,In_4045);
or U330 (N_330,In_2170,In_4462);
nor U331 (N_331,In_2707,In_3815);
or U332 (N_332,In_3411,In_1464);
xnor U333 (N_333,In_1592,In_3957);
nor U334 (N_334,In_2142,In_1841);
nor U335 (N_335,In_4593,In_1135);
and U336 (N_336,In_275,In_3275);
or U337 (N_337,In_952,In_4739);
or U338 (N_338,In_2193,In_3169);
nor U339 (N_339,In_4920,In_2570);
xor U340 (N_340,In_1570,In_327);
nand U341 (N_341,In_3686,In_1794);
nor U342 (N_342,In_52,In_3018);
nand U343 (N_343,In_2894,In_2005);
nand U344 (N_344,In_1160,In_2268);
or U345 (N_345,In_4135,In_4478);
and U346 (N_346,In_3126,In_172);
xnor U347 (N_347,In_2890,In_389);
nand U348 (N_348,In_981,In_242);
and U349 (N_349,In_2254,In_3594);
and U350 (N_350,In_1789,In_945);
nand U351 (N_351,In_3324,In_861);
nand U352 (N_352,In_4337,In_3939);
nor U353 (N_353,In_2491,In_1131);
nor U354 (N_354,In_3007,In_631);
or U355 (N_355,In_2320,In_1641);
xnor U356 (N_356,In_1052,In_3651);
nand U357 (N_357,In_472,In_1534);
or U358 (N_358,In_2054,In_3952);
nand U359 (N_359,In_4417,In_2279);
nand U360 (N_360,In_56,In_2987);
and U361 (N_361,In_4666,In_1522);
or U362 (N_362,In_3814,In_4938);
or U363 (N_363,In_2450,In_2105);
xnor U364 (N_364,In_1432,In_3792);
xnor U365 (N_365,In_1989,In_1653);
or U366 (N_366,In_3649,In_425);
nor U367 (N_367,In_3626,In_1016);
or U368 (N_368,In_114,In_749);
nand U369 (N_369,In_3643,In_4878);
and U370 (N_370,In_4555,In_293);
nor U371 (N_371,In_2228,In_2898);
or U372 (N_372,In_1308,In_2133);
nor U373 (N_373,In_766,In_4873);
xnor U374 (N_374,In_3075,In_1486);
nor U375 (N_375,In_3399,In_3000);
or U376 (N_376,In_2154,In_2378);
and U377 (N_377,In_3519,In_3313);
and U378 (N_378,In_3392,In_2776);
nor U379 (N_379,In_3291,In_3714);
and U380 (N_380,In_4042,In_4379);
and U381 (N_381,In_412,In_1374);
and U382 (N_382,In_4414,In_1759);
xnor U383 (N_383,In_4750,In_1509);
and U384 (N_384,In_748,In_3091);
and U385 (N_385,In_1117,In_4272);
nand U386 (N_386,In_465,In_4869);
nor U387 (N_387,In_333,In_2653);
nand U388 (N_388,In_1443,In_4047);
nand U389 (N_389,In_4071,In_1958);
xor U390 (N_390,In_4551,In_1092);
nand U391 (N_391,In_3326,In_1487);
nor U392 (N_392,In_297,In_3802);
nor U393 (N_393,In_1892,In_632);
xor U394 (N_394,In_1013,In_1804);
or U395 (N_395,In_4989,In_1782);
xnor U396 (N_396,In_3115,In_2118);
nand U397 (N_397,In_4719,In_3797);
xnor U398 (N_398,In_3305,In_1253);
xnor U399 (N_399,In_1210,In_3863);
or U400 (N_400,In_1590,In_3224);
and U401 (N_401,In_4709,In_4019);
or U402 (N_402,In_2758,In_3580);
or U403 (N_403,In_3194,In_4228);
or U404 (N_404,In_1489,In_1325);
or U405 (N_405,In_3008,In_2832);
xnor U406 (N_406,In_423,In_4295);
xnor U407 (N_407,In_3637,In_825);
and U408 (N_408,In_1056,In_4885);
nand U409 (N_409,In_2836,In_4212);
and U410 (N_410,In_469,In_4384);
nor U411 (N_411,In_1019,In_4458);
nand U412 (N_412,In_1084,In_2682);
nand U413 (N_413,In_2906,In_235);
nor U414 (N_414,In_4078,In_3995);
nand U415 (N_415,In_801,In_2160);
nor U416 (N_416,In_4851,In_1071);
and U417 (N_417,In_3972,In_1631);
or U418 (N_418,In_4801,In_1663);
or U419 (N_419,In_177,In_1355);
and U420 (N_420,In_1628,In_2608);
nand U421 (N_421,In_3619,In_3531);
nand U422 (N_422,In_775,In_4215);
nand U423 (N_423,In_3944,In_1655);
nor U424 (N_424,In_4450,In_688);
nand U425 (N_425,In_400,In_1064);
or U426 (N_426,In_3103,In_3791);
and U427 (N_427,In_3524,In_1706);
or U428 (N_428,In_1180,In_2907);
nor U429 (N_429,In_3579,In_4697);
and U430 (N_430,In_2725,In_4426);
nor U431 (N_431,In_4756,In_3131);
nor U432 (N_432,In_187,In_2262);
xor U433 (N_433,In_21,In_2330);
nor U434 (N_434,In_3123,In_4634);
nor U435 (N_435,In_4033,In_3211);
and U436 (N_436,In_84,In_2688);
or U437 (N_437,In_1081,In_1735);
xor U438 (N_438,In_3167,In_4068);
nor U439 (N_439,In_2743,In_969);
nor U440 (N_440,In_4573,In_1147);
xor U441 (N_441,In_3808,In_818);
and U442 (N_442,In_834,In_4672);
nand U443 (N_443,In_1239,In_1102);
and U444 (N_444,In_2136,In_3280);
nand U445 (N_445,In_4330,In_2238);
or U446 (N_446,In_810,In_3236);
and U447 (N_447,In_2539,In_4261);
or U448 (N_448,In_2163,In_1346);
or U449 (N_449,In_4153,In_3442);
or U450 (N_450,In_355,In_139);
xnor U451 (N_451,In_1909,In_1086);
nand U452 (N_452,In_620,In_4211);
nand U453 (N_453,In_4044,In_1383);
nor U454 (N_454,In_4563,In_3540);
and U455 (N_455,In_3858,In_1917);
xnor U456 (N_456,In_1017,In_1388);
nand U457 (N_457,In_1161,In_2990);
nor U458 (N_458,In_984,In_2466);
nor U459 (N_459,In_2401,In_1627);
or U460 (N_460,In_1547,In_4317);
and U461 (N_461,In_3264,In_1290);
nand U462 (N_462,In_2374,In_3270);
nor U463 (N_463,In_2213,In_4880);
nor U464 (N_464,In_1197,In_3337);
and U465 (N_465,In_4298,In_855);
xor U466 (N_466,In_4780,In_4460);
or U467 (N_467,In_2589,In_3953);
and U468 (N_468,In_4436,In_2516);
and U469 (N_469,In_4788,In_3529);
nor U470 (N_470,In_4990,In_379);
nor U471 (N_471,In_2773,In_1494);
xnor U472 (N_472,In_103,In_2966);
or U473 (N_473,In_4451,In_193);
nor U474 (N_474,In_3570,In_2554);
or U475 (N_475,In_2605,In_3074);
nor U476 (N_476,In_4061,In_4300);
nor U477 (N_477,In_3377,In_1890);
nor U478 (N_478,In_3885,In_4341);
nor U479 (N_479,In_4971,In_2956);
nand U480 (N_480,In_98,In_3810);
nor U481 (N_481,In_421,In_2593);
xor U482 (N_482,In_4292,In_3174);
or U483 (N_483,In_1387,In_1227);
or U484 (N_484,In_1817,In_1485);
or U485 (N_485,In_594,In_4931);
nand U486 (N_486,In_2557,In_1575);
or U487 (N_487,In_432,In_1029);
nor U488 (N_488,In_4289,In_2575);
xnor U489 (N_489,In_1898,In_3187);
and U490 (N_490,In_1304,In_784);
nand U491 (N_491,In_342,In_495);
nand U492 (N_492,In_267,In_4094);
xnor U493 (N_493,In_4232,In_1569);
xor U494 (N_494,In_317,In_1242);
nor U495 (N_495,In_742,In_1191);
nand U496 (N_496,In_2880,In_2338);
and U497 (N_497,In_954,In_4140);
and U498 (N_498,In_2574,In_2537);
nor U499 (N_499,In_2346,In_1809);
or U500 (N_500,In_4396,In_3968);
xor U501 (N_501,In_1713,In_2766);
nand U502 (N_502,In_4772,In_1719);
xnor U503 (N_503,In_1429,In_1732);
or U504 (N_504,In_4313,In_1109);
or U505 (N_505,In_1259,In_2333);
and U506 (N_506,In_4675,In_2103);
or U507 (N_507,In_1295,In_1891);
xor U508 (N_508,In_975,In_1611);
or U509 (N_509,In_1236,In_3868);
nand U510 (N_510,In_4633,In_963);
nand U511 (N_511,In_2569,In_451);
and U512 (N_512,In_459,In_3385);
or U513 (N_513,In_1932,In_4491);
or U514 (N_514,In_3537,In_3734);
nor U515 (N_515,In_280,In_3266);
xor U516 (N_516,In_4000,In_1419);
and U517 (N_517,In_2050,In_1311);
nor U518 (N_518,In_850,In_4429);
nor U519 (N_519,In_2546,In_4870);
and U520 (N_520,In_4891,In_1833);
xor U521 (N_521,In_3036,In_1572);
nor U522 (N_522,In_1133,In_2650);
and U523 (N_523,In_1879,In_2048);
and U524 (N_524,In_925,In_300);
nor U525 (N_525,In_932,In_1219);
nand U526 (N_526,In_1589,In_4546);
or U527 (N_527,In_4046,In_2056);
xor U528 (N_528,In_696,In_563);
nand U529 (N_529,In_1282,In_615);
nor U530 (N_530,In_2925,In_1452);
nand U531 (N_531,In_2715,In_4677);
nand U532 (N_532,In_2444,In_4905);
xnor U533 (N_533,In_2463,In_3680);
nand U534 (N_534,In_697,In_1055);
and U535 (N_535,In_926,In_2277);
or U536 (N_536,In_4345,In_3215);
or U537 (N_537,In_3510,In_1170);
or U538 (N_538,In_2151,In_1873);
nand U539 (N_539,In_3740,In_2809);
nand U540 (N_540,In_4609,In_97);
nand U541 (N_541,In_1672,In_3905);
and U542 (N_542,In_1141,In_4737);
nor U543 (N_543,In_4506,In_1500);
nand U544 (N_544,In_2429,In_3659);
nor U545 (N_545,In_1095,In_3813);
nor U546 (N_546,In_1739,In_2280);
xnor U547 (N_547,In_4207,In_560);
nor U548 (N_548,In_1583,In_556);
and U549 (N_549,In_2887,In_3737);
nand U550 (N_550,In_2903,In_4267);
nor U551 (N_551,In_2196,In_2851);
nand U552 (N_552,In_4030,In_1195);
or U553 (N_553,In_3950,In_1559);
or U554 (N_554,In_4476,In_62);
nand U555 (N_555,In_468,In_2422);
or U556 (N_556,In_1128,In_166);
or U557 (N_557,In_4133,In_232);
or U558 (N_558,In_343,In_3909);
nor U559 (N_559,In_3128,In_4804);
nor U560 (N_560,In_2431,In_1847);
xor U561 (N_561,In_1288,In_2326);
xor U562 (N_562,In_3141,In_4049);
nand U563 (N_563,In_100,In_4686);
or U564 (N_564,In_3638,In_185);
nand U565 (N_565,In_28,In_1222);
or U566 (N_566,In_3347,In_43);
nor U567 (N_567,In_3408,In_4698);
nand U568 (N_568,In_1012,In_4565);
xor U569 (N_569,In_705,In_3039);
nand U570 (N_570,In_2949,In_907);
nor U571 (N_571,In_877,In_602);
nor U572 (N_572,In_3440,In_92);
xnor U573 (N_573,In_3982,In_3188);
nor U574 (N_574,In_1212,In_553);
nor U575 (N_575,In_2636,In_2996);
nand U576 (N_576,In_4027,In_1137);
and U577 (N_577,In_1601,In_2398);
nand U578 (N_578,In_2150,In_3355);
nand U579 (N_579,In_3720,In_4560);
nand U580 (N_580,In_4599,In_4293);
and U581 (N_581,In_4684,In_2664);
and U582 (N_582,In_38,In_3751);
nor U583 (N_583,In_4824,In_1318);
xnor U584 (N_584,In_2833,In_4892);
and U585 (N_585,In_453,In_3159);
or U586 (N_586,In_2411,In_2212);
xnor U587 (N_587,In_2547,In_2855);
nand U588 (N_588,In_2360,In_391);
nand U589 (N_589,In_2412,In_1751);
xor U590 (N_590,In_4918,In_1556);
and U591 (N_591,In_4610,In_3573);
nand U592 (N_592,In_3842,In_2913);
or U593 (N_593,In_1238,In_3144);
or U594 (N_594,In_3694,In_884);
xor U595 (N_595,In_4853,In_997);
and U596 (N_596,In_2419,In_3165);
or U597 (N_597,In_2812,In_3568);
and U598 (N_598,In_2615,In_4592);
nand U599 (N_599,In_504,In_3564);
nor U600 (N_600,In_2796,In_730);
xnor U601 (N_601,In_4818,In_4130);
nor U602 (N_602,In_2312,In_1527);
xor U603 (N_603,In_158,In_2509);
or U604 (N_604,In_1348,In_3289);
xnor U605 (N_605,In_93,In_2224);
and U606 (N_606,In_3617,In_2271);
xor U607 (N_607,In_347,In_4612);
and U608 (N_608,In_3946,In_970);
xor U609 (N_609,In_4825,In_428);
and U610 (N_610,In_625,In_528);
xor U611 (N_611,In_2606,In_541);
and U612 (N_612,In_1471,In_4536);
xnor U613 (N_613,In_1829,In_4855);
nor U614 (N_614,In_3623,In_4081);
nor U615 (N_615,In_1978,In_1600);
or U616 (N_616,In_1038,In_427);
nor U617 (N_617,In_1211,In_3170);
or U618 (N_618,In_4585,In_2979);
nand U619 (N_619,In_502,In_1955);
xnor U620 (N_620,In_1882,In_2125);
or U621 (N_621,In_4008,In_4359);
nand U622 (N_622,In_1904,In_3162);
xor U623 (N_623,In_2772,In_1952);
nand U624 (N_624,In_3554,In_446);
or U625 (N_625,In_680,In_761);
xor U626 (N_626,In_4614,In_3718);
or U627 (N_627,In_4724,In_898);
or U628 (N_628,In_3221,In_3733);
nand U629 (N_629,In_778,In_2945);
or U630 (N_630,In_1736,In_2828);
xor U631 (N_631,In_3333,In_848);
nand U632 (N_632,In_1050,In_3627);
xor U633 (N_633,In_2199,In_454);
and U634 (N_634,In_4644,In_746);
and U635 (N_635,In_4111,In_3338);
and U636 (N_636,In_222,In_2049);
and U637 (N_637,In_800,In_2679);
xor U638 (N_638,In_4742,In_4796);
or U639 (N_639,In_1150,In_3916);
nand U640 (N_640,In_2086,In_319);
xor U641 (N_641,In_3150,In_2819);
xor U642 (N_642,In_1949,In_1910);
nand U643 (N_643,In_2716,In_3010);
nand U644 (N_644,In_1075,In_499);
and U645 (N_645,In_3811,In_3653);
or U646 (N_646,In_4860,In_978);
or U647 (N_647,In_3760,In_1042);
and U648 (N_648,In_3647,In_1749);
xor U649 (N_649,In_4158,In_1608);
and U650 (N_650,In_2859,In_1399);
nand U651 (N_651,In_1362,In_878);
nand U652 (N_652,In_4263,In_3851);
and U653 (N_653,In_4721,In_1455);
nand U654 (N_654,In_3222,In_4381);
nor U655 (N_655,In_2905,In_3903);
xnor U656 (N_656,In_1326,In_3606);
nand U657 (N_657,In_3472,In_3757);
nand U658 (N_658,In_972,In_899);
and U659 (N_659,In_651,In_3060);
nor U660 (N_660,In_4364,In_1003);
nand U661 (N_661,In_1912,In_4306);
xnor U662 (N_662,In_2774,In_3522);
and U663 (N_663,In_2623,In_3781);
nor U664 (N_664,In_515,In_449);
or U665 (N_665,In_2603,In_1269);
nand U666 (N_666,In_3879,In_4138);
nor U667 (N_667,In_829,In_2396);
xnor U668 (N_668,In_1930,In_1853);
nor U669 (N_669,In_1907,In_2131);
nand U670 (N_670,In_2560,In_4976);
or U671 (N_671,In_3206,In_4485);
or U672 (N_672,In_3137,In_382);
nor U673 (N_673,In_337,In_648);
nand U674 (N_674,In_4480,In_4586);
xnor U675 (N_675,In_2918,In_1806);
nand U676 (N_676,In_3493,In_1693);
and U677 (N_677,In_2490,In_4674);
and U678 (N_678,In_3153,In_503);
or U679 (N_679,In_1393,In_2864);
nand U680 (N_680,In_2875,In_4362);
xor U681 (N_681,In_17,In_1883);
nor U682 (N_682,In_4389,In_552);
xor U683 (N_683,In_4826,In_4432);
and U684 (N_684,In_3208,In_1336);
xor U685 (N_685,In_2583,In_3112);
or U686 (N_686,In_1594,In_1005);
xor U687 (N_687,In_2214,In_3450);
nor U688 (N_688,In_4441,In_3098);
nor U689 (N_689,In_2625,In_2110);
nand U690 (N_690,In_3492,In_140);
or U691 (N_691,In_2645,In_760);
xnor U692 (N_692,In_534,In_3030);
nor U693 (N_693,In_4760,In_1605);
nor U694 (N_694,In_4496,In_331);
nand U695 (N_695,In_4557,In_4583);
nor U696 (N_696,In_3057,In_685);
xnor U697 (N_697,In_7,In_3025);
and U698 (N_698,In_3889,In_2815);
nand U699 (N_699,In_44,In_2562);
nand U700 (N_700,In_2404,In_756);
and U701 (N_701,In_950,In_161);
nand U702 (N_702,In_2545,In_335);
nand U703 (N_703,In_3945,In_4696);
or U704 (N_704,In_66,In_3940);
nor U705 (N_705,In_4722,In_4370);
nor U706 (N_706,In_1705,In_3448);
nand U707 (N_707,In_1057,In_1692);
nor U708 (N_708,In_3654,In_3300);
nor U709 (N_709,In_4735,In_4181);
xnor U710 (N_710,In_1926,In_4213);
nor U711 (N_711,In_1350,In_637);
xnor U712 (N_712,In_2789,In_1054);
and U713 (N_713,In_1561,In_1938);
or U714 (N_714,In_1331,In_621);
nand U715 (N_715,In_4255,In_4385);
nand U716 (N_716,In_4344,In_4558);
nand U717 (N_717,In_1010,In_2886);
or U718 (N_718,In_2436,In_2739);
nor U719 (N_719,In_768,In_3139);
and U720 (N_720,In_2055,In_489);
or U721 (N_721,In_3743,In_3615);
or U722 (N_722,In_3943,In_2973);
nor U723 (N_723,In_2553,In_2259);
nand U724 (N_724,In_4968,In_4257);
nand U725 (N_725,In_4499,In_4716);
and U726 (N_726,In_3223,In_1769);
or U727 (N_727,In_1372,In_3700);
nand U728 (N_728,In_1149,In_3920);
nand U729 (N_729,In_4116,In_1647);
nor U730 (N_730,In_1157,In_4805);
nor U731 (N_731,In_2243,In_543);
and U732 (N_732,In_3622,In_2730);
xor U733 (N_733,In_262,In_3919);
and U734 (N_734,In_1869,In_254);
or U735 (N_735,In_3559,In_1156);
nand U736 (N_736,In_1737,In_2255);
or U737 (N_737,In_4287,In_3839);
xnor U738 (N_738,In_3855,In_484);
or U739 (N_739,In_104,In_4650);
nand U740 (N_740,In_3308,In_269);
or U741 (N_741,In_894,In_3992);
nand U742 (N_742,In_1680,In_4911);
xnor U743 (N_743,In_4055,In_1317);
or U744 (N_744,In_4425,In_3897);
nand U745 (N_745,In_2995,In_4494);
nand U746 (N_746,In_491,In_4608);
nor U747 (N_747,In_1948,In_1824);
nor U748 (N_748,In_4687,In_2462);
and U749 (N_749,In_211,In_383);
and U750 (N_750,In_2610,In_1367);
nand U751 (N_751,In_1787,In_458);
or U752 (N_752,In_226,In_3732);
or U753 (N_753,In_554,In_2174);
xnor U754 (N_754,In_46,In_3753);
xnor U755 (N_755,In_4368,In_53);
or U756 (N_756,In_1696,In_3665);
xnor U757 (N_757,In_3014,In_4163);
xor U758 (N_758,In_3706,In_4881);
xnor U759 (N_759,In_3132,In_2221);
and U760 (N_760,In_1134,In_2854);
nor U761 (N_761,In_244,In_4605);
nor U762 (N_762,In_872,In_1785);
and U763 (N_763,In_1863,In_2807);
nor U764 (N_764,In_13,In_2594);
and U765 (N_765,In_311,In_1002);
xor U766 (N_766,In_361,In_3561);
xor U767 (N_767,In_3864,In_1107);
nor U768 (N_768,In_2649,In_3847);
or U769 (N_769,In_2514,In_3716);
nand U770 (N_770,In_3599,In_1685);
xnor U771 (N_771,In_3332,In_3421);
or U772 (N_772,In_3460,In_3661);
or U773 (N_773,In_2720,In_2385);
nand U774 (N_774,In_212,In_2286);
nand U775 (N_775,In_658,In_2447);
nor U776 (N_776,In_2335,In_3849);
and U777 (N_777,In_3658,In_1524);
or U778 (N_778,In_4972,In_57);
nand U779 (N_779,In_4797,In_3040);
nor U780 (N_780,In_442,In_3259);
and U781 (N_781,In_3396,In_2117);
nor U782 (N_782,In_2406,In_1264);
xor U783 (N_783,In_3521,In_4912);
and U784 (N_784,In_3157,In_4264);
or U785 (N_785,In_2197,In_846);
and U786 (N_786,In_3790,In_687);
nand U787 (N_787,In_1020,In_305);
nor U788 (N_788,In_4050,In_1790);
xor U789 (N_789,In_12,In_3690);
xnor U790 (N_790,In_4122,In_1368);
and U791 (N_791,In_3394,In_1422);
or U792 (N_792,In_2029,In_4074);
xnor U793 (N_793,In_526,In_2508);
nor U794 (N_794,In_833,In_2904);
or U795 (N_795,In_1660,In_802);
nor U796 (N_796,In_2034,In_4052);
and U797 (N_797,In_1023,In_4146);
or U798 (N_798,In_3361,In_3081);
nor U799 (N_799,In_1985,In_3624);
xor U800 (N_800,In_1553,In_4635);
and U801 (N_801,In_441,In_11);
xnor U802 (N_802,In_3587,In_2970);
nand U803 (N_803,In_3756,In_4240);
xor U804 (N_804,In_1831,In_14);
and U805 (N_805,In_4884,In_702);
nor U806 (N_806,In_4925,In_4431);
nand U807 (N_807,In_1762,In_1577);
or U808 (N_808,In_199,In_1122);
nor U809 (N_809,In_2181,In_329);
and U810 (N_810,In_1154,In_3311);
xor U811 (N_811,In_2345,In_763);
nand U812 (N_812,In_4022,In_4831);
and U813 (N_813,In_1168,In_605);
and U814 (N_814,In_4519,In_1139);
nand U815 (N_815,In_3175,In_1151);
nor U816 (N_816,In_1097,In_4366);
and U817 (N_817,In_4623,In_2270);
xnor U818 (N_818,In_2962,In_4538);
xor U819 (N_819,In_1511,In_3671);
xnor U820 (N_820,In_1565,In_2985);
and U821 (N_821,In_904,In_3901);
nor U822 (N_822,In_2737,In_883);
and U823 (N_823,In_616,In_3181);
xor U824 (N_824,In_2805,In_3741);
or U825 (N_825,In_2511,In_2010);
or U826 (N_826,In_1169,In_315);
xnor U827 (N_827,In_793,In_2997);
nor U828 (N_828,In_2535,In_2745);
xor U829 (N_829,In_523,In_889);
or U830 (N_830,In_1037,In_1939);
xor U831 (N_831,In_2916,In_1624);
nor U832 (N_832,In_73,In_4437);
and U833 (N_833,In_1576,In_4245);
or U834 (N_834,In_3350,In_4390);
xor U835 (N_835,In_4508,In_4901);
nor U836 (N_836,In_603,In_1498);
or U837 (N_837,In_1423,In_3104);
or U838 (N_838,In_1320,In_4256);
or U839 (N_839,In_1252,In_452);
and U840 (N_840,In_299,In_4201);
xnor U841 (N_841,In_1726,In_1741);
nand U842 (N_842,In_1903,In_49);
xnor U843 (N_843,In_2158,In_3993);
or U844 (N_844,In_3687,In_3990);
nand U845 (N_845,In_1456,In_171);
nand U846 (N_846,In_4067,In_2210);
and U847 (N_847,In_4559,In_2402);
and U848 (N_848,In_3583,In_1878);
xor U849 (N_849,In_600,In_2663);
nor U850 (N_850,In_1519,In_3436);
nor U851 (N_851,In_2172,In_4965);
nand U852 (N_852,In_4467,In_1481);
nor U853 (N_853,In_2953,In_1992);
and U854 (N_854,In_1695,In_3890);
or U855 (N_855,In_22,In_4405);
and U856 (N_856,In_3246,In_1229);
xnor U857 (N_857,In_2157,In_2140);
nor U858 (N_858,In_1578,In_4334);
or U859 (N_859,In_1793,In_3189);
nor U860 (N_860,In_3048,In_2523);
nor U861 (N_861,In_3099,In_3071);
nand U862 (N_862,In_2713,In_4139);
and U863 (N_863,In_3731,In_2276);
nor U864 (N_864,In_3357,In_4703);
nor U865 (N_865,In_2495,In_220);
or U866 (N_866,In_259,In_982);
xnor U867 (N_867,In_4303,In_1603);
and U868 (N_868,In_838,In_4607);
xor U869 (N_869,In_206,In_2536);
and U870 (N_870,In_2324,In_2355);
xnor U871 (N_871,In_597,In_4572);
or U872 (N_872,In_4148,In_4461);
nand U873 (N_873,In_2659,In_911);
xnor U874 (N_874,In_4637,In_119);
or U875 (N_875,In_4062,In_1262);
or U876 (N_876,In_4895,In_4890);
nand U877 (N_877,In_1047,In_3290);
and U878 (N_878,In_2147,In_3190);
nor U879 (N_879,In_1072,In_3838);
or U880 (N_880,In_4323,In_1484);
xor U881 (N_881,In_3837,In_91);
nand U882 (N_882,In_4333,In_2227);
nor U883 (N_883,In_1586,In_2219);
nor U884 (N_884,In_1755,In_325);
or U885 (N_885,In_1024,In_4840);
xnor U886 (N_886,In_1746,In_2467);
nand U887 (N_887,In_405,In_295);
and U888 (N_888,In_2129,In_2504);
nand U889 (N_889,In_393,In_1225);
nor U890 (N_890,In_1682,In_1062);
nand U891 (N_891,In_3681,In_1531);
nor U892 (N_892,In_4353,In_3682);
nand U893 (N_893,In_4930,In_887);
and U894 (N_894,In_4717,In_2332);
nor U895 (N_895,In_3886,In_909);
and U896 (N_896,In_902,In_2051);
nand U897 (N_897,In_3590,In_4427);
and U898 (N_898,In_2765,In_1971);
or U899 (N_899,In_546,In_1526);
nand U900 (N_900,In_759,In_221);
and U901 (N_901,In_4921,In_4400);
and U902 (N_902,In_2860,In_1887);
or U903 (N_903,In_1690,In_1811);
xnor U904 (N_904,In_4455,In_1204);
nor U905 (N_905,In_213,In_3752);
and U906 (N_906,In_3958,In_1356);
nor U907 (N_907,In_366,In_4848);
nand U908 (N_908,In_4076,In_542);
or U909 (N_909,In_2563,In_3376);
nor U910 (N_910,In_471,In_2137);
and U911 (N_911,In_2630,In_4168);
nor U912 (N_912,In_4524,In_843);
xnor U913 (N_913,In_1712,In_194);
nor U914 (N_914,In_2201,In_384);
nor U915 (N_915,In_4693,In_3125);
and U916 (N_916,In_1402,In_1514);
nand U917 (N_917,In_2770,In_2842);
and U918 (N_918,In_1287,In_4770);
nand U919 (N_919,In_4800,In_1363);
nand U920 (N_920,In_4100,In_1330);
xor U921 (N_921,In_1199,In_2291);
and U922 (N_922,In_3117,In_1192);
and U923 (N_923,In_360,In_4850);
nor U924 (N_924,In_3517,In_1707);
xnor U925 (N_925,In_339,In_3871);
nor U926 (N_926,In_4619,In_0);
nor U927 (N_927,In_2306,In_4090);
nor U928 (N_928,In_3371,In_493);
nor U929 (N_929,In_2620,In_3004);
and U930 (N_930,In_968,In_1474);
or U931 (N_931,In_1637,In_2524);
xnor U932 (N_932,In_866,In_2712);
or U933 (N_933,In_2223,In_783);
nor U934 (N_934,In_3829,In_2944);
nor U935 (N_935,In_720,In_2393);
and U936 (N_936,In_87,In_3981);
and U937 (N_937,In_3899,In_3534);
nor U938 (N_938,In_1397,In_4967);
and U939 (N_939,In_4142,In_2100);
or U940 (N_940,In_228,In_1360);
xnor U941 (N_941,In_1345,In_4807);
nand U942 (N_942,In_4617,In_4785);
xnor U943 (N_943,In_2409,In_1579);
nor U944 (N_944,In_2933,In_3245);
nand U945 (N_945,In_96,In_1001);
and U946 (N_946,In_3575,In_3597);
and U947 (N_947,In_3974,In_473);
xor U948 (N_948,In_1061,In_3015);
or U949 (N_949,In_2671,In_2343);
and U950 (N_950,In_3873,In_4128);
and U951 (N_951,In_72,In_4058);
xnor U952 (N_952,In_4244,In_2708);
nand U953 (N_953,In_664,In_4898);
nor U954 (N_954,In_4339,In_2233);
xor U955 (N_955,In_2315,In_921);
or U956 (N_956,In_4723,In_4652);
xor U957 (N_957,In_3341,In_601);
xor U958 (N_958,In_396,In_4421);
nor U959 (N_959,In_2204,In_4618);
nand U960 (N_960,In_1965,In_753);
xnor U961 (N_961,In_3629,In_706);
xor U962 (N_962,In_3596,In_2769);
or U963 (N_963,In_4280,In_1571);
xor U964 (N_964,In_463,In_1400);
nor U965 (N_965,In_1962,In_770);
and U966 (N_966,In_918,In_2258);
and U967 (N_967,In_341,In_3755);
or U968 (N_968,In_1625,In_998);
nand U969 (N_969,In_3675,In_4397);
and U970 (N_970,In_3547,In_2239);
nor U971 (N_971,In_415,In_3730);
nor U972 (N_972,In_993,In_946);
nor U973 (N_973,In_4239,In_1312);
or U974 (N_974,In_1412,In_3155);
xor U975 (N_975,In_2784,In_4057);
xnor U976 (N_976,In_3011,In_4075);
nor U977 (N_977,In_976,In_668);
or U978 (N_978,In_1000,In_4016);
and U979 (N_979,In_3961,In_2579);
xnor U980 (N_980,In_3976,In_3506);
xor U981 (N_981,In_431,In_3464);
nor U982 (N_982,In_4301,In_660);
xnor U983 (N_983,In_4879,In_1966);
xnor U984 (N_984,In_4034,In_2376);
nand U985 (N_985,In_3907,In_1004);
nand U986 (N_986,In_3331,In_15);
and U987 (N_987,In_1778,In_4986);
and U988 (N_988,In_4171,In_3565);
nand U989 (N_989,In_2510,In_25);
xnor U990 (N_990,In_147,In_3532);
nor U991 (N_991,In_617,In_223);
or U992 (N_992,In_2313,In_4227);
xor U993 (N_993,In_2037,In_3465);
nor U994 (N_994,In_3348,In_2867);
and U995 (N_995,In_2400,In_4129);
nor U996 (N_996,In_4708,In_1563);
or U997 (N_997,In_2445,In_561);
nor U998 (N_998,In_130,In_2629);
nor U999 (N_999,In_674,In_4907);
nor U1000 (N_1000,In_169,In_1473);
nor U1001 (N_1001,In_2926,In_4942);
or U1002 (N_1002,In_2818,In_4667);
or U1003 (N_1003,In_3567,In_2287);
and U1004 (N_1004,In_2921,In_2);
nor U1005 (N_1005,N_36,In_4616);
nand U1006 (N_1006,In_4836,In_3758);
and U1007 (N_1007,N_93,In_80);
and U1008 (N_1008,N_304,In_3298);
and U1009 (N_1009,In_910,In_157);
xor U1010 (N_1010,In_4273,In_809);
nor U1011 (N_1011,In_2571,In_4615);
xnor U1012 (N_1012,In_248,N_150);
nand U1013 (N_1013,In_2171,In_390);
nand U1014 (N_1014,In_257,N_219);
and U1015 (N_1015,In_2901,In_3676);
nand U1016 (N_1016,In_3317,In_985);
xnor U1017 (N_1017,In_1314,In_251);
nand U1018 (N_1018,In_2717,In_4516);
or U1019 (N_1019,In_1463,N_509);
or U1020 (N_1020,In_4628,In_40);
nand U1021 (N_1021,In_3998,In_1599);
and U1022 (N_1022,N_232,N_170);
xnor U1023 (N_1023,In_2071,N_588);
nand U1024 (N_1024,In_2735,In_4992);
nor U1025 (N_1025,In_37,N_596);
and U1026 (N_1026,In_133,In_2043);
nor U1027 (N_1027,N_985,In_2980);
and U1028 (N_1028,In_2135,In_3955);
nor U1029 (N_1029,In_4479,N_130);
and U1030 (N_1030,In_1366,N_397);
and U1031 (N_1031,In_4286,In_4229);
and U1032 (N_1032,In_3135,In_4182);
or U1033 (N_1033,In_2325,In_1428);
nand U1034 (N_1034,In_3870,In_2845);
or U1035 (N_1035,In_392,N_652);
nand U1036 (N_1036,In_3817,N_377);
xnor U1037 (N_1037,N_936,N_40);
nor U1038 (N_1038,In_3345,In_2395);
nor U1039 (N_1039,In_3928,In_1205);
xnor U1040 (N_1040,In_4754,N_518);
nand U1041 (N_1041,In_2816,N_66);
nand U1042 (N_1042,In_2430,In_1848);
and U1043 (N_1043,In_4728,N_503);
nor U1044 (N_1044,In_318,In_942);
and U1045 (N_1045,In_1391,In_3768);
or U1046 (N_1046,In_4304,In_3409);
or U1047 (N_1047,N_745,In_2781);
nand U1048 (N_1048,In_2643,In_3454);
xnor U1049 (N_1049,In_1548,In_4574);
and U1050 (N_1050,N_716,In_4622);
nand U1051 (N_1051,In_4793,In_2438);
nand U1052 (N_1052,In_4434,In_2381);
or U1053 (N_1053,In_4690,In_845);
xor U1054 (N_1054,N_584,N_783);
xnor U1055 (N_1055,In_4039,In_3378);
and U1056 (N_1056,In_4579,In_1268);
or U1057 (N_1057,In_538,In_1420);
xor U1058 (N_1058,In_522,In_1715);
nand U1059 (N_1059,N_784,In_2189);
xnor U1060 (N_1060,In_4743,N_822);
xnor U1061 (N_1061,In_1596,In_2667);
xnor U1062 (N_1062,In_1028,In_437);
nor U1063 (N_1063,In_1816,In_3261);
and U1064 (N_1064,In_3021,In_4010);
nand U1065 (N_1065,In_3461,In_3552);
and U1066 (N_1066,In_1792,In_947);
or U1067 (N_1067,In_3527,In_955);
or U1068 (N_1068,In_3563,In_871);
and U1069 (N_1069,N_780,In_35);
nor U1070 (N_1070,In_4332,N_340);
and U1071 (N_1071,In_2012,In_2651);
nor U1072 (N_1072,In_4041,In_518);
nor U1073 (N_1073,In_2727,In_1073);
or U1074 (N_1074,In_4525,In_1096);
nor U1075 (N_1075,N_676,In_1629);
or U1076 (N_1076,In_3397,In_4443);
or U1077 (N_1077,In_3749,In_2024);
nand U1078 (N_1078,N_81,In_3954);
or U1079 (N_1079,In_3930,N_83);
or U1080 (N_1080,In_2443,In_2634);
xor U1081 (N_1081,In_2319,N_544);
or U1082 (N_1082,In_1937,In_1609);
or U1083 (N_1083,In_4254,N_342);
xor U1084 (N_1084,In_2066,N_711);
nand U1085 (N_1085,In_3428,N_424);
and U1086 (N_1086,In_1777,In_3748);
nor U1087 (N_1087,In_2492,N_611);
nand U1088 (N_1088,In_1450,In_2942);
and U1089 (N_1089,N_71,In_3297);
nor U1090 (N_1090,In_4113,In_4252);
nor U1091 (N_1091,N_31,In_2230);
and U1092 (N_1092,In_3987,In_966);
nand U1093 (N_1093,N_436,In_3507);
and U1094 (N_1094,In_2141,In_3193);
and U1095 (N_1095,N_447,In_183);
or U1096 (N_1096,In_863,In_3457);
and U1097 (N_1097,In_24,In_4375);
or U1098 (N_1098,In_1702,In_3403);
and U1099 (N_1099,In_991,In_32);
or U1100 (N_1100,In_3848,In_2471);
nor U1101 (N_1101,In_3231,N_577);
xor U1102 (N_1102,In_2247,In_3854);
or U1103 (N_1103,N_963,N_568);
and U1104 (N_1104,In_512,N_924);
or U1105 (N_1105,N_344,In_234);
nor U1106 (N_1106,In_2637,In_3602);
xor U1107 (N_1107,In_3032,In_2008);
nand U1108 (N_1108,In_1510,In_385);
nand U1109 (N_1109,In_2094,N_486);
or U1110 (N_1110,In_3217,In_3200);
xnor U1111 (N_1111,In_1720,In_1543);
xor U1112 (N_1112,In_2923,N_521);
or U1113 (N_1113,In_413,In_3869);
or U1114 (N_1114,N_760,In_3241);
nand U1115 (N_1115,In_703,N_367);
nor U1116 (N_1116,In_1099,In_1986);
and U1117 (N_1117,In_4278,In_2797);
or U1118 (N_1118,In_1658,In_4086);
nand U1119 (N_1119,In_1045,N_838);
and U1120 (N_1120,In_4678,In_827);
or U1121 (N_1121,In_3875,In_3459);
xnor U1122 (N_1122,In_3108,In_3097);
nor U1123 (N_1123,In_151,In_209);
nor U1124 (N_1124,In_1775,In_3677);
or U1125 (N_1125,In_1711,N_755);
or U1126 (N_1126,In_835,In_3111);
nand U1127 (N_1127,In_1501,In_1752);
or U1128 (N_1128,In_3292,In_2299);
nand U1129 (N_1129,In_1552,In_2001);
xor U1130 (N_1130,In_4284,In_2798);
and U1131 (N_1131,In_638,In_4815);
nor U1132 (N_1132,In_1453,In_1068);
or U1133 (N_1133,In_4024,In_3318);
xor U1134 (N_1134,In_1982,In_3610);
xnor U1135 (N_1135,N_478,In_4069);
nor U1136 (N_1136,N_747,In_4629);
or U1137 (N_1137,In_1181,N_288);
and U1138 (N_1138,In_4088,In_4066);
xnor U1139 (N_1139,In_1700,N_912);
or U1140 (N_1140,In_3695,In_582);
and U1141 (N_1141,In_2759,In_773);
or U1142 (N_1142,N_921,In_3230);
xor U1143 (N_1143,In_496,N_981);
nand U1144 (N_1144,N_782,N_119);
nand U1145 (N_1145,N_623,N_636);
or U1146 (N_1146,In_4852,In_1036);
nand U1147 (N_1147,In_2211,In_681);
and U1148 (N_1148,N_79,N_395);
nand U1149 (N_1149,N_257,In_1819);
nor U1150 (N_1150,In_3389,In_578);
nand U1151 (N_1151,In_2683,N_870);
nor U1152 (N_1152,N_634,In_83);
xnor U1153 (N_1153,In_3260,In_3513);
xnor U1154 (N_1154,In_2755,N_998);
nand U1155 (N_1155,In_1158,In_159);
or U1156 (N_1156,N_319,N_691);
or U1157 (N_1157,In_2184,N_99);
and U1158 (N_1158,In_4445,N_554);
and U1159 (N_1159,In_979,In_1914);
or U1160 (N_1160,N_394,N_741);
and U1161 (N_1161,In_198,In_2591);
nor U1162 (N_1162,In_470,N_821);
nand U1163 (N_1163,N_212,In_3986);
and U1164 (N_1164,In_246,N_149);
nand U1165 (N_1165,In_271,In_2588);
xor U1166 (N_1166,In_1856,In_85);
or U1167 (N_1167,In_2304,In_1077);
xnor U1168 (N_1168,In_4060,In_1091);
xnor U1169 (N_1169,In_3366,In_16);
nand U1170 (N_1170,In_2915,N_899);
nand U1171 (N_1171,N_529,In_959);
nand U1172 (N_1172,N_686,In_3555);
xnor U1173 (N_1173,In_4464,In_3836);
or U1174 (N_1174,N_768,In_312);
and U1175 (N_1175,In_1106,In_1354);
nor U1176 (N_1176,In_3922,In_840);
nor U1177 (N_1177,N_559,In_4408);
or U1178 (N_1178,N_997,In_1973);
nor U1179 (N_1179,In_3678,In_3477);
nor U1180 (N_1180,In_1634,In_4556);
and U1181 (N_1181,In_4983,N_409);
nand U1182 (N_1182,N_903,In_1676);
nand U1183 (N_1183,In_2616,In_1564);
xor U1184 (N_1184,N_837,In_4695);
nand U1185 (N_1185,In_2661,In_1606);
and U1186 (N_1186,In_590,In_1503);
or U1187 (N_1187,In_377,In_3252);
nand U1188 (N_1188,In_3455,In_2967);
nand U1189 (N_1189,In_3989,In_2296);
xor U1190 (N_1190,In_168,In_700);
or U1191 (N_1191,In_4957,In_2099);
nand U1192 (N_1192,In_1309,N_507);
and U1193 (N_1193,In_3228,In_403);
nor U1194 (N_1194,In_1307,In_498);
nand U1195 (N_1195,N_391,N_914);
nor U1196 (N_1196,In_4963,In_4369);
and U1197 (N_1197,In_4193,In_48);
or U1198 (N_1198,N_364,In_1332);
nor U1199 (N_1199,In_245,In_4335);
nand U1200 (N_1200,In_3069,In_3003);
xnor U1201 (N_1201,In_2297,In_2485);
xor U1202 (N_1202,N_531,N_773);
and U1203 (N_1203,In_3328,In_654);
and U1204 (N_1204,In_1554,N_289);
nand U1205 (N_1205,In_1281,In_3553);
and U1206 (N_1206,In_3023,N_879);
and U1207 (N_1207,In_4954,In_1414);
and U1208 (N_1208,N_139,In_2841);
or U1209 (N_1209,N_496,In_2900);
nor U1210 (N_1210,N_449,In_2097);
or U1211 (N_1211,N_729,In_4092);
nand U1212 (N_1212,N_13,In_281);
or U1213 (N_1213,In_2052,N_311);
nand U1214 (N_1214,N_242,In_4899);
or U1215 (N_1215,In_1298,N_254);
and U1216 (N_1216,In_370,In_2366);
xor U1217 (N_1217,In_1927,In_3214);
xor U1218 (N_1218,N_147,In_4492);
xor U1219 (N_1219,In_1358,N_67);
or U1220 (N_1220,In_2585,N_58);
nor U1221 (N_1221,In_4856,N_667);
nor U1222 (N_1222,In_940,In_2027);
or U1223 (N_1223,N_762,In_4236);
nand U1224 (N_1224,In_3084,N_802);
xor U1225 (N_1225,In_129,N_546);
nand U1226 (N_1226,In_4655,In_709);
and U1227 (N_1227,In_1271,In_4729);
and U1228 (N_1228,In_1929,In_4875);
and U1229 (N_1229,N_572,In_4064);
nor U1230 (N_1230,In_4994,N_980);
or U1231 (N_1231,N_512,In_121);
nor U1232 (N_1232,In_2959,In_4706);
xor U1233 (N_1233,In_3642,In_2285);
and U1234 (N_1234,In_1970,In_4999);
and U1235 (N_1235,N_993,In_4004);
nor U1236 (N_1236,N_37,In_1142);
nor U1237 (N_1237,In_728,In_2790);
and U1238 (N_1238,In_2020,In_2321);
xor U1239 (N_1239,In_1528,In_1263);
nor U1240 (N_1240,In_2256,N_506);
nand U1241 (N_1241,In_2017,In_4002);
and U1242 (N_1242,N_348,In_399);
or U1243 (N_1243,In_3859,In_608);
nand U1244 (N_1244,N_934,N_883);
or U1245 (N_1245,In_4382,N_245);
nor U1246 (N_1246,In_3207,In_4471);
xor U1247 (N_1247,N_179,In_265);
or U1248 (N_1248,In_1027,In_2122);
xnor U1249 (N_1249,N_157,In_214);
nor U1250 (N_1250,In_4096,In_2014);
nand U1251 (N_1251,In_2162,In_4281);
or U1252 (N_1252,In_3835,In_2046);
nor U1253 (N_1253,In_285,In_2977);
nor U1254 (N_1254,In_4844,In_3393);
and U1255 (N_1255,In_2336,In_4713);
nand U1256 (N_1256,N_378,In_562);
nand U1257 (N_1257,In_1802,In_3729);
or U1258 (N_1258,N_967,In_4119);
nor U1259 (N_1259,N_396,In_995);
xor U1260 (N_1260,In_4838,In_4718);
xor U1261 (N_1261,In_2520,In_3204);
xnor U1262 (N_1262,In_2123,In_1686);
nor U1263 (N_1263,In_3353,In_2685);
xor U1264 (N_1264,In_3630,In_3701);
xnor U1265 (N_1265,In_309,In_302);
or U1266 (N_1266,In_639,N_573);
nand U1267 (N_1267,In_63,In_132);
or U1268 (N_1268,In_1815,In_568);
nor U1269 (N_1269,In_675,N_677);
or U1270 (N_1270,In_1280,N_556);
nand U1271 (N_1271,In_4758,In_2091);
and U1272 (N_1272,In_3445,In_3511);
nor U1273 (N_1273,In_1457,N_468);
nand U1274 (N_1274,In_805,In_4611);
nand U1275 (N_1275,In_138,In_4098);
nand U1276 (N_1276,N_454,N_632);
nor U1277 (N_1277,In_1981,N_330);
xor U1278 (N_1278,In_450,N_648);
or U1279 (N_1279,In_448,In_2722);
or U1280 (N_1280,N_666,In_2803);
xor U1281 (N_1281,N_333,In_2578);
and U1282 (N_1282,N_585,In_4151);
and U1283 (N_1283,In_1551,In_3545);
nand U1284 (N_1284,N_795,In_3476);
nor U1285 (N_1285,In_2640,N_646);
xnor U1286 (N_1286,N_829,In_4321);
or U1287 (N_1287,In_4183,In_4909);
nor U1288 (N_1288,In_394,In_2518);
and U1289 (N_1289,N_864,N_3);
xnor U1290 (N_1290,In_4679,In_2357);
nor U1291 (N_1291,In_481,In_4285);
and U1292 (N_1292,In_4018,In_4886);
or U1293 (N_1293,N_547,In_3395);
nor U1294 (N_1294,In_3800,N_180);
nand U1295 (N_1295,In_1476,N_142);
nor U1296 (N_1296,In_250,In_1251);
and U1297 (N_1297,N_917,In_445);
xnor U1298 (N_1298,In_3900,In_3914);
xnor U1299 (N_1299,In_1144,N_299);
and U1300 (N_1300,N_826,N_558);
or U1301 (N_1301,In_4529,In_4186);
xnor U1302 (N_1302,In_3054,N_194);
or U1303 (N_1303,In_1276,In_628);
and U1304 (N_1304,In_1381,N_498);
nand U1305 (N_1305,N_766,N_471);
nand U1306 (N_1306,In_1956,In_321);
nor U1307 (N_1307,In_1698,In_422);
nor U1308 (N_1308,In_4059,In_2519);
or U1309 (N_1309,In_2607,In_3360);
nand U1310 (N_1310,N_417,In_4404);
or U1311 (N_1311,In_3765,N_110);
or U1312 (N_1312,N_48,In_1060);
or U1313 (N_1313,In_402,In_1226);
nand U1314 (N_1314,In_3013,N_199);
or U1315 (N_1315,In_1983,In_4162);
xnor U1316 (N_1316,N_959,In_4038);
nor U1317 (N_1317,In_852,N_443);
nor U1318 (N_1318,In_613,In_941);
nand U1319 (N_1319,In_1493,N_842);
nor U1320 (N_1320,In_3806,In_1370);
nand U1321 (N_1321,N_225,In_4808);
nor U1322 (N_1322,N_128,N_904);
xnor U1323 (N_1323,In_4720,In_2496);
and U1324 (N_1324,In_1976,In_3059);
xor U1325 (N_1325,N_670,In_4026);
or U1326 (N_1326,In_3711,In_1742);
or U1327 (N_1327,In_4562,In_3180);
and U1328 (N_1328,In_4367,In_2359);
or U1329 (N_1329,In_4318,In_3016);
nand U1330 (N_1330,N_891,In_3685);
nand U1331 (N_1331,N_308,In_2470);
xnor U1332 (N_1332,In_4646,In_3866);
xnor U1333 (N_1333,In_439,N_950);
nand U1334 (N_1334,N_520,N_790);
nor U1335 (N_1335,In_3826,In_2657);
nand U1336 (N_1336,In_606,In_701);
or U1337 (N_1337,In_2994,N_616);
nand U1338 (N_1338,In_1604,In_869);
and U1339 (N_1339,In_10,In_2806);
nand U1340 (N_1340,In_4025,In_2477);
xnor U1341 (N_1341,In_3789,In_583);
xor U1342 (N_1342,In_4520,In_1011);
and U1343 (N_1343,In_1392,In_4358);
or U1344 (N_1344,In_1591,In_1417);
nand U1345 (N_1345,N_203,In_630);
and U1346 (N_1346,In_676,N_76);
xor U1347 (N_1347,In_2542,In_1537);
nand U1348 (N_1348,In_3463,In_3149);
nand U1349 (N_1349,N_707,In_3799);
nand U1350 (N_1350,In_1729,N_514);
and U1351 (N_1351,In_1717,N_960);
and U1352 (N_1352,In_3603,N_484);
nand U1353 (N_1353,N_316,In_719);
and U1354 (N_1354,In_4416,N_606);
or U1355 (N_1355,In_3055,In_3965);
xnor U1356 (N_1356,In_2061,In_4837);
and U1357 (N_1357,In_186,In_2107);
or U1358 (N_1358,N_132,In_4939);
and U1359 (N_1359,In_2232,In_3546);
and U1360 (N_1360,In_4392,N_739);
nor U1361 (N_1361,In_1825,In_2408);
or U1362 (N_1362,In_1065,In_2389);
and U1363 (N_1363,In_1889,In_4145);
and U1364 (N_1364,In_4077,In_4578);
nand U1365 (N_1365,In_1477,In_2253);
and U1366 (N_1366,In_596,In_2220);
and U1367 (N_1367,In_71,In_1854);
nand U1368 (N_1368,In_3005,In_2928);
nand U1369 (N_1369,In_623,N_201);
and U1370 (N_1370,In_4996,In_401);
nor U1371 (N_1371,In_2175,In_4734);
and U1372 (N_1372,In_1832,N_858);
nor U1373 (N_1373,In_2192,In_3778);
nand U1374 (N_1374,In_1296,In_3161);
nor U1375 (N_1375,In_2870,In_4247);
nor U1376 (N_1376,In_4597,In_1861);
or U1377 (N_1377,In_569,N_896);
and U1378 (N_1378,N_690,In_2205);
or U1379 (N_1379,In_2823,N_28);
or U1380 (N_1380,In_4121,In_733);
nand U1381 (N_1381,In_2248,In_1646);
and U1382 (N_1382,In_4326,N_86);
or U1383 (N_1383,In_2274,In_2072);
nand U1384 (N_1384,N_174,In_3490);
nor U1385 (N_1385,In_2164,In_897);
or U1386 (N_1386,In_2173,In_4778);
or U1387 (N_1387,In_2622,In_3276);
or U1388 (N_1388,N_236,N_714);
nor U1389 (N_1389,In_659,N_810);
nand U1390 (N_1390,In_1132,In_679);
nand U1391 (N_1391,In_4843,In_4157);
or U1392 (N_1392,In_3413,In_3535);
or U1393 (N_1393,N_307,In_1300);
nor U1394 (N_1394,In_4156,N_416);
and U1395 (N_1395,In_1858,In_1597);
or U1396 (N_1396,In_4951,In_3247);
or U1397 (N_1397,In_1207,In_3970);
nor U1398 (N_1398,In_3844,N_947);
or U1399 (N_1399,In_4564,In_836);
and U1400 (N_1400,In_4982,In_3592);
and U1401 (N_1401,In_4007,N_737);
nand U1402 (N_1402,N_926,In_497);
and U1403 (N_1403,In_2468,In_4645);
xnor U1404 (N_1404,N_976,In_1885);
nor U1405 (N_1405,N_151,In_4020);
and U1406 (N_1406,In_916,In_813);
nand U1407 (N_1407,In_1951,In_917);
xnor U1408 (N_1408,In_4580,In_3340);
and U1409 (N_1409,In_1469,In_3911);
nor U1410 (N_1410,In_4218,In_3793);
and U1411 (N_1411,In_4639,In_233);
or U1412 (N_1412,In_4747,N_840);
nor U1413 (N_1413,In_110,N_705);
or U1414 (N_1414,N_94,N_765);
xor U1415 (N_1415,In_4966,In_2302);
nand U1416 (N_1416,In_4446,In_3002);
nand U1417 (N_1417,In_924,N_731);
nor U1418 (N_1418,In_1125,N_155);
xor U1419 (N_1419,In_1213,N_393);
xor U1420 (N_1420,N_607,In_1727);
xor U1421 (N_1421,In_795,In_4108);
or U1422 (N_1422,In_1415,In_1850);
and U1423 (N_1423,N_587,In_3717);
xor U1424 (N_1424,N_723,In_2592);
nand U1425 (N_1425,In_2309,In_1175);
and U1426 (N_1426,N_165,In_3949);
xnor U1427 (N_1427,N_181,In_4505);
and U1428 (N_1428,In_508,In_3523);
nand U1429 (N_1429,In_4777,In_3904);
nand U1430 (N_1430,N_843,N_224);
or U1431 (N_1431,In_1960,In_4320);
xnor U1432 (N_1432,N_948,In_1549);
nand U1433 (N_1433,N_622,In_200);
or U1434 (N_1434,N_730,In_1088);
and U1435 (N_1435,In_3582,In_2742);
nor U1436 (N_1436,In_2244,In_2550);
nand U1437 (N_1437,In_4430,In_1895);
nor U1438 (N_1438,In_1622,In_663);
or U1439 (N_1439,In_238,In_36);
and U1440 (N_1440,In_460,In_3229);
nand U1441 (N_1441,In_433,N_645);
or U1442 (N_1442,N_75,In_824);
nand U1443 (N_1443,In_1386,In_4589);
or U1444 (N_1444,In_4176,N_470);
and U1445 (N_1445,In_324,N_931);
xor U1446 (N_1446,In_3834,In_3244);
xor U1447 (N_1447,In_1285,In_1665);
and U1448 (N_1448,In_576,In_440);
and U1449 (N_1449,In_4694,N_426);
or U1450 (N_1450,In_1803,In_3636);
nor U1451 (N_1451,N_649,In_2250);
nor U1452 (N_1452,In_544,In_3370);
xnor U1453 (N_1453,In_3160,In_162);
nand U1454 (N_1454,N_474,N_354);
and U1455 (N_1455,In_796,In_2927);
and U1456 (N_1456,N_152,In_782);
nand U1457 (N_1457,In_4897,In_4226);
and U1458 (N_1458,N_902,In_635);
nor U1459 (N_1459,In_2838,In_4829);
nand U1460 (N_1460,N_261,In_1094);
and U1461 (N_1461,In_4949,N_639);
nor U1462 (N_1462,In_3896,In_488);
nor U1463 (N_1463,In_1277,N_408);
or U1464 (N_1464,In_2968,In_2308);
or U1465 (N_1465,In_3284,In_1796);
or U1466 (N_1466,In_2484,In_943);
xnor U1467 (N_1467,In_1233,In_2454);
xnor U1468 (N_1468,In_3881,In_2225);
and U1469 (N_1469,In_831,In_4459);
or U1470 (N_1470,In_4265,In_1083);
nand U1471 (N_1471,In_973,In_1979);
nor U1472 (N_1472,In_367,In_117);
nand U1473 (N_1473,In_4262,N_504);
xnor U1474 (N_1474,In_74,In_1265);
or U1475 (N_1475,N_148,N_104);
or U1476 (N_1476,In_1619,In_1733);
nor U1477 (N_1477,In_634,In_381);
nand U1478 (N_1478,In_3020,N_265);
and U1479 (N_1479,In_812,In_494);
nor U1480 (N_1480,In_938,In_1562);
or U1481 (N_1481,In_517,N_186);
or U1482 (N_1482,N_953,In_999);
nor U1483 (N_1483,N_665,In_2754);
xor U1484 (N_1484,In_1768,In_3285);
or U1485 (N_1485,In_1515,In_2793);
and U1486 (N_1486,In_4762,N_365);
or U1487 (N_1487,In_971,In_3860);
xnor U1488 (N_1488,In_170,In_3410);
xor U1489 (N_1489,N_290,In_1327);
and U1490 (N_1490,In_1967,In_3975);
nor U1491 (N_1491,In_3240,N_562);
and U1492 (N_1492,In_643,In_2882);
and U1493 (N_1493,In_1774,N_258);
or U1494 (N_1494,In_3578,In_4647);
and U1495 (N_1495,N_193,In_4243);
xnor U1496 (N_1496,In_816,In_3035);
nand U1497 (N_1497,N_875,In_671);
nand U1498 (N_1498,In_3467,In_4322);
xor U1499 (N_1499,In_2740,N_384);
nand U1500 (N_1500,N_405,In_1826);
nor U1501 (N_1501,In_1928,In_537);
and U1502 (N_1502,N_599,In_3558);
or U1503 (N_1503,In_3631,N_517);
or U1504 (N_1504,N_785,In_1689);
and U1505 (N_1505,N_410,In_3556);
xnor U1506 (N_1506,N_602,In_3983);
nor U1507 (N_1507,In_1209,In_2760);
nand U1508 (N_1508,In_2695,N_266);
or U1509 (N_1509,N_123,N_673);
and U1510 (N_1510,In_4601,In_2917);
and U1511 (N_1511,In_4685,In_1176);
or U1512 (N_1512,In_3581,In_2045);
nor U1513 (N_1513,In_386,In_4624);
or U1514 (N_1514,In_501,In_4406);
xor U1515 (N_1515,In_2126,In_2924);
nand U1516 (N_1516,In_1860,N_250);
nor U1517 (N_1517,N_510,N_414);
nor U1518 (N_1518,In_1461,In_2292);
and U1519 (N_1519,In_1389,In_4545);
nor U1520 (N_1520,In_644,In_1146);
nand U1521 (N_1521,In_2965,N_566);
and U1522 (N_1522,N_429,In_882);
xor U1523 (N_1523,In_4356,In_2113);
and U1524 (N_1524,In_3807,In_588);
nor U1525 (N_1525,N_640,In_4533);
xor U1526 (N_1526,N_863,In_1080);
xor U1527 (N_1527,In_4103,In_2098);
and U1528 (N_1528,N_360,In_4682);
nand U1529 (N_1529,In_3667,In_4125);
or U1530 (N_1530,In_4845,In_2597);
or U1531 (N_1531,N_73,In_4547);
xor U1532 (N_1532,In_1006,In_189);
nor U1533 (N_1533,In_3105,In_710);
nand U1534 (N_1534,N_19,In_994);
nor U1535 (N_1535,N_418,In_713);
xnor U1536 (N_1536,N_35,In_3043);
nand U1537 (N_1537,In_1946,In_3312);
and U1538 (N_1538,In_1842,In_4509);
and U1539 (N_1539,N_56,In_3841);
nand U1540 (N_1540,In_2564,In_3456);
and U1541 (N_1541,In_4587,In_131);
and U1542 (N_1542,In_3140,N_725);
xor U1543 (N_1543,In_3648,In_3274);
xor U1544 (N_1544,In_1969,In_2863);
nand U1545 (N_1545,N_33,In_298);
nand U1546 (N_1546,In_4109,N_630);
and U1547 (N_1547,In_88,In_939);
and U1548 (N_1548,In_4861,N_594);
and U1549 (N_1549,In_3012,In_3483);
xnor U1550 (N_1550,In_3935,N_476);
nor U1551 (N_1551,In_529,N_7);
xor U1552 (N_1552,In_3942,In_2612);
xor U1553 (N_1553,In_3213,In_4028);
and U1554 (N_1554,N_657,In_3888);
and U1555 (N_1555,In_1786,N_275);
nand U1556 (N_1556,In_4202,N_469);
or U1557 (N_1557,In_1866,N_50);
xnor U1558 (N_1558,In_134,In_3106);
xor U1559 (N_1559,N_539,In_1550);
nand U1560 (N_1560,In_4412,In_3113);
and U1561 (N_1561,In_2459,In_2465);
nor U1562 (N_1562,In_4712,In_3613);
and U1563 (N_1563,In_3249,In_9);
and U1564 (N_1564,N_336,N_803);
and U1565 (N_1565,In_3469,In_4465);
nand U1566 (N_1566,In_4420,In_2372);
nand U1567 (N_1567,In_956,N_264);
or U1568 (N_1568,N_823,In_682);
and U1569 (N_1569,N_911,In_1808);
nand U1570 (N_1570,N_732,In_2689);
nor U1571 (N_1571,In_2128,In_673);
and U1572 (N_1572,In_1516,N_116);
nand U1573 (N_1573,In_2053,In_365);
or U1574 (N_1574,In_461,N_283);
and U1575 (N_1575,N_996,In_2111);
xor U1576 (N_1576,In_692,In_270);
and U1577 (N_1577,In_2435,In_624);
nand U1578 (N_1578,N_597,In_1540);
nand U1579 (N_1579,In_3452,In_2405);
xnor U1580 (N_1580,In_3795,N_746);
xnor U1581 (N_1581,In_1410,In_3843);
nor U1582 (N_1582,In_2595,In_1920);
or U1583 (N_1583,In_1260,In_1661);
or U1584 (N_1584,In_4632,In_2721);
nor U1585 (N_1585,In_3295,In_3572);
xnor U1586 (N_1586,N_98,In_888);
xor U1587 (N_1587,N_990,In_4235);
and U1588 (N_1588,In_2930,N_695);
nor U1589 (N_1589,In_988,In_1201);
xor U1590 (N_1590,In_1044,In_2804);
nand U1591 (N_1591,In_4123,In_4924);
nor U1592 (N_1592,In_3391,In_2399);
or U1593 (N_1593,N_215,In_3096);
xor U1594 (N_1594,In_3424,In_4568);
xor U1595 (N_1595,In_3679,N_533);
or U1596 (N_1596,N_804,In_1416);
xnor U1597 (N_1597,In_2628,In_2032);
nor U1598 (N_1598,N_816,N_681);
or U1599 (N_1599,In_2040,In_64);
nand U1600 (N_1600,In_2567,In_3321);
nor U1601 (N_1601,In_208,In_4962);
and U1602 (N_1602,In_1536,N_708);
nor U1603 (N_1603,N_222,In_3414);
xor U1604 (N_1604,In_4648,N_332);
nor U1605 (N_1605,In_4504,In_3022);
nand U1606 (N_1606,In_2340,N_781);
nand U1607 (N_1607,In_3857,In_2572);
or U1608 (N_1608,In_4401,In_4689);
or U1609 (N_1609,N_682,In_1538);
nand U1610 (N_1610,In_127,In_2869);
xor U1611 (N_1611,N_975,In_4641);
nand U1612 (N_1612,In_1919,In_740);
nand U1613 (N_1613,In_1467,In_2092);
and U1614 (N_1614,N_184,In_2779);
nand U1615 (N_1615,In_3745,In_1014);
or U1616 (N_1616,In_55,In_3883);
or U1617 (N_1617,In_3322,In_1830);
nand U1618 (N_1618,In_3614,In_3319);
nor U1619 (N_1619,N_624,In_3142);
nand U1620 (N_1620,In_4540,In_2351);
and U1621 (N_1621,N_43,In_3267);
or U1622 (N_1622,N_309,N_713);
or U1623 (N_1623,N_125,In_4846);
and U1624 (N_1624,In_1364,In_4023);
nand U1625 (N_1625,N_834,In_3713);
xnor U1626 (N_1626,In_3702,In_3805);
and U1627 (N_1627,N_890,In_3819);
xnor U1628 (N_1628,In_407,In_1744);
xnor U1629 (N_1629,In_4338,N_920);
nand U1630 (N_1630,In_2472,N_233);
nand U1631 (N_1631,In_3708,In_3915);
nand U1632 (N_1632,In_1517,N_989);
nand U1633 (N_1633,In_3689,In_4596);
or U1634 (N_1634,In_1722,In_2190);
and U1635 (N_1635,In_1460,In_4582);
nor U1636 (N_1636,N_575,In_524);
or U1637 (N_1637,In_1896,In_3533);
and U1638 (N_1638,In_2245,In_4948);
and U1639 (N_1639,In_4584,In_3382);
or U1640 (N_1640,In_1659,In_3474);
nand U1641 (N_1641,N_463,In_1357);
and U1642 (N_1642,In_1918,In_4683);
nor U1643 (N_1643,In_1394,N_861);
nor U1644 (N_1644,In_2390,N_617);
or U1645 (N_1645,N_905,In_195);
and U1646 (N_1646,In_2738,N_228);
and U1647 (N_1647,N_548,N_763);
nor U1648 (N_1648,In_1814,In_4487);
nand U1649 (N_1649,In_4771,In_2101);
or U1650 (N_1650,In_4154,In_1623);
or U1651 (N_1651,In_847,In_1079);
nor U1652 (N_1652,N_560,In_3574);
and U1653 (N_1653,In_1669,In_2526);
and U1654 (N_1654,In_2464,In_2417);
nand U1655 (N_1655,In_2428,N_272);
nand U1656 (N_1656,In_252,In_2382);
or U1657 (N_1657,In_1250,In_4365);
xor U1658 (N_1658,In_2919,In_1026);
xor U1659 (N_1659,In_2041,In_611);
xnor U1660 (N_1660,In_411,In_577);
nor U1661 (N_1661,In_4131,In_757);
or U1662 (N_1662,N_793,In_372);
nand U1663 (N_1663,In_4782,In_776);
and U1664 (N_1664,In_4513,In_215);
and U1665 (N_1665,In_106,In_1492);
nor U1666 (N_1666,In_3435,In_2696);
xor U1667 (N_1667,In_4383,In_4160);
and U1668 (N_1668,In_1980,In_3420);
xor U1669 (N_1669,In_649,In_718);
xor U1670 (N_1670,In_4640,In_2584);
or U1671 (N_1671,In_3874,In_4311);
and U1672 (N_1672,In_4453,In_4798);
or U1673 (N_1673,In_353,In_4175);
nor U1674 (N_1674,In_4775,In_2260);
xnor U1675 (N_1675,In_2350,In_2746);
or U1676 (N_1676,In_2517,In_4241);
or U1677 (N_1677,N_318,In_4127);
and U1678 (N_1678,N_277,In_1820);
and U1679 (N_1679,In_4208,In_820);
and U1680 (N_1680,In_2839,In_3422);
nand U1681 (N_1681,N_335,N_145);
nand U1682 (N_1682,In_3198,In_2893);
and U1683 (N_1683,In_4219,N_525);
or U1684 (N_1684,In_2347,In_4791);
and U1685 (N_1685,In_2912,In_1836);
nand U1686 (N_1686,In_2750,In_376);
or U1687 (N_1687,In_2505,In_336);
nand U1688 (N_1688,In_3372,In_4120);
or U1689 (N_1689,In_684,N_315);
nand U1690 (N_1690,In_2433,In_2473);
nor U1691 (N_1691,In_4015,N_115);
xor U1692 (N_1692,In_1642,In_3609);
nand U1693 (N_1693,In_4932,N_129);
nor U1694 (N_1694,N_187,In_3584);
nand U1695 (N_1695,In_1258,In_1651);
nor U1696 (N_1696,N_633,In_3618);
or U1697 (N_1697,In_2935,In_4266);
and U1698 (N_1698,In_20,In_4776);
nand U1699 (N_1699,N_994,N_255);
or U1700 (N_1700,In_1283,In_3635);
or U1701 (N_1701,In_3912,In_2448);
or U1702 (N_1702,In_3234,In_3077);
or U1703 (N_1703,N_208,In_2316);
nor U1704 (N_1704,N_6,In_3390);
nor U1705 (N_1705,In_913,N_992);
xor U1706 (N_1706,N_361,N_592);
nor U1707 (N_1707,N_831,In_276);
xnor U1708 (N_1708,N_349,In_933);
or U1709 (N_1709,N_664,In_294);
and U1710 (N_1710,N_805,In_3400);
and U1711 (N_1711,In_4566,In_4732);
xnor U1712 (N_1712,N_852,In_2992);
xor U1713 (N_1713,In_3342,In_2609);
nor U1714 (N_1714,N_446,In_2365);
xor U1715 (N_1715,In_478,N_300);
nand U1716 (N_1716,In_1677,N_329);
or U1717 (N_1717,In_1179,In_3404);
nand U1718 (N_1718,In_1688,In_2426);
nand U1719 (N_1719,In_1630,In_2352);
or U1720 (N_1720,In_2734,N_860);
xnor U1721 (N_1721,In_47,In_1043);
xnor U1722 (N_1722,N_452,In_4497);
nand U1723 (N_1723,In_4799,In_2850);
and U1724 (N_1724,N_522,In_3354);
xor U1725 (N_1725,N_684,N_90);
xnor U1726 (N_1726,In_4161,In_3049);
or U1727 (N_1727,In_1436,N_366);
xor U1728 (N_1728,N_256,N_352);
nand U1729 (N_1729,In_29,N_549);
xor U1730 (N_1730,In_2058,In_3185);
or U1731 (N_1731,N_800,In_1532);
xor U1732 (N_1732,In_3767,In_3947);
and U1733 (N_1733,In_2206,In_4764);
or U1734 (N_1734,In_1272,In_4248);
xor U1735 (N_1735,In_4606,In_937);
and U1736 (N_1736,In_3831,In_3562);
nand U1737 (N_1737,N_857,In_430);
and U1738 (N_1738,In_2108,N_302);
nand U1739 (N_1739,N_919,N_744);
xnor U1740 (N_1740,In_842,N_724);
or U1741 (N_1741,In_3569,In_1165);
or U1742 (N_1742,N_526,In_3779);
nand U1743 (N_1743,In_178,In_4813);
nand U1744 (N_1744,In_739,In_1194);
nor U1745 (N_1745,In_4859,In_4590);
xnor U1746 (N_1746,In_2573,In_2413);
nand U1747 (N_1747,N_39,In_2881);
nor U1748 (N_1748,N_295,In_2999);
and U1749 (N_1749,In_3576,In_2234);
or U1750 (N_1750,In_2991,In_4554);
nor U1751 (N_1751,In_1448,N_830);
xor U1752 (N_1752,N_983,N_398);
xnor U1753 (N_1753,In_263,In_1313);
xor U1754 (N_1754,In_1143,In_3664);
or U1755 (N_1755,In_2581,In_4037);
or U1756 (N_1756,In_65,In_3101);
or U1757 (N_1757,In_2853,N_877);
nor U1758 (N_1758,In_4029,In_571);
nor U1759 (N_1759,In_4388,In_4253);
or U1760 (N_1760,N_238,In_1316);
nand U1761 (N_1761,N_642,In_4507);
and U1762 (N_1762,In_645,In_1921);
xor U1763 (N_1763,In_3906,In_2544);
nor U1764 (N_1764,In_4725,In_4475);
nor U1765 (N_1765,N_34,In_1687);
or U1766 (N_1766,In_1520,In_656);
nand U1767 (N_1767,In_4926,In_2177);
xnor U1768 (N_1768,In_3772,In_2549);
xor U1769 (N_1769,N_578,In_4082);
or U1770 (N_1770,In_3127,In_3750);
nor U1771 (N_1771,In_2070,N_370);
xor U1772 (N_1772,In_3898,N_728);
and U1773 (N_1773,In_2821,In_4056);
or U1774 (N_1774,In_58,N_422);
xor U1775 (N_1775,In_1678,In_3484);
nand U1776 (N_1776,In_804,In_1953);
or U1777 (N_1777,N_751,In_4834);
nand U1778 (N_1778,In_4117,N_15);
xor U1779 (N_1779,In_3344,In_3001);
and U1780 (N_1780,In_2115,In_196);
or U1781 (N_1781,N_900,In_3499);
and U1782 (N_1782,N_227,In_1449);
nand U1783 (N_1783,In_3646,In_3375);
nor U1784 (N_1784,In_572,In_2846);
xnor U1785 (N_1785,In_4091,In_4553);
nand U1786 (N_1786,In_4980,In_1105);
and U1787 (N_1787,In_2425,In_3967);
nor U1788 (N_1788,In_4576,In_1846);
nor U1789 (N_1789,In_744,N_687);
or U1790 (N_1790,N_376,In_2947);
and U1791 (N_1791,In_1539,In_886);
or U1792 (N_1792,N_656,In_1943);
nor U1793 (N_1793,In_2479,In_1445);
nor U1794 (N_1794,N_528,N_167);
or U1795 (N_1795,In_3076,N_490);
or U1796 (N_1796,N_812,In_2503);
nand U1797 (N_1797,N_701,N_101);
nand U1798 (N_1798,N_710,In_2694);
nand U1799 (N_1799,In_2543,In_667);
xnor U1800 (N_1800,In_960,N_347);
xnor U1801 (N_1801,N_248,In_1478);
nor U1802 (N_1802,In_3894,In_2002);
nand U1803 (N_1803,In_745,In_181);
and U1804 (N_1804,In_3887,In_3656);
and U1805 (N_1805,In_832,In_598);
and U1806 (N_1806,In_4297,N_609);
and U1807 (N_1807,In_3094,In_1936);
and U1808 (N_1808,N_479,N_767);
or U1809 (N_1809,In_2824,In_3367);
nand U1810 (N_1810,In_3655,In_3959);
and U1811 (N_1811,N_579,N_445);
xnor U1812 (N_1812,In_711,In_3612);
nor U1813 (N_1813,N_570,In_2087);
nand U1814 (N_1814,In_1612,In_2613);
or U1815 (N_1815,N_412,N_259);
nor U1816 (N_1816,In_1266,In_2060);
and U1817 (N_1817,N_564,In_2452);
and U1818 (N_1818,In_2424,In_2814);
nand U1819 (N_1819,In_240,In_1409);
and U1820 (N_1820,In_2635,In_3053);
xnor U1821 (N_1821,N_962,In_2783);
xor U1822 (N_1822,In_4613,In_3759);
nand U1823 (N_1823,N_565,In_3744);
and U1824 (N_1824,In_3853,N_433);
nand U1825 (N_1825,In_146,In_2513);
nand U1826 (N_1826,In_587,In_116);
xnor U1827 (N_1827,N_23,In_2369);
nand U1828 (N_1828,In_2751,In_1231);
nand U1829 (N_1829,In_4809,N_106);
xor U1830 (N_1830,In_492,In_2675);
xnor U1831 (N_1831,In_1908,N_495);
or U1832 (N_1832,N_96,N_127);
nor U1833 (N_1833,N_788,N_759);
xnor U1834 (N_1834,In_3473,In_1795);
nand U1835 (N_1835,In_1502,In_205);
nor U1836 (N_1836,N_855,In_4474);
and U1837 (N_1837,In_3801,N_462);
or U1838 (N_1838,In_1584,N_721);
or U1839 (N_1839,N_345,In_2540);
and U1840 (N_1840,N_661,In_3114);
nor U1841 (N_1841,In_1944,In_2699);
xnor U1842 (N_1842,In_474,N_957);
nand U1843 (N_1843,In_4946,In_1289);
nor U1844 (N_1844,N_389,In_4343);
or U1845 (N_1845,In_4093,In_3257);
nor U1846 (N_1846,N_162,In_3310);
and U1847 (N_1847,In_2799,In_3721);
and U1848 (N_1848,In_1721,In_3929);
xor U1849 (N_1849,In_3988,In_4084);
xor U1850 (N_1850,In_3538,N_608);
nor U1851 (N_1851,N_274,N_97);
xor U1852 (N_1852,In_2726,In_86);
and U1853 (N_1853,In_1760,N_240);
xor U1854 (N_1854,In_722,In_4231);
or U1855 (N_1855,In_2387,In_1648);
xnor U1856 (N_1856,In_1876,N_114);
nand U1857 (N_1857,In_2646,In_1404);
and U1858 (N_1858,In_3303,N_441);
nand U1859 (N_1859,In_1337,In_2862);
or U1860 (N_1860,In_3846,In_2194);
xor U1861 (N_1861,In_1593,In_4448);
and U1862 (N_1862,N_698,In_3548);
nor U1863 (N_1863,In_2478,N_859);
xor U1864 (N_1864,In_2678,In_4537);
xnor U1865 (N_1865,N_87,In_2794);
and U1866 (N_1866,In_150,N_743);
nor U1867 (N_1867,In_1699,In_1812);
and U1868 (N_1868,In_1030,In_4670);
and U1869 (N_1869,In_912,In_3334);
or U1870 (N_1870,In_4380,In_774);
or U1871 (N_1871,In_4410,N_249);
or U1872 (N_1872,In_3299,In_4350);
or U1873 (N_1873,In_1654,In_841);
and U1874 (N_1874,In_1294,In_3458);
nand U1875 (N_1875,In_2075,In_2525);
nor U1876 (N_1876,In_4224,In_2529);
and U1877 (N_1877,In_3166,In_3495);
or U1878 (N_1878,In_4903,N_21);
nor U1879 (N_1879,In_4676,In_4288);
or U1880 (N_1880,In_4187,In_3272);
nand U1881 (N_1881,In_356,N_968);
or U1882 (N_1882,In_2506,In_3064);
or U1883 (N_1883,In_105,In_4857);
xnor U1884 (N_1884,In_4319,In_2498);
or U1885 (N_1885,In_4209,In_203);
and U1886 (N_1886,N_488,In_3158);
and U1887 (N_1887,N_668,In_1454);
and U1888 (N_1888,In_4688,N_278);
xor U1889 (N_1889,N_92,N_271);
nand U1890 (N_1890,N_466,In_1615);
and U1891 (N_1891,In_2078,In_3173);
xor U1892 (N_1892,In_4820,In_622);
xnor U1893 (N_1893,N_183,N_625);
nand U1894 (N_1894,In_4828,In_4087);
xnor U1895 (N_1895,In_1913,N_813);
nor U1896 (N_1896,In_2733,N_444);
and U1897 (N_1897,In_570,In_3219);
xor U1898 (N_1898,In_2031,In_3588);
nand U1899 (N_1899,In_426,In_2481);
xor U1900 (N_1900,In_2420,In_3645);
xnor U1901 (N_1901,N_613,In_896);
nor U1902 (N_1902,In_4251,In_2577);
nor U1903 (N_1903,In_3960,N_658);
and U1904 (N_1904,In_3288,In_1857);
xnor U1905 (N_1905,In_2368,In_4210);
nor U1906 (N_1906,In_4065,In_2895);
and U1907 (N_1907,In_694,In_1087);
nand U1908 (N_1908,In_2600,N_631);
nor U1909 (N_1909,In_691,In_665);
nor U1910 (N_1910,In_4447,In_1138);
nor U1911 (N_1911,In_256,In_2458);
or U1912 (N_1912,In_3462,N_778);
nand U1913 (N_1913,In_3938,N_662);
xor U1914 (N_1914,N_794,In_368);
and U1915 (N_1915,N_866,In_1870);
nand U1916 (N_1916,In_3316,In_81);
nand U1917 (N_1917,In_3195,N_820);
nor U1918 (N_1918,In_2179,N_74);
xnor U1919 (N_1919,In_3736,In_1103);
and U1920 (N_1920,N_282,In_539);
nor U1921 (N_1921,In_2096,In_4868);
nor U1922 (N_1922,In_476,In_2042);
or U1923 (N_1923,N_650,In_2283);
nor U1924 (N_1924,In_1136,In_1334);
nand U1925 (N_1925,N_873,In_2156);
xor U1926 (N_1926,In_2674,N_126);
xor U1927 (N_1927,In_1216,In_4011);
nor U1928 (N_1928,In_2655,In_2931);
xnor U1929 (N_1929,N_103,N_51);
nand U1930 (N_1930,In_527,In_4012);
nor U1931 (N_1931,In_655,In_4786);
or U1932 (N_1932,In_4115,In_1246);
nand U1933 (N_1933,N_943,In_2442);
or U1934 (N_1934,In_3498,In_467);
nor U1935 (N_1935,In_122,In_647);
nand U1936 (N_1936,In_2356,In_980);
nand U1937 (N_1937,N_419,In_201);
nor U1938 (N_1938,In_320,In_4484);
or U1939 (N_1939,In_2474,In_2825);
xor U1940 (N_1940,In_1488,In_4656);
nand U1941 (N_1941,In_2009,N_693);
or U1942 (N_1942,N_221,In_4987);
and U1943 (N_1943,N_182,In_962);
nand U1944 (N_1944,In_1754,N_638);
and U1945 (N_1945,In_1587,N_815);
xnor U1946 (N_1946,N_253,In_2780);
xor U1947 (N_1947,In_3650,N_176);
nor U1948 (N_1948,N_709,N_679);
or U1949 (N_1949,In_247,In_243);
xnor U1950 (N_1950,In_260,In_1171);
and U1951 (N_1951,In_4501,In_1761);
and U1952 (N_1952,In_4542,In_2461);
or U1953 (N_1953,In_4489,N_941);
nand U1954 (N_1954,In_4331,N_29);
or U1955 (N_1955,In_2028,In_4360);
and U1956 (N_1956,In_1256,In_936);
nand U1957 (N_1957,In_636,N_369);
or U1958 (N_1958,In_4167,In_4541);
and U1959 (N_1959,In_4933,N_748);
nand U1960 (N_1960,In_4936,N_872);
nor U1961 (N_1961,In_306,In_922);
nand U1962 (N_1962,N_825,In_525);
or U1963 (N_1963,In_137,In_409);
xnor U1964 (N_1964,N_519,In_4296);
or U1965 (N_1965,N_995,In_4952);
and U1966 (N_1966,N_453,N_346);
or U1967 (N_1967,In_184,In_3607);
or U1968 (N_1968,In_2499,N_647);
and U1969 (N_1969,In_2515,N_404);
nor U1970 (N_1970,In_1818,In_1580);
and U1971 (N_1971,In_3984,In_704);
nor U1972 (N_1972,In_4442,In_304);
nand U1973 (N_1973,In_2534,In_520);
nor U1974 (N_1974,In_3192,In_395);
or U1975 (N_1975,N_535,In_4781);
and U1976 (N_1976,In_3956,In_2884);
nor U1977 (N_1977,In_777,In_1375);
nand U1978 (N_1978,N_703,N_351);
xnor U1979 (N_1979,In_1302,In_4919);
xnor U1980 (N_1980,In_2723,In_4214);
or U1981 (N_1981,In_890,In_1497);
and U1982 (N_1982,In_3037,N_442);
nand U1983 (N_1983,In_2380,N_493);
or U1984 (N_1984,In_3090,In_4974);
nand U1985 (N_1985,In_76,In_1293);
nand U1986 (N_1986,In_1343,In_3764);
nand U1987 (N_1987,In_2166,In_2030);
xnor U1988 (N_1988,In_1206,N_915);
or U1989 (N_1989,In_4488,N_545);
nand U1990 (N_1990,N_534,In_4625);
xnor U1991 (N_1991,In_3425,N_68);
or U1992 (N_1992,In_3381,In_4230);
or U1993 (N_1993,In_1644,N_263);
nor U1994 (N_1994,In_3433,N_669);
xnor U1995 (N_1995,In_986,N_536);
nor U1996 (N_1996,In_1673,In_1581);
nor U1997 (N_1997,In_217,In_3611);
xor U1998 (N_1998,In_2339,In_2891);
nor U1999 (N_1999,In_1441,In_2834);
or U2000 (N_2000,In_1224,In_4398);
or U2001 (N_2001,In_885,In_4290);
nor U2002 (N_2002,N_1497,N_1843);
xnor U2003 (N_2003,N_154,In_2263);
nor U2004 (N_2004,In_857,N_1634);
or U2005 (N_2005,In_4468,N_1260);
or U2006 (N_2006,In_4051,N_1992);
or U2007 (N_2007,N_1079,In_752);
or U2008 (N_2008,N_143,In_3314);
nand U2009 (N_2009,In_4733,In_229);
nor U2010 (N_2010,In_4997,N_1706);
nand U2011 (N_2011,In_2943,In_4415);
nor U2012 (N_2012,In_2972,N_1209);
nor U2013 (N_2013,In_2951,In_715);
nand U2014 (N_2014,In_3182,In_2961);
or U2015 (N_2015,N_1722,In_873);
or U2016 (N_2016,In_2929,In_4469);
nor U2017 (N_2017,In_4943,N_1445);
xnor U2018 (N_2018,In_650,In_585);
xnor U2019 (N_2019,In_3343,In_3600);
nor U2020 (N_2020,In_4841,In_2134);
or U2021 (N_2021,N_1013,N_334);
and U2022 (N_2022,N_867,In_3163);
nor U2023 (N_2023,N_1395,In_4711);
xor U2024 (N_2024,N_1515,N_1425);
xnor U2025 (N_2025,In_2958,N_1169);
xor U2026 (N_2026,In_3725,In_2632);
nor U2027 (N_2027,N_432,N_1017);
xnor U2028 (N_2028,N_966,In_1639);
or U2029 (N_2029,N_1977,N_402);
and U2030 (N_2030,N_1826,In_3449);
nor U2031 (N_2031,N_502,In_595);
nor U2032 (N_2032,In_3951,N_1314);
or U2033 (N_2033,N_234,N_38);
xnor U2034 (N_2034,In_1671,N_551);
and U2035 (N_2035,N_84,In_1821);
and U2036 (N_2036,N_1704,In_3212);
nor U2037 (N_2037,N_1778,N_754);
nand U2038 (N_2038,In_1865,N_1066);
xor U2039 (N_2039,In_4761,N_358);
and U2040 (N_2040,In_39,In_2706);
nor U2041 (N_2041,In_4166,In_2222);
and U2042 (N_2042,N_1245,In_686);
xnor U2043 (N_2043,In_160,N_160);
nand U2044 (N_2044,In_1758,N_979);
or U2045 (N_2045,N_1712,In_4463);
and U2046 (N_2046,N_1254,In_1049);
nor U2047 (N_2047,N_1422,In_1491);
nand U2048 (N_2048,In_3832,In_3122);
xnor U2049 (N_2049,In_1110,In_3560);
nand U2050 (N_2050,In_2621,N_1660);
xor U2051 (N_2051,In_2844,N_53);
nand U2052 (N_2052,In_2394,N_1285);
xnor U2053 (N_2053,In_2067,In_2619);
xnor U2054 (N_2054,N_589,In_2782);
or U2055 (N_2055,In_3148,N_325);
nor U2056 (N_2056,N_1355,N_696);
xnor U2057 (N_2057,N_1407,N_1959);
xnor U2058 (N_2058,In_1684,N_1063);
nor U2059 (N_2059,N_886,N_55);
nand U2060 (N_2060,In_1667,N_827);
nand U2061 (N_2061,N_761,N_1705);
nand U2062 (N_2062,N_301,N_1647);
nand U2063 (N_2063,N_550,In_2801);
nor U2064 (N_2064,N_1539,In_436);
nand U2065 (N_2065,In_1950,N_218);
nand U2066 (N_2066,In_3503,N_1791);
and U2067 (N_2067,In_101,N_1136);
and U2068 (N_2068,N_1755,N_437);
and U2069 (N_2069,N_47,N_1218);
or U2070 (N_2070,N_1760,N_321);
or U2071 (N_2071,In_2731,N_100);
and U2072 (N_2072,In_2680,N_320);
nor U2073 (N_2073,In_2033,In_2026);
and U2074 (N_2074,In_4449,In_3589);
nor U2075 (N_2075,N_1085,N_1385);
and U2076 (N_2076,N_1200,In_314);
xnor U2077 (N_2077,N_1562,N_1543);
nor U2078 (N_2078,N_1906,In_1506);
xor U2079 (N_2079,N_1077,In_273);
nand U2080 (N_2080,N_1431,N_1989);
nand U2081 (N_2081,In_4823,N_1917);
nand U2082 (N_2082,In_819,N_1646);
and U2083 (N_2083,N_937,In_3910);
nor U2084 (N_2084,N_598,N_969);
xnor U2085 (N_2085,In_1116,N_1616);
or U2086 (N_2086,N_1321,In_3197);
and U2087 (N_2087,N_769,N_89);
or U2088 (N_2088,N_1239,In_1574);
or U2089 (N_2089,In_3301,In_2138);
or U2090 (N_2090,N_1093,In_274);
or U2091 (N_2091,In_2004,In_2022);
and U2092 (N_2092,In_4923,In_4327);
nand U2093 (N_2093,In_3416,N_1740);
or U2094 (N_2094,N_487,In_2681);
and U2095 (N_2095,N_1389,In_2626);
xor U2096 (N_2096,N_1728,In_398);
and U2097 (N_2097,In_1275,N_1192);
nand U2098 (N_2098,In_3323,In_3278);
nor U2099 (N_2099,N_1251,N_1969);
nor U2100 (N_2100,In_3539,N_1953);
nor U2101 (N_2101,N_874,N_343);
and U2102 (N_2102,N_1341,In_862);
xor U2103 (N_2103,In_3673,N_1583);
nand U2104 (N_2104,In_2116,In_2120);
nor U2105 (N_2105,N_1006,In_3315);
xor U2106 (N_2106,In_4402,N_1867);
nor U2107 (N_2107,N_1481,N_1398);
nor U2108 (N_2108,In_1617,In_3092);
xnor U2109 (N_2109,N_1749,In_1613);
xnor U2110 (N_2110,N_1584,In_350);
nor U2111 (N_2111,In_4833,In_2236);
nand U2112 (N_2112,N_1488,In_1254);
nor U2113 (N_2113,In_18,In_1541);
xor U2114 (N_2114,In_2974,N_1860);
or U2115 (N_2115,N_1159,In_1544);
nor U2116 (N_2116,N_1866,N_1080);
nand U2117 (N_2117,In_3330,N_1919);
or U2118 (N_2118,N_1292,In_923);
or U2119 (N_2119,In_3083,N_1930);
xor U2120 (N_2120,N_846,In_787);
xor U2121 (N_2121,In_2273,In_1482);
or U2122 (N_2122,N_1530,N_16);
xor U2123 (N_2123,In_4189,In_727);
nand U2124 (N_2124,N_1384,N_1101);
xor U2125 (N_2125,N_1976,N_1465);
nor U2126 (N_2126,In_1776,In_3339);
xnor U2127 (N_2127,In_1851,In_1349);
or U2128 (N_2128,N_935,In_1270);
or U2129 (N_2129,N_1480,In_1813);
and U2130 (N_2130,N_61,N_1912);
nor U2131 (N_2131,N_1566,N_267);
nand U2132 (N_2132,N_1994,N_583);
and U2133 (N_2133,In_754,N_1148);
nor U2134 (N_2134,N_1560,N_1027);
nor U2135 (N_2135,N_1614,In_4900);
or U2136 (N_2136,N_1761,N_987);
xor U2137 (N_2137,In_8,In_4928);
and U2138 (N_2138,N_1713,N_1520);
and U2139 (N_2139,N_1262,N_494);
nand U2140 (N_2140,In_3489,N_1296);
xnor U2141 (N_2141,In_514,In_4744);
or U2142 (N_2142,N_1776,N_1138);
nand U2143 (N_2143,In_2705,In_41);
and U2144 (N_2144,N_1880,N_482);
nor U2145 (N_2145,N_1030,In_771);
or U2146 (N_2146,N_322,In_2764);
nand U2147 (N_2147,N_1650,N_1940);
nor U2148 (N_2148,In_1100,N_381);
and U2149 (N_2149,In_163,N_901);
xnor U2150 (N_2150,N_175,In_2808);
nand U2151 (N_2151,N_371,N_1436);
nand U2152 (N_2152,N_1405,In_4534);
nor U2153 (N_2153,In_4847,In_4642);
nand U2154 (N_2154,N_591,N_1454);
nand U2155 (N_2155,In_1424,In_4376);
nand U2156 (N_2156,In_3451,In_4315);
nor U2157 (N_2157,N_399,In_870);
xnor U2158 (N_2158,In_4657,In_2079);
xor U2159 (N_2159,In_173,In_126);
xor U2160 (N_2160,In_323,In_3821);
and U2161 (N_2161,In_3431,N_618);
nor U2162 (N_2162,N_1765,N_1362);
nor U2163 (N_2163,In_530,In_781);
and U2164 (N_2164,In_1670,N_1388);
nand U2165 (N_2165,In_4377,N_1591);
nand U2166 (N_2166,In_3738,In_1297);
xor U2167 (N_2167,In_2861,N_1001);
nand U2168 (N_2168,N_719,N_971);
xnor U2169 (N_2169,N_1009,N_1931);
or U2170 (N_2170,In_1274,N_1112);
or U2171 (N_2171,N_1598,N_226);
xnor U2172 (N_2172,N_483,N_102);
and U2173 (N_2173,N_1268,In_2251);
xnor U2174 (N_2174,N_952,N_1466);
nor U2175 (N_2175,N_1391,N_1582);
xnor U2176 (N_2176,N_700,In_1763);
nor U2177 (N_2177,In_2124,N_1684);
or U2178 (N_2178,N_1835,N_824);
nor U2179 (N_2179,N_796,In_1178);
xor U2180 (N_2180,N_516,In_3816);
or U2181 (N_2181,N_1375,N_1152);
and U2182 (N_2182,In_466,In_1022);
nand U2183 (N_2183,In_927,N_1430);
and U2184 (N_2184,In_2827,N_383);
and U2185 (N_2185,In_148,N_1475);
nor U2186 (N_2186,In_3203,In_1435);
nor U2187 (N_2187,In_3979,In_4745);
nand U2188 (N_2188,In_1196,N_1683);
and U2189 (N_2189,In_1379,N_1226);
nand U2190 (N_2190,N_1350,In_4079);
xor U2191 (N_2191,N_1911,N_216);
or U2192 (N_2192,In_141,In_2802);
xor U2193 (N_2193,N_1164,N_1211);
xor U2194 (N_2194,In_2203,N_1746);
nor U2195 (N_2195,N_819,In_1406);
nand U2196 (N_2196,N_298,N_341);
and U2197 (N_2197,In_3256,N_492);
or U2198 (N_2198,In_4200,N_1916);
or U2199 (N_2199,In_4569,N_1386);
or U2200 (N_2200,In_197,N_1419);
or U2201 (N_2201,In_4021,In_3062);
or U2202 (N_2202,In_580,In_1991);
or U2203 (N_2203,N_923,N_1575);
xnor U2204 (N_2204,In_4347,In_3502);
nor U2205 (N_2205,In_4638,In_1339);
and U2206 (N_2206,In_3727,In_2269);
or U2207 (N_2207,In_406,N_949);
nor U2208 (N_2208,In_237,N_626);
nor U2209 (N_2209,In_3586,In_3501);
nand U2210 (N_2210,In_1101,N_1204);
and U2211 (N_2211,In_3481,In_3937);
or U2212 (N_2212,In_2437,In_1126);
nand U2213 (N_2213,In_4969,In_4522);
or U2214 (N_2214,N_1711,N_312);
or U2215 (N_2215,In_1545,In_1573);
and U2216 (N_2216,N_1411,N_758);
xnor U2217 (N_2217,In_59,N_702);
nand U2218 (N_2218,In_3296,In_607);
xor U2219 (N_2219,In_2813,N_1811);
xnor U2220 (N_2220,In_4896,N_303);
nor U2221 (N_2221,In_1111,N_1656);
or U2222 (N_2222,In_2551,N_1118);
or U2223 (N_2223,N_511,In_2216);
and U2224 (N_2224,In_1996,In_4054);
and U2225 (N_2225,In_2633,N_111);
xnor U2226 (N_2226,In_3120,N_610);
and U2227 (N_2227,In_4876,In_3070);
or U2228 (N_2228,N_323,In_2093);
nor U2229 (N_2229,In_3087,N_1392);
nand U2230 (N_2230,In_1845,In_3439);
xor U2231 (N_2231,In_4973,In_4393);
xnor U2232 (N_2232,In_974,N_603);
and U2233 (N_2233,N_60,In_2795);
or U2234 (N_2234,N_604,N_1965);
nor U2235 (N_2235,In_1187,In_357);
or U2236 (N_2236,In_2323,N_1939);
nand U2237 (N_2237,N_1752,In_1301);
nand U2238 (N_2238,N_1549,N_1351);
xnor U2239 (N_2239,In_2364,N_324);
and U2240 (N_2240,In_2538,N_1998);
xor U2241 (N_2241,In_176,In_3666);
nand U2242 (N_2242,N_1220,N_1470);
or U2243 (N_2243,In_876,In_3891);
nor U2244 (N_2244,N_1198,N_1443);
or U2245 (N_2245,N_1179,In_2753);
nor U2246 (N_2246,N_359,In_1459);
nor U2247 (N_2247,N_1837,N_475);
xnor U2248 (N_2248,In_3608,In_359);
xor U2249 (N_2249,N_764,N_72);
or U2250 (N_2250,N_229,In_2018);
xor U2251 (N_2251,In_2038,N_1067);
or U2252 (N_2252,In_3453,N_467);
xnor U2253 (N_2253,N_1674,In_1113);
or U2254 (N_2254,In_867,N_1876);
nor U2255 (N_2255,In_1942,In_2084);
nand U2256 (N_2256,In_815,N_1247);
and U2257 (N_2257,In_4959,In_1184);
xor U2258 (N_2258,In_619,In_1421);
xor U2259 (N_2259,N_27,In_3852);
nand U2260 (N_2260,N_1952,In_3683);
and U2261 (N_2261,N_1346,N_1955);
and U2262 (N_2262,N_1123,In_4944);
and U2263 (N_2263,N_1799,In_2198);
xor U2264 (N_2264,In_1306,N_1460);
nand U2265 (N_2265,N_1895,N_1521);
or U2266 (N_2266,In_1800,In_953);
and U2267 (N_2267,N_1213,In_1555);
or U2268 (N_2268,N_355,In_1167);
and U2269 (N_2269,N_1182,In_1021);
and U2270 (N_2270,N_1212,N_464);
nor U2271 (N_2271,In_2719,In_2301);
and U2272 (N_2272,In_1675,N_641);
or U2273 (N_2273,N_124,In_736);
xnor U2274 (N_2274,In_3827,In_2687);
or U2275 (N_2275,N_1933,In_3405);
xnor U2276 (N_2276,In_1234,N_689);
xor U2277 (N_2277,In_2541,In_45);
or U2278 (N_2278,N_1408,In_2275);
xnor U2279 (N_2279,In_2358,N_1918);
and U2280 (N_2280,In_788,In_4704);
xnor U2281 (N_2281,N_1259,In_3991);
nand U2282 (N_2282,N_472,In_1643);
xnor U2283 (N_2283,N_1222,N_1439);
nor U2284 (N_2284,N_1000,In_4539);
nand U2285 (N_2285,In_2011,In_4602);
and U2286 (N_2286,N_1231,N_108);
nand U2287 (N_2287,In_3833,In_4604);
xnor U2288 (N_2288,In_2648,N_1119);
xnor U2289 (N_2289,In_1957,N_1897);
and U2290 (N_2290,N_1495,In_4766);
or U2291 (N_2291,In_4661,N_1461);
and U2292 (N_2292,In_1632,In_4073);
nand U2293 (N_2293,N_1023,N_1418);
nor U2294 (N_2294,In_4170,N_1588);
nor U2295 (N_2295,In_4514,In_2371);
or U2296 (N_2296,In_3183,In_4195);
or U2297 (N_2297,N_1622,In_2015);
nand U2298 (N_2298,N_1358,N_1675);
xor U2299 (N_2299,N_1892,N_1950);
nor U2300 (N_2300,N_2,N_52);
and U2301 (N_2301,N_508,N_1637);
and U2302 (N_2302,N_246,In_2191);
nand U2303 (N_2303,In_4486,N_1004);
and U2304 (N_2304,In_4204,N_1537);
and U2305 (N_2305,N_1854,N_163);
nand U2306 (N_2306,In_3209,In_928);
and U2307 (N_2307,N_1464,In_1984);
nor U2308 (N_2308,In_283,In_2314);
nor U2309 (N_2309,In_4439,N_1215);
nand U2310 (N_2310,N_1738,N_1730);
nor U2311 (N_2311,In_2451,In_4032);
nand U2312 (N_2312,In_1240,In_4621);
xnor U2313 (N_2313,In_272,N_69);
xnor U2314 (N_2314,In_4197,N_1196);
xnor U2315 (N_2315,In_4934,N_1289);
and U2316 (N_2316,In_4874,N_1774);
xor U2317 (N_2317,N_284,N_1781);
and U2318 (N_2318,N_1783,In_1278);
and U2319 (N_2319,N_1810,In_4922);
xor U2320 (N_2320,N_1636,In_3362);
or U2321 (N_2321,N_1682,In_2180);
or U2322 (N_2322,N_1687,N_1579);
nor U2323 (N_2323,N_1010,N_1265);
or U2324 (N_2324,N_1472,In_4669);
nor U2325 (N_2325,In_3412,In_1221);
and U2326 (N_2326,In_1941,N_423);
and U2327 (N_2327,N_1991,In_4155);
nand U2328 (N_2328,N_1168,N_1036);
and U2329 (N_2329,In_3543,N_386);
nand U2330 (N_2330,N_1847,In_2920);
xnor U2331 (N_2331,N_1455,N_1451);
and U2332 (N_2332,In_1255,In_2295);
nor U2333 (N_2333,In_1323,N_247);
and U2334 (N_2334,In_2310,N_801);
or U2335 (N_2335,N_1404,In_1620);
and U2336 (N_2336,In_1875,In_1859);
nor U2337 (N_2337,N_1485,In_4950);
or U2338 (N_2338,N_1668,N_1850);
and U2339 (N_2339,N_1894,N_1029);
nor U2340 (N_2340,N_1035,In_1709);
nand U2341 (N_2341,In_4308,N_1437);
and U2342 (N_2342,In_3387,In_4752);
nor U2343 (N_2343,In_4205,N_1872);
nand U2344 (N_2344,N_1663,N_1197);
and U2345 (N_2345,N_651,In_352);
or U2346 (N_2346,N_85,N_141);
nor U2347 (N_2347,N_956,In_3604);
and U2348 (N_2348,N_1459,N_832);
or U2349 (N_2349,N_1373,N_9);
nor U2350 (N_2350,N_1050,N_1324);
and U2351 (N_2351,In_3526,N_1559);
or U2352 (N_2352,In_1093,In_2085);
and U2353 (N_2353,N_1891,N_291);
and U2354 (N_2354,N_1564,In_2521);
nor U2355 (N_2355,In_3777,In_2989);
and U2356 (N_2356,In_4324,In_3253);
nand U2357 (N_2357,In_1902,N_881);
and U2358 (N_2358,N_1606,In_3138);
nor U2359 (N_2359,N_136,N_1294);
nand U2360 (N_2360,N_1046,N_1482);
nor U2361 (N_2361,N_1555,In_1361);
and U2362 (N_2362,In_290,In_1267);
nand U2363 (N_2363,In_3688,In_708);
and U2364 (N_2364,N_736,N_451);
nor U2365 (N_2365,N_895,In_1053);
nand U2366 (N_2366,N_356,In_3147);
or U2367 (N_2367,In_2982,In_3512);
nand U2368 (N_2368,In_4221,In_4527);
xnor U2369 (N_2369,In_1738,In_2983);
and U2370 (N_2370,N_1686,N_1840);
xnor U2371 (N_2371,N_1553,N_1626);
or U2372 (N_2372,N_1874,In_919);
xnor U2373 (N_2373,N_1817,N_1946);
xor U2374 (N_2374,N_505,N_1185);
nor U2375 (N_2375,In_3644,In_477);
nor U2376 (N_2376,N_285,In_2215);
xnor U2377 (N_2377,N_1057,N_1848);
or U2378 (N_2378,N_1904,In_291);
nor U2379 (N_2379,N_1428,N_1261);
nand U2380 (N_2380,In_2829,N_717);
xnor U2381 (N_2381,N_1763,In_2349);
nor U2382 (N_2382,N_1217,In_2946);
nand U2383 (N_2383,In_772,In_860);
or U2384 (N_2384,In_1567,N_1089);
and U2385 (N_2385,N_1764,In_3402);
xor U2386 (N_2386,In_2692,N_230);
nand U2387 (N_2387,N_1069,In_4663);
or U2388 (N_2388,N_1631,N_1468);
xnor U2389 (N_2389,N_1941,N_379);
and U2390 (N_2390,N_1337,N_1525);
xnor U2391 (N_2391,In_591,In_4769);
nand U2392 (N_2392,N_1161,N_1467);
and U2393 (N_2393,N_1267,In_1322);
xor U2394 (N_2394,In_3585,In_30);
or U2395 (N_2395,N_1238,In_2502);
or U2396 (N_2396,In_3595,In_3325);
and U2397 (N_2397,In_4085,N_455);
nand U2398 (N_2398,In_207,N_1723);
xnor U2399 (N_2399,N_619,In_4794);
nand U2400 (N_2400,N_1055,In_4053);
or U2401 (N_2401,N_974,N_204);
and U2402 (N_2402,In_762,In_3707);
nor U2403 (N_2403,N_133,N_1277);
and U2404 (N_2404,N_553,N_1178);
and U2405 (N_2405,N_1898,In_661);
nor U2406 (N_2406,N_1597,In_4089);
nand U2407 (N_2407,N_1508,In_4822);
xor U2408 (N_2408,N_1383,N_1527);
nand U2409 (N_2409,In_1163,In_2457);
xor U2410 (N_2410,N_552,In_1855);
nand U2411 (N_2411,N_675,In_2639);
nor U2412 (N_2412,N_206,N_1073);
nor U2413 (N_2413,In_1483,N_1381);
and U2414 (N_2414,In_2362,N_1469);
xnor U2415 (N_2415,N_387,In_2872);
nor U2416 (N_2416,In_2057,N_24);
xnor U2417 (N_2417,In_2710,In_4970);
or U2418 (N_2418,In_4104,In_3320);
nand U2419 (N_2419,In_3763,In_1931);
or U2420 (N_2420,N_1975,N_1900);
xnor U2421 (N_2421,N_1410,In_4985);
or U2422 (N_2422,N_153,N_927);
and U2423 (N_2423,N_1456,N_1863);
xor U2424 (N_2424,In_1881,In_4329);
xnor U2425 (N_2425,N_940,In_3633);
xor U2426 (N_2426,In_2848,In_3923);
nor U2427 (N_2427,In_3818,In_4741);
xor U2428 (N_2428,N_1697,In_2527);
and U2429 (N_2429,N_1661,In_2161);
nor U2430 (N_2430,N_235,In_4152);
nor U2431 (N_2431,In_2892,In_750);
xor U2432 (N_2432,In_4309,N_1972);
nand U2433 (N_2433,In_1338,In_920);
nand U2434 (N_2434,N_1170,In_1007);
nor U2435 (N_2435,In_3009,In_4511);
nand U2436 (N_2436,N_853,N_1709);
nor U2437 (N_2437,In_1198,In_2068);
nor U2438 (N_2438,In_2976,N_909);
nor U2439 (N_2439,N_1233,In_3095);
and U2440 (N_2440,N_1114,In_3996);
or U2441 (N_2441,N_1323,N_456);
or U2442 (N_2442,In_2439,In_3672);
nor U2443 (N_2443,In_1924,In_2494);
and U2444 (N_2444,N_10,N_434);
xnor U2445 (N_2445,N_1556,N_1534);
and U2446 (N_2446,N_1082,N_146);
nand U2447 (N_2447,N_1271,N_1281);
and U2448 (N_2448,N_297,N_1804);
nor U2449 (N_2449,In_136,N_1621);
nand U2450 (N_2450,In_2497,N_327);
xnor U2451 (N_2451,N_1025,In_255);
nand U2452 (N_2452,N_1715,N_605);
or U2453 (N_2453,N_1869,In_175);
or U2454 (N_2454,N_757,N_1102);
nor U2455 (N_2455,N_1855,In_738);
or U2456 (N_2456,N_1581,In_3771);
nand U2457 (N_2457,N_1227,In_4664);
nand U2458 (N_2458,N_540,In_3882);
nand U2459 (N_2459,In_2732,In_2342);
and U2460 (N_2460,In_1468,In_4665);
and U2461 (N_2461,In_3093,N_1914);
nor U2462 (N_2462,In_990,N_91);
or U2463 (N_2463,N_1394,N_1762);
xnor U2464 (N_2464,N_1571,N_1278);
or U2465 (N_2465,In_4854,In_6);
and U2466 (N_2466,In_737,N_1990);
and U2467 (N_2467,N_14,In_51);
or U2468 (N_2468,N_339,In_4456);
nand U2469 (N_2469,In_811,In_1418);
nand U2470 (N_2470,In_1513,N_1087);
and U2471 (N_2471,In_1241,In_1035);
xnor U2472 (N_2472,N_1978,N_211);
nand U2473 (N_2473,In_726,In_915);
nor U2474 (N_2474,In_2747,In_3762);
and U2475 (N_2475,N_1845,In_948);
nor U2476 (N_2476,In_4570,In_4351);
xor U2477 (N_2477,In_4681,In_3352);
or U2478 (N_2478,In_3769,In_3151);
xor U2479 (N_2479,In_2035,In_1299);
and U2480 (N_2480,N_1165,In_2582);
and U2481 (N_2481,In_351,N_1157);
nor U2482 (N_2482,N_1708,N_1970);
nand U2483 (N_2483,N_933,In_3056);
nand U2484 (N_2484,N_1429,In_4374);
xor U2485 (N_2485,N_1172,In_2978);
nor U2486 (N_2486,N_63,In_3566);
and U2487 (N_2487,N_972,In_1766);
or U2488 (N_2488,N_1945,In_2704);
xnor U2489 (N_2489,In_155,In_1868);
xnor U2490 (N_2490,In_1214,N_986);
xnor U2491 (N_2491,In_3980,N_1105);
or U2492 (N_2492,In_2290,In_1114);
or U2493 (N_2493,N_1115,In_533);
nand U2494 (N_2494,N_78,N_1852);
or U2495 (N_2495,In_4668,N_884);
xnor U2496 (N_2496,N_1971,N_1532);
nand U2497 (N_2497,N_1298,In_2558);
and U2498 (N_2498,N_1693,N_1458);
and U2499 (N_2499,N_1979,N_185);
and U2500 (N_2500,N_1049,N_1028);
and U2501 (N_2501,N_168,N_172);
xor U2502 (N_2502,N_542,In_287);
nor U2503 (N_2503,In_3426,N_1827);
nor U2504 (N_2504,In_3709,In_4126);
or U2505 (N_2505,N_1100,N_1328);
nor U2506 (N_2506,N_749,In_266);
nor U2507 (N_2507,In_3632,In_1972);
nor U2508 (N_2508,N_1615,N_251);
and U2509 (N_2509,N_1580,N_1166);
or U2510 (N_2510,In_2684,N_970);
xnor U2511 (N_2511,N_1059,N_1828);
xnor U2512 (N_2512,In_3171,In_268);
nand U2513 (N_2513,N_1889,N_1618);
and U2514 (N_2514,In_1783,In_2998);
or U2515 (N_2515,N_1305,N_159);
and U2516 (N_2516,In_2178,N_0);
or U2517 (N_2517,N_787,N_41);
xnor U2518 (N_2518,In_2857,N_984);
xor U2519 (N_2519,In_4600,N_1493);
nand U2520 (N_2520,N_1716,In_113);
xor U2521 (N_2521,In_2552,In_4493);
and U2522 (N_2522,N_480,N_310);
xor U2523 (N_2523,N_1356,In_1390);
xor U2524 (N_2524,In_3356,N_286);
and U2525 (N_2525,In_1090,N_1075);
nor U2526 (N_2526,N_1147,N_1927);
xnor U2527 (N_2527,N_1011,N_1691);
or U2528 (N_2528,N_833,N_1453);
or U2529 (N_2529,In_416,In_1595);
nand U2530 (N_2530,In_4865,In_4830);
and U2531 (N_2531,N_678,N_1974);
or U2532 (N_2532,In_2183,In_548);
or U2533 (N_2533,In_4035,N_1542);
nor U2534 (N_2534,In_1922,In_2159);
nand U2535 (N_2535,In_4814,In_3079);
and U2536 (N_2536,In_695,In_165);
nand U2537 (N_2537,In_2596,In_859);
nand U2538 (N_2538,In_3129,N_1297);
nor U2539 (N_2539,N_1890,In_1823);
xnor U2540 (N_2540,In_2391,N_1293);
nor U2541 (N_2541,N_1187,N_1370);
nand U2542 (N_2542,N_1244,In_3783);
or U2543 (N_2543,N_913,N_1415);
nand U2544 (N_2544,N_1070,N_854);
xor U2545 (N_2545,N_1768,In_4937);
xor U2546 (N_2546,In_1347,N_1664);
nand U2547 (N_2547,N_954,In_2000);
and U2548 (N_2548,N_1331,N_1343);
or U2549 (N_2549,In_2388,N_1772);
nand U2550 (N_2550,In_3351,In_1530);
and U2551 (N_2551,In_4164,N_1985);
or U2552 (N_2552,In_1884,In_1512);
and U2553 (N_2553,N_326,In_4225);
nor U2554 (N_2554,In_3052,N_1357);
nand U2555 (N_2555,N_30,In_4188);
or U2556 (N_2556,In_1153,In_1708);
or U2557 (N_2557,In_4433,N_1246);
nand U2558 (N_2558,In_2284,In_1193);
nor U2559 (N_2559,In_2047,In_2003);
or U2560 (N_2560,In_2460,N_1864);
or U2561 (N_2561,In_457,In_3423);
and U2562 (N_2562,In_1877,In_599);
or U2563 (N_2563,In_1041,N_350);
and U2564 (N_2564,N_659,N_1002);
or U2565 (N_2565,N_742,N_1071);
nor U2566 (N_2566,In_4517,In_3329);
or U2567 (N_2567,In_4753,In_2941);
nor U2568 (N_2568,In_2533,N_601);
xnor U2569 (N_2569,In_3364,In_4352);
nor U2570 (N_2570,N_1750,N_1737);
nor U2571 (N_2571,N_1273,N_1748);
and U2572 (N_2572,N_835,In_779);
xor U2573 (N_2573,In_1697,In_1508);
nand U2574 (N_2574,N_1039,N_171);
and U2575 (N_2575,N_1679,N_1506);
and U2576 (N_2576,N_1753,In_67);
xnor U2577 (N_2577,N_1401,In_2440);
nand U2578 (N_2578,N_1449,N_1478);
xor U2579 (N_2579,N_1125,N_1150);
nand U2580 (N_2580,N_1505,N_1899);
nand U2581 (N_2581,N_1756,In_565);
xnor U2582 (N_2582,N_1139,N_1249);
and U2583 (N_2583,In_3917,In_1743);
xnor U2584 (N_2584,In_2267,In_2278);
xnor U2585 (N_2585,In_424,In_1916);
or U2586 (N_2586,N_808,N_22);
and U2587 (N_2587,In_3086,N_1317);
nand U2588 (N_2588,N_1842,N_1380);
nand U2589 (N_2589,In_822,N_1685);
or U2590 (N_2590,N_1951,N_156);
nand U2591 (N_2591,N_955,In_2019);
nand U2592 (N_2592,N_220,N_1836);
nor U2593 (N_2593,In_2729,In_455);
or U2594 (N_2594,In_1340,In_3479);
and U2595 (N_2595,N_1483,In_4591);
and U2596 (N_2596,N_293,N_1264);
nor U2597 (N_2597,N_694,N_1669);
nand U2598 (N_2598,In_4727,N_1541);
nand U2599 (N_2599,N_1423,In_1867);
xnor U2600 (N_2600,N_1657,In_4423);
nor U2601 (N_2601,N_489,In_3089);
nor U2602 (N_2602,In_4357,N_134);
or U2603 (N_2603,In_2293,In_4258);
xor U2604 (N_2604,In_2403,In_1714);
nand U2605 (N_2605,In_2528,N_252);
and U2606 (N_2606,N_1625,In_751);
nand U2607 (N_2607,N_1382,In_780);
or U2608 (N_2608,N_1736,In_4095);
nand U2609 (N_2609,In_2642,N_241);
nor U2610 (N_2610,In_4283,N_1725);
nand U2611 (N_2611,N_1037,In_1446);
xnor U2612 (N_2612,N_885,In_1753);
and U2613 (N_2613,N_1645,In_4871);
and U2614 (N_2614,In_2768,N_1773);
or U2615 (N_2615,N_1286,N_1270);
xor U2616 (N_2616,In_3202,N_1361);
nor U2617 (N_2617,In_2736,In_1118);
and U2618 (N_2618,In_4787,In_3823);
xor U2619 (N_2619,N_1742,In_747);
nor U2620 (N_2620,In_2888,N_363);
nand U2621 (N_2621,N_499,In_723);
xnor U2622 (N_2622,In_3497,N_1548);
nand U2623 (N_2623,In_2155,N_501);
nand U2624 (N_2624,N_1619,In_108);
and U2625 (N_2625,In_219,N_1325);
nand U2626 (N_2626,N_107,N_18);
nor U2627 (N_2627,In_1657,In_89);
xnor U2628 (N_2628,In_3383,N_543);
or U2629 (N_2629,N_1016,N_1417);
nand U2630 (N_2630,In_1351,N_1090);
nor U2631 (N_2631,N_862,In_3061);
or U2632 (N_2632,N_929,In_957);
and U2633 (N_2633,In_3346,N_1558);
or U2634 (N_2634,In_4913,N_1003);
xor U2635 (N_2635,N_1219,N_571);
nand U2636 (N_2636,N_1516,In_224);
nand U2637 (N_2637,N_1021,N_718);
nand U2638 (N_2638,In_1959,N_1720);
xnor U2639 (N_2639,In_823,N_362);
and U2640 (N_2640,N_223,In_2095);
xor U2641 (N_2641,N_1526,N_77);
nor U2642 (N_2642,N_999,In_2363);
or U2643 (N_2643,N_191,N_214);
xor U2644 (N_2644,In_2993,N_1096);
or U2645 (N_2645,N_1241,In_3058);
nand U2646 (N_2646,N_897,In_4740);
nor U2647 (N_2647,In_4910,N_1528);
or U2648 (N_2648,N_1031,In_142);
or U2649 (N_2649,N_1104,N_775);
and U2650 (N_2650,N_1144,In_3109);
or U2651 (N_2651,In_1378,N_1607);
or U2652 (N_2652,N_158,In_1864);
xor U2653 (N_2653,N_296,N_1958);
and U2654 (N_2654,In_1791,N_1909);
nand U2655 (N_2655,N_655,In_3130);
nor U2656 (N_2656,In_1947,N_635);
xor U2657 (N_2657,In_4817,N_1610);
nor U2658 (N_2658,N_1665,N_1177);
and U2659 (N_2659,N_1928,In_4419);
or U2660 (N_2660,In_4746,In_4150);
or U2661 (N_2661,In_1382,N_1908);
or U2662 (N_2662,In_303,In_1662);
nand U2663 (N_2663,In_4726,N_735);
and U2664 (N_2664,In_3598,In_3045);
and U2665 (N_2665,In_1458,In_1810);
nor U2666 (N_2666,N_1648,In_4960);
nor U2667 (N_2667,N_1308,N_368);
xor U2668 (N_2668,N_1142,In_3121);
xnor U2669 (N_2669,N_1873,In_4413);
xor U2670 (N_2670,N_841,N_1338);
nand U2671 (N_2671,N_653,N_1967);
nand U2672 (N_2672,N_1427,N_1288);
nand U2673 (N_2673,In_550,In_3220);
xor U2674 (N_2674,In_3265,In_1728);
nor U2675 (N_2675,N_663,N_582);
nor U2676 (N_2676,N_477,In_1245);
xnor U2677 (N_2677,In_4512,In_3812);
nand U2678 (N_2678,In_1112,In_1899);
and U2679 (N_2679,N_294,N_590);
or U2680 (N_2680,In_1679,In_2896);
and U2681 (N_2681,In_380,In_2007);
and U2682 (N_2682,N_1462,In_4991);
nand U2683 (N_2683,In_905,In_799);
nand U2684 (N_2684,N_1186,N_1412);
xor U2685 (N_2685,In_1009,N_699);
and U2686 (N_2686,N_1500,N_1595);
nand U2687 (N_2687,N_1106,N_1007);
or U2688 (N_2688,N_807,N_244);
xor U2689 (N_2689,N_1544,N_1739);
or U2690 (N_2690,In_3485,N_1201);
and U2691 (N_2691,N_1496,In_2910);
xor U2692 (N_2692,In_1140,N_109);
xor U2693 (N_2693,In_3470,In_2698);
and U2694 (N_2694,N_1690,In_1935);
and U2695 (N_2695,In_4399,N_1053);
or U2696 (N_2696,In_4409,N_1232);
xnor U2697 (N_2697,N_1300,In_1668);
or U2698 (N_2698,In_4101,N_1770);
nor U2699 (N_2699,N_1586,N_1365);
xor U2700 (N_2700,N_1224,N_1888);
or U2701 (N_2701,In_2565,In_4147);
xnor U2702 (N_2702,N_593,In_1964);
or U2703 (N_2703,N_916,In_1525);
and U2704 (N_2704,In_1740,In_4550);
nor U2705 (N_2705,In_1104,N_1859);
nor U2706 (N_2706,In_2073,N_1949);
nor U2707 (N_2707,N_1932,In_3398);
nand U2708 (N_2708,N_177,In_3178);
nor U2709 (N_2709,N_1514,In_3722);
nand U2710 (N_2710,N_1256,In_3867);
and U2711 (N_2711,N_1141,N_715);
and U2712 (N_2712,In_4714,N_1696);
nand U2713 (N_2713,N_1015,In_589);
or U2714 (N_2714,In_3282,N_1371);
xor U2715 (N_2715,N_1809,N_1176);
xor U2716 (N_2716,N_1137,N_513);
nor U2717 (N_2717,N_1628,N_1);
nand U2718 (N_2718,In_278,N_1507);
or U2719 (N_2719,In_3997,In_3024);
or U2720 (N_2720,In_344,N_1043);
xnor U2721 (N_2721,In_26,N_1272);
xnor U2722 (N_2722,In_3258,N_1915);
or U2723 (N_2723,In_798,In_191);
or U2724 (N_2724,In_358,N_1574);
or U2725 (N_2725,N_1886,N_1962);
xnor U2726 (N_2726,N_1963,N_753);
nand U2727 (N_2727,In_4340,N_279);
and U2728 (N_2728,In_1321,In_1683);
or U2729 (N_2729,N_1377,N_1019);
or U2730 (N_2730,In_1872,In_1747);
xnor U2731 (N_2731,In_3444,In_1934);
or U2732 (N_2732,N_1189,N_752);
or U2733 (N_2733,In_2627,In_4528);
and U2734 (N_2734,In_2771,In_3746);
xor U2735 (N_2735,N_1326,N_400);
xnor U2736 (N_2736,In_931,N_1807);
and U2737 (N_2737,N_600,In_483);
xnor U2738 (N_2738,N_1569,N_1446);
xor U2739 (N_2739,In_125,In_1480);
nor U2740 (N_2740,In_2914,N_1352);
xor U2741 (N_2741,In_2530,N_401);
nor U2742 (N_2742,In_1292,In_1650);
nor U2743 (N_2743,In_3365,In_1504);
xor U2744 (N_2744,N_1858,N_1632);
and U2745 (N_2745,In_375,In_2341);
and U2746 (N_2746,In_2778,N_1191);
nand U2747 (N_2747,N_1523,In_3963);
nand U2748 (N_2748,N_1140,In_3309);
and U2749 (N_2749,N_1083,N_450);
nand U2750 (N_2750,N_1345,N_1120);
and U2751 (N_2751,In_4883,N_1258);
and U2752 (N_2752,N_1937,In_284);
nand U2753 (N_2753,N_1074,In_4544);
or U2754 (N_2754,N_1617,In_2246);
nand U2755 (N_2755,N_581,In_2877);
nand U2756 (N_2756,N_1364,N_1964);
xor U2757 (N_2757,N_1195,In_2076);
nand U2758 (N_2758,In_4457,In_4177);
nand U2759 (N_2759,In_3369,In_4371);
and U2760 (N_2760,In_3865,N_1426);
xor U2761 (N_2761,In_2724,N_734);
and U2762 (N_2762,In_112,In_4889);
nand U2763 (N_2763,In_2586,In_4490);
nand U2764 (N_2764,N_54,In_4036);
or U2765 (N_2765,N_1202,N_481);
nor U2766 (N_2766,In_3964,In_1993);
and U2767 (N_2767,N_907,In_2453);
nor U2768 (N_2768,N_1434,In_3571);
nand U2769 (N_2769,In_397,In_4792);
nor U2770 (N_2770,In_1189,N_925);
nand U2771 (N_2771,In_2149,In_3742);
nor U2772 (N_2772,N_1276,In_4598);
nand U2773 (N_2773,N_269,In_3210);
nor U2774 (N_2774,N_1033,In_837);
nor U2775 (N_2775,N_1879,In_2456);
nor U2776 (N_2776,In_3374,N_1655);
or U2777 (N_2777,In_3136,In_90);
or U2778 (N_2778,In_903,In_4386);
xnor U2779 (N_2779,N_1275,N_1790);
nand U2780 (N_2780,In_3824,In_4510);
xnor U2781 (N_2781,In_2083,N_458);
and U2782 (N_2782,In_2167,N_1813);
or U2783 (N_2783,In_1731,N_1995);
nor U2784 (N_2784,N_1524,N_580);
xor U2785 (N_2785,N_1825,N_537);
or U2786 (N_2786,In_4518,N_420);
and U2787 (N_2787,N_1747,N_1639);
and U2788 (N_2788,N_231,In_764);
or U2789 (N_2789,N_1163,N_5);
nand U2790 (N_2790,In_1701,N_1966);
and U2791 (N_2791,N_11,N_674);
or U2792 (N_2792,N_105,In_900);
nor U2793 (N_2793,N_1390,N_1092);
xnor U2794 (N_2794,In_1411,N_660);
or U2795 (N_2795,In_2264,In_3447);
nor U2796 (N_2796,N_1585,In_3443);
nand U2797 (N_2797,N_189,In_3042);
and U2798 (N_2798,N_1681,In_2647);
xor U2799 (N_2799,In_1636,N_1721);
or U2800 (N_2800,N_1047,N_1076);
xnor U2801 (N_2801,N_1316,In_935);
or U2802 (N_2802,In_4355,N_615);
or U2803 (N_2803,In_3726,In_3530);
nor U2804 (N_2804,In_3380,In_1303);
xor U2805 (N_2805,In_410,N_1424);
xor U2806 (N_2806,In_1475,In_879);
nand U2807 (N_2807,N_1127,In_1365);
xor U2808 (N_2808,N_1733,In_1704);
or U2809 (N_2809,In_1,N_1576);
or U2810 (N_2810,In_4549,N_871);
xor U2811 (N_2811,In_3927,N_1041);
xor U2812 (N_2812,N_1203,N_1214);
nor U2813 (N_2813,N_1862,In_2229);
or U2814 (N_2814,In_1208,N_770);
xor U2815 (N_2815,N_847,N_1938);
xnor U2816 (N_2816,N_1567,N_1578);
xnor U2817 (N_2817,In_1495,In_3359);
and U2818 (N_2818,N_1190,In_2373);
or U2819 (N_2819,In_4277,N_1926);
nor U2820 (N_2820,In_1582,N_213);
nand U2821 (N_2821,N_1921,In_4132);
nand U2822 (N_2822,In_4915,N_353);
nand U2823 (N_2823,In_1123,N_1414);
or U2824 (N_2824,In_893,N_791);
nand U2825 (N_2825,N_1968,N_1406);
xnor U2826 (N_2826,In_3697,N_1519);
nor U2827 (N_2827,N_135,In_3494);
xnor U2828 (N_2828,N_1143,In_438);
and U2829 (N_2829,In_683,N_628);
or U2830 (N_2830,In_1408,N_1599);
nor U2831 (N_2831,In_2611,N_1934);
xor U2832 (N_2832,In_1405,In_3384);
or U2833 (N_2833,N_1235,N_1920);
and U2834 (N_2834,In_310,In_725);
xnor U2835 (N_2835,N_460,In_2059);
and U2836 (N_2836,In_509,In_1040);
xor U2837 (N_2837,In_3286,N_893);
xnor U2838 (N_2838,N_425,N_317);
nor U2839 (N_2839,In_3418,N_465);
or U2840 (N_2840,N_209,In_1888);
nand U2841 (N_2841,In_3926,N_733);
nand U2842 (N_2842,In_3263,N_849);
nand U2843 (N_2843,In_4141,In_1129);
and U2844 (N_2844,N_435,In_4768);
and U2845 (N_2845,In_4291,In_735);
and U2846 (N_2846,N_439,N_1536);
and U2847 (N_2847,In_549,N_614);
or U2848 (N_2848,In_2489,In_485);
nand U2849 (N_2849,In_4631,In_1063);
xnor U2850 (N_2850,In_4198,N_260);
nor U2851 (N_2851,N_806,N_1820);
or U2852 (N_2852,In_1034,In_1764);
nand U2853 (N_2853,In_4206,N_268);
or U2854 (N_2854,N_541,N_811);
nor U2855 (N_2855,In_2785,N_1551);
and U2856 (N_2856,N_59,In_1961);
nor U2857 (N_2857,In_4730,N_497);
nand U2858 (N_2858,N_1754,N_1432);
nand U2859 (N_2859,N_1240,In_2487);
and U2860 (N_2860,N_1330,In_2109);
xor U2861 (N_2861,In_2691,In_657);
and U2862 (N_2862,N_1335,N_1734);
nor U2863 (N_2863,N_1831,In_4165);
and U2864 (N_2864,N_415,In_4354);
and U2865 (N_2865,In_4275,In_99);
xnor U2866 (N_2866,N_1068,In_593);
and U2867 (N_2867,In_729,In_1235);
xnor U2868 (N_2868,In_2102,In_2418);
xnor U2869 (N_2869,N_1922,N_270);
or U2870 (N_2870,N_1794,N_64);
nand U2871 (N_2871,In_1664,In_19);
or U2872 (N_2872,N_173,N_1183);
and U2873 (N_2873,N_1484,In_2971);
nand U2874 (N_2874,N_1344,In_1046);
xor U2875 (N_2875,In_2476,In_1975);
nor U2876 (N_2876,N_1777,N_906);
and U2877 (N_2877,N_207,In_4523);
xor U2878 (N_2878,In_4978,In_4660);
xnor U2879 (N_2879,In_3427,N_1091);
xnor U2880 (N_2880,N_1857,N_26);
or U2881 (N_2881,In_1546,In_2434);
xor U2882 (N_2882,In_1433,N_1376);
xor U2883 (N_2883,N_1283,N_1318);
or U2884 (N_2884,In_716,In_2148);
xnor U2885 (N_2885,In_1098,N_1589);
xnor U2886 (N_2886,N_262,In_4105);
nor U2887 (N_2887,N_1098,N_1984);
or U2888 (N_2888,In_2964,N_1547);
xor U2889 (N_2889,In_1217,In_1342);
and U2890 (N_2890,N_1925,N_1757);
nor U2891 (N_2891,In_4070,N_1981);
and U2892 (N_2892,N_375,N_1780);
nor U2893 (N_2893,In_2955,N_1111);
or U2894 (N_2894,N_1741,In_4424);
xnor U2895 (N_2895,In_42,In_1626);
xor U2896 (N_2896,N_1688,In_4995);
nor U2897 (N_2897,N_1905,In_1341);
nor U2898 (N_2898,In_1999,In_4106);
xor U2899 (N_2899,N_1342,In_2354);
or U2900 (N_2900,N_1363,In_296);
or U2901 (N_2901,In_3047,In_4953);
nor U2902 (N_2902,In_4902,N_1116);
nor U2903 (N_2903,N_982,In_3031);
xnor U2904 (N_2904,In_3893,In_672);
xor U2905 (N_2905,N_1444,N_372);
or U2906 (N_2906,N_1779,N_1605);
nor U2907 (N_2907,In_629,N_1552);
and U2908 (N_2908,In_989,N_792);
and U2909 (N_2909,In_4237,N_1128);
xnor U2910 (N_2910,In_2441,N_1703);
nor U2911 (N_2911,N_1596,N_706);
nor U2912 (N_2912,N_382,N_1570);
or U2913 (N_2913,In_3172,In_3496);
nor U2914 (N_2914,In_3551,N_117);
and U2915 (N_2915,N_1789,N_1107);
xor U2916 (N_2916,N_113,In_2153);
or U2917 (N_2917,N_1194,N_1601);
or U2918 (N_2918,N_880,N_1158);
xnor U2919 (N_2919,In_1172,In_289);
nand U2920 (N_2920,In_586,In_3146);
nor U2921 (N_2921,N_1490,N_12);
and U2922 (N_2922,N_1448,N_1263);
and U2923 (N_2923,In_31,N_629);
and U2924 (N_2924,In_61,In_3417);
xor U2925 (N_2925,N_1870,N_1996);
or U2926 (N_2926,N_771,N_1957);
or U2927 (N_2927,N_688,In_4699);
xor U2928 (N_2928,In_853,N_1884);
nand U2929 (N_2929,In_3785,N_407);
or U2930 (N_2930,In_618,N_958);
or U2931 (N_2931,In_1618,N_817);
or U2932 (N_2932,In_2874,In_2817);
nor U2933 (N_2933,N_1563,N_814);
xnor U2934 (N_2934,In_662,In_3196);
and U2935 (N_2935,N_1727,In_4651);
nor U2936 (N_2936,N_80,In_4191);
or U2937 (N_2937,N_413,In_4014);
nor U2938 (N_2938,N_1184,In_3508);
nor U2939 (N_2939,N_865,N_178);
nor U2940 (N_2940,In_4336,N_1109);
or U2941 (N_2941,N_1099,N_876);
nor U2942 (N_2942,N_828,N_964);
and U2943 (N_2943,N_1311,N_411);
nor U2944 (N_2944,N_273,In_1403);
nor U2945 (N_2945,N_1907,In_2249);
or U2946 (N_2946,N_1048,In_2631);
nand U2947 (N_2947,In_2062,N_1399);
or U2948 (N_2948,In_1148,N_1154);
and U2949 (N_2949,In_2114,In_1694);
xnor U2950 (N_2950,N_198,N_1788);
or U2951 (N_2951,In_3724,In_4473);
or U2952 (N_2952,N_1044,N_1509);
nand U2953 (N_2953,N_888,N_1061);
nand U2954 (N_2954,N_1902,In_2146);
nand U2955 (N_2955,In_3505,In_3932);
nor U2956 (N_2956,In_4194,In_2119);
or U2957 (N_2957,N_637,In_2748);
or U2958 (N_2958,In_3478,N_672);
nand U2959 (N_2959,In_4958,In_408);
nand U2960 (N_2960,In_2130,In_2081);
or U2961 (N_2961,In_2044,N_1554);
and U2962 (N_2962,In_1353,N_1603);
or U2963 (N_2963,In_2911,N_1421);
or U2964 (N_2964,N_1121,N_1769);
nand U2965 (N_2965,In_1827,N_1206);
nand U2966 (N_2966,N_621,In_4867);
xnor U2967 (N_2967,In_1838,In_807);
xnor U2968 (N_2968,In_1610,N_1667);
nand U2969 (N_2969,In_2614,N_1269);
or U2970 (N_2970,N_928,In_4530);
nor U2971 (N_2971,N_1242,In_3591);
nor U2972 (N_2972,In_4849,N_1225);
xor U2973 (N_2973,N_1349,In_3770);
or U2974 (N_2974,In_3046,In_2693);
nand U2975 (N_2975,In_3825,N_388);
xnor U2976 (N_2976,N_557,N_1875);
xnor U2977 (N_2977,In_604,N_440);
or U2978 (N_2978,N_280,N_1883);
and U2979 (N_2979,N_1529,N_799);
nand U2980 (N_2980,In_107,N_1710);
and U2981 (N_2981,In_786,N_1644);
nand U2982 (N_2982,N_1903,N_1024);
xor U2983 (N_2983,In_3784,N_1751);
xnor U2984 (N_2984,N_1042,N_1255);
or U2985 (N_2985,N_1208,N_1162);
nand U2986 (N_2986,In_364,N_1402);
and U2987 (N_2987,N_1052,N_1237);
xnor U2988 (N_2988,In_4784,In_2837);
xnor U2989 (N_2989,In_4839,N_1374);
nor U2990 (N_2990,In_95,N_942);
nor U2991 (N_2991,In_1376,In_1505);
or U2992 (N_2992,N_137,In_814);
nor U2993 (N_2993,N_1018,N_1379);
or U2994 (N_2994,In_4955,In_3670);
nand U2995 (N_2995,In_2327,N_1856);
nor U2996 (N_2996,In_1542,In_1425);
xor U2997 (N_2997,N_1173,In_4521);
nor U2998 (N_2998,N_1279,N_1306);
xnor U2999 (N_2999,N_1122,In_149);
and U3000 (N_3000,In_5,In_1507);
or U3001 (N_3001,N_2348,In_3368);
and U3002 (N_3002,N_2571,In_3828);
xor U3003 (N_3003,N_1492,In_279);
nand U3004 (N_3004,In_1413,N_2457);
and U3005 (N_3005,N_2525,N_2379);
xnor U3006 (N_3006,N_1701,N_1732);
or U3007 (N_3007,N_2291,N_200);
or U3008 (N_3008,N_2324,N_2236);
xor U3009 (N_3009,N_2371,N_2798);
nand U3010 (N_3010,N_2906,N_774);
or U3011 (N_3011,N_704,In_1954);
or U3012 (N_3012,In_4438,N_2569);
and U3013 (N_3013,N_1815,N_2508);
xor U3014 (N_3014,N_2141,N_685);
and U3015 (N_3015,N_2862,In_2690);
nand U3016 (N_3016,In_326,N_2676);
nor U3017 (N_3017,N_2474,N_1193);
and U3018 (N_3018,N_740,N_2750);
or U3019 (N_3019,N_1814,In_856);
nor U3020 (N_3020,N_2488,N_2231);
nand U3021 (N_3021,N_2456,N_1689);
xor U3022 (N_3022,N_2184,N_2596);
nor U3023 (N_3023,N_2229,N_2036);
xor U3024 (N_3024,In_2446,N_2622);
nor U3025 (N_3025,In_3544,In_475);
nand U3026 (N_3026,In_3235,N_1816);
and U3027 (N_3027,N_2493,N_2182);
nand U3028 (N_3028,N_2900,N_2955);
or U3029 (N_3029,N_1387,In_821);
nand U3030 (N_3030,In_3652,N_2514);
xnor U3031 (N_3031,N_2331,N_2953);
nand U3032 (N_3032,In_4222,In_3415);
and U3033 (N_3033,In_1218,N_2113);
and U3034 (N_3034,N_2605,In_4391);
or U3035 (N_3035,N_1771,N_2185);
xnor U3036 (N_3036,N_2385,In_3616);
xor U3037 (N_3037,In_4945,N_2986);
or U3038 (N_3038,N_1699,N_2061);
nor U3039 (N_3039,N_2322,N_2151);
and U3040 (N_3040,N_2561,In_230);
nor U3041 (N_3041,N_2226,N_1366);
nand U3042 (N_3042,In_1228,N_1327);
xnor U3043 (N_3043,In_3251,N_2096);
nor U3044 (N_3044,In_4894,N_2294);
and U3045 (N_3045,N_2360,N_2079);
or U3046 (N_3046,In_2741,N_2806);
nor U3047 (N_3047,N_1347,N_1315);
xnor U3048 (N_3048,N_2347,N_2355);
nor U3049 (N_3049,N_2237,N_2188);
nor U3050 (N_3050,N_1248,N_2031);
and U3051 (N_3051,In_1933,N_2176);
nor U3052 (N_3052,N_1303,N_2729);
nor U3053 (N_3053,In_4893,N_2833);
nand U3054 (N_3054,N_2694,N_2942);
or U3055 (N_3055,N_1290,N_1797);
nand U3056 (N_3056,N_1097,N_2252);
or U3057 (N_3057,N_2821,N_932);
or U3058 (N_3058,In_2202,N_683);
and U3059 (N_3059,In_1773,N_2118);
and U3060 (N_3060,N_4,N_939);
and U3061 (N_3061,N_1322,N_2746);
and U3062 (N_3062,In_731,N_2111);
or U3063 (N_3063,N_1504,In_4917);
xor U3064 (N_3064,N_1887,In_1666);
nand U3065 (N_3065,N_2850,N_2894);
xor U3066 (N_3066,N_2831,N_2937);
and U3067 (N_3067,N_2202,N_2603);
or U3068 (N_3068,In_23,In_4348);
xor U3069 (N_3069,N_1620,In_3692);
xor U3070 (N_3070,In_4143,N_2480);
nand U3071 (N_3071,N_2004,N_2243);
and U3072 (N_3072,N_1367,N_2238);
xor U3073 (N_3073,In_875,N_197);
xor U3074 (N_3074,N_2144,N_2087);
nand U3075 (N_3075,N_2179,In_2407);
or U3076 (N_3076,In_3026,N_2645);
and U3077 (N_3077,N_2242,N_1149);
nand U3078 (N_3078,N_2208,In_2878);
and U3079 (N_3079,N_977,In_3237);
or U3080 (N_3080,N_1997,In_3068);
nor U3081 (N_3081,N_2044,In_4470);
or U3082 (N_3082,In_4581,N_2146);
or U3083 (N_3083,In_1640,N_2829);
xor U3084 (N_3084,N_779,N_2939);
nor U3085 (N_3085,N_17,In_4342);
nand U3086 (N_3086,N_2918,In_2090);
or U3087 (N_3087,In_4535,In_4302);
or U3088 (N_3088,N_1672,N_2993);
xnor U3089 (N_3089,N_1767,In_429);
nor U3090 (N_3090,N_2931,N_2957);
xnor U3091 (N_3091,In_4246,N_2784);
nor U3092 (N_3092,N_1072,N_2781);
xor U3093 (N_3093,N_2930,In_2240);
or U3094 (N_3094,In_3179,N_756);
and U3095 (N_3095,N_2470,In_2761);
and U3096 (N_3096,N_2110,N_431);
and U3097 (N_3097,N_2532,N_2015);
xor U3098 (N_3098,N_1378,N_2726);
xnor U3099 (N_3099,N_1942,In_765);
or U3100 (N_3100,N_2374,In_1305);
nor U3101 (N_3101,N_2914,N_1108);
nand U3102 (N_3102,N_2544,N_2977);
nor U3103 (N_3103,N_1171,N_2984);
or U3104 (N_3104,N_2919,In_3705);
nor U3105 (N_3105,N_1400,N_2978);
and U3106 (N_3106,N_2548,N_2203);
xnor U3107 (N_3107,N_1457,N_2905);
and U3108 (N_3108,N_1611,N_2206);
nand U3109 (N_3109,N_726,N_1302);
nand U3110 (N_3110,N_1174,N_2895);
nand U3111 (N_3111,N_1339,N_2691);
and U3112 (N_3112,N_1435,In_1237);
and U3113 (N_3113,N_2777,In_1074);
nand U3114 (N_3114,N_2414,N_2359);
or U3115 (N_3115,N_2134,N_2462);
xnor U3116 (N_3116,N_1846,N_2663);
xnor U3117 (N_3117,N_1499,In_4118);
xnor U3118 (N_3118,In_2089,N_2736);
and U3119 (N_3119,N_2126,N_1538);
and U3120 (N_3120,In_4418,N_1878);
nor U3121 (N_3121,N_2556,N_2879);
and U3122 (N_3122,N_2306,In_2714);
or U3123 (N_3123,In_1395,N_2416);
or U3124 (N_3124,N_2099,In_1185);
nor U3125 (N_3125,N_1792,N_2178);
xor U3126 (N_3126,N_2059,In_261);
nor U3127 (N_3127,N_2839,N_2244);
nand U3128 (N_3128,N_2959,N_2510);
or U3129 (N_3129,N_1805,N_2365);
nand U3130 (N_3130,N_2021,N_898);
nor U3131 (N_3131,N_2912,N_2199);
xor U3132 (N_3132,In_4680,N_2521);
xor U3133 (N_3133,In_4819,N_2787);
xor U3134 (N_3134,N_2153,N_1960);
nor U3135 (N_3135,N_2090,N_1731);
nor U3136 (N_3136,N_2800,N_380);
and U3137 (N_3137,N_2686,N_2799);
xnor U3138 (N_3138,N_2366,N_2629);
xor U3139 (N_3139,N_2539,N_2408);
xnor U3140 (N_3140,N_2450,N_2007);
xor U3141 (N_3141,In_689,N_2803);
or U3142 (N_3142,N_1929,N_1502);
nand U3143 (N_3143,N_2092,N_2611);
nand U3144 (N_3144,In_371,N_2357);
and U3145 (N_3145,N_1032,N_1056);
or U3146 (N_3146,N_2171,N_2391);
xor U3147 (N_3147,N_2191,N_2034);
nand U3148 (N_3148,N_1662,N_1221);
or U3149 (N_3149,N_2852,N_2297);
xnor U3150 (N_3150,N_2704,In_2756);
and U3151 (N_3151,N_2923,In_111);
nor U3152 (N_3152,N_2884,N_2478);
or U3153 (N_3153,N_1986,In_4626);
nand U3154 (N_3154,In_75,N_2681);
and U3155 (N_3155,N_2173,N_1333);
xor U3156 (N_3156,N_2782,In_4941);
nand U3157 (N_3157,N_2765,N_2965);
nand U3158 (N_3158,In_264,In_1220);
or U3159 (N_3159,N_1849,N_1823);
xnor U3160 (N_3160,N_2362,N_2672);
nor U3161 (N_3161,N_2116,N_2692);
and U3162 (N_3162,N_2473,N_1517);
and U3163 (N_3163,N_2254,N_2811);
xor U3164 (N_3164,N_57,N_8);
xor U3165 (N_3165,N_2094,In_2700);
nand U3166 (N_3166,N_237,N_2752);
nand U3167 (N_3167,N_2519,In_2936);
or U3168 (N_3168,In_1230,N_2251);
nand U3169 (N_3169,N_1452,N_2938);
and U3170 (N_3170,N_1329,In_4234);
nor U3171 (N_3171,In_3621,N_818);
nor U3172 (N_3172,N_1447,In_1032);
xnor U3173 (N_3173,N_2209,N_2581);
nor U3174 (N_3174,N_2886,N_2926);
nor U3175 (N_3175,N_2382,N_2258);
nor U3176 (N_3176,In_241,N_2721);
nand U3177 (N_3177,N_2792,N_2017);
nand U3178 (N_3178,N_2133,N_164);
or U3179 (N_3179,N_2654,N_1812);
nand U3180 (N_3180,N_2716,In_1897);
xnor U3181 (N_3181,N_1947,N_1759);
xor U3182 (N_3182,N_2971,N_2861);
and U3183 (N_3183,N_2985,N_2815);
nor U3184 (N_3184,N_2341,In_2195);
and U3185 (N_3185,N_1800,N_2644);
nor U3186 (N_3186,In_2200,N_2816);
and U3187 (N_3187,N_2826,In_4395);
and U3188 (N_3188,N_2342,N_563);
or U3189 (N_3189,N_2838,In_3803);
nor U3190 (N_3190,In_3388,N_2910);
nor U3191 (N_3191,N_2696,N_2313);
xor U3192 (N_3192,N_946,N_2896);
nor U3193 (N_3193,In_1145,N_292);
or U3194 (N_3194,N_2353,In_123);
and U3195 (N_3195,N_1565,N_643);
or U3196 (N_3196,N_2597,N_2832);
xor U3197 (N_3197,N_2709,N_2076);
nand U3198 (N_3198,N_1808,N_2817);
nor U3199 (N_3199,N_2275,N_2125);
or U3200 (N_3200,N_1086,In_2065);
and U3201 (N_3201,N_2536,N_2990);
xnor U3202 (N_3202,N_889,N_2227);
or U3203 (N_3203,In_1018,In_2077);
or U3204 (N_3204,N_2309,N_2602);
and U3205 (N_3205,In_2143,N_2628);
xnor U3206 (N_3206,In_4110,N_2310);
or U3207 (N_3207,In_646,N_2557);
or U3208 (N_3208,N_1360,N_2776);
xnor U3209 (N_3209,N_2738,N_188);
or U3210 (N_3210,N_2327,In_3933);
nand U3211 (N_3211,In_2548,N_1413);
xnor U3212 (N_3212,N_2925,N_2170);
or U3213 (N_3213,N_2156,In_2656);
xor U3214 (N_3214,N_2066,N_2160);
or U3215 (N_3215,N_2717,In_3168);
nor U3216 (N_3216,N_2859,N_2128);
and U3217 (N_3217,N_1729,N_1474);
or U3218 (N_3218,N_2995,N_2697);
and U3219 (N_3219,In_1871,In_521);
xor U3220 (N_3220,N_2162,N_1658);
and U3221 (N_3221,N_2135,N_2876);
and U3222 (N_3222,N_1677,In_3205);
nor U3223 (N_3223,N_2454,N_1501);
or U3224 (N_3224,N_2865,N_878);
and U3225 (N_3225,N_2576,In_2885);
nand U3226 (N_3226,N_2551,N_697);
nor U3227 (N_3227,In_1968,In_3124);
xor U3228 (N_3228,N_1640,In_2392);
xor U3229 (N_3229,In_3050,N_2403);
or U3230 (N_3230,In_4748,N_2659);
nand U3231 (N_3231,N_1822,N_2875);
nor U3232 (N_3232,N_2642,N_473);
nand U3233 (N_3233,N_2565,N_2293);
and U3234 (N_3234,In_3116,In_3620);
nor U3235 (N_3235,N_448,N_2713);
nor U3236 (N_3236,N_1282,N_2235);
xnor U3237 (N_3237,N_1320,N_2946);
or U3238 (N_3238,N_2677,N_2883);
nor U3239 (N_3239,In_444,N_1084);
or U3240 (N_3240,N_2277,In_699);
and U3241 (N_3241,N_2468,N_786);
nand U3242 (N_3242,N_2661,N_2268);
nor U3243 (N_3243,N_1726,N_2624);
nand U3244 (N_3244,N_2169,N_2073);
or U3245 (N_3245,N_2741,N_427);
nor U3246 (N_3246,N_2880,In_3549);
or U3247 (N_3247,N_2751,N_2409);
xnor U3248 (N_3248,N_2507,In_1598);
nand U3249 (N_3249,In_2168,N_373);
and U3250 (N_3250,N_1635,N_2728);
nor U3251 (N_3251,N_2584,N_2288);
xor U3252 (N_3252,N_140,N_2680);
and U3253 (N_3253,N_1652,In_109);
nand U3254 (N_3254,In_4864,N_2836);
nor U3255 (N_3255,In_4691,N_2108);
xnor U3256 (N_3256,N_527,N_1295);
nor U3257 (N_3257,N_2214,In_462);
and U3258 (N_3258,In_4866,N_1861);
xnor U3259 (N_3259,N_1113,N_1471);
xnor U3260 (N_3260,N_2014,In_2969);
xor U3261 (N_3261,In_3918,N_1511);
xor U3262 (N_3262,In_1159,In_3199);
or U3263 (N_3263,N_1348,N_1393);
xor U3264 (N_3264,N_2845,N_2593);
or U3265 (N_3265,N_2973,N_720);
or U3266 (N_3266,In_4984,N_2068);
nor U3267 (N_3267,In_3921,In_2475);
or U3268 (N_3268,N_2786,N_2037);
nand U3269 (N_3269,In_1533,N_2404);
nand U3270 (N_3270,In_1750,N_1936);
nor U3271 (N_3271,N_2049,In_797);
nand U3272 (N_3272,N_2967,N_2406);
nor U3273 (N_3273,N_2830,N_1250);
xnor U3274 (N_3274,N_2762,In_4707);
nand U3275 (N_3275,N_45,In_374);
xor U3276 (N_3276,In_653,N_2701);
xnor U3277 (N_3277,N_2030,N_2350);
and U3278 (N_3278,N_1369,N_2870);
nor U3279 (N_3279,In_4372,N_120);
or U3280 (N_3280,N_1561,N_2345);
xor U3281 (N_3281,N_2996,In_3051);
and U3282 (N_3282,N_2748,N_2055);
nand U3283 (N_3283,N_314,N_2158);
nor U3284 (N_3284,N_2361,N_2944);
nand U3285 (N_3285,N_2956,N_32);
xor U3286 (N_3286,N_2853,In_567);
xor U3287 (N_3287,N_2326,N_2020);
xor U3288 (N_3288,N_2490,N_2881);
or U3289 (N_3289,N_1821,In_2231);
and U3290 (N_3290,N_2755,N_2384);
nor U3291 (N_3291,N_118,N_2444);
and U3292 (N_3292,In_1344,N_2774);
xnor U3293 (N_3293,N_1442,N_1956);
xor U3294 (N_3294,N_2769,N_2949);
and U3295 (N_3295,N_2065,N_2107);
and U3296 (N_3296,N_2579,N_2898);
nor U3297 (N_3297,N_2432,N_2196);
nor U3298 (N_3298,N_2148,N_2181);
nor U3299 (N_3299,N_2968,N_2506);
nand U3300 (N_3300,N_406,N_2215);
and U3301 (N_3301,In_614,N_2766);
and U3302 (N_3302,N_1234,N_2212);
or U3303 (N_3303,N_2767,N_313);
and U3304 (N_3304,N_1510,In_3931);
or U3305 (N_3305,N_2377,In_225);
xor U3306 (N_3306,N_2641,N_2482);
and U3307 (N_3307,N_2280,N_2705);
xnor U3308 (N_3308,N_2868,N_1801);
or U3309 (N_3309,N_390,N_2623);
or U3310 (N_3310,N_2608,N_2916);
nor U3311 (N_3311,N_2523,N_738);
nor U3312 (N_3312,N_459,N_2335);
and U3313 (N_3313,N_2131,N_2303);
or U3314 (N_3314,N_2813,N_524);
or U3315 (N_3315,N_2999,In_3557);
and U3316 (N_3316,In_4217,N_2352);
xor U3317 (N_3317,N_2289,N_644);
or U3318 (N_3318,N_2970,In_102);
nor U3319 (N_3319,N_2877,N_2056);
xnor U3320 (N_3320,N_2662,N_2230);
or U3321 (N_3321,N_2234,N_82);
and U3322 (N_3322,N_65,In_3102);
and U3323 (N_3323,N_2591,In_4040);
nor U3324 (N_3324,In_3691,N_2533);
nand U3325 (N_3325,N_2458,N_1673);
nand U3326 (N_3326,N_2009,N_1913);
nor U3327 (N_3327,In_4806,N_2735);
or U3328 (N_3328,In_4001,N_281);
and U3329 (N_3329,N_2285,N_2143);
nor U3330 (N_3330,In_3073,N_1653);
and U3331 (N_3331,In_1069,N_2329);
or U3332 (N_3332,N_2594,In_1431);
nand U3333 (N_3333,N_2370,N_671);
xor U3334 (N_3334,In_1261,N_2976);
or U3335 (N_3335,N_2583,In_4268);
nor U3336 (N_3336,N_2878,N_2262);
or U3337 (N_3337,N_2632,N_2563);
xnor U3338 (N_3338,N_2820,N_1638);
and U3339 (N_3339,N_2987,N_2617);
and U3340 (N_3340,N_961,N_2019);
or U3341 (N_3341,N_1332,N_2139);
nor U3342 (N_3342,N_2424,N_2290);
and U3343 (N_3343,In_4472,N_1629);
xor U3344 (N_3344,N_2292,N_2867);
and U3345 (N_3345,N_1040,N_2566);
and U3346 (N_3346,N_1284,N_2438);
xor U3347 (N_3347,N_965,In_3668);
nand U3348 (N_3348,N_1557,N_144);
xnor U3349 (N_3349,In_1602,N_2412);
or U3350 (N_3350,N_2211,In_1369);
nand U3351 (N_3351,N_2189,N_1735);
or U3352 (N_3352,N_1353,N_2513);
nand U3353 (N_3353,N_2940,In_3775);
nor U3354 (N_3354,N_1633,In_3430);
xnor U3355 (N_3355,N_2001,In_3605);
nand U3356 (N_3356,In_864,N_2270);
xnor U3357 (N_3357,In_3856,N_2530);
nand U3358 (N_3358,N_2032,N_2527);
nor U3359 (N_3359,N_2464,N_2785);
or U3360 (N_3360,In_4114,N_1540);
and U3361 (N_3361,N_1593,N_2657);
and U3362 (N_3362,In_2370,N_2587);
nand U3363 (N_3363,N_457,N_2026);
or U3364 (N_3364,In_2063,N_2604);
xor U3365 (N_3365,N_2130,N_2607);
xnor U3366 (N_3366,In_2868,N_2295);
xnor U3367 (N_3367,In_4877,In_3227);
xor U3368 (N_3368,In_4827,N_2340);
or U3369 (N_3369,N_2627,N_1546);
or U3370 (N_3370,In_2493,N_2541);
nand U3371 (N_3371,N_1882,N_2770);
or U3372 (N_3372,N_1834,In_4561);
nand U3373 (N_3373,N_1627,N_421);
or U3374 (N_3374,N_908,N_2402);
or U3375 (N_3375,N_2674,N_1440);
nand U3376 (N_3376,N_2653,N_2463);
nand U3377 (N_3377,N_2682,N_1051);
xor U3378 (N_3378,N_2000,N_1973);
nand U3379 (N_3379,N_2369,N_121);
nand U3380 (N_3380,N_195,N_62);
or U3381 (N_3381,N_2504,In_2383);
nand U3382 (N_3382,N_1531,N_2712);
nand U3383 (N_3383,N_2201,N_2660);
nand U3384 (N_3384,N_2471,N_848);
and U3385 (N_3385,N_2964,In_4620);
and U3386 (N_3386,N_2219,In_145);
and U3387 (N_3387,N_2025,N_1901);
xnor U3388 (N_3388,N_777,N_2947);
or U3389 (N_3389,N_1117,N_722);
or U3390 (N_3390,N_2119,N_2520);
nand U3391 (N_3391,N_1700,N_1868);
nor U3392 (N_3392,In_3038,In_3438);
nor U3393 (N_3393,N_612,N_2749);
xor U3394 (N_3394,N_1160,In_4927);
or U3395 (N_3395,N_1910,N_2304);
nand U3396 (N_3396,N_2643,N_2543);
nand U3397 (N_3397,In_3971,N_2103);
xnor U3398 (N_3398,In_575,N_2351);
or U3399 (N_3399,N_2398,In_3699);
nor U3400 (N_3400,In_4567,N_2667);
nor U3401 (N_3401,N_1503,In_4552);
nand U3402 (N_3402,N_88,N_2844);
nor U3403 (N_3403,N_2502,In_4299);
or U3404 (N_3404,N_2452,N_1252);
or U3405 (N_3405,N_1124,N_2442);
nand U3406 (N_3406,N_2824,N_1983);
and U3407 (N_3407,N_2932,N_1954);
xor U3408 (N_3408,N_2546,N_2887);
or U3409 (N_3409,In_2786,In_1291);
nand U3410 (N_3410,In_2654,N_217);
or U3411 (N_3411,N_2278,N_2070);
or U3412 (N_3412,N_2373,In_70);
nor U3413 (N_3413,N_1416,N_2739);
or U3414 (N_3414,In_1039,In_1756);
nand U3415 (N_3415,In_4003,N_2724);
and U3416 (N_3416,In_434,N_2180);
and U3417 (N_3417,N_2969,N_1806);
xnor U3418 (N_3418,N_1012,In_4795);
nor U3419 (N_3419,N_1795,N_2006);
or U3420 (N_3420,N_2319,N_2210);
or U3421 (N_3421,N_2592,N_1604);
and U3422 (N_3422,N_2899,N_438);
or U3423 (N_3423,N_2166,In_4588);
and U3424 (N_3424,N_2650,N_2220);
or U3425 (N_3425,N_1641,In_1988);
nor U3426 (N_3426,N_2305,In_551);
nand U3427 (N_3427,N_1034,N_2072);
or U3428 (N_3428,N_190,N_1498);
nor U3429 (N_3429,In_2576,N_2423);
nor U3430 (N_3430,N_844,In_4842);
nand U3431 (N_3431,N_1291,N_2547);
or U3432 (N_3432,N_2613,N_2841);
xnor U3433 (N_3433,N_2866,N_2354);
or U3434 (N_3434,N_2333,N_627);
or U3435 (N_3435,N_1786,N_2028);
nor U3436 (N_3436,N_1396,N_2102);
nor U3437 (N_3437,N_973,N_1590);
xnor U3438 (N_3438,N_2420,In_1977);
nor U3439 (N_3439,N_2933,In_4705);
xnor U3440 (N_3440,N_1336,N_2666);
nor U3441 (N_3441,N_2197,N_2979);
xnor U3442 (N_3442,N_2318,N_1146);
nand U3443 (N_3443,N_2085,N_2198);
nor U3444 (N_3444,In_1008,N_2731);
xor U3445 (N_3445,N_2630,N_2451);
xor U3446 (N_3446,N_2554,N_1830);
nor U3447 (N_3447,N_2764,N_2634);
nor U3448 (N_3448,N_2796,In_1652);
or U3449 (N_3449,N_2733,N_2276);
and U3450 (N_3450,N_1666,N_776);
nand U3451 (N_3451,N_2747,N_1678);
nand U3452 (N_3452,N_2515,N_2024);
and U3453 (N_3453,N_2687,In_1286);
xnor U3454 (N_3454,In_1284,N_2847);
xnor U3455 (N_3455,N_1135,N_2152);
and U3456 (N_3456,N_2086,N_1094);
xor U3457 (N_3457,N_2619,N_2038);
and U3458 (N_3458,N_2725,N_1229);
nor U3459 (N_3459,N_2834,N_2395);
and U3460 (N_3460,In_4821,In_4271);
or U3461 (N_3461,N_1844,In_1249);
or U3462 (N_3462,N_809,In_332);
nand U3463 (N_3463,N_1851,In_1108);
nand U3464 (N_3464,N_2418,N_1078);
xor U3465 (N_3465,N_2714,N_2187);
and U3466 (N_3466,N_1766,N_2901);
xor U3467 (N_3467,In_3279,N_1287);
and U3468 (N_3468,N_1745,In_2121);
xnor U3469 (N_3469,N_1167,N_1839);
nor U3470 (N_3470,N_2590,N_576);
or U3471 (N_3471,In_3475,In_4654);
and U3472 (N_3472,N_2194,N_2435);
nor U3473 (N_3473,N_1719,N_894);
or U3474 (N_3474,N_2511,In_388);
nor U3475 (N_3475,N_2400,N_2793);
and U3476 (N_3476,N_2337,In_987);
nor U3477 (N_3477,In_2986,In_4515);
nand U3478 (N_3478,N_2047,N_2903);
nor U3479 (N_3479,In_456,N_2339);
nand U3480 (N_3480,N_1207,In_532);
nor U3481 (N_3481,N_2380,N_2753);
nand U3482 (N_3482,N_1340,N_2497);
nand U3483 (N_3483,N_1487,N_2027);
nand U3484 (N_3484,N_2720,In_4013);
nor U3485 (N_3485,N_2598,N_2757);
or U3486 (N_3486,In_3628,In_1407);
or U3487 (N_3487,In_1466,N_1110);
nor U3488 (N_3488,N_2496,N_2963);
xnor U3489 (N_3489,In_3488,N_2387);
nor U3490 (N_3490,N_2794,N_574);
or U3491 (N_3491,N_2129,In_34);
xnor U3492 (N_3492,N_1060,N_2429);
xor U3493 (N_3493,N_1280,N_1829);
and U3494 (N_3494,In_3504,In_4373);
nor U3495 (N_3495,N_1743,N_2531);
and U3496 (N_3496,N_2323,N_2088);
xor U3497 (N_3497,N_485,N_1491);
nand U3498 (N_3498,N_845,N_2837);
xnor U3499 (N_3499,N_1307,In_1518);
nand U3500 (N_3500,N_2484,N_1518);
and U3501 (N_3501,N_2935,N_2069);
or U3502 (N_3502,N_2742,N_2849);
or U3503 (N_3503,N_2316,In_156);
nand U3504 (N_3504,N_1572,N_2213);
nor U3505 (N_3505,N_2240,N_2282);
and U3506 (N_3506,N_1714,N_2860);
xnor U3507 (N_3507,N_2936,N_2740);
nor U3508 (N_3508,N_2419,N_2149);
or U3509 (N_3509,In_1828,In_2377);
xor U3510 (N_3510,N_2616,In_633);
and U3511 (N_3511,In_1439,N_2042);
xnor U3512 (N_3512,N_1354,In_3892);
nor U3513 (N_3513,N_2958,N_1210);
xor U3514 (N_3514,In_2669,In_891);
nand U3515 (N_3515,N_2105,In_152);
and U3516 (N_3516,N_2114,N_2512);
xor U3517 (N_3517,In_2337,In_1130);
xor U3518 (N_3518,In_540,N_2248);
nor U3519 (N_3519,N_2274,N_1062);
xor U3520 (N_3520,N_2023,N_2997);
xor U3521 (N_3521,In_54,N_680);
or U3522 (N_3522,In_3242,N_1153);
nand U3523 (N_3523,N_2320,N_2772);
or U3524 (N_3524,N_70,In_1674);
nor U3525 (N_3525,N_1463,N_2051);
or U3526 (N_3526,N_2271,N_2161);
nand U3527 (N_3527,N_2582,N_2904);
and U3528 (N_3528,N_2658,N_2568);
nand U3529 (N_3529,N_1132,N_1243);
nor U3530 (N_3530,N_869,N_1131);
nor U3531 (N_3531,N_2467,In_3085);
xnor U3532 (N_3532,N_2425,In_4269);
xnor U3533 (N_3533,In_4812,N_2410);
xnor U3534 (N_3534,In_4242,N_166);
or U3535 (N_3535,In_641,In_4975);
and U3536 (N_3536,N_2960,N_2328);
xnor U3537 (N_3537,In_3710,N_2018);
xnor U3538 (N_3538,In_363,N_2981);
and U3539 (N_3539,N_2296,N_1216);
nor U3540 (N_3540,N_2364,N_882);
nor U3541 (N_3541,N_2225,N_2228);
nand U3542 (N_3542,N_1228,N_930);
and U3543 (N_3543,N_798,N_2863);
and U3544 (N_3544,In_1997,In_373);
nand U3545 (N_3545,In_3233,N_2550);
nand U3546 (N_3546,N_1654,N_1473);
nor U3547 (N_3547,In_2344,N_2703);
nand U3548 (N_3548,N_2980,In_1479);
and U3549 (N_3549,N_2801,N_2163);
nor U3550 (N_3550,N_2908,In_4603);
and U3551 (N_3551,In_513,N_1309);
xnor U3552 (N_3552,N_1782,In_1987);
xnor U3553 (N_3553,N_2789,N_2609);
nor U3554 (N_3554,N_2706,In_2307);
nor U3555 (N_3555,N_2437,N_2168);
nand U3556 (N_3556,N_1841,N_586);
and U3557 (N_3557,N_169,In_906);
or U3558 (N_3558,N_138,N_2190);
or U3559 (N_3559,In_2261,N_2871);
nor U3560 (N_3560,N_1438,N_1486);
nand U3561 (N_3561,N_2719,N_2651);
xor U3562 (N_3562,In_519,N_161);
or U3563 (N_3563,In_486,N_2455);
and U3564 (N_3564,In_2871,N_2314);
and U3565 (N_3565,N_2578,N_2636);
or U3566 (N_3566,N_2635,N_2445);
xor U3567 (N_3567,N_1257,N_2638);
or U3568 (N_3568,In_2763,In_4124);
nand U3569 (N_3569,N_2810,N_2138);
nand U3570 (N_3570,N_2889,In_2415);
xor U3571 (N_3571,N_2892,N_1476);
and U3572 (N_3572,N_2555,N_1982);
nor U3573 (N_3573,N_2501,N_331);
nand U3574 (N_3574,N_1045,In_2432);
xnor U3575 (N_3575,N_2601,In_190);
xor U3576 (N_3576,N_2489,N_1999);
nand U3577 (N_3577,N_1961,In_3152);
or U3578 (N_3578,N_2443,N_2417);
or U3579 (N_3579,In_640,N_2759);
nor U3580 (N_3580,In_2587,N_1987);
xor U3581 (N_3581,N_2917,N_202);
nor U3582 (N_3582,N_2461,N_2177);
nor U3583 (N_3583,N_2505,In_4940);
or U3584 (N_3584,N_2145,N_2447);
nor U3585 (N_3585,N_2626,N_2155);
and U3586 (N_3586,N_2580,N_1081);
nor U3587 (N_3587,N_1784,N_2648);
nor U3588 (N_3588,N_2612,N_1718);
xor U3589 (N_3589,N_1676,In_1523);
and U3590 (N_3590,N_2553,N_1818);
nor U3591 (N_3591,N_2137,In_3471);
or U3592 (N_3592,N_2902,N_2223);
nand U3593 (N_3593,In_1995,N_2246);
nand U3594 (N_3594,N_2053,N_2893);
or U3595 (N_3595,N_1865,N_2625);
nor U3596 (N_3596,In_418,N_192);
or U3597 (N_3597,N_2476,N_2106);
nor U3598 (N_3598,N_1188,N_2760);
and U3599 (N_3599,N_1223,In_2701);
or U3600 (N_3600,In_4495,N_850);
or U3601 (N_3601,N_2495,N_2913);
nor U3602 (N_3602,N_2945,N_2008);
and U3603 (N_3603,N_2983,N_2952);
nand U3604 (N_3604,N_2710,N_2640);
or U3605 (N_3605,N_1651,N_1433);
and U3606 (N_3606,N_2427,N_2874);
and U3607 (N_3607,N_2991,N_515);
nand U3608 (N_3608,N_1568,N_2950);
xor U3609 (N_3609,N_2961,N_2734);
nand U3610 (N_3610,N_2207,N_2778);
xor U3611 (N_3611,In_4276,N_338);
nand U3612 (N_3612,N_2469,In_2483);
nor U3613 (N_3613,N_2545,N_2054);
and U3614 (N_3614,N_2487,N_2929);
nor U3615 (N_3615,N_2122,N_2909);
and U3616 (N_3616,N_2698,N_2503);
nor U3617 (N_3617,N_988,In_3255);
nor U3618 (N_3618,N_1943,In_4906);
nor U3619 (N_3619,In_182,In_2144);
xnor U3620 (N_3620,N_2029,In_3804);
xor U3621 (N_3621,N_305,In_1248);
xnor U3622 (N_3622,N_1885,N_2279);
nor U3623 (N_3623,N_2057,N_2250);
and U3624 (N_3624,N_2922,N_2315);
nand U3625 (N_3625,N_2494,N_2711);
xor U3626 (N_3626,In_1923,N_1871);
nand U3627 (N_3627,N_2994,N_2221);
and U3628 (N_3628,N_2312,N_2039);
nand U3629 (N_3629,In_292,N_2195);
and U3630 (N_3630,N_2064,In_3065);
or U3631 (N_3631,N_1005,In_2658);
nor U3632 (N_3632,In_340,N_2574);
nor U3633 (N_3633,N_2012,N_2528);
nor U3634 (N_3634,N_1304,N_1602);
and U3635 (N_3635,N_2095,N_1573);
nand U3636 (N_3636,N_2091,N_2637);
nor U3637 (N_3637,N_2301,In_1200);
nor U3638 (N_3638,N_2426,In_1568);
or U3639 (N_3639,N_2737,N_131);
nand U3640 (N_3640,N_2097,N_2718);
and U3641 (N_3641,N_1643,N_2273);
xnor U3642 (N_3642,N_727,N_2255);
nand U3643 (N_3643,N_2537,N_2974);
xor U3644 (N_3644,N_1310,N_2620);
and U3645 (N_3645,In_2021,In_4363);
nor U3646 (N_3646,In_3006,N_2193);
and U3647 (N_3647,N_2854,In_1462);
nor U3648 (N_3648,N_2330,N_1299);
xor U3649 (N_3649,N_2773,In_3796);
or U3650 (N_3650,N_2060,In_2744);
and U3651 (N_3651,In_4274,N_1230);
or U3652 (N_3652,N_797,N_2063);
nor U3653 (N_3653,In_3480,In_4981);
xnor U3654 (N_3654,N_2812,N_2606);
nand U3655 (N_3655,In_4858,N_2389);
and U3656 (N_3656,N_2472,N_1600);
xor U3657 (N_3657,In_1051,N_1522);
and U3658 (N_3658,N_2685,In_2176);
xnor U3659 (N_3659,N_1026,N_1609);
xnor U3660 (N_3660,N_2308,In_874);
or U3661 (N_3661,N_2695,N_1372);
nand U3662 (N_3662,N_2093,N_2205);
nand U3663 (N_3663,N_2647,In_610);
or U3664 (N_3664,N_2283,N_2941);
nor U3665 (N_3665,N_1670,N_2344);
xnor U3666 (N_3666,N_1441,N_2534);
and U3667 (N_3667,N_2265,N_49);
nand U3668 (N_3668,N_2577,N_2430);
xor U3669 (N_3669,N_2529,N_2259);
xor U3670 (N_3670,N_2011,N_2264);
and U3671 (N_3671,N_2656,N_2486);
nor U3672 (N_3672,N_2368,In_1426);
or U3673 (N_3673,N_2575,N_1550);
or U3674 (N_3674,N_2665,N_1649);
nand U3675 (N_3675,N_2392,N_1312);
or U3676 (N_3676,N_951,In_2561);
xnor U3677 (N_3677,In_1770,N_2459);
and U3678 (N_3678,In_4548,N_555);
nand U3679 (N_3679,N_491,In_4702);
or U3680 (N_3680,In_4872,In_3268);
xor U3681 (N_3681,In_1839,N_2869);
xor U3682 (N_3682,N_2121,N_2825);
or U3683 (N_3683,In_3107,N_1724);
xor U3684 (N_3684,N_2460,In_4914);
nor U3685 (N_3685,In_3027,In_4199);
nand U3686 (N_3686,N_2795,N_2082);
nand U3687 (N_3687,In_4361,N_2927);
xor U3688 (N_3688,N_287,In_2348);
or U3689 (N_3689,In_2328,N_2943);
nor U3690 (N_3690,In_2665,N_2522);
or U3691 (N_3691,In_1607,In_4190);
or U3692 (N_3692,In_1862,In_4174);
and U3693 (N_3693,In_3363,N_1785);
nor U3694 (N_3694,N_1397,In_2840);
nand U3695 (N_3695,In_2311,In_2852);
and U3696 (N_3696,N_25,N_2302);
or U3697 (N_3697,N_2517,In_992);
xor U3698 (N_3698,N_2924,N_2715);
xor U3699 (N_3699,N_2723,N_2071);
or U3700 (N_3700,In_3041,In_865);
nand U3701 (N_3701,In_2566,N_2589);
and U3702 (N_3702,N_2754,N_403);
nor U3703 (N_3703,N_1155,N_2649);
nor U3704 (N_3704,N_2802,N_276);
nand U3705 (N_3705,In_3432,N_2257);
and U3706 (N_3706,N_2267,N_2897);
xor U3707 (N_3707,N_2518,N_2127);
nand U3708 (N_3708,In_4444,In_1066);
xor U3709 (N_3709,N_2346,N_1692);
or U3710 (N_3710,In_1058,N_44);
or U3711 (N_3711,N_2157,N_2048);
and U3712 (N_3712,N_1896,N_2390);
or U3713 (N_3713,N_1301,In_2410);
nand U3714 (N_3714,N_1608,N_2167);
xnor U3715 (N_3715,N_1199,In_3238);
xnor U3716 (N_3716,N_2679,N_1359);
nand U3717 (N_3717,N_2002,In_4882);
xor U3718 (N_3718,N_2491,N_2332);
xnor U3719 (N_3719,N_1512,In_3872);
and U3720 (N_3720,In_1328,N_2975);
or U3721 (N_3721,N_868,N_2077);
and U3722 (N_3722,N_2245,N_2101);
xor U3723 (N_3723,N_2763,N_1266);
xnor U3724 (N_3724,N_122,N_2954);
and U3725 (N_3725,N_2396,N_2807);
nor U3726 (N_3726,N_2123,In_4627);
nand U3727 (N_3727,N_2192,N_2851);
nor U3728 (N_3728,N_2669,In_734);
or U3729 (N_3729,N_1253,N_2858);
or U3730 (N_3730,In_2602,N_2075);
nand U3731 (N_3731,In_2638,N_2440);
or U3732 (N_3732,N_2074,N_922);
or U3733 (N_3733,In_1182,N_2084);
nor U3734 (N_3734,N_839,N_239);
xor U3735 (N_3735,N_2768,N_2745);
nor U3736 (N_3736,N_2453,N_2828);
nor U3737 (N_3737,In_346,N_2040);
nand U3738 (N_3738,N_2052,N_2120);
nand U3739 (N_3739,In_4314,In_1223);
or U3740 (N_3740,In_1401,N_2013);
nand U3741 (N_3741,N_2835,In_785);
nand U3742 (N_3742,N_2538,N_2165);
nor U3743 (N_3743,In_3985,N_2439);
or U3744 (N_3744,N_2689,In_4);
and U3745 (N_3745,N_2485,N_567);
nor U3746 (N_3746,N_2857,N_2664);
nor U3747 (N_3747,N_2422,N_1642);
xor U3748 (N_3748,N_1988,In_1784);
and U3749 (N_3749,N_2411,N_430);
xor U3750 (N_3750,In_135,N_1923);
nor U3751 (N_3751,N_2562,N_2610);
nand U3752 (N_3752,N_2045,N_2222);
xor U3753 (N_3753,N_1014,In_2331);
xor U3754 (N_3754,N_1924,N_2989);
nand U3755 (N_3755,N_2224,In_1078);
nor U3756 (N_3756,In_3406,In_2791);
and U3757 (N_3757,N_910,N_1513);
xnor U3758 (N_3758,N_1151,N_1533);
nor U3759 (N_3759,N_2558,N_1695);
nor U3760 (N_3760,N_2393,N_2272);
nand U3761 (N_3761,In_4203,N_2915);
and U3762 (N_3762,N_2043,N_2790);
nand U3763 (N_3763,N_385,In_2379);
xor U3764 (N_3764,N_2343,N_2394);
xor U3765 (N_3765,N_1613,N_2140);
nand U3766 (N_3766,In_2088,N_1065);
xnor U3767 (N_3767,N_1707,N_2200);
xor U3768 (N_3768,In_743,N_2311);
or U3769 (N_3769,N_1236,N_20);
or U3770 (N_3770,N_2567,In_1874);
and U3771 (N_3771,N_2239,In_531);
or U3772 (N_3772,In_3861,N_2287);
nand U3773 (N_3773,N_2022,N_945);
nand U3774 (N_3774,N_1717,N_2124);
xnor U3775 (N_3775,In_4250,N_2805);
xor U3776 (N_3776,N_2564,In_3072);
and U3777 (N_3777,In_3862,N_2281);
nand U3778 (N_3778,N_530,N_2465);
and U3779 (N_3779,In_1718,N_1274);
or U3780 (N_3780,N_2998,N_918);
and U3781 (N_3781,N_2891,N_2646);
or U3782 (N_3782,N_2154,N_2599);
xor U3783 (N_3783,N_569,N_2100);
xor U3784 (N_3784,N_2150,N_1594);
nor U3785 (N_3785,In_2899,N_836);
xor U3786 (N_3786,N_2992,N_2041);
or U3787 (N_3787,N_2109,In_2728);
or U3788 (N_3788,N_1129,N_1838);
and U3789 (N_3789,N_2062,N_2683);
nor U3790 (N_3790,N_2372,N_1134);
or U3791 (N_3791,N_2848,N_2572);
or U3792 (N_3792,In_4216,N_2475);
and U3793 (N_3793,N_2573,In_2865);
nor U3794 (N_3794,N_2588,N_1145);
nor U3795 (N_3795,In_3486,N_2819);
xor U3796 (N_3796,N_1450,In_1788);
and U3797 (N_3797,N_2982,In_3936);
xnor U3798 (N_3798,N_2407,N_500);
xnor U3799 (N_3799,N_2299,N_2621);
nand U3800 (N_3800,In_3273,N_2560);
or U3801 (N_3801,In_3386,N_2298);
and U3802 (N_3802,N_2050,N_2436);
or U3803 (N_3803,N_2334,In_2023);
nand U3804 (N_3804,N_2951,N_1420);
nor U3805 (N_3805,In_983,N_654);
xnor U3806 (N_3806,In_1745,N_1008);
nand U3807 (N_3807,In_4816,N_2921);
or U3808 (N_3808,In_2822,In_3100);
xnor U3809 (N_3809,N_1744,In_479);
nor U3810 (N_3810,In_2512,In_2265);
nor U3811 (N_3811,N_2864,N_1935);
xnor U3812 (N_3812,N_2855,N_1694);
nor U3813 (N_3813,N_2559,In_2367);
xnor U3814 (N_3814,In_2670,N_1612);
xnor U3815 (N_3815,N_2671,N_2399);
xor U3816 (N_3816,N_1409,N_1630);
or U3817 (N_3817,N_1993,N_2081);
and U3818 (N_3818,In_118,N_2492);
or U3819 (N_3819,N_2183,In_1186);
nor U3820 (N_3820,In_3663,N_1881);
or U3821 (N_3821,N_2397,In_558);
nand U3822 (N_3822,N_2499,N_2241);
nand U3823 (N_3823,In_1781,In_2709);
nor U3824 (N_3824,N_2448,N_1775);
nand U3825 (N_3825,In_4789,In_1772);
xnor U3826 (N_3826,N_2758,In_3999);
or U3827 (N_3827,In_1067,N_1787);
nor U3828 (N_3828,N_2585,In_1994);
nor U3829 (N_3829,In_1177,N_2083);
and U3830 (N_3830,In_4005,N_750);
and U3831 (N_3831,N_2172,N_2358);
nand U3832 (N_3832,N_2827,N_2888);
xor U3833 (N_3833,N_1479,N_2089);
nand U3834 (N_3834,In_3446,N_2673);
nand U3835 (N_3835,N_428,In_3262);
nand U3836 (N_3836,N_2174,In_929);
nor U3837 (N_3837,N_851,In_573);
nand U3838 (N_3838,N_2668,N_2540);
nand U3839 (N_3839,N_2232,N_887);
nand U3840 (N_3840,In_3066,N_2552);
and U3841 (N_3841,N_2433,N_2614);
nand U3842 (N_3842,In_2954,In_3029);
xnor U3843 (N_3843,N_1058,In_1990);
nand U3844 (N_3844,N_2732,N_2633);
nand U3845 (N_3845,N_595,N_461);
nor U3846 (N_3846,N_1535,In_2353);
and U3847 (N_3847,N_978,N_1126);
and U3848 (N_3848,N_2386,N_2349);
nor U3849 (N_3849,N_1022,N_2256);
and U3850 (N_3850,In_1616,N_2132);
and U3851 (N_3851,N_2966,In_511);
nor U3852 (N_3852,N_374,N_1659);
xor U3853 (N_3853,N_2325,N_2035);
nand U3854 (N_3854,In_4658,N_938);
xor U3855 (N_3855,In_794,N_2744);
nand U3856 (N_3856,In_2082,N_2481);
or U3857 (N_3857,N_2449,N_1671);
and U3858 (N_3858,N_2542,In_2384);
or U3859 (N_3859,N_2775,N_1680);
nand U3860 (N_3860,N_1489,N_2707);
nor U3861 (N_3861,In_4048,N_856);
nor U3862 (N_3862,In_4503,N_2136);
and U3863 (N_3863,In_3913,N_2284);
nand U3864 (N_3864,N_2756,N_2856);
and U3865 (N_3865,N_1088,N_1156);
or U3866 (N_3866,N_2843,N_2500);
nor U3867 (N_3867,In_2469,In_308);
or U3868 (N_3868,In_1835,In_2800);
nand U3869 (N_3869,In_2697,N_2804);
and U3870 (N_3870,N_620,N_2317);
nand U3871 (N_3871,N_2117,N_2788);
and U3872 (N_3872,N_2595,N_523);
and U3873 (N_3873,N_196,N_210);
and U3874 (N_3874,In_378,N_2046);
nor U3875 (N_3875,N_2367,N_2067);
or U3876 (N_3876,In_3349,N_1095);
xor U3877 (N_3877,In_33,N_306);
or U3878 (N_3878,N_2010,In_4149);
and U3879 (N_3879,N_2249,N_2840);
or U3880 (N_3880,In_2876,N_712);
nor U3881 (N_3881,N_1494,In_2858);
xnor U3882 (N_3882,N_2376,N_2142);
nor U3883 (N_3883,In_3509,N_2600);
or U3884 (N_3884,N_2631,N_1819);
nand U3885 (N_3885,N_2690,N_1802);
nand U3886 (N_3886,In_3281,N_2016);
xnor U3887 (N_3887,In_3525,In_4017);
and U3888 (N_3888,In_3669,N_2727);
nor U3889 (N_3889,N_2684,N_2693);
xnor U3890 (N_3890,N_2928,N_2300);
and U3891 (N_3891,N_2247,N_2675);
nor U3892 (N_3892,N_2217,N_772);
and U3893 (N_3893,N_2233,In_2252);
nor U3894 (N_3894,N_2962,In_2106);
and U3895 (N_3895,N_2972,In_3304);
or U3896 (N_3896,In_806,N_2336);
or U3897 (N_3897,N_1796,In_3306);
or U3898 (N_3898,N_2286,N_944);
and U3899 (N_3899,N_2615,N_2948);
nand U3900 (N_3900,N_2428,N_2783);
nor U3901 (N_3901,In_1115,N_2375);
and U3902 (N_3902,In_3528,N_1853);
or U3903 (N_3903,N_2771,N_2509);
nand U3904 (N_3904,N_2269,N_1824);
nor U3905 (N_3905,In_2169,N_1205);
nand U3906 (N_3906,N_2431,N_357);
nor U3907 (N_3907,In_3401,N_2186);
nor U3908 (N_3908,N_2524,N_2260);
nand U3909 (N_3909,In_609,N_2890);
nor U3910 (N_3910,N_2818,N_2033);
or U3911 (N_3911,N_2934,N_46);
or U3912 (N_3912,N_2761,In_1444);
xor U3913 (N_3913,N_2112,N_2526);
and U3914 (N_3914,In_4736,N_2413);
xnor U3915 (N_3915,N_1587,N_1133);
and U3916 (N_3916,In_3625,N_2401);
or U3917 (N_3917,N_2791,N_2261);
nor U3918 (N_3918,In_4862,N_2164);
or U3919 (N_3919,N_2655,N_538);
and U3920 (N_3920,N_2003,In_1352);
nand U3921 (N_3921,N_2873,N_2907);
or U3922 (N_3922,N_2688,N_1103);
or U3923 (N_3923,N_2988,N_1980);
and U3924 (N_3924,N_2307,In_3941);
and U3925 (N_3925,N_1893,N_1403);
and U3926 (N_3926,In_3017,N_2253);
xor U3927 (N_3927,N_2466,In_3254);
and U3928 (N_3928,N_2115,N_1334);
or U3929 (N_3929,In_3754,In_4659);
nand U3930 (N_3930,N_2263,In_2938);
xor U3931 (N_3931,N_532,In_4249);
or U3932 (N_3932,N_2441,N_2381);
and U3933 (N_3933,N_1477,N_2477);
xnor U3934 (N_3934,N_2809,N_95);
xnor U3935 (N_3935,N_2479,N_1054);
nor U3936 (N_3936,N_2434,N_2814);
nor U3937 (N_3937,N_2872,N_205);
nor U3938 (N_3938,In_2673,N_2885);
nand U3939 (N_3939,N_2216,In_741);
nand U3940 (N_3940,N_1877,N_2356);
and U3941 (N_3941,N_991,N_1624);
xor U3942 (N_3942,N_42,N_1798);
nor U3943 (N_3943,N_1758,N_1180);
and U3944 (N_3944,In_3287,N_2415);
nor U3945 (N_3945,In_2500,N_2498);
nand U3946 (N_3946,N_1130,N_2378);
xnor U3947 (N_3947,N_2920,N_2058);
and U3948 (N_3948,N_1319,In_3088);
and U3949 (N_3949,N_2797,N_2483);
or U3950 (N_3950,N_2678,In_4435);
or U3951 (N_3951,N_337,N_1623);
and U3952 (N_3952,N_2846,N_2702);
and U3953 (N_3953,In_4279,In_154);
or U3954 (N_3954,N_2730,N_2421);
and U3955 (N_3955,In_2288,N_2405);
and U3956 (N_3956,N_789,In_2208);
or U3957 (N_3957,N_243,N_561);
nand U3958 (N_3958,N_2321,N_2779);
and U3959 (N_3959,N_1592,In_2305);
and U3960 (N_3960,In_2820,In_4159);
nand U3961 (N_3961,N_112,In_4169);
or U3962 (N_3962,In_4349,N_2570);
xnor U3963 (N_3963,In_82,In_1529);
nor U3964 (N_3964,N_2266,In_1901);
and U3965 (N_3965,N_2743,N_2670);
or U3966 (N_3966,N_1064,N_1803);
xor U3967 (N_3967,N_2098,N_1181);
nor U3968 (N_3968,N_2078,N_2204);
nor U3969 (N_3969,N_1175,N_2363);
or U3970 (N_3970,N_2652,N_1944);
nor U3971 (N_3971,In_3684,N_1698);
nand U3972 (N_3972,N_1948,In_3601);
nor U3973 (N_3973,In_1359,N_2383);
xnor U3974 (N_3974,N_2708,N_2080);
or U3975 (N_3975,In_4543,N_1368);
or U3976 (N_3976,N_2549,N_1702);
xnor U3977 (N_3977,N_892,N_2535);
or U3978 (N_3978,N_1038,N_2388);
nor U3979 (N_3979,N_2175,N_2808);
and U3980 (N_3980,In_2835,N_2446);
or U3981 (N_3981,In_3336,N_2618);
and U3982 (N_3982,N_2823,N_1313);
or U3983 (N_3983,N_2639,N_2842);
xor U3984 (N_3984,N_2104,N_2699);
or U3985 (N_3985,N_2338,In_4394);
xor U3986 (N_3986,N_2147,N_1545);
xor U3987 (N_3987,N_692,N_2722);
xor U3988 (N_3988,N_2586,N_328);
xor U3989 (N_3989,N_1577,In_4220);
or U3990 (N_3990,N_1832,In_4715);
nand U3991 (N_3991,N_2218,N_1793);
nand U3992 (N_3992,In_1963,N_2516);
and U3993 (N_3993,In_3703,N_2882);
nor U3994 (N_3994,N_2700,N_2780);
or U3995 (N_3995,N_1020,In_3243);
and U3996 (N_3996,N_2822,N_1833);
or U3997 (N_3997,N_2911,In_1033);
nand U3998 (N_3998,N_2159,N_392);
nand U3999 (N_3999,In_2036,N_2005);
nand U4000 (N_4000,N_3479,N_3769);
nor U4001 (N_4001,N_3786,N_3173);
nor U4002 (N_4002,N_3324,N_3216);
nand U4003 (N_4003,N_3808,N_3162);
nor U4004 (N_4004,N_3567,N_3950);
nand U4005 (N_4005,N_3291,N_3500);
xnor U4006 (N_4006,N_3093,N_3636);
xor U4007 (N_4007,N_3067,N_3775);
nor U4008 (N_4008,N_3704,N_3174);
or U4009 (N_4009,N_3123,N_3319);
nor U4010 (N_4010,N_3825,N_3459);
or U4011 (N_4011,N_3360,N_3321);
and U4012 (N_4012,N_3794,N_3272);
and U4013 (N_4013,N_3647,N_3311);
xnor U4014 (N_4014,N_3768,N_3401);
and U4015 (N_4015,N_3962,N_3638);
and U4016 (N_4016,N_3664,N_3457);
nor U4017 (N_4017,N_3629,N_3493);
nand U4018 (N_4018,N_3005,N_3804);
or U4019 (N_4019,N_3037,N_3721);
or U4020 (N_4020,N_3663,N_3908);
and U4021 (N_4021,N_3259,N_3778);
xor U4022 (N_4022,N_3016,N_3247);
nor U4023 (N_4023,N_3284,N_3235);
and U4024 (N_4024,N_3084,N_3336);
or U4025 (N_4025,N_3572,N_3119);
xnor U4026 (N_4026,N_3575,N_3211);
or U4027 (N_4027,N_3810,N_3449);
nand U4028 (N_4028,N_3683,N_3850);
or U4029 (N_4029,N_3275,N_3024);
nand U4030 (N_4030,N_3831,N_3858);
nor U4031 (N_4031,N_3818,N_3377);
and U4032 (N_4032,N_3608,N_3928);
nor U4033 (N_4033,N_3489,N_3674);
and U4034 (N_4034,N_3602,N_3759);
or U4035 (N_4035,N_3732,N_3548);
or U4036 (N_4036,N_3588,N_3849);
nand U4037 (N_4037,N_3237,N_3913);
or U4038 (N_4038,N_3670,N_3862);
nand U4039 (N_4039,N_3814,N_3028);
xor U4040 (N_4040,N_3957,N_3737);
and U4041 (N_4041,N_3731,N_3342);
and U4042 (N_4042,N_3081,N_3780);
nand U4043 (N_4043,N_3581,N_3551);
xor U4044 (N_4044,N_3085,N_3458);
or U4045 (N_4045,N_3148,N_3512);
xnor U4046 (N_4046,N_3365,N_3313);
or U4047 (N_4047,N_3337,N_3533);
and U4048 (N_4048,N_3203,N_3022);
nor U4049 (N_4049,N_3919,N_3982);
nor U4050 (N_4050,N_3451,N_3792);
and U4051 (N_4051,N_3529,N_3442);
or U4052 (N_4052,N_3215,N_3745);
xor U4053 (N_4053,N_3589,N_3438);
xor U4054 (N_4054,N_3556,N_3104);
xor U4055 (N_4055,N_3565,N_3899);
or U4056 (N_4056,N_3357,N_3115);
or U4057 (N_4057,N_3487,N_3332);
and U4058 (N_4058,N_3640,N_3349);
nor U4059 (N_4059,N_3511,N_3419);
nor U4060 (N_4060,N_3662,N_3325);
nand U4061 (N_4061,N_3273,N_3008);
xnor U4062 (N_4062,N_3131,N_3201);
nand U4063 (N_4063,N_3117,N_3777);
nor U4064 (N_4064,N_3530,N_3111);
nor U4065 (N_4065,N_3723,N_3931);
or U4066 (N_4066,N_3010,N_3498);
and U4067 (N_4067,N_3783,N_3985);
or U4068 (N_4068,N_3169,N_3813);
xnor U4069 (N_4069,N_3524,N_3754);
nor U4070 (N_4070,N_3803,N_3582);
or U4071 (N_4071,N_3776,N_3748);
nor U4072 (N_4072,N_3616,N_3964);
and U4073 (N_4073,N_3716,N_3279);
xor U4074 (N_4074,N_3323,N_3209);
or U4075 (N_4075,N_3452,N_3920);
xnor U4076 (N_4076,N_3274,N_3376);
nand U4077 (N_4077,N_3897,N_3064);
nor U4078 (N_4078,N_3988,N_3916);
nor U4079 (N_4079,N_3242,N_3822);
or U4080 (N_4080,N_3651,N_3128);
and U4081 (N_4081,N_3220,N_3422);
and U4082 (N_4082,N_3281,N_3735);
or U4083 (N_4083,N_3027,N_3513);
and U4084 (N_4084,N_3655,N_3143);
nand U4085 (N_4085,N_3806,N_3091);
nor U4086 (N_4086,N_3253,N_3348);
and U4087 (N_4087,N_3222,N_3437);
xnor U4088 (N_4088,N_3309,N_3439);
nand U4089 (N_4089,N_3627,N_3074);
xnor U4090 (N_4090,N_3878,N_3961);
or U4091 (N_4091,N_3755,N_3947);
nand U4092 (N_4092,N_3254,N_3331);
or U4093 (N_4093,N_3155,N_3066);
xor U4094 (N_4094,N_3076,N_3391);
xor U4095 (N_4095,N_3416,N_3300);
or U4096 (N_4096,N_3503,N_3884);
nand U4097 (N_4097,N_3047,N_3502);
and U4098 (N_4098,N_3694,N_3466);
nand U4099 (N_4099,N_3105,N_3743);
and U4100 (N_4100,N_3612,N_3264);
or U4101 (N_4101,N_3396,N_3531);
xor U4102 (N_4102,N_3346,N_3573);
xnor U4103 (N_4103,N_3139,N_3369);
nor U4104 (N_4104,N_3527,N_3427);
nor U4105 (N_4105,N_3007,N_3987);
xnor U4106 (N_4106,N_3374,N_3764);
and U4107 (N_4107,N_3303,N_3089);
xnor U4108 (N_4108,N_3102,N_3477);
nor U4109 (N_4109,N_3017,N_3326);
and U4110 (N_4110,N_3137,N_3302);
nand U4111 (N_4111,N_3939,N_3127);
nand U4112 (N_4112,N_3577,N_3560);
or U4113 (N_4113,N_3000,N_3989);
and U4114 (N_4114,N_3191,N_3960);
and U4115 (N_4115,N_3568,N_3952);
nor U4116 (N_4116,N_3366,N_3249);
or U4117 (N_4117,N_3358,N_3684);
nor U4118 (N_4118,N_3620,N_3590);
and U4119 (N_4119,N_3494,N_3842);
and U4120 (N_4120,N_3317,N_3853);
xor U4121 (N_4121,N_3854,N_3070);
or U4122 (N_4122,N_3465,N_3993);
or U4123 (N_4123,N_3713,N_3157);
xor U4124 (N_4124,N_3368,N_3834);
and U4125 (N_4125,N_3221,N_3001);
nand U4126 (N_4126,N_3386,N_3545);
xor U4127 (N_4127,N_3048,N_3659);
or U4128 (N_4128,N_3763,N_3671);
or U4129 (N_4129,N_3888,N_3866);
or U4130 (N_4130,N_3844,N_3189);
or U4131 (N_4131,N_3447,N_3969);
nor U4132 (N_4132,N_3845,N_3030);
or U4133 (N_4133,N_3676,N_3370);
nand U4134 (N_4134,N_3911,N_3433);
nor U4135 (N_4135,N_3474,N_3891);
nor U4136 (N_4136,N_3399,N_3648);
or U4137 (N_4137,N_3823,N_3009);
and U4138 (N_4138,N_3518,N_3885);
xor U4139 (N_4139,N_3910,N_3921);
and U4140 (N_4140,N_3902,N_3553);
or U4141 (N_4141,N_3956,N_3226);
nor U4142 (N_4142,N_3877,N_3395);
xnor U4143 (N_4143,N_3562,N_3953);
nor U4144 (N_4144,N_3795,N_3923);
xor U4145 (N_4145,N_3506,N_3967);
and U4146 (N_4146,N_3815,N_3948);
and U4147 (N_4147,N_3637,N_3519);
xor U4148 (N_4148,N_3618,N_3793);
nor U4149 (N_4149,N_3043,N_3855);
and U4150 (N_4150,N_3132,N_3029);
nor U4151 (N_4151,N_3287,N_3430);
nor U4152 (N_4152,N_3686,N_3238);
nor U4153 (N_4153,N_3765,N_3943);
nor U4154 (N_4154,N_3178,N_3955);
and U4155 (N_4155,N_3444,N_3271);
and U4156 (N_4156,N_3784,N_3478);
and U4157 (N_4157,N_3860,N_3975);
and U4158 (N_4158,N_3431,N_3425);
and U4159 (N_4159,N_3999,N_3796);
xor U4160 (N_4160,N_3270,N_3603);
xnor U4161 (N_4161,N_3062,N_3224);
nand U4162 (N_4162,N_3516,N_3470);
nor U4163 (N_4163,N_3187,N_3023);
or U4164 (N_4164,N_3100,N_3693);
nor U4165 (N_4165,N_3387,N_3817);
nor U4166 (N_4166,N_3420,N_3078);
xnor U4167 (N_4167,N_3320,N_3382);
xnor U4168 (N_4168,N_3175,N_3669);
or U4169 (N_4169,N_3484,N_3625);
nand U4170 (N_4170,N_3918,N_3690);
xnor U4171 (N_4171,N_3994,N_3383);
nor U4172 (N_4172,N_3464,N_3381);
xor U4173 (N_4173,N_3068,N_3244);
xnor U4174 (N_4174,N_3171,N_3836);
and U4175 (N_4175,N_3140,N_3103);
xnor U4176 (N_4176,N_3549,N_3504);
nor U4177 (N_4177,N_3257,N_3747);
and U4178 (N_4178,N_3838,N_3014);
or U4179 (N_4179,N_3329,N_3473);
and U4180 (N_4180,N_3712,N_3557);
nor U4181 (N_4181,N_3979,N_3894);
xnor U4182 (N_4182,N_3547,N_3392);
or U4183 (N_4183,N_3801,N_3604);
and U4184 (N_4184,N_3497,N_3176);
and U4185 (N_4185,N_3371,N_3056);
or U4186 (N_4186,N_3893,N_3065);
and U4187 (N_4187,N_3012,N_3402);
nor U4188 (N_4188,N_3871,N_3697);
xor U4189 (N_4189,N_3340,N_3650);
xor U4190 (N_4190,N_3632,N_3297);
nand U4191 (N_4191,N_3197,N_3865);
nor U4192 (N_4192,N_3060,N_3592);
or U4193 (N_4193,N_3058,N_3811);
nand U4194 (N_4194,N_3821,N_3248);
nor U4195 (N_4195,N_3886,N_3977);
xor U4196 (N_4196,N_3744,N_3408);
xnor U4197 (N_4197,N_3196,N_3681);
and U4198 (N_4198,N_3398,N_3312);
or U4199 (N_4199,N_3002,N_3296);
nand U4200 (N_4200,N_3614,N_3841);
nand U4201 (N_4201,N_3976,N_3901);
xor U4202 (N_4202,N_3996,N_3316);
xnor U4203 (N_4203,N_3193,N_3350);
nand U4204 (N_4204,N_3772,N_3734);
nor U4205 (N_4205,N_3574,N_3424);
nand U4206 (N_4206,N_3586,N_3071);
nand U4207 (N_4207,N_3134,N_3032);
nand U4208 (N_4208,N_3468,N_3345);
or U4209 (N_4209,N_3940,N_3631);
nand U4210 (N_4210,N_3829,N_3040);
and U4211 (N_4211,N_3812,N_3781);
or U4212 (N_4212,N_3266,N_3053);
and U4213 (N_4213,N_3657,N_3179);
xnor U4214 (N_4214,N_3426,N_3252);
nor U4215 (N_4215,N_3613,N_3034);
nor U4216 (N_4216,N_3429,N_3159);
xnor U4217 (N_4217,N_3990,N_3546);
nor U4218 (N_4218,N_3643,N_3958);
or U4219 (N_4219,N_3409,N_3846);
xor U4220 (N_4220,N_3537,N_3243);
xnor U4221 (N_4221,N_3073,N_3021);
nor U4222 (N_4222,N_3630,N_3403);
nor U4223 (N_4223,N_3144,N_3523);
xnor U4224 (N_4224,N_3949,N_3766);
and U4225 (N_4225,N_3944,N_3660);
and U4226 (N_4226,N_3268,N_3917);
nor U4227 (N_4227,N_3805,N_3550);
xor U4228 (N_4228,N_3185,N_3749);
xnor U4229 (N_4229,N_3757,N_3057);
xnor U4230 (N_4230,N_3970,N_3767);
xnor U4231 (N_4231,N_3199,N_3959);
nand U4232 (N_4232,N_3857,N_3455);
and U4233 (N_4233,N_3339,N_3079);
xor U4234 (N_4234,N_3699,N_3276);
or U4235 (N_4235,N_3868,N_3318);
xor U4236 (N_4236,N_3026,N_3265);
nand U4237 (N_4237,N_3267,N_3039);
or U4238 (N_4238,N_3698,N_3789);
xnor U4239 (N_4239,N_3033,N_3837);
nand U4240 (N_4240,N_3843,N_3475);
or U4241 (N_4241,N_3869,N_3397);
nand U4242 (N_4242,N_3384,N_3307);
or U4243 (N_4243,N_3232,N_3156);
nand U4244 (N_4244,N_3328,N_3063);
nand U4245 (N_4245,N_3535,N_3004);
nand U4246 (N_4246,N_3106,N_3668);
nand U4247 (N_4247,N_3750,N_3285);
nor U4248 (N_4248,N_3025,N_3986);
and U4249 (N_4249,N_3968,N_3110);
xor U4250 (N_4250,N_3367,N_3052);
nor U4251 (N_4251,N_3709,N_3710);
and U4252 (N_4252,N_3622,N_3725);
or U4253 (N_4253,N_3832,N_3875);
and U4254 (N_4254,N_3770,N_3413);
xor U4255 (N_4255,N_3042,N_3239);
nor U4256 (N_4256,N_3405,N_3649);
xnor U4257 (N_4257,N_3501,N_3212);
or U4258 (N_4258,N_3330,N_3347);
nor U4259 (N_4259,N_3544,N_3003);
and U4260 (N_4260,N_3483,N_3564);
and U4261 (N_4261,N_3467,N_3802);
or U4262 (N_4262,N_3116,N_3540);
or U4263 (N_4263,N_3998,N_3543);
or U4264 (N_4264,N_3966,N_3675);
or U4265 (N_4265,N_3055,N_3163);
nor U4266 (N_4266,N_3788,N_3210);
xnor U4267 (N_4267,N_3705,N_3020);
or U4268 (N_4268,N_3509,N_3870);
nor U4269 (N_4269,N_3359,N_3799);
nor U4270 (N_4270,N_3656,N_3180);
nor U4271 (N_4271,N_3739,N_3161);
or U4272 (N_4272,N_3751,N_3092);
nor U4273 (N_4273,N_3114,N_3299);
nor U4274 (N_4274,N_3454,N_3703);
and U4275 (N_4275,N_3372,N_3536);
nand U4276 (N_4276,N_3354,N_3691);
nand U4277 (N_4277,N_3192,N_3972);
or U4278 (N_4278,N_3135,N_3482);
and U4279 (N_4279,N_3086,N_3121);
nand U4280 (N_4280,N_3375,N_3492);
or U4281 (N_4281,N_3202,N_3214);
nor U4282 (N_4282,N_3490,N_3661);
nand U4283 (N_4283,N_3819,N_3905);
or U4284 (N_4284,N_3771,N_3720);
nor U4285 (N_4285,N_3672,N_3130);
xnor U4286 (N_4286,N_3715,N_3665);
nand U4287 (N_4287,N_3292,N_3652);
or U4288 (N_4288,N_3898,N_3120);
xnor U4289 (N_4289,N_3400,N_3282);
nand U4290 (N_4290,N_3892,N_3122);
and U4291 (N_4291,N_3621,N_3798);
or U4292 (N_4292,N_3390,N_3234);
nor U4293 (N_4293,N_3532,N_3246);
nor U4294 (N_4294,N_3418,N_3283);
or U4295 (N_4295,N_3142,N_3099);
xnor U4296 (N_4296,N_3044,N_3785);
nand U4297 (N_4297,N_3054,N_3436);
xnor U4298 (N_4298,N_3059,N_3797);
nand U4299 (N_4299,N_3515,N_3118);
nor U4300 (N_4300,N_3194,N_3230);
nor U4301 (N_4301,N_3667,N_3486);
xnor U4302 (N_4302,N_3445,N_3205);
or U4303 (N_4303,N_3847,N_3356);
nor U4304 (N_4304,N_3035,N_3840);
and U4305 (N_4305,N_3554,N_3983);
and U4306 (N_4306,N_3889,N_3411);
nor U4307 (N_4307,N_3415,N_3166);
and U4308 (N_4308,N_3929,N_3733);
and U4309 (N_4309,N_3261,N_3521);
nor U4310 (N_4310,N_3149,N_3742);
xor U4311 (N_4311,N_3634,N_3154);
nor U4312 (N_4312,N_3423,N_3965);
nor U4313 (N_4313,N_3606,N_3177);
or U4314 (N_4314,N_3774,N_3096);
nand U4315 (N_4315,N_3779,N_3200);
nor U4316 (N_4316,N_3217,N_3666);
or U4317 (N_4317,N_3295,N_3938);
nand U4318 (N_4318,N_3343,N_3941);
nor U4319 (N_4319,N_3679,N_3628);
or U4320 (N_4320,N_3633,N_3380);
or U4321 (N_4321,N_3700,N_3088);
and U4322 (N_4322,N_3787,N_3204);
or U4323 (N_4323,N_3236,N_3167);
xnor U4324 (N_4324,N_3126,N_3213);
or U4325 (N_4325,N_3828,N_3900);
nor U4326 (N_4326,N_3926,N_3315);
nand U4327 (N_4327,N_3355,N_3584);
xor U4328 (N_4328,N_3288,N_3927);
or U4329 (N_4329,N_3914,N_3930);
nand U4330 (N_4330,N_3496,N_3555);
nand U4331 (N_4331,N_3946,N_3434);
nand U4332 (N_4332,N_3251,N_3839);
and U4333 (N_4333,N_3587,N_3394);
xor U4334 (N_4334,N_3514,N_3463);
xnor U4335 (N_4335,N_3626,N_3129);
xnor U4336 (N_4336,N_3019,N_3364);
or U4337 (N_4337,N_3097,N_3756);
nor U4338 (N_4338,N_3980,N_3476);
and U4339 (N_4339,N_3136,N_3873);
or U4340 (N_4340,N_3228,N_3183);
nor U4341 (N_4341,N_3726,N_3605);
or U4342 (N_4342,N_3108,N_3680);
nand U4343 (N_4343,N_3450,N_3225);
nor U4344 (N_4344,N_3414,N_3864);
xnor U4345 (N_4345,N_3800,N_3168);
nand U4346 (N_4346,N_3534,N_3015);
or U4347 (N_4347,N_3717,N_3006);
and U4348 (N_4348,N_3038,N_3113);
and U4349 (N_4349,N_3233,N_3441);
xor U4350 (N_4350,N_3353,N_3881);
or U4351 (N_4351,N_3685,N_3673);
nand U4352 (N_4352,N_3170,N_3491);
nand U4353 (N_4353,N_3827,N_3701);
nor U4354 (N_4354,N_3256,N_3566);
and U4355 (N_4355,N_3761,N_3301);
and U4356 (N_4356,N_3147,N_3984);
or U4357 (N_4357,N_3125,N_3526);
and U4358 (N_4358,N_3576,N_3945);
nand U4359 (N_4359,N_3051,N_3925);
nand U4360 (N_4360,N_3080,N_3609);
xor U4361 (N_4361,N_3903,N_3936);
nor U4362 (N_4362,N_3098,N_3883);
nor U4363 (N_4363,N_3453,N_3896);
and U4364 (N_4364,N_3522,N_3188);
and U4365 (N_4365,N_3727,N_3207);
or U4366 (N_4366,N_3443,N_3255);
xnor U4367 (N_4367,N_3508,N_3682);
or U4368 (N_4368,N_3379,N_3830);
nand U4369 (N_4369,N_3992,N_3389);
nand U4370 (N_4370,N_3981,N_3654);
and U4371 (N_4371,N_3245,N_3488);
and U4372 (N_4372,N_3714,N_3623);
nor U4373 (N_4373,N_3362,N_3934);
or U4374 (N_4374,N_3876,N_3031);
nor U4375 (N_4375,N_3820,N_3542);
and U4376 (N_4376,N_3525,N_3141);
nor U4377 (N_4377,N_3569,N_3752);
xnor U4378 (N_4378,N_3791,N_3646);
nor U4379 (N_4379,N_3250,N_3421);
and U4380 (N_4380,N_3240,N_3932);
and U4381 (N_4381,N_3760,N_3594);
xnor U4382 (N_4382,N_3585,N_3190);
xnor U4383 (N_4383,N_3909,N_3707);
nand U4384 (N_4384,N_3971,N_3593);
xnor U4385 (N_4385,N_3075,N_3570);
nor U4386 (N_4386,N_3809,N_3890);
nor U4387 (N_4387,N_3195,N_3013);
nand U4388 (N_4388,N_3198,N_3229);
nor U4389 (N_4389,N_3107,N_3924);
xnor U4390 (N_4390,N_3472,N_3124);
or U4391 (N_4391,N_3915,N_3677);
and U4392 (N_4392,N_3112,N_3528);
xor U4393 (N_4393,N_3363,N_3305);
xnor U4394 (N_4394,N_3880,N_3327);
nor U4395 (N_4395,N_3824,N_3578);
nor U4396 (N_4396,N_3186,N_3077);
xnor U4397 (N_4397,N_3995,N_3101);
nand U4398 (N_4398,N_3378,N_3728);
xnor U4399 (N_4399,N_3160,N_3231);
nor U4400 (N_4400,N_3887,N_3635);
and U4401 (N_4401,N_3872,N_3306);
xor U4402 (N_4402,N_3719,N_3471);
xnor U4403 (N_4403,N_3942,N_3294);
nor U4404 (N_4404,N_3617,N_3746);
or U4405 (N_4405,N_3644,N_3485);
and U4406 (N_4406,N_3507,N_3262);
and U4407 (N_4407,N_3158,N_3417);
nand U4408 (N_4408,N_3373,N_3645);
nor U4409 (N_4409,N_3615,N_3184);
nor U4410 (N_4410,N_3642,N_3041);
or U4411 (N_4411,N_3895,N_3807);
xor U4412 (N_4412,N_3410,N_3597);
and U4413 (N_4413,N_3729,N_3595);
xnor U4414 (N_4414,N_3208,N_3706);
or U4415 (N_4415,N_3773,N_3352);
nand U4416 (N_4416,N_3607,N_3428);
nor U4417 (N_4417,N_3835,N_3338);
and U4418 (N_4418,N_3481,N_3722);
nand U4419 (N_4419,N_3753,N_3904);
nand U4420 (N_4420,N_3152,N_3061);
nand U4421 (N_4421,N_3954,N_3385);
xor U4422 (N_4422,N_3462,N_3935);
xor U4423 (N_4423,N_3510,N_3172);
and U4424 (N_4424,N_3738,N_3182);
or U4425 (N_4425,N_3580,N_3310);
nor U4426 (N_4426,N_3145,N_3393);
or U4427 (N_4427,N_3624,N_3861);
xor U4428 (N_4428,N_3882,N_3571);
or U4429 (N_4429,N_3598,N_3388);
or U4430 (N_4430,N_3552,N_3499);
xor U4431 (N_4431,N_3011,N_3090);
or U4432 (N_4432,N_3322,N_3790);
and U4433 (N_4433,N_3460,N_3639);
xor U4434 (N_4434,N_3083,N_3146);
or U4435 (N_4435,N_3351,N_3610);
nand U4436 (N_4436,N_3541,N_3298);
and U4437 (N_4437,N_3469,N_3448);
nor U4438 (N_4438,N_3561,N_3308);
and U4439 (N_4439,N_3708,N_3702);
and U4440 (N_4440,N_3539,N_3906);
nand U4441 (N_4441,N_3933,N_3289);
nand U4442 (N_4442,N_3018,N_3583);
nand U4443 (N_4443,N_3361,N_3069);
nand U4444 (N_4444,N_3973,N_3711);
or U4445 (N_4445,N_3658,N_3730);
or U4446 (N_4446,N_3688,N_3563);
nor U4447 (N_4447,N_3951,N_3596);
nor U4448 (N_4448,N_3335,N_3852);
nor U4449 (N_4449,N_3689,N_3782);
xor U4450 (N_4450,N_3461,N_3874);
xor U4451 (N_4451,N_3559,N_3741);
or U4452 (N_4452,N_3082,N_3599);
nor U4453 (N_4453,N_3260,N_3095);
and U4454 (N_4454,N_3072,N_3206);
xnor U4455 (N_4455,N_3278,N_3558);
or U4456 (N_4456,N_3520,N_3258);
and U4457 (N_4457,N_3695,N_3263);
or U4458 (N_4458,N_3591,N_3718);
or U4459 (N_4459,N_3867,N_3412);
nand U4460 (N_4460,N_3133,N_3138);
or U4461 (N_4461,N_3109,N_3181);
nand U4462 (N_4462,N_3280,N_3611);
or U4463 (N_4463,N_3050,N_3241);
nand U4464 (N_4464,N_3164,N_3692);
and U4465 (N_4465,N_3762,N_3087);
or U4466 (N_4466,N_3227,N_3696);
and U4467 (N_4467,N_3601,N_3495);
or U4468 (N_4468,N_3304,N_3736);
nand U4469 (N_4469,N_3922,N_3094);
nand U4470 (N_4470,N_3406,N_3407);
nand U4471 (N_4471,N_3991,N_3153);
xnor U4472 (N_4472,N_3334,N_3974);
or U4473 (N_4473,N_3937,N_3833);
and U4474 (N_4474,N_3269,N_3277);
nor U4475 (N_4475,N_3912,N_3600);
and U4476 (N_4476,N_3907,N_3879);
nor U4477 (N_4477,N_3446,N_3333);
nand U4478 (N_4478,N_3440,N_3435);
xor U4479 (N_4479,N_3740,N_3859);
and U4480 (N_4480,N_3505,N_3619);
and U4481 (N_4481,N_3165,N_3286);
nand U4482 (N_4482,N_3219,N_3978);
or U4483 (N_4483,N_3314,N_3724);
or U4484 (N_4484,N_3579,N_3046);
xor U4485 (N_4485,N_3963,N_3150);
and U4486 (N_4486,N_3456,N_3290);
nor U4487 (N_4487,N_3223,N_3863);
or U4488 (N_4488,N_3848,N_3049);
xnor U4489 (N_4489,N_3480,N_3856);
nor U4490 (N_4490,N_3758,N_3641);
xor U4491 (N_4491,N_3826,N_3653);
or U4492 (N_4492,N_3293,N_3538);
and U4493 (N_4493,N_3404,N_3851);
and U4494 (N_4494,N_3687,N_3341);
or U4495 (N_4495,N_3816,N_3036);
xnor U4496 (N_4496,N_3517,N_3678);
nor U4497 (N_4497,N_3045,N_3344);
xnor U4498 (N_4498,N_3218,N_3997);
and U4499 (N_4499,N_3432,N_3151);
nand U4500 (N_4500,N_3237,N_3551);
and U4501 (N_4501,N_3640,N_3503);
nand U4502 (N_4502,N_3437,N_3067);
and U4503 (N_4503,N_3277,N_3095);
and U4504 (N_4504,N_3138,N_3317);
nand U4505 (N_4505,N_3286,N_3556);
and U4506 (N_4506,N_3105,N_3830);
and U4507 (N_4507,N_3800,N_3877);
or U4508 (N_4508,N_3713,N_3961);
nand U4509 (N_4509,N_3016,N_3714);
nand U4510 (N_4510,N_3545,N_3278);
and U4511 (N_4511,N_3142,N_3306);
or U4512 (N_4512,N_3828,N_3415);
or U4513 (N_4513,N_3445,N_3309);
xnor U4514 (N_4514,N_3737,N_3693);
xnor U4515 (N_4515,N_3530,N_3859);
or U4516 (N_4516,N_3050,N_3924);
xor U4517 (N_4517,N_3668,N_3216);
and U4518 (N_4518,N_3876,N_3305);
and U4519 (N_4519,N_3685,N_3765);
and U4520 (N_4520,N_3292,N_3103);
or U4521 (N_4521,N_3417,N_3192);
nand U4522 (N_4522,N_3601,N_3932);
nor U4523 (N_4523,N_3968,N_3671);
xnor U4524 (N_4524,N_3955,N_3444);
nand U4525 (N_4525,N_3906,N_3322);
and U4526 (N_4526,N_3179,N_3369);
and U4527 (N_4527,N_3259,N_3935);
or U4528 (N_4528,N_3337,N_3982);
nand U4529 (N_4529,N_3311,N_3388);
nand U4530 (N_4530,N_3822,N_3924);
xor U4531 (N_4531,N_3958,N_3357);
nand U4532 (N_4532,N_3801,N_3507);
and U4533 (N_4533,N_3092,N_3986);
or U4534 (N_4534,N_3204,N_3094);
and U4535 (N_4535,N_3582,N_3471);
xnor U4536 (N_4536,N_3817,N_3713);
and U4537 (N_4537,N_3013,N_3851);
xnor U4538 (N_4538,N_3370,N_3098);
xnor U4539 (N_4539,N_3538,N_3646);
nor U4540 (N_4540,N_3548,N_3456);
nor U4541 (N_4541,N_3603,N_3093);
nand U4542 (N_4542,N_3966,N_3968);
or U4543 (N_4543,N_3597,N_3362);
or U4544 (N_4544,N_3786,N_3136);
and U4545 (N_4545,N_3760,N_3851);
and U4546 (N_4546,N_3263,N_3775);
and U4547 (N_4547,N_3986,N_3918);
nand U4548 (N_4548,N_3028,N_3899);
nor U4549 (N_4549,N_3937,N_3080);
xor U4550 (N_4550,N_3770,N_3800);
nand U4551 (N_4551,N_3544,N_3301);
nand U4552 (N_4552,N_3379,N_3339);
xnor U4553 (N_4553,N_3457,N_3142);
nand U4554 (N_4554,N_3750,N_3667);
nor U4555 (N_4555,N_3077,N_3207);
and U4556 (N_4556,N_3588,N_3567);
nor U4557 (N_4557,N_3157,N_3462);
xor U4558 (N_4558,N_3314,N_3841);
nor U4559 (N_4559,N_3102,N_3439);
xnor U4560 (N_4560,N_3875,N_3291);
and U4561 (N_4561,N_3081,N_3904);
nand U4562 (N_4562,N_3819,N_3912);
or U4563 (N_4563,N_3289,N_3640);
nor U4564 (N_4564,N_3107,N_3660);
and U4565 (N_4565,N_3204,N_3386);
xnor U4566 (N_4566,N_3280,N_3728);
xor U4567 (N_4567,N_3686,N_3998);
and U4568 (N_4568,N_3074,N_3112);
and U4569 (N_4569,N_3549,N_3063);
nor U4570 (N_4570,N_3019,N_3784);
nand U4571 (N_4571,N_3813,N_3779);
and U4572 (N_4572,N_3175,N_3761);
xor U4573 (N_4573,N_3530,N_3689);
nor U4574 (N_4574,N_3313,N_3706);
and U4575 (N_4575,N_3915,N_3776);
nand U4576 (N_4576,N_3992,N_3483);
nand U4577 (N_4577,N_3072,N_3893);
nor U4578 (N_4578,N_3426,N_3363);
and U4579 (N_4579,N_3094,N_3943);
nand U4580 (N_4580,N_3875,N_3659);
xnor U4581 (N_4581,N_3110,N_3750);
nor U4582 (N_4582,N_3855,N_3845);
xor U4583 (N_4583,N_3894,N_3208);
xor U4584 (N_4584,N_3763,N_3824);
and U4585 (N_4585,N_3408,N_3561);
xor U4586 (N_4586,N_3665,N_3969);
nand U4587 (N_4587,N_3262,N_3190);
nand U4588 (N_4588,N_3405,N_3222);
and U4589 (N_4589,N_3920,N_3945);
nor U4590 (N_4590,N_3059,N_3457);
and U4591 (N_4591,N_3602,N_3925);
or U4592 (N_4592,N_3276,N_3977);
xor U4593 (N_4593,N_3464,N_3516);
xnor U4594 (N_4594,N_3257,N_3888);
nor U4595 (N_4595,N_3865,N_3235);
and U4596 (N_4596,N_3101,N_3549);
nor U4597 (N_4597,N_3238,N_3269);
or U4598 (N_4598,N_3431,N_3459);
xnor U4599 (N_4599,N_3404,N_3049);
nor U4600 (N_4600,N_3811,N_3966);
or U4601 (N_4601,N_3541,N_3046);
and U4602 (N_4602,N_3354,N_3536);
nor U4603 (N_4603,N_3548,N_3682);
or U4604 (N_4604,N_3919,N_3140);
or U4605 (N_4605,N_3138,N_3758);
nor U4606 (N_4606,N_3034,N_3212);
nand U4607 (N_4607,N_3956,N_3463);
nor U4608 (N_4608,N_3279,N_3029);
nor U4609 (N_4609,N_3406,N_3375);
or U4610 (N_4610,N_3676,N_3965);
xnor U4611 (N_4611,N_3105,N_3467);
xnor U4612 (N_4612,N_3149,N_3746);
or U4613 (N_4613,N_3304,N_3894);
nand U4614 (N_4614,N_3279,N_3744);
or U4615 (N_4615,N_3450,N_3905);
nor U4616 (N_4616,N_3291,N_3263);
or U4617 (N_4617,N_3704,N_3208);
or U4618 (N_4618,N_3646,N_3904);
and U4619 (N_4619,N_3168,N_3546);
nor U4620 (N_4620,N_3154,N_3060);
or U4621 (N_4621,N_3185,N_3419);
or U4622 (N_4622,N_3968,N_3167);
xnor U4623 (N_4623,N_3689,N_3892);
nor U4624 (N_4624,N_3082,N_3701);
nor U4625 (N_4625,N_3490,N_3646);
and U4626 (N_4626,N_3560,N_3542);
or U4627 (N_4627,N_3187,N_3370);
xor U4628 (N_4628,N_3760,N_3206);
xnor U4629 (N_4629,N_3985,N_3841);
nand U4630 (N_4630,N_3825,N_3294);
or U4631 (N_4631,N_3669,N_3339);
or U4632 (N_4632,N_3839,N_3693);
and U4633 (N_4633,N_3396,N_3835);
or U4634 (N_4634,N_3727,N_3473);
xor U4635 (N_4635,N_3992,N_3941);
or U4636 (N_4636,N_3711,N_3263);
nand U4637 (N_4637,N_3975,N_3555);
nand U4638 (N_4638,N_3593,N_3342);
xor U4639 (N_4639,N_3157,N_3750);
xnor U4640 (N_4640,N_3437,N_3745);
xnor U4641 (N_4641,N_3372,N_3547);
or U4642 (N_4642,N_3460,N_3768);
nand U4643 (N_4643,N_3058,N_3377);
or U4644 (N_4644,N_3770,N_3849);
xor U4645 (N_4645,N_3958,N_3483);
or U4646 (N_4646,N_3873,N_3878);
xnor U4647 (N_4647,N_3522,N_3504);
and U4648 (N_4648,N_3268,N_3603);
or U4649 (N_4649,N_3041,N_3447);
nor U4650 (N_4650,N_3546,N_3886);
or U4651 (N_4651,N_3214,N_3101);
or U4652 (N_4652,N_3049,N_3445);
xor U4653 (N_4653,N_3290,N_3538);
or U4654 (N_4654,N_3130,N_3169);
xor U4655 (N_4655,N_3520,N_3725);
nand U4656 (N_4656,N_3700,N_3471);
and U4657 (N_4657,N_3483,N_3818);
nor U4658 (N_4658,N_3409,N_3962);
or U4659 (N_4659,N_3663,N_3766);
or U4660 (N_4660,N_3729,N_3012);
xor U4661 (N_4661,N_3439,N_3057);
nor U4662 (N_4662,N_3659,N_3685);
xor U4663 (N_4663,N_3482,N_3370);
or U4664 (N_4664,N_3381,N_3886);
xor U4665 (N_4665,N_3411,N_3242);
nor U4666 (N_4666,N_3244,N_3021);
or U4667 (N_4667,N_3274,N_3162);
nand U4668 (N_4668,N_3716,N_3036);
xnor U4669 (N_4669,N_3721,N_3459);
and U4670 (N_4670,N_3767,N_3059);
or U4671 (N_4671,N_3127,N_3934);
nand U4672 (N_4672,N_3080,N_3362);
nand U4673 (N_4673,N_3977,N_3750);
and U4674 (N_4674,N_3509,N_3907);
nor U4675 (N_4675,N_3519,N_3817);
and U4676 (N_4676,N_3789,N_3727);
and U4677 (N_4677,N_3176,N_3755);
xor U4678 (N_4678,N_3999,N_3057);
nor U4679 (N_4679,N_3143,N_3691);
nand U4680 (N_4680,N_3232,N_3910);
and U4681 (N_4681,N_3473,N_3734);
and U4682 (N_4682,N_3420,N_3768);
or U4683 (N_4683,N_3193,N_3274);
or U4684 (N_4684,N_3019,N_3343);
nor U4685 (N_4685,N_3670,N_3100);
nand U4686 (N_4686,N_3852,N_3025);
or U4687 (N_4687,N_3474,N_3074);
nand U4688 (N_4688,N_3115,N_3602);
or U4689 (N_4689,N_3788,N_3868);
nand U4690 (N_4690,N_3977,N_3423);
and U4691 (N_4691,N_3311,N_3216);
and U4692 (N_4692,N_3959,N_3647);
xor U4693 (N_4693,N_3515,N_3617);
nand U4694 (N_4694,N_3876,N_3811);
xnor U4695 (N_4695,N_3247,N_3239);
xnor U4696 (N_4696,N_3001,N_3979);
and U4697 (N_4697,N_3999,N_3727);
and U4698 (N_4698,N_3190,N_3634);
nand U4699 (N_4699,N_3593,N_3325);
nand U4700 (N_4700,N_3525,N_3020);
and U4701 (N_4701,N_3013,N_3820);
xor U4702 (N_4702,N_3381,N_3467);
xor U4703 (N_4703,N_3534,N_3295);
nand U4704 (N_4704,N_3445,N_3717);
and U4705 (N_4705,N_3591,N_3537);
and U4706 (N_4706,N_3368,N_3614);
nand U4707 (N_4707,N_3590,N_3125);
nand U4708 (N_4708,N_3689,N_3548);
nand U4709 (N_4709,N_3772,N_3248);
xnor U4710 (N_4710,N_3110,N_3727);
xnor U4711 (N_4711,N_3434,N_3424);
and U4712 (N_4712,N_3754,N_3976);
and U4713 (N_4713,N_3154,N_3175);
xnor U4714 (N_4714,N_3303,N_3839);
nand U4715 (N_4715,N_3391,N_3849);
nand U4716 (N_4716,N_3896,N_3227);
or U4717 (N_4717,N_3493,N_3055);
or U4718 (N_4718,N_3255,N_3839);
xor U4719 (N_4719,N_3363,N_3629);
xor U4720 (N_4720,N_3754,N_3442);
or U4721 (N_4721,N_3618,N_3624);
and U4722 (N_4722,N_3668,N_3441);
nand U4723 (N_4723,N_3836,N_3616);
nand U4724 (N_4724,N_3424,N_3351);
and U4725 (N_4725,N_3007,N_3932);
xor U4726 (N_4726,N_3279,N_3759);
xor U4727 (N_4727,N_3474,N_3476);
or U4728 (N_4728,N_3202,N_3444);
and U4729 (N_4729,N_3954,N_3452);
nand U4730 (N_4730,N_3927,N_3372);
nor U4731 (N_4731,N_3436,N_3337);
or U4732 (N_4732,N_3376,N_3168);
nand U4733 (N_4733,N_3055,N_3110);
xor U4734 (N_4734,N_3015,N_3777);
and U4735 (N_4735,N_3128,N_3049);
nor U4736 (N_4736,N_3237,N_3969);
or U4737 (N_4737,N_3063,N_3828);
and U4738 (N_4738,N_3679,N_3457);
or U4739 (N_4739,N_3258,N_3274);
nand U4740 (N_4740,N_3136,N_3359);
or U4741 (N_4741,N_3837,N_3957);
nand U4742 (N_4742,N_3583,N_3827);
nor U4743 (N_4743,N_3890,N_3869);
and U4744 (N_4744,N_3830,N_3529);
and U4745 (N_4745,N_3313,N_3643);
xor U4746 (N_4746,N_3005,N_3938);
and U4747 (N_4747,N_3319,N_3585);
xor U4748 (N_4748,N_3078,N_3940);
or U4749 (N_4749,N_3400,N_3264);
nand U4750 (N_4750,N_3416,N_3119);
or U4751 (N_4751,N_3806,N_3328);
or U4752 (N_4752,N_3313,N_3390);
or U4753 (N_4753,N_3096,N_3612);
xor U4754 (N_4754,N_3440,N_3380);
xnor U4755 (N_4755,N_3097,N_3179);
nand U4756 (N_4756,N_3333,N_3938);
and U4757 (N_4757,N_3422,N_3900);
nand U4758 (N_4758,N_3511,N_3969);
nand U4759 (N_4759,N_3399,N_3190);
or U4760 (N_4760,N_3659,N_3226);
xnor U4761 (N_4761,N_3422,N_3152);
or U4762 (N_4762,N_3264,N_3825);
xor U4763 (N_4763,N_3385,N_3260);
xor U4764 (N_4764,N_3620,N_3201);
or U4765 (N_4765,N_3087,N_3646);
and U4766 (N_4766,N_3242,N_3745);
nor U4767 (N_4767,N_3638,N_3412);
xnor U4768 (N_4768,N_3514,N_3948);
and U4769 (N_4769,N_3530,N_3843);
xor U4770 (N_4770,N_3019,N_3779);
and U4771 (N_4771,N_3364,N_3805);
and U4772 (N_4772,N_3153,N_3270);
nand U4773 (N_4773,N_3956,N_3868);
nand U4774 (N_4774,N_3746,N_3252);
nor U4775 (N_4775,N_3630,N_3035);
or U4776 (N_4776,N_3196,N_3932);
or U4777 (N_4777,N_3714,N_3433);
and U4778 (N_4778,N_3434,N_3659);
and U4779 (N_4779,N_3053,N_3270);
or U4780 (N_4780,N_3246,N_3707);
or U4781 (N_4781,N_3230,N_3692);
and U4782 (N_4782,N_3764,N_3328);
nor U4783 (N_4783,N_3413,N_3014);
or U4784 (N_4784,N_3455,N_3079);
nand U4785 (N_4785,N_3087,N_3862);
nor U4786 (N_4786,N_3365,N_3461);
or U4787 (N_4787,N_3400,N_3088);
xnor U4788 (N_4788,N_3992,N_3321);
nand U4789 (N_4789,N_3093,N_3730);
and U4790 (N_4790,N_3305,N_3553);
and U4791 (N_4791,N_3758,N_3339);
xor U4792 (N_4792,N_3165,N_3171);
xor U4793 (N_4793,N_3720,N_3293);
and U4794 (N_4794,N_3363,N_3999);
nor U4795 (N_4795,N_3944,N_3010);
and U4796 (N_4796,N_3055,N_3540);
and U4797 (N_4797,N_3382,N_3316);
nand U4798 (N_4798,N_3478,N_3461);
or U4799 (N_4799,N_3852,N_3224);
nor U4800 (N_4800,N_3100,N_3264);
or U4801 (N_4801,N_3769,N_3003);
xor U4802 (N_4802,N_3872,N_3723);
nand U4803 (N_4803,N_3046,N_3734);
nor U4804 (N_4804,N_3192,N_3830);
or U4805 (N_4805,N_3168,N_3112);
and U4806 (N_4806,N_3357,N_3166);
nor U4807 (N_4807,N_3272,N_3630);
or U4808 (N_4808,N_3165,N_3814);
and U4809 (N_4809,N_3428,N_3800);
or U4810 (N_4810,N_3676,N_3938);
or U4811 (N_4811,N_3517,N_3316);
nor U4812 (N_4812,N_3941,N_3409);
xor U4813 (N_4813,N_3919,N_3968);
and U4814 (N_4814,N_3475,N_3337);
or U4815 (N_4815,N_3655,N_3715);
or U4816 (N_4816,N_3078,N_3532);
and U4817 (N_4817,N_3858,N_3802);
nor U4818 (N_4818,N_3465,N_3662);
or U4819 (N_4819,N_3859,N_3945);
and U4820 (N_4820,N_3927,N_3688);
xor U4821 (N_4821,N_3210,N_3198);
nor U4822 (N_4822,N_3743,N_3407);
xor U4823 (N_4823,N_3728,N_3927);
or U4824 (N_4824,N_3220,N_3001);
nor U4825 (N_4825,N_3654,N_3435);
and U4826 (N_4826,N_3076,N_3339);
and U4827 (N_4827,N_3861,N_3137);
xor U4828 (N_4828,N_3329,N_3557);
nand U4829 (N_4829,N_3737,N_3884);
xnor U4830 (N_4830,N_3150,N_3189);
xnor U4831 (N_4831,N_3550,N_3943);
xnor U4832 (N_4832,N_3774,N_3355);
and U4833 (N_4833,N_3913,N_3513);
xor U4834 (N_4834,N_3701,N_3975);
nand U4835 (N_4835,N_3665,N_3985);
nand U4836 (N_4836,N_3199,N_3680);
nand U4837 (N_4837,N_3193,N_3130);
or U4838 (N_4838,N_3771,N_3702);
xor U4839 (N_4839,N_3973,N_3563);
or U4840 (N_4840,N_3363,N_3272);
xor U4841 (N_4841,N_3361,N_3851);
and U4842 (N_4842,N_3384,N_3700);
and U4843 (N_4843,N_3771,N_3011);
nand U4844 (N_4844,N_3663,N_3440);
or U4845 (N_4845,N_3127,N_3977);
and U4846 (N_4846,N_3802,N_3132);
xor U4847 (N_4847,N_3152,N_3506);
nand U4848 (N_4848,N_3278,N_3335);
or U4849 (N_4849,N_3038,N_3385);
and U4850 (N_4850,N_3743,N_3468);
or U4851 (N_4851,N_3670,N_3011);
or U4852 (N_4852,N_3279,N_3462);
nor U4853 (N_4853,N_3107,N_3802);
or U4854 (N_4854,N_3945,N_3514);
xnor U4855 (N_4855,N_3932,N_3350);
nor U4856 (N_4856,N_3543,N_3821);
and U4857 (N_4857,N_3245,N_3351);
nor U4858 (N_4858,N_3801,N_3083);
xor U4859 (N_4859,N_3743,N_3907);
nor U4860 (N_4860,N_3619,N_3740);
xor U4861 (N_4861,N_3396,N_3268);
nor U4862 (N_4862,N_3181,N_3384);
nor U4863 (N_4863,N_3780,N_3646);
or U4864 (N_4864,N_3230,N_3114);
nand U4865 (N_4865,N_3867,N_3944);
or U4866 (N_4866,N_3046,N_3808);
or U4867 (N_4867,N_3723,N_3533);
and U4868 (N_4868,N_3831,N_3778);
xnor U4869 (N_4869,N_3940,N_3515);
or U4870 (N_4870,N_3019,N_3601);
and U4871 (N_4871,N_3390,N_3161);
xnor U4872 (N_4872,N_3902,N_3602);
nand U4873 (N_4873,N_3152,N_3184);
xnor U4874 (N_4874,N_3907,N_3931);
or U4875 (N_4875,N_3692,N_3313);
xor U4876 (N_4876,N_3223,N_3292);
nor U4877 (N_4877,N_3766,N_3535);
and U4878 (N_4878,N_3720,N_3696);
and U4879 (N_4879,N_3960,N_3617);
or U4880 (N_4880,N_3226,N_3609);
nor U4881 (N_4881,N_3349,N_3504);
nor U4882 (N_4882,N_3588,N_3597);
nand U4883 (N_4883,N_3703,N_3639);
nor U4884 (N_4884,N_3436,N_3510);
nor U4885 (N_4885,N_3305,N_3104);
nor U4886 (N_4886,N_3920,N_3022);
or U4887 (N_4887,N_3252,N_3878);
and U4888 (N_4888,N_3032,N_3430);
xor U4889 (N_4889,N_3315,N_3317);
nand U4890 (N_4890,N_3930,N_3676);
or U4891 (N_4891,N_3340,N_3388);
xor U4892 (N_4892,N_3441,N_3463);
nand U4893 (N_4893,N_3347,N_3025);
xnor U4894 (N_4894,N_3659,N_3212);
or U4895 (N_4895,N_3752,N_3166);
nor U4896 (N_4896,N_3527,N_3775);
nor U4897 (N_4897,N_3334,N_3129);
nand U4898 (N_4898,N_3471,N_3404);
nor U4899 (N_4899,N_3206,N_3699);
xor U4900 (N_4900,N_3196,N_3395);
or U4901 (N_4901,N_3498,N_3254);
xor U4902 (N_4902,N_3342,N_3130);
and U4903 (N_4903,N_3126,N_3681);
xnor U4904 (N_4904,N_3046,N_3175);
or U4905 (N_4905,N_3669,N_3521);
and U4906 (N_4906,N_3115,N_3014);
nor U4907 (N_4907,N_3199,N_3678);
xor U4908 (N_4908,N_3400,N_3460);
nand U4909 (N_4909,N_3832,N_3867);
or U4910 (N_4910,N_3156,N_3647);
xor U4911 (N_4911,N_3218,N_3527);
nor U4912 (N_4912,N_3997,N_3149);
and U4913 (N_4913,N_3675,N_3468);
nor U4914 (N_4914,N_3737,N_3245);
and U4915 (N_4915,N_3040,N_3213);
nor U4916 (N_4916,N_3025,N_3776);
nand U4917 (N_4917,N_3916,N_3046);
nor U4918 (N_4918,N_3387,N_3318);
xor U4919 (N_4919,N_3982,N_3299);
and U4920 (N_4920,N_3221,N_3487);
or U4921 (N_4921,N_3906,N_3267);
nand U4922 (N_4922,N_3236,N_3610);
and U4923 (N_4923,N_3842,N_3617);
nor U4924 (N_4924,N_3005,N_3341);
and U4925 (N_4925,N_3613,N_3459);
nand U4926 (N_4926,N_3611,N_3578);
nor U4927 (N_4927,N_3371,N_3573);
xor U4928 (N_4928,N_3646,N_3944);
and U4929 (N_4929,N_3367,N_3398);
nor U4930 (N_4930,N_3923,N_3532);
and U4931 (N_4931,N_3597,N_3492);
nand U4932 (N_4932,N_3353,N_3718);
nor U4933 (N_4933,N_3044,N_3731);
and U4934 (N_4934,N_3889,N_3703);
nor U4935 (N_4935,N_3013,N_3778);
nor U4936 (N_4936,N_3411,N_3003);
nor U4937 (N_4937,N_3289,N_3231);
and U4938 (N_4938,N_3094,N_3147);
xnor U4939 (N_4939,N_3237,N_3750);
nand U4940 (N_4940,N_3115,N_3406);
nor U4941 (N_4941,N_3209,N_3684);
nor U4942 (N_4942,N_3015,N_3227);
xor U4943 (N_4943,N_3677,N_3635);
nand U4944 (N_4944,N_3285,N_3386);
xor U4945 (N_4945,N_3271,N_3717);
nand U4946 (N_4946,N_3677,N_3132);
and U4947 (N_4947,N_3779,N_3310);
and U4948 (N_4948,N_3371,N_3798);
nand U4949 (N_4949,N_3871,N_3913);
or U4950 (N_4950,N_3463,N_3506);
and U4951 (N_4951,N_3837,N_3590);
nand U4952 (N_4952,N_3326,N_3458);
xor U4953 (N_4953,N_3233,N_3684);
xor U4954 (N_4954,N_3079,N_3701);
or U4955 (N_4955,N_3661,N_3525);
and U4956 (N_4956,N_3952,N_3979);
nand U4957 (N_4957,N_3320,N_3984);
nor U4958 (N_4958,N_3766,N_3920);
and U4959 (N_4959,N_3865,N_3654);
nand U4960 (N_4960,N_3720,N_3313);
or U4961 (N_4961,N_3782,N_3425);
nor U4962 (N_4962,N_3114,N_3333);
or U4963 (N_4963,N_3043,N_3697);
xnor U4964 (N_4964,N_3257,N_3337);
and U4965 (N_4965,N_3593,N_3337);
xor U4966 (N_4966,N_3059,N_3152);
nor U4967 (N_4967,N_3960,N_3070);
nor U4968 (N_4968,N_3592,N_3179);
nand U4969 (N_4969,N_3344,N_3938);
xnor U4970 (N_4970,N_3638,N_3760);
or U4971 (N_4971,N_3742,N_3052);
and U4972 (N_4972,N_3949,N_3425);
or U4973 (N_4973,N_3476,N_3129);
xor U4974 (N_4974,N_3727,N_3107);
and U4975 (N_4975,N_3146,N_3378);
xor U4976 (N_4976,N_3420,N_3456);
nand U4977 (N_4977,N_3245,N_3083);
nor U4978 (N_4978,N_3573,N_3548);
nand U4979 (N_4979,N_3944,N_3215);
nor U4980 (N_4980,N_3530,N_3298);
nand U4981 (N_4981,N_3581,N_3297);
nor U4982 (N_4982,N_3809,N_3657);
or U4983 (N_4983,N_3317,N_3829);
or U4984 (N_4984,N_3620,N_3606);
or U4985 (N_4985,N_3620,N_3051);
xnor U4986 (N_4986,N_3994,N_3583);
and U4987 (N_4987,N_3104,N_3919);
nand U4988 (N_4988,N_3552,N_3721);
or U4989 (N_4989,N_3857,N_3707);
nor U4990 (N_4990,N_3736,N_3324);
and U4991 (N_4991,N_3543,N_3209);
nand U4992 (N_4992,N_3514,N_3623);
and U4993 (N_4993,N_3491,N_3641);
or U4994 (N_4994,N_3827,N_3835);
xnor U4995 (N_4995,N_3921,N_3945);
nor U4996 (N_4996,N_3113,N_3093);
and U4997 (N_4997,N_3156,N_3997);
and U4998 (N_4998,N_3487,N_3472);
xor U4999 (N_4999,N_3038,N_3217);
or U5000 (N_5000,N_4404,N_4216);
xnor U5001 (N_5001,N_4407,N_4171);
or U5002 (N_5002,N_4324,N_4303);
or U5003 (N_5003,N_4277,N_4594);
xor U5004 (N_5004,N_4622,N_4565);
nor U5005 (N_5005,N_4109,N_4624);
nand U5006 (N_5006,N_4557,N_4647);
nor U5007 (N_5007,N_4527,N_4447);
or U5008 (N_5008,N_4217,N_4950);
nor U5009 (N_5009,N_4784,N_4777);
and U5010 (N_5010,N_4202,N_4646);
nor U5011 (N_5011,N_4899,N_4966);
and U5012 (N_5012,N_4639,N_4862);
nor U5013 (N_5013,N_4045,N_4379);
xnor U5014 (N_5014,N_4755,N_4246);
xnor U5015 (N_5015,N_4026,N_4485);
nor U5016 (N_5016,N_4805,N_4143);
or U5017 (N_5017,N_4386,N_4947);
nand U5018 (N_5018,N_4403,N_4849);
nand U5019 (N_5019,N_4429,N_4833);
xnor U5020 (N_5020,N_4186,N_4920);
nand U5021 (N_5021,N_4278,N_4825);
xnor U5022 (N_5022,N_4121,N_4590);
and U5023 (N_5023,N_4494,N_4205);
xor U5024 (N_5024,N_4453,N_4891);
xnor U5025 (N_5025,N_4270,N_4348);
and U5026 (N_5026,N_4089,N_4929);
and U5027 (N_5027,N_4400,N_4921);
or U5028 (N_5028,N_4712,N_4612);
nand U5029 (N_5029,N_4293,N_4911);
or U5030 (N_5030,N_4245,N_4084);
xor U5031 (N_5031,N_4812,N_4537);
nor U5032 (N_5032,N_4504,N_4123);
or U5033 (N_5033,N_4025,N_4066);
and U5034 (N_5034,N_4640,N_4840);
nor U5035 (N_5035,N_4038,N_4550);
xor U5036 (N_5036,N_4676,N_4809);
and U5037 (N_5037,N_4832,N_4895);
and U5038 (N_5038,N_4319,N_4868);
nor U5039 (N_5039,N_4092,N_4057);
and U5040 (N_5040,N_4367,N_4304);
nand U5041 (N_5041,N_4659,N_4352);
and U5042 (N_5042,N_4432,N_4964);
or U5043 (N_5043,N_4918,N_4154);
nand U5044 (N_5044,N_4933,N_4359);
or U5045 (N_5045,N_4110,N_4059);
and U5046 (N_5046,N_4545,N_4573);
nor U5047 (N_5047,N_4002,N_4489);
nor U5048 (N_5048,N_4028,N_4309);
nor U5049 (N_5049,N_4714,N_4015);
xnor U5050 (N_5050,N_4466,N_4415);
and U5051 (N_5051,N_4881,N_4859);
and U5052 (N_5052,N_4741,N_4175);
nand U5053 (N_5053,N_4495,N_4405);
or U5054 (N_5054,N_4905,N_4858);
xnor U5055 (N_5055,N_4004,N_4611);
nand U5056 (N_5056,N_4915,N_4155);
nand U5057 (N_5057,N_4876,N_4433);
nand U5058 (N_5058,N_4830,N_4315);
and U5059 (N_5059,N_4468,N_4042);
nand U5060 (N_5060,N_4981,N_4364);
and U5061 (N_5061,N_4816,N_4526);
and U5062 (N_5062,N_4257,N_4783);
and U5063 (N_5063,N_4681,N_4058);
nand U5064 (N_5064,N_4987,N_4397);
nor U5065 (N_5065,N_4283,N_4888);
nor U5066 (N_5066,N_4112,N_4148);
nor U5067 (N_5067,N_4363,N_4074);
and U5068 (N_5068,N_4749,N_4583);
xnor U5069 (N_5069,N_4725,N_4700);
xor U5070 (N_5070,N_4321,N_4962);
or U5071 (N_5071,N_4541,N_4815);
nand U5072 (N_5072,N_4563,N_4197);
nand U5073 (N_5073,N_4423,N_4383);
nor U5074 (N_5074,N_4484,N_4803);
xor U5075 (N_5075,N_4238,N_4976);
and U5076 (N_5076,N_4705,N_4768);
and U5077 (N_5077,N_4422,N_4795);
xor U5078 (N_5078,N_4625,N_4836);
xor U5079 (N_5079,N_4663,N_4446);
nor U5080 (N_5080,N_4075,N_4022);
nand U5081 (N_5081,N_4445,N_4956);
nand U5082 (N_5082,N_4564,N_4952);
nand U5083 (N_5083,N_4491,N_4736);
nand U5084 (N_5084,N_4419,N_4431);
nor U5085 (N_5085,N_4925,N_4726);
nor U5086 (N_5086,N_4276,N_4691);
nand U5087 (N_5087,N_4016,N_4299);
or U5088 (N_5088,N_4522,N_4680);
xor U5089 (N_5089,N_4193,N_4543);
and U5090 (N_5090,N_4596,N_4050);
xor U5091 (N_5091,N_4924,N_4312);
nor U5092 (N_5092,N_4887,N_4693);
nand U5093 (N_5093,N_4538,N_4243);
and U5094 (N_5094,N_4571,N_4737);
nor U5095 (N_5095,N_4280,N_4141);
nor U5096 (N_5096,N_4720,N_4983);
or U5097 (N_5097,N_4591,N_4452);
or U5098 (N_5098,N_4461,N_4560);
and U5099 (N_5099,N_4880,N_4839);
and U5100 (N_5100,N_4290,N_4052);
nand U5101 (N_5101,N_4247,N_4963);
and U5102 (N_5102,N_4988,N_4917);
xnor U5103 (N_5103,N_4626,N_4508);
and U5104 (N_5104,N_4706,N_4487);
nand U5105 (N_5105,N_4576,N_4451);
or U5106 (N_5106,N_4150,N_4204);
nand U5107 (N_5107,N_4584,N_4307);
nor U5108 (N_5108,N_4636,N_4819);
or U5109 (N_5109,N_4081,N_4256);
nor U5110 (N_5110,N_4023,N_4960);
xor U5111 (N_5111,N_4475,N_4394);
nor U5112 (N_5112,N_4398,N_4345);
nand U5113 (N_5113,N_4160,N_4897);
or U5114 (N_5114,N_4107,N_4046);
nand U5115 (N_5115,N_4845,N_4174);
and U5116 (N_5116,N_4606,N_4989);
or U5117 (N_5117,N_4800,N_4692);
and U5118 (N_5118,N_4592,N_4686);
and U5119 (N_5119,N_4203,N_4993);
or U5120 (N_5120,N_4296,N_4757);
nand U5121 (N_5121,N_4234,N_4972);
nand U5122 (N_5122,N_4406,N_4745);
or U5123 (N_5123,N_4566,N_4472);
nand U5124 (N_5124,N_4613,N_4088);
and U5125 (N_5125,N_4501,N_4418);
or U5126 (N_5126,N_4834,N_4514);
or U5127 (N_5127,N_4284,N_4267);
and U5128 (N_5128,N_4699,N_4281);
xnor U5129 (N_5129,N_4380,N_4331);
and U5130 (N_5130,N_4879,N_4984);
xor U5131 (N_5131,N_4698,N_4717);
nor U5132 (N_5132,N_4060,N_4730);
or U5133 (N_5133,N_4619,N_4817);
nand U5134 (N_5134,N_4532,N_4497);
xnor U5135 (N_5135,N_4076,N_4306);
or U5136 (N_5136,N_4311,N_4582);
xor U5137 (N_5137,N_4655,N_4765);
nor U5138 (N_5138,N_4941,N_4579);
or U5139 (N_5139,N_4609,N_4152);
or U5140 (N_5140,N_4439,N_4629);
or U5141 (N_5141,N_4919,N_4213);
and U5142 (N_5142,N_4697,N_4760);
or U5143 (N_5143,N_4673,N_4971);
nor U5144 (N_5144,N_4551,N_4580);
nand U5145 (N_5145,N_4967,N_4793);
or U5146 (N_5146,N_4827,N_4035);
xnor U5147 (N_5147,N_4739,N_4190);
nor U5148 (N_5148,N_4512,N_4926);
xor U5149 (N_5149,N_4722,N_4430);
nor U5150 (N_5150,N_4965,N_4562);
xnor U5151 (N_5151,N_4530,N_4601);
nand U5152 (N_5152,N_4464,N_4511);
or U5153 (N_5153,N_4649,N_4342);
nand U5154 (N_5154,N_4934,N_4027);
or U5155 (N_5155,N_4417,N_4391);
nand U5156 (N_5156,N_4347,N_4250);
nor U5157 (N_5157,N_4008,N_4214);
nor U5158 (N_5158,N_4269,N_4224);
and U5159 (N_5159,N_4172,N_4199);
nor U5160 (N_5160,N_4457,N_4033);
nand U5161 (N_5161,N_4240,N_4212);
nor U5162 (N_5162,N_4223,N_4441);
and U5163 (N_5163,N_4338,N_4413);
nand U5164 (N_5164,N_4638,N_4863);
xnor U5165 (N_5165,N_4648,N_4598);
or U5166 (N_5166,N_4853,N_4944);
nor U5167 (N_5167,N_4158,N_4883);
nand U5168 (N_5168,N_4374,N_4589);
xor U5169 (N_5169,N_4228,N_4835);
nor U5170 (N_5170,N_4436,N_4847);
and U5171 (N_5171,N_4822,N_4116);
nor U5172 (N_5172,N_4523,N_4569);
or U5173 (N_5173,N_4459,N_4137);
nor U5174 (N_5174,N_4130,N_4738);
or U5175 (N_5175,N_4753,N_4288);
nand U5176 (N_5176,N_4043,N_4393);
or U5177 (N_5177,N_4420,N_4115);
nand U5178 (N_5178,N_4310,N_4103);
nor U5179 (N_5179,N_4802,N_4011);
nand U5180 (N_5180,N_4159,N_4305);
nor U5181 (N_5181,N_4382,N_4533);
xor U5182 (N_5182,N_4361,N_4558);
or U5183 (N_5183,N_4239,N_4469);
and U5184 (N_5184,N_4916,N_4664);
nor U5185 (N_5185,N_4292,N_4279);
xor U5186 (N_5186,N_4961,N_4326);
nand U5187 (N_5187,N_4282,N_4156);
and U5188 (N_5188,N_4785,N_4470);
and U5189 (N_5189,N_4080,N_4334);
and U5190 (N_5190,N_4848,N_4180);
nor U5191 (N_5191,N_4260,N_4861);
nand U5192 (N_5192,N_4255,N_4153);
xnor U5193 (N_5193,N_4544,N_4442);
and U5194 (N_5194,N_4774,N_4034);
nand U5195 (N_5195,N_4806,N_4846);
nor U5196 (N_5196,N_4721,N_4837);
nand U5197 (N_5197,N_4724,N_4164);
nand U5198 (N_5198,N_4631,N_4670);
nand U5199 (N_5199,N_4574,N_4012);
nand U5200 (N_5200,N_4192,N_4053);
nor U5201 (N_5201,N_4854,N_4796);
or U5202 (N_5202,N_4824,N_4614);
and U5203 (N_5203,N_4426,N_4873);
nor U5204 (N_5204,N_4906,N_4411);
or U5205 (N_5205,N_4082,N_4781);
or U5206 (N_5206,N_4792,N_4652);
nor U5207 (N_5207,N_4097,N_4914);
and U5208 (N_5208,N_4465,N_4069);
xor U5209 (N_5209,N_4946,N_4608);
nand U5210 (N_5210,N_4503,N_4684);
or U5211 (N_5211,N_4567,N_4384);
nor U5212 (N_5212,N_4675,N_4857);
or U5213 (N_5213,N_4500,N_4460);
or U5214 (N_5214,N_4340,N_4823);
and U5215 (N_5215,N_4227,N_4799);
xor U5216 (N_5216,N_4658,N_4147);
nor U5217 (N_5217,N_4617,N_4593);
or U5218 (N_5218,N_4764,N_4923);
and U5219 (N_5219,N_4392,N_4065);
and U5220 (N_5220,N_4300,N_4264);
or U5221 (N_5221,N_4645,N_4759);
and U5222 (N_5222,N_4553,N_4351);
nor U5223 (N_5223,N_4395,N_4808);
nand U5224 (N_5224,N_4168,N_4492);
or U5225 (N_5225,N_4030,N_4695);
nand U5226 (N_5226,N_4992,N_4024);
nor U5227 (N_5227,N_4323,N_4685);
nand U5228 (N_5228,N_4371,N_4597);
xor U5229 (N_5229,N_4463,N_4129);
nand U5230 (N_5230,N_4937,N_4689);
or U5231 (N_5231,N_4122,N_4478);
and U5232 (N_5232,N_4587,N_4274);
xor U5233 (N_5233,N_4729,N_4126);
nor U5234 (N_5234,N_4173,N_4241);
or U5235 (N_5235,N_4771,N_4661);
xor U5236 (N_5236,N_4818,N_4077);
nor U5237 (N_5237,N_4235,N_4095);
xor U5238 (N_5238,N_4249,N_4373);
xor U5239 (N_5239,N_4874,N_4878);
nor U5240 (N_5240,N_4385,N_4814);
or U5241 (N_5241,N_4935,N_4268);
or U5242 (N_5242,N_4291,N_4546);
xnor U5243 (N_5243,N_4146,N_4448);
nor U5244 (N_5244,N_4473,N_4029);
nor U5245 (N_5245,N_4958,N_4525);
or U5246 (N_5246,N_4682,N_4266);
or U5247 (N_5247,N_4851,N_4585);
nor U5248 (N_5248,N_4886,N_4510);
nand U5249 (N_5249,N_4826,N_4850);
xor U5250 (N_5250,N_4940,N_4272);
or U5251 (N_5251,N_4237,N_4618);
or U5252 (N_5252,N_4009,N_4285);
xnor U5253 (N_5253,N_4506,N_4376);
and U5254 (N_5254,N_4381,N_4099);
xor U5255 (N_5255,N_4225,N_4101);
xnor U5256 (N_5256,N_4534,N_4360);
nand U5257 (N_5257,N_4339,N_4356);
or U5258 (N_5258,N_4434,N_4054);
xor U5259 (N_5259,N_4125,N_4995);
and U5260 (N_5260,N_4632,N_4021);
xnor U5261 (N_5261,N_4210,N_4020);
nor U5262 (N_5262,N_4317,N_4456);
and U5263 (N_5263,N_4061,N_4633);
or U5264 (N_5264,N_4111,N_4201);
or U5265 (N_5265,N_4810,N_4733);
xor U5266 (N_5266,N_4412,N_4913);
xnor U5267 (N_5267,N_4807,N_4620);
xnor U5268 (N_5268,N_4083,N_4410);
and U5269 (N_5269,N_4734,N_4483);
nor U5270 (N_5270,N_4679,N_4196);
and U5271 (N_5271,N_4656,N_4499);
nor U5272 (N_5272,N_4337,N_4261);
nor U5273 (N_5273,N_4704,N_4780);
or U5274 (N_5274,N_4586,N_4747);
nor U5275 (N_5275,N_4665,N_4390);
xor U5276 (N_5276,N_4073,N_4401);
xor U5277 (N_5277,N_4302,N_4801);
xor U5278 (N_5278,N_4041,N_4672);
xor U5279 (N_5279,N_4488,N_4108);
nand U5280 (N_5280,N_4355,N_4377);
xor U5281 (N_5281,N_4170,N_4643);
nand U5282 (N_5282,N_4513,N_4654);
nor U5283 (N_5283,N_4169,N_4762);
xnor U5284 (N_5284,N_4683,N_4006);
nand U5285 (N_5285,N_4751,N_4554);
or U5286 (N_5286,N_4408,N_4010);
nor U5287 (N_5287,N_4071,N_4973);
xor U5288 (N_5288,N_4754,N_4570);
nor U5289 (N_5289,N_4273,N_4841);
nor U5290 (N_5290,N_4969,N_4328);
nor U5291 (N_5291,N_4948,N_4875);
or U5292 (N_5292,N_4427,N_4908);
nor U5293 (N_5293,N_4336,N_4215);
nand U5294 (N_5294,N_4229,N_4098);
xnor U5295 (N_5295,N_4425,N_4068);
and U5296 (N_5296,N_4329,N_4298);
nand U5297 (N_5297,N_4767,N_4718);
and U5298 (N_5298,N_4939,N_4909);
nor U5299 (N_5299,N_4630,N_4669);
and U5300 (N_5300,N_4896,N_4244);
nor U5301 (N_5301,N_4572,N_4040);
xnor U5302 (N_5302,N_4829,N_4894);
nand U5303 (N_5303,N_4157,N_4182);
nor U5304 (N_5304,N_4438,N_4688);
nand U5305 (N_5305,N_4974,N_4135);
nor U5306 (N_5306,N_4927,N_4756);
nor U5307 (N_5307,N_4232,N_4703);
and U5308 (N_5308,N_4831,N_4744);
xnor U5309 (N_5309,N_4637,N_4555);
and U5310 (N_5310,N_4540,N_4788);
nand U5311 (N_5311,N_4758,N_4467);
xnor U5312 (N_5312,N_4177,N_4687);
xor U5313 (N_5313,N_4713,N_4354);
or U5314 (N_5314,N_4561,N_4287);
or U5315 (N_5315,N_4165,N_4389);
xnor U5316 (N_5316,N_4662,N_4271);
nand U5317 (N_5317,N_4674,N_4871);
xnor U5318 (N_5318,N_4102,N_4221);
and U5319 (N_5319,N_4322,N_4610);
and U5320 (N_5320,N_4838,N_4032);
nor U5321 (N_5321,N_4399,N_4211);
and U5322 (N_5322,N_4294,N_4772);
and U5323 (N_5323,N_4366,N_4440);
xor U5324 (N_5324,N_4922,N_4127);
and U5325 (N_5325,N_4458,N_4134);
and U5326 (N_5326,N_4036,N_4671);
nor U5327 (N_5327,N_4031,N_4607);
nand U5328 (N_5328,N_4388,N_4990);
and U5329 (N_5329,N_4435,N_4140);
and U5330 (N_5330,N_4362,N_4761);
nand U5331 (N_5331,N_4517,N_4798);
nor U5332 (N_5332,N_4275,N_4811);
xnor U5333 (N_5333,N_4890,N_4051);
nor U5334 (N_5334,N_4982,N_4396);
or U5335 (N_5335,N_4930,N_4943);
nand U5336 (N_5336,N_4444,N_4144);
or U5337 (N_5337,N_4450,N_4124);
nor U5338 (N_5338,N_4820,N_4748);
or U5339 (N_5339,N_4437,N_4200);
nor U5340 (N_5340,N_4657,N_4220);
and U5341 (N_5341,N_4365,N_4882);
or U5342 (N_5342,N_4120,N_4368);
or U5343 (N_5343,N_4536,N_4163);
and U5344 (N_5344,N_4602,N_4480);
or U5345 (N_5345,N_4262,N_4867);
and U5346 (N_5346,N_4207,N_4870);
xor U5347 (N_5347,N_4013,N_4524);
or U5348 (N_5348,N_4454,N_4605);
or U5349 (N_5349,N_4114,N_4001);
nand U5350 (N_5350,N_4954,N_4251);
nor U5351 (N_5351,N_4105,N_4991);
nor U5352 (N_5352,N_4330,N_4770);
or U5353 (N_5353,N_4968,N_4666);
and U5354 (N_5354,N_4949,N_4953);
xor U5355 (N_5355,N_4660,N_4194);
and U5356 (N_5356,N_4187,N_4138);
and U5357 (N_5357,N_4320,N_4118);
nand U5358 (N_5358,N_4865,N_4327);
nand U5359 (N_5359,N_4372,N_4106);
xor U5360 (N_5360,N_4634,N_4219);
and U5361 (N_5361,N_4715,N_4149);
nor U5362 (N_5362,N_4615,N_4603);
nor U5363 (N_5363,N_4975,N_4778);
and U5364 (N_5364,N_4344,N_4980);
nand U5365 (N_5365,N_4094,N_4653);
and U5366 (N_5366,N_4222,N_4297);
xnor U5367 (N_5367,N_4860,N_4252);
and U5368 (N_5368,N_4498,N_4167);
xor U5369 (N_5369,N_4804,N_4998);
nand U5370 (N_5370,N_4142,N_4677);
nor U5371 (N_5371,N_4064,N_4719);
nand U5372 (N_5372,N_4085,N_4985);
xnor U5373 (N_5373,N_4507,N_4628);
nor U5374 (N_5374,N_4341,N_4047);
nor U5375 (N_5375,N_4486,N_4242);
and U5376 (N_5376,N_4369,N_4039);
nor U5377 (N_5377,N_4017,N_4635);
and U5378 (N_5378,N_4402,N_4902);
and U5379 (N_5379,N_4178,N_4308);
and U5380 (N_5380,N_4353,N_4893);
or U5381 (N_5381,N_4938,N_4575);
or U5382 (N_5382,N_4889,N_4179);
nand U5383 (N_5383,N_4481,N_4387);
and U5384 (N_5384,N_4707,N_4236);
nand U5385 (N_5385,N_4014,N_4866);
and U5386 (N_5386,N_4037,N_4132);
nor U5387 (N_5387,N_4185,N_4462);
and U5388 (N_5388,N_4195,N_4184);
or U5389 (N_5389,N_4740,N_4313);
and U5390 (N_5390,N_4056,N_4230);
nor U5391 (N_5391,N_4128,N_4782);
xor U5392 (N_5392,N_4421,N_4723);
xnor U5393 (N_5393,N_4790,N_4710);
and U5394 (N_5394,N_4455,N_4568);
nor U5395 (N_5395,N_4977,N_4789);
or U5396 (N_5396,N_4959,N_4424);
nor U5397 (N_5397,N_4623,N_4139);
and U5398 (N_5398,N_4496,N_4335);
xnor U5399 (N_5399,N_4951,N_4086);
xnor U5400 (N_5400,N_4314,N_4901);
nor U5401 (N_5401,N_4932,N_4233);
nor U5402 (N_5402,N_4333,N_4477);
xnor U5403 (N_5403,N_4955,N_4884);
and U5404 (N_5404,N_4779,N_4316);
nand U5405 (N_5405,N_4520,N_4078);
and U5406 (N_5406,N_4642,N_4869);
xor U5407 (N_5407,N_4588,N_4581);
or U5408 (N_5408,N_4189,N_4957);
and U5409 (N_5409,N_4709,N_4048);
nand U5410 (N_5410,N_4842,N_4482);
and U5411 (N_5411,N_4070,N_4100);
nor U5412 (N_5412,N_4518,N_4117);
nor U5413 (N_5413,N_4528,N_4728);
nor U5414 (N_5414,N_4776,N_4090);
and U5415 (N_5415,N_4191,N_4005);
or U5416 (N_5416,N_4375,N_4821);
xnor U5417 (N_5417,N_4794,N_4539);
or U5418 (N_5418,N_4621,N_4119);
nand U5419 (N_5419,N_4515,N_4079);
nand U5420 (N_5420,N_4254,N_4828);
or U5421 (N_5421,N_4742,N_4295);
xor U5422 (N_5422,N_4253,N_4378);
or U5423 (N_5423,N_4529,N_4265);
nand U5424 (N_5424,N_4750,N_4556);
and U5425 (N_5425,N_4996,N_4667);
xor U5426 (N_5426,N_4549,N_4516);
xnor U5427 (N_5427,N_4131,N_4797);
nand U5428 (N_5428,N_4490,N_4161);
or U5429 (N_5429,N_4259,N_4735);
and U5430 (N_5430,N_4502,N_4509);
and U5431 (N_5431,N_4904,N_4521);
and U5432 (N_5432,N_4209,N_4151);
and U5433 (N_5433,N_4994,N_4578);
xor U5434 (N_5434,N_4535,N_4852);
xor U5435 (N_5435,N_4104,N_4018);
xnor U5436 (N_5436,N_4711,N_4844);
or U5437 (N_5437,N_4176,N_4049);
and U5438 (N_5438,N_4616,N_4595);
xor U5439 (N_5439,N_4651,N_4231);
and U5440 (N_5440,N_4763,N_4542);
nand U5441 (N_5441,N_4443,N_4072);
and U5442 (N_5442,N_4218,N_4289);
nor U5443 (N_5443,N_4900,N_4096);
and U5444 (N_5444,N_4258,N_4206);
nor U5445 (N_5445,N_4449,N_4007);
xor U5446 (N_5446,N_4577,N_4226);
nand U5447 (N_5447,N_4349,N_4208);
nor U5448 (N_5448,N_4248,N_4903);
or U5449 (N_5449,N_4000,N_4731);
or U5450 (N_5450,N_4505,N_4343);
xor U5451 (N_5451,N_4787,N_4732);
nor U5452 (N_5452,N_4864,N_4727);
xnor U5453 (N_5453,N_4766,N_4198);
nand U5454 (N_5454,N_4936,N_4907);
nand U5455 (N_5455,N_4559,N_4087);
xor U5456 (N_5456,N_4414,N_4696);
xnor U5457 (N_5457,N_4892,N_4773);
nand U5458 (N_5458,N_4062,N_4346);
nand U5459 (N_5459,N_4332,N_4548);
xor U5460 (N_5460,N_4743,N_4769);
or U5461 (N_5461,N_4428,N_4912);
or U5462 (N_5462,N_4843,N_4350);
nand U5463 (N_5463,N_4690,N_4519);
nand U5464 (N_5464,N_4650,N_4701);
nand U5465 (N_5465,N_4286,N_4325);
or U5466 (N_5466,N_4409,N_4370);
nand U5467 (N_5467,N_4627,N_4694);
nor U5468 (N_5468,N_4970,N_4063);
nand U5469 (N_5469,N_4928,N_4945);
nor U5470 (N_5470,N_4877,N_4145);
nor U5471 (N_5471,N_4746,N_4856);
or U5472 (N_5472,N_4872,N_4986);
nand U5473 (N_5473,N_4318,N_4855);
xor U5474 (N_5474,N_4188,N_4416);
or U5475 (N_5475,N_4067,N_4166);
and U5476 (N_5476,N_4604,N_4133);
nand U5477 (N_5477,N_4479,N_4471);
nand U5478 (N_5478,N_4600,N_4716);
and U5479 (N_5479,N_4357,N_4910);
nor U5480 (N_5480,N_4997,N_4183);
or U5481 (N_5481,N_4552,N_4474);
or U5482 (N_5482,N_4885,N_4931);
or U5483 (N_5483,N_4942,N_4786);
nor U5484 (N_5484,N_4044,N_4547);
xnor U5485 (N_5485,N_4668,N_4708);
xor U5486 (N_5486,N_4702,N_4476);
and U5487 (N_5487,N_4813,N_4791);
xor U5488 (N_5488,N_4599,N_4136);
nor U5489 (N_5489,N_4493,N_4775);
xor U5490 (N_5490,N_4091,N_4003);
nor U5491 (N_5491,N_4181,N_4301);
xnor U5492 (N_5492,N_4093,N_4641);
nand U5493 (N_5493,N_4644,N_4019);
and U5494 (N_5494,N_4752,N_4531);
nand U5495 (N_5495,N_4898,N_4113);
and U5496 (N_5496,N_4358,N_4055);
nand U5497 (N_5497,N_4999,N_4678);
nand U5498 (N_5498,N_4162,N_4979);
nor U5499 (N_5499,N_4263,N_4978);
nand U5500 (N_5500,N_4595,N_4698);
nor U5501 (N_5501,N_4039,N_4735);
and U5502 (N_5502,N_4464,N_4841);
and U5503 (N_5503,N_4008,N_4834);
nand U5504 (N_5504,N_4038,N_4880);
nor U5505 (N_5505,N_4277,N_4218);
nand U5506 (N_5506,N_4111,N_4682);
nand U5507 (N_5507,N_4780,N_4874);
nor U5508 (N_5508,N_4687,N_4658);
xnor U5509 (N_5509,N_4543,N_4423);
nor U5510 (N_5510,N_4547,N_4218);
nor U5511 (N_5511,N_4352,N_4330);
or U5512 (N_5512,N_4567,N_4806);
xor U5513 (N_5513,N_4031,N_4173);
or U5514 (N_5514,N_4721,N_4359);
xor U5515 (N_5515,N_4558,N_4118);
and U5516 (N_5516,N_4498,N_4795);
and U5517 (N_5517,N_4480,N_4040);
nand U5518 (N_5518,N_4000,N_4610);
nand U5519 (N_5519,N_4124,N_4912);
or U5520 (N_5520,N_4658,N_4391);
and U5521 (N_5521,N_4319,N_4415);
and U5522 (N_5522,N_4725,N_4401);
or U5523 (N_5523,N_4360,N_4773);
and U5524 (N_5524,N_4522,N_4569);
and U5525 (N_5525,N_4868,N_4445);
nand U5526 (N_5526,N_4251,N_4212);
nor U5527 (N_5527,N_4189,N_4089);
or U5528 (N_5528,N_4363,N_4274);
xor U5529 (N_5529,N_4078,N_4580);
or U5530 (N_5530,N_4765,N_4868);
and U5531 (N_5531,N_4927,N_4526);
nand U5532 (N_5532,N_4866,N_4962);
xnor U5533 (N_5533,N_4744,N_4105);
nand U5534 (N_5534,N_4104,N_4558);
nand U5535 (N_5535,N_4122,N_4568);
xor U5536 (N_5536,N_4168,N_4748);
nor U5537 (N_5537,N_4022,N_4872);
nor U5538 (N_5538,N_4402,N_4166);
nand U5539 (N_5539,N_4253,N_4732);
xnor U5540 (N_5540,N_4141,N_4395);
nand U5541 (N_5541,N_4145,N_4710);
nand U5542 (N_5542,N_4462,N_4573);
nor U5543 (N_5543,N_4661,N_4139);
or U5544 (N_5544,N_4894,N_4517);
nor U5545 (N_5545,N_4789,N_4669);
and U5546 (N_5546,N_4000,N_4746);
xnor U5547 (N_5547,N_4065,N_4393);
or U5548 (N_5548,N_4304,N_4018);
xnor U5549 (N_5549,N_4362,N_4077);
xnor U5550 (N_5550,N_4690,N_4513);
and U5551 (N_5551,N_4897,N_4106);
nor U5552 (N_5552,N_4394,N_4956);
xnor U5553 (N_5553,N_4945,N_4099);
and U5554 (N_5554,N_4989,N_4973);
nand U5555 (N_5555,N_4258,N_4040);
or U5556 (N_5556,N_4683,N_4181);
xnor U5557 (N_5557,N_4048,N_4654);
or U5558 (N_5558,N_4616,N_4104);
nand U5559 (N_5559,N_4210,N_4028);
or U5560 (N_5560,N_4022,N_4099);
xnor U5561 (N_5561,N_4921,N_4801);
nor U5562 (N_5562,N_4162,N_4172);
nand U5563 (N_5563,N_4703,N_4800);
and U5564 (N_5564,N_4175,N_4133);
nor U5565 (N_5565,N_4150,N_4014);
or U5566 (N_5566,N_4129,N_4893);
xor U5567 (N_5567,N_4850,N_4233);
xnor U5568 (N_5568,N_4718,N_4696);
nor U5569 (N_5569,N_4631,N_4674);
and U5570 (N_5570,N_4598,N_4232);
xnor U5571 (N_5571,N_4242,N_4352);
and U5572 (N_5572,N_4228,N_4219);
or U5573 (N_5573,N_4133,N_4370);
nor U5574 (N_5574,N_4813,N_4999);
nor U5575 (N_5575,N_4484,N_4263);
nand U5576 (N_5576,N_4955,N_4038);
xor U5577 (N_5577,N_4177,N_4452);
xnor U5578 (N_5578,N_4215,N_4555);
nor U5579 (N_5579,N_4377,N_4023);
or U5580 (N_5580,N_4579,N_4914);
nand U5581 (N_5581,N_4085,N_4057);
xor U5582 (N_5582,N_4532,N_4879);
or U5583 (N_5583,N_4135,N_4575);
xor U5584 (N_5584,N_4694,N_4664);
nand U5585 (N_5585,N_4949,N_4202);
nand U5586 (N_5586,N_4307,N_4018);
nand U5587 (N_5587,N_4169,N_4147);
nand U5588 (N_5588,N_4647,N_4166);
nor U5589 (N_5589,N_4326,N_4013);
xor U5590 (N_5590,N_4629,N_4282);
xnor U5591 (N_5591,N_4758,N_4559);
or U5592 (N_5592,N_4873,N_4565);
or U5593 (N_5593,N_4789,N_4323);
xnor U5594 (N_5594,N_4294,N_4390);
nor U5595 (N_5595,N_4157,N_4836);
xor U5596 (N_5596,N_4993,N_4536);
and U5597 (N_5597,N_4823,N_4714);
or U5598 (N_5598,N_4268,N_4265);
or U5599 (N_5599,N_4299,N_4738);
or U5600 (N_5600,N_4303,N_4087);
nand U5601 (N_5601,N_4840,N_4812);
nand U5602 (N_5602,N_4569,N_4207);
xor U5603 (N_5603,N_4321,N_4172);
nand U5604 (N_5604,N_4168,N_4981);
and U5605 (N_5605,N_4634,N_4591);
or U5606 (N_5606,N_4519,N_4990);
xnor U5607 (N_5607,N_4510,N_4010);
nor U5608 (N_5608,N_4186,N_4226);
or U5609 (N_5609,N_4607,N_4561);
xnor U5610 (N_5610,N_4324,N_4071);
nor U5611 (N_5611,N_4647,N_4452);
xor U5612 (N_5612,N_4601,N_4261);
and U5613 (N_5613,N_4500,N_4417);
or U5614 (N_5614,N_4315,N_4753);
nor U5615 (N_5615,N_4095,N_4420);
and U5616 (N_5616,N_4557,N_4241);
nand U5617 (N_5617,N_4343,N_4340);
nand U5618 (N_5618,N_4499,N_4411);
nand U5619 (N_5619,N_4099,N_4387);
or U5620 (N_5620,N_4994,N_4628);
nand U5621 (N_5621,N_4037,N_4593);
nand U5622 (N_5622,N_4990,N_4030);
nor U5623 (N_5623,N_4451,N_4146);
and U5624 (N_5624,N_4109,N_4513);
nor U5625 (N_5625,N_4861,N_4715);
and U5626 (N_5626,N_4014,N_4846);
and U5627 (N_5627,N_4694,N_4805);
xnor U5628 (N_5628,N_4090,N_4411);
xnor U5629 (N_5629,N_4213,N_4029);
xor U5630 (N_5630,N_4582,N_4102);
and U5631 (N_5631,N_4030,N_4156);
nor U5632 (N_5632,N_4134,N_4393);
and U5633 (N_5633,N_4739,N_4356);
or U5634 (N_5634,N_4204,N_4482);
xnor U5635 (N_5635,N_4972,N_4192);
nand U5636 (N_5636,N_4065,N_4090);
or U5637 (N_5637,N_4436,N_4574);
xor U5638 (N_5638,N_4004,N_4091);
and U5639 (N_5639,N_4561,N_4302);
and U5640 (N_5640,N_4899,N_4906);
or U5641 (N_5641,N_4800,N_4048);
nor U5642 (N_5642,N_4132,N_4855);
nand U5643 (N_5643,N_4763,N_4397);
xnor U5644 (N_5644,N_4436,N_4494);
xor U5645 (N_5645,N_4722,N_4877);
nand U5646 (N_5646,N_4668,N_4302);
nor U5647 (N_5647,N_4419,N_4398);
nor U5648 (N_5648,N_4880,N_4177);
xor U5649 (N_5649,N_4410,N_4583);
nor U5650 (N_5650,N_4097,N_4897);
and U5651 (N_5651,N_4118,N_4925);
or U5652 (N_5652,N_4947,N_4850);
nor U5653 (N_5653,N_4595,N_4704);
and U5654 (N_5654,N_4941,N_4477);
nor U5655 (N_5655,N_4169,N_4506);
xnor U5656 (N_5656,N_4954,N_4667);
nand U5657 (N_5657,N_4431,N_4985);
nor U5658 (N_5658,N_4062,N_4185);
nand U5659 (N_5659,N_4948,N_4586);
nor U5660 (N_5660,N_4862,N_4554);
nand U5661 (N_5661,N_4394,N_4863);
xnor U5662 (N_5662,N_4932,N_4410);
nor U5663 (N_5663,N_4460,N_4914);
nor U5664 (N_5664,N_4943,N_4732);
nand U5665 (N_5665,N_4225,N_4994);
or U5666 (N_5666,N_4890,N_4958);
nand U5667 (N_5667,N_4630,N_4401);
nor U5668 (N_5668,N_4917,N_4914);
nor U5669 (N_5669,N_4895,N_4422);
and U5670 (N_5670,N_4294,N_4658);
nor U5671 (N_5671,N_4495,N_4260);
and U5672 (N_5672,N_4408,N_4368);
nor U5673 (N_5673,N_4448,N_4737);
nand U5674 (N_5674,N_4581,N_4723);
xor U5675 (N_5675,N_4963,N_4353);
xor U5676 (N_5676,N_4829,N_4364);
xor U5677 (N_5677,N_4836,N_4543);
or U5678 (N_5678,N_4949,N_4704);
nor U5679 (N_5679,N_4767,N_4443);
nand U5680 (N_5680,N_4395,N_4109);
and U5681 (N_5681,N_4406,N_4694);
or U5682 (N_5682,N_4673,N_4682);
nor U5683 (N_5683,N_4301,N_4110);
nand U5684 (N_5684,N_4948,N_4140);
nor U5685 (N_5685,N_4413,N_4398);
nor U5686 (N_5686,N_4023,N_4256);
or U5687 (N_5687,N_4222,N_4457);
and U5688 (N_5688,N_4431,N_4176);
or U5689 (N_5689,N_4666,N_4199);
nand U5690 (N_5690,N_4958,N_4377);
nor U5691 (N_5691,N_4897,N_4764);
nor U5692 (N_5692,N_4207,N_4738);
or U5693 (N_5693,N_4296,N_4585);
nor U5694 (N_5694,N_4963,N_4186);
nand U5695 (N_5695,N_4360,N_4218);
xnor U5696 (N_5696,N_4917,N_4746);
nand U5697 (N_5697,N_4699,N_4763);
and U5698 (N_5698,N_4854,N_4991);
or U5699 (N_5699,N_4739,N_4803);
or U5700 (N_5700,N_4970,N_4803);
and U5701 (N_5701,N_4291,N_4320);
and U5702 (N_5702,N_4098,N_4633);
nand U5703 (N_5703,N_4578,N_4517);
and U5704 (N_5704,N_4861,N_4993);
and U5705 (N_5705,N_4104,N_4284);
nand U5706 (N_5706,N_4732,N_4239);
and U5707 (N_5707,N_4990,N_4802);
or U5708 (N_5708,N_4922,N_4889);
or U5709 (N_5709,N_4927,N_4830);
nor U5710 (N_5710,N_4626,N_4248);
xnor U5711 (N_5711,N_4971,N_4152);
nor U5712 (N_5712,N_4924,N_4223);
or U5713 (N_5713,N_4384,N_4064);
or U5714 (N_5714,N_4930,N_4919);
nand U5715 (N_5715,N_4957,N_4726);
nor U5716 (N_5716,N_4387,N_4143);
nand U5717 (N_5717,N_4984,N_4590);
and U5718 (N_5718,N_4834,N_4074);
xnor U5719 (N_5719,N_4382,N_4558);
or U5720 (N_5720,N_4483,N_4565);
or U5721 (N_5721,N_4031,N_4028);
and U5722 (N_5722,N_4462,N_4018);
nand U5723 (N_5723,N_4231,N_4946);
nor U5724 (N_5724,N_4762,N_4037);
xnor U5725 (N_5725,N_4245,N_4658);
nor U5726 (N_5726,N_4625,N_4650);
xnor U5727 (N_5727,N_4421,N_4464);
xor U5728 (N_5728,N_4189,N_4888);
nor U5729 (N_5729,N_4919,N_4017);
xnor U5730 (N_5730,N_4206,N_4334);
or U5731 (N_5731,N_4432,N_4268);
or U5732 (N_5732,N_4223,N_4992);
nor U5733 (N_5733,N_4089,N_4236);
and U5734 (N_5734,N_4878,N_4322);
nand U5735 (N_5735,N_4811,N_4036);
nor U5736 (N_5736,N_4540,N_4503);
nand U5737 (N_5737,N_4763,N_4799);
nand U5738 (N_5738,N_4948,N_4137);
xor U5739 (N_5739,N_4085,N_4919);
xor U5740 (N_5740,N_4244,N_4226);
xor U5741 (N_5741,N_4488,N_4874);
nor U5742 (N_5742,N_4080,N_4062);
xor U5743 (N_5743,N_4492,N_4706);
nor U5744 (N_5744,N_4208,N_4523);
nand U5745 (N_5745,N_4181,N_4896);
nand U5746 (N_5746,N_4164,N_4669);
or U5747 (N_5747,N_4084,N_4375);
nor U5748 (N_5748,N_4532,N_4538);
or U5749 (N_5749,N_4795,N_4393);
and U5750 (N_5750,N_4521,N_4944);
nor U5751 (N_5751,N_4610,N_4121);
and U5752 (N_5752,N_4124,N_4664);
xnor U5753 (N_5753,N_4055,N_4314);
nor U5754 (N_5754,N_4399,N_4690);
nand U5755 (N_5755,N_4149,N_4609);
or U5756 (N_5756,N_4883,N_4169);
or U5757 (N_5757,N_4411,N_4944);
nand U5758 (N_5758,N_4510,N_4250);
nor U5759 (N_5759,N_4319,N_4085);
nand U5760 (N_5760,N_4003,N_4800);
xor U5761 (N_5761,N_4691,N_4966);
nor U5762 (N_5762,N_4434,N_4991);
xor U5763 (N_5763,N_4908,N_4288);
or U5764 (N_5764,N_4584,N_4168);
or U5765 (N_5765,N_4409,N_4154);
and U5766 (N_5766,N_4951,N_4548);
or U5767 (N_5767,N_4535,N_4038);
xor U5768 (N_5768,N_4791,N_4638);
and U5769 (N_5769,N_4102,N_4657);
and U5770 (N_5770,N_4831,N_4948);
xor U5771 (N_5771,N_4820,N_4640);
xor U5772 (N_5772,N_4627,N_4390);
or U5773 (N_5773,N_4437,N_4569);
or U5774 (N_5774,N_4526,N_4271);
or U5775 (N_5775,N_4915,N_4502);
nand U5776 (N_5776,N_4710,N_4446);
nand U5777 (N_5777,N_4785,N_4583);
nor U5778 (N_5778,N_4093,N_4106);
nor U5779 (N_5779,N_4351,N_4963);
nor U5780 (N_5780,N_4012,N_4389);
xor U5781 (N_5781,N_4566,N_4271);
and U5782 (N_5782,N_4143,N_4385);
nor U5783 (N_5783,N_4957,N_4204);
nor U5784 (N_5784,N_4041,N_4469);
xnor U5785 (N_5785,N_4063,N_4234);
and U5786 (N_5786,N_4295,N_4170);
and U5787 (N_5787,N_4200,N_4397);
xor U5788 (N_5788,N_4594,N_4655);
xnor U5789 (N_5789,N_4939,N_4625);
and U5790 (N_5790,N_4087,N_4258);
nor U5791 (N_5791,N_4122,N_4045);
nor U5792 (N_5792,N_4781,N_4273);
nor U5793 (N_5793,N_4624,N_4202);
xor U5794 (N_5794,N_4461,N_4046);
nand U5795 (N_5795,N_4567,N_4399);
or U5796 (N_5796,N_4435,N_4212);
nand U5797 (N_5797,N_4837,N_4132);
xor U5798 (N_5798,N_4287,N_4328);
and U5799 (N_5799,N_4807,N_4704);
nor U5800 (N_5800,N_4037,N_4806);
xor U5801 (N_5801,N_4288,N_4473);
xnor U5802 (N_5802,N_4751,N_4090);
xnor U5803 (N_5803,N_4500,N_4900);
nor U5804 (N_5804,N_4373,N_4559);
nand U5805 (N_5805,N_4243,N_4286);
and U5806 (N_5806,N_4467,N_4594);
nand U5807 (N_5807,N_4548,N_4296);
nand U5808 (N_5808,N_4674,N_4630);
xnor U5809 (N_5809,N_4018,N_4030);
nand U5810 (N_5810,N_4639,N_4519);
nand U5811 (N_5811,N_4118,N_4204);
xnor U5812 (N_5812,N_4340,N_4055);
and U5813 (N_5813,N_4852,N_4181);
xnor U5814 (N_5814,N_4626,N_4381);
nand U5815 (N_5815,N_4286,N_4497);
or U5816 (N_5816,N_4914,N_4959);
xnor U5817 (N_5817,N_4373,N_4653);
and U5818 (N_5818,N_4602,N_4814);
nor U5819 (N_5819,N_4916,N_4136);
and U5820 (N_5820,N_4029,N_4767);
and U5821 (N_5821,N_4173,N_4136);
nor U5822 (N_5822,N_4274,N_4376);
nor U5823 (N_5823,N_4333,N_4398);
or U5824 (N_5824,N_4511,N_4050);
nand U5825 (N_5825,N_4467,N_4046);
nand U5826 (N_5826,N_4897,N_4328);
or U5827 (N_5827,N_4282,N_4744);
xor U5828 (N_5828,N_4330,N_4520);
nor U5829 (N_5829,N_4324,N_4905);
and U5830 (N_5830,N_4672,N_4738);
nand U5831 (N_5831,N_4337,N_4119);
or U5832 (N_5832,N_4210,N_4266);
or U5833 (N_5833,N_4446,N_4373);
and U5834 (N_5834,N_4768,N_4269);
or U5835 (N_5835,N_4297,N_4790);
xor U5836 (N_5836,N_4989,N_4453);
nor U5837 (N_5837,N_4373,N_4094);
or U5838 (N_5838,N_4128,N_4859);
nor U5839 (N_5839,N_4068,N_4605);
or U5840 (N_5840,N_4709,N_4220);
nand U5841 (N_5841,N_4048,N_4517);
nand U5842 (N_5842,N_4403,N_4468);
or U5843 (N_5843,N_4138,N_4207);
xor U5844 (N_5844,N_4120,N_4853);
or U5845 (N_5845,N_4271,N_4757);
and U5846 (N_5846,N_4436,N_4676);
or U5847 (N_5847,N_4038,N_4834);
nand U5848 (N_5848,N_4862,N_4041);
and U5849 (N_5849,N_4537,N_4650);
and U5850 (N_5850,N_4276,N_4903);
and U5851 (N_5851,N_4629,N_4579);
nor U5852 (N_5852,N_4125,N_4518);
or U5853 (N_5853,N_4662,N_4230);
xor U5854 (N_5854,N_4461,N_4790);
xnor U5855 (N_5855,N_4386,N_4744);
or U5856 (N_5856,N_4386,N_4992);
nor U5857 (N_5857,N_4169,N_4862);
nor U5858 (N_5858,N_4044,N_4996);
and U5859 (N_5859,N_4748,N_4412);
and U5860 (N_5860,N_4146,N_4579);
and U5861 (N_5861,N_4883,N_4748);
nand U5862 (N_5862,N_4478,N_4040);
and U5863 (N_5863,N_4493,N_4934);
xnor U5864 (N_5864,N_4386,N_4085);
and U5865 (N_5865,N_4764,N_4547);
nand U5866 (N_5866,N_4867,N_4256);
nand U5867 (N_5867,N_4608,N_4596);
nand U5868 (N_5868,N_4015,N_4014);
xnor U5869 (N_5869,N_4753,N_4242);
and U5870 (N_5870,N_4698,N_4490);
nand U5871 (N_5871,N_4794,N_4420);
nor U5872 (N_5872,N_4480,N_4719);
and U5873 (N_5873,N_4057,N_4497);
and U5874 (N_5874,N_4538,N_4306);
or U5875 (N_5875,N_4627,N_4805);
nand U5876 (N_5876,N_4058,N_4360);
or U5877 (N_5877,N_4613,N_4371);
or U5878 (N_5878,N_4776,N_4388);
nand U5879 (N_5879,N_4158,N_4760);
or U5880 (N_5880,N_4269,N_4100);
nand U5881 (N_5881,N_4060,N_4677);
nor U5882 (N_5882,N_4708,N_4719);
nor U5883 (N_5883,N_4431,N_4757);
and U5884 (N_5884,N_4275,N_4368);
nor U5885 (N_5885,N_4303,N_4835);
or U5886 (N_5886,N_4802,N_4393);
nand U5887 (N_5887,N_4555,N_4964);
nor U5888 (N_5888,N_4733,N_4232);
nand U5889 (N_5889,N_4395,N_4305);
and U5890 (N_5890,N_4165,N_4527);
xnor U5891 (N_5891,N_4924,N_4975);
nor U5892 (N_5892,N_4433,N_4029);
nand U5893 (N_5893,N_4983,N_4828);
or U5894 (N_5894,N_4858,N_4783);
or U5895 (N_5895,N_4379,N_4031);
nor U5896 (N_5896,N_4455,N_4298);
or U5897 (N_5897,N_4258,N_4946);
or U5898 (N_5898,N_4760,N_4050);
or U5899 (N_5899,N_4215,N_4668);
nor U5900 (N_5900,N_4838,N_4377);
nand U5901 (N_5901,N_4382,N_4209);
nand U5902 (N_5902,N_4225,N_4656);
nand U5903 (N_5903,N_4260,N_4041);
nand U5904 (N_5904,N_4249,N_4399);
nor U5905 (N_5905,N_4880,N_4028);
and U5906 (N_5906,N_4709,N_4337);
xnor U5907 (N_5907,N_4217,N_4369);
nand U5908 (N_5908,N_4267,N_4610);
nand U5909 (N_5909,N_4011,N_4203);
or U5910 (N_5910,N_4458,N_4332);
nand U5911 (N_5911,N_4377,N_4135);
and U5912 (N_5912,N_4401,N_4271);
and U5913 (N_5913,N_4294,N_4225);
nor U5914 (N_5914,N_4953,N_4326);
xor U5915 (N_5915,N_4484,N_4008);
nand U5916 (N_5916,N_4771,N_4110);
nor U5917 (N_5917,N_4695,N_4918);
nand U5918 (N_5918,N_4349,N_4345);
nor U5919 (N_5919,N_4401,N_4636);
xnor U5920 (N_5920,N_4488,N_4827);
and U5921 (N_5921,N_4996,N_4679);
nand U5922 (N_5922,N_4088,N_4038);
or U5923 (N_5923,N_4337,N_4759);
xnor U5924 (N_5924,N_4142,N_4683);
nor U5925 (N_5925,N_4711,N_4845);
nor U5926 (N_5926,N_4760,N_4067);
and U5927 (N_5927,N_4420,N_4736);
nand U5928 (N_5928,N_4958,N_4765);
nor U5929 (N_5929,N_4065,N_4416);
xor U5930 (N_5930,N_4453,N_4630);
nand U5931 (N_5931,N_4062,N_4193);
nor U5932 (N_5932,N_4795,N_4707);
nand U5933 (N_5933,N_4069,N_4509);
xnor U5934 (N_5934,N_4585,N_4467);
nor U5935 (N_5935,N_4561,N_4132);
or U5936 (N_5936,N_4094,N_4581);
xor U5937 (N_5937,N_4302,N_4144);
nor U5938 (N_5938,N_4614,N_4586);
nand U5939 (N_5939,N_4084,N_4527);
xnor U5940 (N_5940,N_4651,N_4149);
or U5941 (N_5941,N_4868,N_4793);
xnor U5942 (N_5942,N_4835,N_4944);
nand U5943 (N_5943,N_4528,N_4370);
nor U5944 (N_5944,N_4266,N_4426);
nand U5945 (N_5945,N_4605,N_4707);
or U5946 (N_5946,N_4355,N_4553);
nor U5947 (N_5947,N_4449,N_4348);
or U5948 (N_5948,N_4814,N_4774);
nand U5949 (N_5949,N_4271,N_4269);
or U5950 (N_5950,N_4376,N_4026);
nor U5951 (N_5951,N_4723,N_4736);
and U5952 (N_5952,N_4379,N_4475);
or U5953 (N_5953,N_4910,N_4655);
xor U5954 (N_5954,N_4654,N_4234);
nand U5955 (N_5955,N_4921,N_4479);
and U5956 (N_5956,N_4834,N_4344);
nor U5957 (N_5957,N_4756,N_4650);
xnor U5958 (N_5958,N_4034,N_4184);
nor U5959 (N_5959,N_4266,N_4980);
xor U5960 (N_5960,N_4729,N_4984);
and U5961 (N_5961,N_4245,N_4833);
and U5962 (N_5962,N_4093,N_4736);
and U5963 (N_5963,N_4253,N_4712);
nand U5964 (N_5964,N_4848,N_4131);
nand U5965 (N_5965,N_4806,N_4990);
nor U5966 (N_5966,N_4326,N_4889);
nor U5967 (N_5967,N_4254,N_4900);
and U5968 (N_5968,N_4140,N_4408);
and U5969 (N_5969,N_4053,N_4368);
nand U5970 (N_5970,N_4779,N_4482);
and U5971 (N_5971,N_4782,N_4340);
or U5972 (N_5972,N_4942,N_4127);
xor U5973 (N_5973,N_4184,N_4275);
nand U5974 (N_5974,N_4055,N_4293);
nand U5975 (N_5975,N_4042,N_4680);
or U5976 (N_5976,N_4300,N_4261);
xnor U5977 (N_5977,N_4884,N_4463);
nor U5978 (N_5978,N_4553,N_4158);
xnor U5979 (N_5979,N_4930,N_4934);
and U5980 (N_5980,N_4042,N_4907);
or U5981 (N_5981,N_4034,N_4606);
xor U5982 (N_5982,N_4086,N_4637);
nor U5983 (N_5983,N_4418,N_4881);
xnor U5984 (N_5984,N_4456,N_4243);
and U5985 (N_5985,N_4179,N_4578);
and U5986 (N_5986,N_4365,N_4292);
xor U5987 (N_5987,N_4297,N_4174);
and U5988 (N_5988,N_4164,N_4928);
and U5989 (N_5989,N_4275,N_4307);
or U5990 (N_5990,N_4184,N_4608);
or U5991 (N_5991,N_4321,N_4903);
nor U5992 (N_5992,N_4967,N_4285);
nand U5993 (N_5993,N_4045,N_4143);
and U5994 (N_5994,N_4984,N_4835);
xnor U5995 (N_5995,N_4954,N_4492);
and U5996 (N_5996,N_4058,N_4996);
and U5997 (N_5997,N_4862,N_4519);
xnor U5998 (N_5998,N_4274,N_4914);
xnor U5999 (N_5999,N_4049,N_4266);
and U6000 (N_6000,N_5034,N_5962);
xor U6001 (N_6001,N_5727,N_5688);
and U6002 (N_6002,N_5801,N_5771);
nor U6003 (N_6003,N_5265,N_5552);
or U6004 (N_6004,N_5492,N_5024);
xor U6005 (N_6005,N_5021,N_5286);
xnor U6006 (N_6006,N_5385,N_5884);
or U6007 (N_6007,N_5025,N_5754);
nor U6008 (N_6008,N_5347,N_5646);
or U6009 (N_6009,N_5732,N_5082);
nand U6010 (N_6010,N_5847,N_5791);
nor U6011 (N_6011,N_5018,N_5151);
or U6012 (N_6012,N_5364,N_5616);
xnor U6013 (N_6013,N_5127,N_5147);
nor U6014 (N_6014,N_5271,N_5993);
nand U6015 (N_6015,N_5348,N_5572);
or U6016 (N_6016,N_5504,N_5963);
xnor U6017 (N_6017,N_5096,N_5189);
xor U6018 (N_6018,N_5695,N_5242);
xnor U6019 (N_6019,N_5674,N_5063);
nor U6020 (N_6020,N_5078,N_5828);
and U6021 (N_6021,N_5359,N_5883);
xnor U6022 (N_6022,N_5533,N_5457);
or U6023 (N_6023,N_5879,N_5972);
and U6024 (N_6024,N_5991,N_5509);
and U6025 (N_6025,N_5800,N_5042);
or U6026 (N_6026,N_5454,N_5167);
and U6027 (N_6027,N_5470,N_5876);
xnor U6028 (N_6028,N_5463,N_5448);
xnor U6029 (N_6029,N_5611,N_5916);
nor U6030 (N_6030,N_5798,N_5396);
or U6031 (N_6031,N_5226,N_5164);
nor U6032 (N_6032,N_5440,N_5925);
and U6033 (N_6033,N_5994,N_5829);
nor U6034 (N_6034,N_5941,N_5651);
nor U6035 (N_6035,N_5569,N_5842);
nor U6036 (N_6036,N_5395,N_5686);
and U6037 (N_6037,N_5355,N_5642);
nand U6038 (N_6038,N_5554,N_5239);
or U6039 (N_6039,N_5205,N_5526);
nand U6040 (N_6040,N_5425,N_5679);
or U6041 (N_6041,N_5669,N_5843);
or U6042 (N_6042,N_5822,N_5356);
nor U6043 (N_6043,N_5452,N_5950);
nand U6044 (N_6044,N_5817,N_5826);
nor U6045 (N_6045,N_5442,N_5146);
and U6046 (N_6046,N_5134,N_5767);
xnor U6047 (N_6047,N_5224,N_5917);
nand U6048 (N_6048,N_5989,N_5525);
nand U6049 (N_6049,N_5091,N_5506);
nand U6050 (N_6050,N_5550,N_5543);
nand U6051 (N_6051,N_5663,N_5183);
nor U6052 (N_6052,N_5320,N_5805);
nand U6053 (N_6053,N_5423,N_5712);
and U6054 (N_6054,N_5198,N_5468);
or U6055 (N_6055,N_5045,N_5460);
or U6056 (N_6056,N_5904,N_5176);
or U6057 (N_6057,N_5584,N_5105);
xor U6058 (N_6058,N_5296,N_5580);
and U6059 (N_6059,N_5621,N_5086);
or U6060 (N_6060,N_5092,N_5330);
nor U6061 (N_6061,N_5726,N_5048);
and U6062 (N_6062,N_5590,N_5441);
or U6063 (N_6063,N_5041,N_5603);
xor U6064 (N_6064,N_5053,N_5627);
or U6065 (N_6065,N_5786,N_5598);
nand U6066 (N_6066,N_5974,N_5629);
or U6067 (N_6067,N_5586,N_5599);
xor U6068 (N_6068,N_5277,N_5612);
xnor U6069 (N_6069,N_5938,N_5957);
xor U6070 (N_6070,N_5606,N_5336);
nand U6071 (N_6071,N_5966,N_5403);
xor U6072 (N_6072,N_5520,N_5943);
and U6073 (N_6073,N_5417,N_5834);
nor U6074 (N_6074,N_5303,N_5148);
or U6075 (N_6075,N_5382,N_5353);
xor U6076 (N_6076,N_5668,N_5722);
and U6077 (N_6077,N_5389,N_5664);
xor U6078 (N_6078,N_5307,N_5793);
nor U6079 (N_6079,N_5539,N_5778);
nor U6080 (N_6080,N_5536,N_5282);
nand U6081 (N_6081,N_5777,N_5190);
nor U6082 (N_6082,N_5420,N_5749);
xor U6083 (N_6083,N_5772,N_5229);
and U6084 (N_6084,N_5773,N_5225);
and U6085 (N_6085,N_5819,N_5243);
xor U6086 (N_6086,N_5683,N_5415);
nand U6087 (N_6087,N_5581,N_5267);
nand U6088 (N_6088,N_5233,N_5115);
or U6089 (N_6089,N_5033,N_5366);
nand U6090 (N_6090,N_5371,N_5909);
and U6091 (N_6091,N_5593,N_5835);
and U6092 (N_6092,N_5076,N_5394);
nand U6093 (N_6093,N_5751,N_5634);
xor U6094 (N_6094,N_5792,N_5367);
nand U6095 (N_6095,N_5212,N_5874);
xnor U6096 (N_6096,N_5799,N_5142);
nand U6097 (N_6097,N_5975,N_5133);
and U6098 (N_6098,N_5971,N_5781);
and U6099 (N_6099,N_5535,N_5764);
nand U6100 (N_6100,N_5861,N_5928);
nor U6101 (N_6101,N_5338,N_5335);
or U6102 (N_6102,N_5859,N_5156);
nor U6103 (N_6103,N_5545,N_5266);
and U6104 (N_6104,N_5108,N_5854);
or U6105 (N_6105,N_5221,N_5062);
nor U6106 (N_6106,N_5649,N_5685);
xnor U6107 (N_6107,N_5517,N_5121);
xnor U6108 (N_6108,N_5191,N_5731);
nor U6109 (N_6109,N_5272,N_5245);
nor U6110 (N_6110,N_5377,N_5787);
nor U6111 (N_6111,N_5428,N_5459);
or U6112 (N_6112,N_5057,N_5852);
nand U6113 (N_6113,N_5345,N_5500);
nor U6114 (N_6114,N_5085,N_5630);
xnor U6115 (N_6115,N_5215,N_5472);
nand U6116 (N_6116,N_5788,N_5940);
nand U6117 (N_6117,N_5703,N_5114);
nor U6118 (N_6118,N_5900,N_5295);
nor U6119 (N_6119,N_5376,N_5275);
and U6120 (N_6120,N_5650,N_5476);
xnor U6121 (N_6121,N_5565,N_5163);
or U6122 (N_6122,N_5567,N_5093);
and U6123 (N_6123,N_5583,N_5182);
or U6124 (N_6124,N_5639,N_5564);
xor U6125 (N_6125,N_5813,N_5160);
nand U6126 (N_6126,N_5246,N_5313);
and U6127 (N_6127,N_5387,N_5125);
or U6128 (N_6128,N_5138,N_5723);
xor U6129 (N_6129,N_5869,N_5162);
or U6130 (N_6130,N_5112,N_5426);
nand U6131 (N_6131,N_5103,N_5432);
nor U6132 (N_6132,N_5809,N_5628);
xor U6133 (N_6133,N_5109,N_5578);
nor U6134 (N_6134,N_5770,N_5740);
nor U6135 (N_6135,N_5064,N_5475);
nand U6136 (N_6136,N_5661,N_5568);
or U6137 (N_6137,N_5942,N_5481);
nor U6138 (N_6138,N_5269,N_5720);
and U6139 (N_6139,N_5849,N_5635);
and U6140 (N_6140,N_5766,N_5036);
or U6141 (N_6141,N_5206,N_5231);
xnor U6142 (N_6142,N_5002,N_5696);
nand U6143 (N_6143,N_5370,N_5692);
nor U6144 (N_6144,N_5824,N_5424);
nand U6145 (N_6145,N_5549,N_5633);
nand U6146 (N_6146,N_5363,N_5278);
nor U6147 (N_6147,N_5181,N_5038);
xnor U6148 (N_6148,N_5710,N_5193);
nor U6149 (N_6149,N_5840,N_5706);
nand U6150 (N_6150,N_5268,N_5238);
xnor U6151 (N_6151,N_5083,N_5640);
nand U6152 (N_6152,N_5050,N_5850);
nand U6153 (N_6153,N_5073,N_5736);
and U6154 (N_6154,N_5281,N_5742);
nand U6155 (N_6155,N_5702,N_5136);
nand U6156 (N_6156,N_5982,N_5297);
xor U6157 (N_6157,N_5592,N_5241);
and U6158 (N_6158,N_5340,N_5744);
and U6159 (N_6159,N_5293,N_5891);
and U6160 (N_6160,N_5285,N_5289);
or U6161 (N_6161,N_5375,N_5131);
xor U6162 (N_6162,N_5350,N_5343);
or U6163 (N_6163,N_5218,N_5524);
or U6164 (N_6164,N_5204,N_5645);
nor U6165 (N_6165,N_5422,N_5689);
and U6166 (N_6166,N_5935,N_5124);
nor U6167 (N_6167,N_5899,N_5489);
nand U6168 (N_6168,N_5601,N_5166);
or U6169 (N_6169,N_5066,N_5965);
nand U6170 (N_6170,N_5806,N_5625);
nand U6171 (N_6171,N_5930,N_5381);
xnor U6172 (N_6172,N_5737,N_5538);
or U6173 (N_6173,N_5283,N_5264);
xor U6174 (N_6174,N_5200,N_5249);
xnor U6175 (N_6175,N_5230,N_5017);
nand U6176 (N_6176,N_5467,N_5469);
nand U6177 (N_6177,N_5986,N_5914);
and U6178 (N_6178,N_5069,N_5179);
or U6179 (N_6179,N_5889,N_5443);
and U6180 (N_6180,N_5790,N_5450);
nand U6181 (N_6181,N_5043,N_5833);
nand U6182 (N_6182,N_5969,N_5956);
xnor U6183 (N_6183,N_5429,N_5310);
or U6184 (N_6184,N_5372,N_5028);
nor U6185 (N_6185,N_5318,N_5309);
nor U6186 (N_6186,N_5122,N_5352);
xor U6187 (N_6187,N_5911,N_5001);
nor U6188 (N_6188,N_5358,N_5201);
xor U6189 (N_6189,N_5090,N_5258);
and U6190 (N_6190,N_5923,N_5701);
and U6191 (N_6191,N_5551,N_5186);
nand U6192 (N_6192,N_5102,N_5088);
nor U6193 (N_6193,N_5211,N_5287);
and U6194 (N_6194,N_5743,N_5814);
or U6195 (N_6195,N_5576,N_5292);
nor U6196 (N_6196,N_5818,N_5919);
nand U6197 (N_6197,N_5810,N_5161);
xor U6198 (N_6198,N_5501,N_5519);
nand U6199 (N_6199,N_5208,N_5841);
nand U6200 (N_6200,N_5071,N_5838);
and U6201 (N_6201,N_5217,N_5196);
nor U6202 (N_6202,N_5721,N_5011);
and U6203 (N_6203,N_5404,N_5939);
and U6204 (N_6204,N_5312,N_5715);
nor U6205 (N_6205,N_5279,N_5080);
nor U6206 (N_6206,N_5557,N_5753);
xnor U6207 (N_6207,N_5298,N_5158);
xnor U6208 (N_6208,N_5321,N_5037);
and U6209 (N_6209,N_5747,N_5487);
xor U6210 (N_6210,N_5046,N_5110);
and U6211 (N_6211,N_5014,N_5780);
nand U6212 (N_6212,N_5708,N_5479);
nand U6213 (N_6213,N_5860,N_5739);
nor U6214 (N_6214,N_5932,N_5153);
xnor U6215 (N_6215,N_5416,N_5301);
xnor U6216 (N_6216,N_5027,N_5608);
and U6217 (N_6217,N_5623,N_5734);
nand U6218 (N_6218,N_5199,N_5234);
or U6219 (N_6219,N_5529,N_5169);
or U6220 (N_6220,N_5261,N_5155);
xor U6221 (N_6221,N_5290,N_5738);
nor U6222 (N_6222,N_5380,N_5936);
nor U6223 (N_6223,N_5390,N_5180);
and U6224 (N_6224,N_5613,N_5253);
and U6225 (N_6225,N_5713,N_5111);
nor U6226 (N_6226,N_5979,N_5887);
xnor U6227 (N_6227,N_5931,N_5202);
and U6228 (N_6228,N_5259,N_5354);
nand U6229 (N_6229,N_5797,N_5273);
and U6230 (N_6230,N_5893,N_5728);
or U6231 (N_6231,N_5302,N_5100);
or U6232 (N_6232,N_5015,N_5362);
xnor U6233 (N_6233,N_5074,N_5845);
and U6234 (N_6234,N_5653,N_5832);
xor U6235 (N_6235,N_5216,N_5300);
nand U6236 (N_6236,N_5915,N_5735);
nor U6237 (N_6237,N_5808,N_5398);
and U6238 (N_6238,N_5958,N_5471);
nand U6239 (N_6239,N_5383,N_5905);
nor U6240 (N_6240,N_5903,N_5856);
nand U6241 (N_6241,N_5756,N_5049);
or U6242 (N_6242,N_5837,N_5368);
or U6243 (N_6243,N_5405,N_5369);
and U6244 (N_6244,N_5433,N_5748);
nor U6245 (N_6245,N_5349,N_5502);
and U6246 (N_6246,N_5528,N_5174);
and U6247 (N_6247,N_5484,N_5126);
nor U6248 (N_6248,N_5235,N_5591);
nor U6249 (N_6249,N_5937,N_5711);
nor U6250 (N_6250,N_5908,N_5888);
xnor U6251 (N_6251,N_5673,N_5906);
nor U6252 (N_6252,N_5351,N_5365);
xor U6253 (N_6253,N_5563,N_5816);
xor U6254 (N_6254,N_5513,N_5473);
or U6255 (N_6255,N_5830,N_5435);
nor U6256 (N_6256,N_5339,N_5836);
nand U6257 (N_6257,N_5719,N_5907);
or U6258 (N_6258,N_5388,N_5516);
nor U6259 (N_6259,N_5095,N_5141);
or U6260 (N_6260,N_5152,N_5707);
xor U6261 (N_6261,N_5803,N_5746);
nand U6262 (N_6262,N_5718,N_5776);
nor U6263 (N_6263,N_5026,N_5980);
nand U6264 (N_6264,N_5288,N_5408);
nand U6265 (N_6265,N_5765,N_5761);
xor U6266 (N_6266,N_5948,N_5760);
and U6267 (N_6267,N_5056,N_5401);
or U6268 (N_6268,N_5610,N_5544);
xnor U6269 (N_6269,N_5047,N_5973);
nor U6270 (N_6270,N_5030,N_5665);
and U6271 (N_6271,N_5863,N_5944);
or U6272 (N_6272,N_5392,N_5522);
nor U6273 (N_6273,N_5400,N_5490);
nand U6274 (N_6274,N_5699,N_5750);
xor U6275 (N_6275,N_5546,N_5219);
nand U6276 (N_6276,N_5600,N_5494);
and U6277 (N_6277,N_5412,N_5276);
and U6278 (N_6278,N_5004,N_5990);
or U6279 (N_6279,N_5391,N_5007);
or U6280 (N_6280,N_5117,N_5924);
and U6281 (N_6281,N_5755,N_5065);
or U6282 (N_6282,N_5588,N_5875);
and U6283 (N_6283,N_5029,N_5060);
and U6284 (N_6284,N_5120,N_5531);
or U6285 (N_6285,N_5260,N_5143);
xor U6286 (N_6286,N_5055,N_5514);
xnor U6287 (N_6287,N_5573,N_5019);
nand U6288 (N_6288,N_5725,N_5556);
nand U6289 (N_6289,N_5137,N_5717);
nor U6290 (N_6290,N_5676,N_5058);
nand U6291 (N_6291,N_5192,N_5465);
or U6292 (N_6292,N_5154,N_5178);
and U6293 (N_6293,N_5762,N_5223);
nand U6294 (N_6294,N_5051,N_5327);
and U6295 (N_6295,N_5763,N_5427);
xor U6296 (N_6296,N_5220,N_5537);
and U6297 (N_6297,N_5970,N_5698);
xnor U6298 (N_6298,N_5173,N_5342);
xnor U6299 (N_6299,N_5729,N_5263);
and U6300 (N_6300,N_5107,N_5857);
and U6301 (N_6301,N_5248,N_5308);
xnor U6302 (N_6302,N_5922,N_5988);
nand U6303 (N_6303,N_5855,N_5194);
xor U6304 (N_6304,N_5040,N_5687);
and U6305 (N_6305,N_5684,N_5784);
and U6306 (N_6306,N_5150,N_5254);
or U6307 (N_6307,N_5123,N_5605);
nand U6308 (N_6308,N_5885,N_5532);
or U6309 (N_6309,N_5437,N_5961);
or U6310 (N_6310,N_5654,N_5682);
and U6311 (N_6311,N_5839,N_5553);
nand U6312 (N_6312,N_5118,N_5009);
nor U6313 (N_6313,N_5119,N_5631);
xor U6314 (N_6314,N_5411,N_5992);
and U6315 (N_6315,N_5305,N_5172);
nand U6316 (N_6316,N_5329,N_5068);
and U6317 (N_6317,N_5087,N_5977);
xnor U6318 (N_6318,N_5304,N_5324);
or U6319 (N_6319,N_5759,N_5099);
xnor U6320 (N_6320,N_5256,N_5149);
or U6321 (N_6321,N_5474,N_5694);
or U6322 (N_6322,N_5769,N_5185);
or U6323 (N_6323,N_5555,N_5116);
nand U6324 (N_6324,N_5171,N_5414);
xnor U6325 (N_6325,N_5890,N_5913);
xor U6326 (N_6326,N_5848,N_5785);
and U6327 (N_6327,N_5745,N_5097);
or U6328 (N_6328,N_5602,N_5491);
nand U6329 (N_6329,N_5498,N_5831);
nor U6330 (N_6330,N_5807,N_5378);
xnor U6331 (N_6331,N_5020,N_5503);
nor U6332 (N_6332,N_5976,N_5978);
xnor U6333 (N_6333,N_5579,N_5796);
nand U6334 (N_6334,N_5952,N_5059);
xnor U6335 (N_6335,N_5130,N_5637);
xor U6336 (N_6336,N_5252,N_5901);
and U6337 (N_6337,N_5098,N_5140);
or U6338 (N_6338,N_5203,N_5228);
or U6339 (N_6339,N_5575,N_5488);
and U6340 (N_6340,N_5455,N_5458);
nand U6341 (N_6341,N_5604,N_5210);
and U6342 (N_6342,N_5315,N_5089);
or U6343 (N_6343,N_5571,N_5968);
nand U6344 (N_6344,N_5862,N_5274);
or U6345 (N_6345,N_5188,N_5559);
nor U6346 (N_6346,N_5132,N_5647);
nand U6347 (N_6347,N_5620,N_5508);
and U6348 (N_6348,N_5644,N_5896);
and U6349 (N_6349,N_5779,N_5912);
or U6350 (N_6350,N_5039,N_5496);
and U6351 (N_6351,N_5827,N_5983);
xnor U6352 (N_6352,N_5951,N_5825);
nand U6353 (N_6353,N_5314,N_5864);
and U6354 (N_6354,N_5566,N_5878);
or U6355 (N_6355,N_5540,N_5758);
or U6356 (N_6356,N_5866,N_5168);
nor U6357 (N_6357,N_5334,N_5407);
nand U6358 (N_6358,N_5462,N_5195);
xnor U6359 (N_6359,N_5733,N_5232);
nand U6360 (N_6360,N_5386,N_5461);
xor U6361 (N_6361,N_5714,N_5270);
and U6362 (N_6362,N_5430,N_5344);
nand U6363 (N_6363,N_5693,N_5477);
nor U6364 (N_6364,N_5445,N_5444);
or U6365 (N_6365,N_5752,N_5657);
xor U6366 (N_6366,N_5548,N_5031);
and U6367 (N_6367,N_5337,N_5022);
or U6368 (N_6368,N_5933,N_5655);
nand U6369 (N_6369,N_5851,N_5811);
nor U6370 (N_6370,N_5280,N_5374);
nand U6371 (N_6371,N_5724,N_5128);
and U6372 (N_6372,N_5618,N_5624);
or U6373 (N_6373,N_5013,N_5902);
and U6374 (N_6374,N_5981,N_5322);
nand U6375 (N_6375,N_5081,N_5177);
and U6376 (N_6376,N_5844,N_5010);
and U6377 (N_6377,N_5691,N_5954);
xnor U6378 (N_6378,N_5678,N_5317);
nand U6379 (N_6379,N_5449,N_5061);
nand U6380 (N_6380,N_5697,N_5871);
nand U6381 (N_6381,N_5257,N_5542);
xor U6382 (N_6382,N_5619,N_5328);
and U6383 (N_6383,N_5789,N_5892);
or U6384 (N_6384,N_5480,N_5333);
and U6385 (N_6385,N_5596,N_5658);
or U6386 (N_6386,N_5486,N_5493);
xnor U6387 (N_6387,N_5521,N_5853);
nor U6388 (N_6388,N_5434,N_5341);
xnor U6389 (N_6389,N_5413,N_5291);
and U6390 (N_6390,N_5570,N_5898);
nor U6391 (N_6391,N_5084,N_5299);
or U6392 (N_6392,N_5464,N_5964);
nor U6393 (N_6393,N_5187,N_5453);
nor U6394 (N_6394,N_5709,N_5595);
xor U6395 (N_6395,N_5802,N_5730);
or U6396 (N_6396,N_5894,N_5794);
xnor U6397 (N_6397,N_5244,N_5373);
or U6398 (N_6398,N_5451,N_5251);
or U6399 (N_6399,N_5774,N_5240);
nor U6400 (N_6400,N_5667,N_5632);
nand U6401 (N_6401,N_5527,N_5886);
nor U6402 (N_6402,N_5577,N_5671);
and U6403 (N_6403,N_5823,N_5466);
and U6404 (N_6404,N_5880,N_5741);
xnor U6405 (N_6405,N_5323,N_5918);
or U6406 (N_6406,N_5873,N_5035);
xor U6407 (N_6407,N_5998,N_5384);
nand U6408 (N_6408,N_5607,N_5804);
and U6409 (N_6409,N_5615,N_5139);
and U6410 (N_6410,N_5512,N_5052);
and U6411 (N_6411,N_5012,N_5659);
xnor U6412 (N_6412,N_5106,N_5070);
xor U6413 (N_6413,N_5626,N_5782);
or U6414 (N_6414,N_5016,N_5237);
and U6415 (N_6415,N_5775,N_5582);
nand U6416 (N_6416,N_5497,N_5757);
and U6417 (N_6417,N_5690,N_5795);
nor U6418 (N_6418,N_5006,N_5431);
or U6419 (N_6419,N_5409,N_5507);
and U6420 (N_6420,N_5032,N_5820);
and U6421 (N_6421,N_5129,N_5929);
and U6422 (N_6422,N_5222,N_5000);
and U6423 (N_6423,N_5705,N_5960);
or U6424 (N_6424,N_5945,N_5947);
xnor U6425 (N_6425,N_5560,N_5700);
nand U6426 (N_6426,N_5648,N_5921);
and U6427 (N_6427,N_5541,N_5585);
or U6428 (N_6428,N_5675,N_5934);
nand U6429 (N_6429,N_5609,N_5574);
nor U6430 (N_6430,N_5159,N_5325);
nand U6431 (N_6431,N_5184,N_5326);
and U6432 (N_6432,N_5589,N_5439);
or U6433 (N_6433,N_5999,N_5868);
nor U6434 (N_6434,N_5145,N_5867);
nand U6435 (N_6435,N_5846,N_5421);
or U6436 (N_6436,N_5558,N_5996);
nand U6437 (N_6437,N_5547,N_5967);
nand U6438 (N_6438,N_5997,N_5144);
nor U6439 (N_6439,N_5670,N_5207);
or U6440 (N_6440,N_5008,N_5495);
and U6441 (N_6441,N_5920,N_5680);
nand U6442 (N_6442,N_5023,N_5227);
or U6443 (N_6443,N_5306,N_5597);
xnor U6444 (N_6444,N_5783,N_5406);
xnor U6445 (N_6445,N_5858,N_5079);
nor U6446 (N_6446,N_5643,N_5067);
nor U6447 (N_6447,N_5331,N_5209);
or U6448 (N_6448,N_5666,N_5077);
or U6449 (N_6449,N_5402,N_5821);
or U6450 (N_6450,N_5101,N_5534);
nor U6451 (N_6451,N_5294,N_5213);
nand U6452 (N_6452,N_5247,N_5870);
nand U6453 (N_6453,N_5446,N_5005);
nor U6454 (N_6454,N_5499,N_5346);
xor U6455 (N_6455,N_5250,N_5872);
nand U6456 (N_6456,N_5987,N_5515);
nand U6457 (N_6457,N_5561,N_5003);
nor U6458 (N_6458,N_5895,N_5418);
and U6459 (N_6459,N_5897,N_5165);
nand U6460 (N_6460,N_5959,N_5946);
or U6461 (N_6461,N_5704,N_5113);
and U6462 (N_6462,N_5478,N_5054);
and U6463 (N_6463,N_5399,N_5438);
or U6464 (N_6464,N_5636,N_5094);
nor U6465 (N_6465,N_5170,N_5436);
nor U6466 (N_6466,N_5638,N_5511);
and U6467 (N_6467,N_5316,N_5660);
xnor U6468 (N_6468,N_5530,N_5410);
or U6469 (N_6469,N_5518,N_5953);
and U6470 (N_6470,N_5510,N_5652);
xnor U6471 (N_6471,N_5236,N_5311);
nand U6472 (N_6472,N_5812,N_5505);
nor U6473 (N_6473,N_5910,N_5984);
nand U6474 (N_6474,N_5768,N_5104);
nor U6475 (N_6475,N_5622,N_5262);
xor U6476 (N_6476,N_5677,N_5360);
xor U6477 (N_6477,N_5447,N_5985);
nor U6478 (N_6478,N_5135,N_5397);
or U6479 (N_6479,N_5815,N_5075);
or U6480 (N_6480,N_5482,N_5485);
nor U6481 (N_6481,N_5617,N_5284);
and U6482 (N_6482,N_5681,N_5662);
or U6483 (N_6483,N_5594,N_5523);
or U6484 (N_6484,N_5044,N_5157);
nand U6485 (N_6485,N_5995,N_5877);
nand U6486 (N_6486,N_5881,N_5175);
nand U6487 (N_6487,N_5927,N_5255);
and U6488 (N_6488,N_5614,N_5656);
nor U6489 (N_6489,N_5072,N_5882);
nor U6490 (N_6490,N_5214,N_5483);
and U6491 (N_6491,N_5587,N_5361);
or U6492 (N_6492,N_5332,N_5672);
xor U6493 (N_6493,N_5379,N_5955);
or U6494 (N_6494,N_5926,N_5419);
and U6495 (N_6495,N_5949,N_5197);
nand U6496 (N_6496,N_5456,N_5319);
nand U6497 (N_6497,N_5641,N_5357);
and U6498 (N_6498,N_5393,N_5716);
and U6499 (N_6499,N_5865,N_5562);
nor U6500 (N_6500,N_5523,N_5713);
xnor U6501 (N_6501,N_5041,N_5425);
and U6502 (N_6502,N_5680,N_5938);
nor U6503 (N_6503,N_5819,N_5583);
and U6504 (N_6504,N_5359,N_5707);
nor U6505 (N_6505,N_5765,N_5588);
xnor U6506 (N_6506,N_5112,N_5502);
and U6507 (N_6507,N_5926,N_5574);
nor U6508 (N_6508,N_5713,N_5426);
xnor U6509 (N_6509,N_5112,N_5275);
nor U6510 (N_6510,N_5052,N_5003);
nor U6511 (N_6511,N_5884,N_5303);
xnor U6512 (N_6512,N_5246,N_5709);
and U6513 (N_6513,N_5717,N_5758);
nand U6514 (N_6514,N_5050,N_5925);
xnor U6515 (N_6515,N_5236,N_5879);
nand U6516 (N_6516,N_5030,N_5371);
and U6517 (N_6517,N_5560,N_5319);
and U6518 (N_6518,N_5815,N_5581);
nor U6519 (N_6519,N_5028,N_5749);
and U6520 (N_6520,N_5032,N_5299);
nor U6521 (N_6521,N_5416,N_5399);
or U6522 (N_6522,N_5088,N_5595);
nor U6523 (N_6523,N_5393,N_5286);
and U6524 (N_6524,N_5799,N_5904);
xor U6525 (N_6525,N_5177,N_5772);
or U6526 (N_6526,N_5880,N_5021);
and U6527 (N_6527,N_5349,N_5223);
and U6528 (N_6528,N_5359,N_5703);
and U6529 (N_6529,N_5192,N_5795);
and U6530 (N_6530,N_5798,N_5180);
nand U6531 (N_6531,N_5985,N_5113);
and U6532 (N_6532,N_5026,N_5718);
and U6533 (N_6533,N_5392,N_5518);
or U6534 (N_6534,N_5434,N_5241);
nand U6535 (N_6535,N_5039,N_5632);
or U6536 (N_6536,N_5068,N_5712);
nand U6537 (N_6537,N_5332,N_5751);
or U6538 (N_6538,N_5991,N_5800);
and U6539 (N_6539,N_5178,N_5346);
nand U6540 (N_6540,N_5415,N_5938);
nand U6541 (N_6541,N_5560,N_5114);
nor U6542 (N_6542,N_5653,N_5135);
xor U6543 (N_6543,N_5146,N_5539);
nor U6544 (N_6544,N_5012,N_5503);
and U6545 (N_6545,N_5430,N_5883);
or U6546 (N_6546,N_5482,N_5579);
nand U6547 (N_6547,N_5235,N_5193);
and U6548 (N_6548,N_5800,N_5436);
nand U6549 (N_6549,N_5132,N_5988);
or U6550 (N_6550,N_5681,N_5020);
nand U6551 (N_6551,N_5215,N_5135);
or U6552 (N_6552,N_5815,N_5206);
and U6553 (N_6553,N_5468,N_5574);
nand U6554 (N_6554,N_5155,N_5714);
and U6555 (N_6555,N_5407,N_5378);
nand U6556 (N_6556,N_5611,N_5887);
nor U6557 (N_6557,N_5097,N_5563);
and U6558 (N_6558,N_5704,N_5224);
xnor U6559 (N_6559,N_5205,N_5884);
and U6560 (N_6560,N_5220,N_5210);
or U6561 (N_6561,N_5858,N_5700);
or U6562 (N_6562,N_5641,N_5556);
and U6563 (N_6563,N_5978,N_5873);
xnor U6564 (N_6564,N_5821,N_5462);
nand U6565 (N_6565,N_5027,N_5365);
nand U6566 (N_6566,N_5537,N_5606);
and U6567 (N_6567,N_5716,N_5876);
or U6568 (N_6568,N_5282,N_5710);
xnor U6569 (N_6569,N_5834,N_5476);
and U6570 (N_6570,N_5140,N_5901);
nand U6571 (N_6571,N_5565,N_5912);
and U6572 (N_6572,N_5450,N_5183);
or U6573 (N_6573,N_5983,N_5437);
and U6574 (N_6574,N_5262,N_5648);
xnor U6575 (N_6575,N_5830,N_5516);
and U6576 (N_6576,N_5350,N_5752);
or U6577 (N_6577,N_5640,N_5108);
and U6578 (N_6578,N_5185,N_5890);
and U6579 (N_6579,N_5381,N_5212);
xnor U6580 (N_6580,N_5886,N_5336);
xnor U6581 (N_6581,N_5939,N_5997);
xor U6582 (N_6582,N_5963,N_5166);
xor U6583 (N_6583,N_5520,N_5811);
xnor U6584 (N_6584,N_5251,N_5854);
nand U6585 (N_6585,N_5714,N_5372);
xnor U6586 (N_6586,N_5293,N_5237);
or U6587 (N_6587,N_5174,N_5123);
and U6588 (N_6588,N_5863,N_5855);
nand U6589 (N_6589,N_5187,N_5742);
nand U6590 (N_6590,N_5950,N_5418);
or U6591 (N_6591,N_5427,N_5610);
or U6592 (N_6592,N_5957,N_5726);
or U6593 (N_6593,N_5142,N_5834);
and U6594 (N_6594,N_5075,N_5885);
nand U6595 (N_6595,N_5763,N_5881);
or U6596 (N_6596,N_5269,N_5369);
nand U6597 (N_6597,N_5330,N_5649);
and U6598 (N_6598,N_5254,N_5099);
or U6599 (N_6599,N_5255,N_5143);
and U6600 (N_6600,N_5782,N_5338);
nand U6601 (N_6601,N_5215,N_5542);
or U6602 (N_6602,N_5672,N_5817);
nand U6603 (N_6603,N_5134,N_5079);
xnor U6604 (N_6604,N_5251,N_5652);
nand U6605 (N_6605,N_5047,N_5684);
nand U6606 (N_6606,N_5477,N_5603);
and U6607 (N_6607,N_5572,N_5749);
xnor U6608 (N_6608,N_5360,N_5991);
xor U6609 (N_6609,N_5558,N_5750);
xor U6610 (N_6610,N_5137,N_5096);
and U6611 (N_6611,N_5875,N_5950);
nand U6612 (N_6612,N_5622,N_5892);
nand U6613 (N_6613,N_5807,N_5085);
nor U6614 (N_6614,N_5121,N_5851);
or U6615 (N_6615,N_5445,N_5063);
and U6616 (N_6616,N_5150,N_5978);
xnor U6617 (N_6617,N_5601,N_5655);
nand U6618 (N_6618,N_5652,N_5744);
and U6619 (N_6619,N_5327,N_5822);
nand U6620 (N_6620,N_5357,N_5073);
xnor U6621 (N_6621,N_5367,N_5172);
and U6622 (N_6622,N_5318,N_5218);
nand U6623 (N_6623,N_5767,N_5133);
and U6624 (N_6624,N_5173,N_5531);
nor U6625 (N_6625,N_5751,N_5398);
or U6626 (N_6626,N_5468,N_5716);
and U6627 (N_6627,N_5674,N_5208);
xor U6628 (N_6628,N_5938,N_5903);
xnor U6629 (N_6629,N_5266,N_5767);
and U6630 (N_6630,N_5045,N_5439);
and U6631 (N_6631,N_5458,N_5226);
or U6632 (N_6632,N_5414,N_5342);
xnor U6633 (N_6633,N_5938,N_5674);
xor U6634 (N_6634,N_5615,N_5512);
xor U6635 (N_6635,N_5408,N_5218);
xnor U6636 (N_6636,N_5404,N_5234);
or U6637 (N_6637,N_5371,N_5943);
or U6638 (N_6638,N_5028,N_5151);
nor U6639 (N_6639,N_5425,N_5016);
nor U6640 (N_6640,N_5188,N_5677);
and U6641 (N_6641,N_5265,N_5671);
or U6642 (N_6642,N_5138,N_5808);
xor U6643 (N_6643,N_5190,N_5095);
nand U6644 (N_6644,N_5755,N_5083);
and U6645 (N_6645,N_5272,N_5702);
nand U6646 (N_6646,N_5880,N_5451);
or U6647 (N_6647,N_5648,N_5979);
or U6648 (N_6648,N_5989,N_5300);
or U6649 (N_6649,N_5235,N_5890);
nand U6650 (N_6650,N_5381,N_5688);
xor U6651 (N_6651,N_5789,N_5032);
nor U6652 (N_6652,N_5643,N_5359);
and U6653 (N_6653,N_5368,N_5892);
or U6654 (N_6654,N_5715,N_5229);
nand U6655 (N_6655,N_5926,N_5181);
nor U6656 (N_6656,N_5724,N_5799);
nor U6657 (N_6657,N_5223,N_5189);
or U6658 (N_6658,N_5840,N_5168);
nor U6659 (N_6659,N_5555,N_5255);
and U6660 (N_6660,N_5098,N_5067);
xnor U6661 (N_6661,N_5675,N_5130);
nand U6662 (N_6662,N_5230,N_5173);
nor U6663 (N_6663,N_5703,N_5354);
nor U6664 (N_6664,N_5904,N_5195);
nor U6665 (N_6665,N_5866,N_5296);
xor U6666 (N_6666,N_5032,N_5324);
nor U6667 (N_6667,N_5410,N_5079);
nor U6668 (N_6668,N_5559,N_5827);
and U6669 (N_6669,N_5605,N_5511);
and U6670 (N_6670,N_5780,N_5072);
xor U6671 (N_6671,N_5339,N_5268);
nor U6672 (N_6672,N_5160,N_5129);
nor U6673 (N_6673,N_5829,N_5862);
or U6674 (N_6674,N_5570,N_5334);
nor U6675 (N_6675,N_5421,N_5892);
or U6676 (N_6676,N_5212,N_5070);
nand U6677 (N_6677,N_5487,N_5885);
and U6678 (N_6678,N_5807,N_5524);
nand U6679 (N_6679,N_5147,N_5837);
xor U6680 (N_6680,N_5709,N_5070);
xnor U6681 (N_6681,N_5051,N_5181);
nor U6682 (N_6682,N_5082,N_5009);
and U6683 (N_6683,N_5959,N_5850);
and U6684 (N_6684,N_5848,N_5953);
nand U6685 (N_6685,N_5418,N_5027);
xnor U6686 (N_6686,N_5029,N_5762);
or U6687 (N_6687,N_5030,N_5785);
or U6688 (N_6688,N_5059,N_5317);
nand U6689 (N_6689,N_5800,N_5503);
xnor U6690 (N_6690,N_5260,N_5788);
and U6691 (N_6691,N_5279,N_5863);
nor U6692 (N_6692,N_5138,N_5689);
or U6693 (N_6693,N_5616,N_5381);
or U6694 (N_6694,N_5122,N_5872);
nand U6695 (N_6695,N_5922,N_5235);
nand U6696 (N_6696,N_5872,N_5715);
or U6697 (N_6697,N_5707,N_5741);
nor U6698 (N_6698,N_5388,N_5274);
xnor U6699 (N_6699,N_5478,N_5232);
and U6700 (N_6700,N_5226,N_5093);
and U6701 (N_6701,N_5253,N_5258);
xor U6702 (N_6702,N_5314,N_5993);
nand U6703 (N_6703,N_5255,N_5528);
or U6704 (N_6704,N_5583,N_5030);
or U6705 (N_6705,N_5892,N_5182);
nand U6706 (N_6706,N_5684,N_5994);
nor U6707 (N_6707,N_5807,N_5028);
nor U6708 (N_6708,N_5783,N_5469);
nand U6709 (N_6709,N_5218,N_5834);
and U6710 (N_6710,N_5748,N_5835);
nor U6711 (N_6711,N_5077,N_5069);
nand U6712 (N_6712,N_5447,N_5402);
nand U6713 (N_6713,N_5876,N_5522);
nand U6714 (N_6714,N_5768,N_5644);
nand U6715 (N_6715,N_5050,N_5512);
and U6716 (N_6716,N_5659,N_5474);
nand U6717 (N_6717,N_5002,N_5544);
or U6718 (N_6718,N_5562,N_5176);
xnor U6719 (N_6719,N_5721,N_5392);
nor U6720 (N_6720,N_5947,N_5865);
or U6721 (N_6721,N_5295,N_5518);
or U6722 (N_6722,N_5641,N_5874);
nor U6723 (N_6723,N_5503,N_5038);
and U6724 (N_6724,N_5233,N_5626);
or U6725 (N_6725,N_5349,N_5817);
nor U6726 (N_6726,N_5325,N_5151);
nand U6727 (N_6727,N_5649,N_5843);
xnor U6728 (N_6728,N_5632,N_5685);
xnor U6729 (N_6729,N_5610,N_5933);
nand U6730 (N_6730,N_5274,N_5969);
xor U6731 (N_6731,N_5983,N_5127);
and U6732 (N_6732,N_5007,N_5211);
nor U6733 (N_6733,N_5695,N_5326);
and U6734 (N_6734,N_5007,N_5891);
or U6735 (N_6735,N_5749,N_5458);
or U6736 (N_6736,N_5903,N_5062);
and U6737 (N_6737,N_5090,N_5471);
and U6738 (N_6738,N_5374,N_5918);
or U6739 (N_6739,N_5445,N_5044);
nor U6740 (N_6740,N_5562,N_5697);
nand U6741 (N_6741,N_5525,N_5166);
nor U6742 (N_6742,N_5332,N_5138);
xor U6743 (N_6743,N_5089,N_5744);
nor U6744 (N_6744,N_5063,N_5323);
nor U6745 (N_6745,N_5803,N_5683);
or U6746 (N_6746,N_5052,N_5226);
nor U6747 (N_6747,N_5102,N_5590);
nand U6748 (N_6748,N_5038,N_5943);
nor U6749 (N_6749,N_5707,N_5713);
nor U6750 (N_6750,N_5924,N_5511);
and U6751 (N_6751,N_5457,N_5042);
nor U6752 (N_6752,N_5879,N_5301);
nand U6753 (N_6753,N_5688,N_5557);
and U6754 (N_6754,N_5613,N_5797);
and U6755 (N_6755,N_5234,N_5167);
xor U6756 (N_6756,N_5241,N_5205);
or U6757 (N_6757,N_5389,N_5649);
or U6758 (N_6758,N_5770,N_5982);
and U6759 (N_6759,N_5365,N_5570);
or U6760 (N_6760,N_5921,N_5789);
or U6761 (N_6761,N_5423,N_5123);
nand U6762 (N_6762,N_5155,N_5278);
xnor U6763 (N_6763,N_5772,N_5076);
xor U6764 (N_6764,N_5355,N_5353);
xor U6765 (N_6765,N_5057,N_5828);
and U6766 (N_6766,N_5237,N_5466);
nor U6767 (N_6767,N_5997,N_5580);
and U6768 (N_6768,N_5648,N_5493);
nand U6769 (N_6769,N_5793,N_5075);
nor U6770 (N_6770,N_5993,N_5441);
nor U6771 (N_6771,N_5663,N_5276);
or U6772 (N_6772,N_5523,N_5667);
and U6773 (N_6773,N_5019,N_5494);
or U6774 (N_6774,N_5731,N_5197);
nor U6775 (N_6775,N_5039,N_5115);
nor U6776 (N_6776,N_5115,N_5945);
and U6777 (N_6777,N_5887,N_5465);
nand U6778 (N_6778,N_5706,N_5761);
or U6779 (N_6779,N_5895,N_5684);
and U6780 (N_6780,N_5327,N_5345);
and U6781 (N_6781,N_5831,N_5236);
xnor U6782 (N_6782,N_5407,N_5056);
or U6783 (N_6783,N_5623,N_5944);
and U6784 (N_6784,N_5626,N_5065);
or U6785 (N_6785,N_5052,N_5765);
xor U6786 (N_6786,N_5993,N_5753);
and U6787 (N_6787,N_5353,N_5891);
and U6788 (N_6788,N_5990,N_5655);
and U6789 (N_6789,N_5883,N_5979);
nor U6790 (N_6790,N_5136,N_5533);
nand U6791 (N_6791,N_5849,N_5766);
and U6792 (N_6792,N_5182,N_5831);
nand U6793 (N_6793,N_5744,N_5255);
or U6794 (N_6794,N_5276,N_5801);
and U6795 (N_6795,N_5580,N_5641);
nand U6796 (N_6796,N_5474,N_5230);
xor U6797 (N_6797,N_5978,N_5908);
and U6798 (N_6798,N_5357,N_5444);
xnor U6799 (N_6799,N_5793,N_5487);
nor U6800 (N_6800,N_5582,N_5310);
and U6801 (N_6801,N_5865,N_5976);
or U6802 (N_6802,N_5135,N_5500);
xnor U6803 (N_6803,N_5912,N_5822);
nand U6804 (N_6804,N_5138,N_5412);
nor U6805 (N_6805,N_5322,N_5540);
nor U6806 (N_6806,N_5565,N_5905);
nor U6807 (N_6807,N_5536,N_5973);
nand U6808 (N_6808,N_5208,N_5617);
nor U6809 (N_6809,N_5467,N_5007);
and U6810 (N_6810,N_5701,N_5642);
xor U6811 (N_6811,N_5158,N_5068);
nand U6812 (N_6812,N_5634,N_5815);
nand U6813 (N_6813,N_5152,N_5816);
and U6814 (N_6814,N_5003,N_5573);
nand U6815 (N_6815,N_5685,N_5983);
or U6816 (N_6816,N_5755,N_5495);
nor U6817 (N_6817,N_5926,N_5995);
nand U6818 (N_6818,N_5626,N_5528);
xnor U6819 (N_6819,N_5304,N_5992);
and U6820 (N_6820,N_5291,N_5358);
or U6821 (N_6821,N_5039,N_5694);
nand U6822 (N_6822,N_5910,N_5364);
and U6823 (N_6823,N_5506,N_5722);
nand U6824 (N_6824,N_5378,N_5770);
and U6825 (N_6825,N_5173,N_5353);
nand U6826 (N_6826,N_5488,N_5454);
or U6827 (N_6827,N_5891,N_5197);
nand U6828 (N_6828,N_5628,N_5952);
or U6829 (N_6829,N_5834,N_5180);
and U6830 (N_6830,N_5753,N_5451);
xnor U6831 (N_6831,N_5111,N_5344);
nor U6832 (N_6832,N_5650,N_5443);
and U6833 (N_6833,N_5497,N_5955);
or U6834 (N_6834,N_5988,N_5230);
nand U6835 (N_6835,N_5096,N_5170);
xor U6836 (N_6836,N_5397,N_5264);
and U6837 (N_6837,N_5761,N_5470);
nor U6838 (N_6838,N_5701,N_5041);
nand U6839 (N_6839,N_5838,N_5165);
xnor U6840 (N_6840,N_5461,N_5767);
nor U6841 (N_6841,N_5661,N_5422);
nand U6842 (N_6842,N_5897,N_5573);
nand U6843 (N_6843,N_5149,N_5689);
or U6844 (N_6844,N_5654,N_5888);
or U6845 (N_6845,N_5403,N_5862);
xor U6846 (N_6846,N_5266,N_5158);
xor U6847 (N_6847,N_5379,N_5752);
and U6848 (N_6848,N_5377,N_5444);
xor U6849 (N_6849,N_5262,N_5428);
or U6850 (N_6850,N_5682,N_5822);
and U6851 (N_6851,N_5291,N_5544);
and U6852 (N_6852,N_5267,N_5130);
and U6853 (N_6853,N_5068,N_5882);
nor U6854 (N_6854,N_5890,N_5918);
nor U6855 (N_6855,N_5763,N_5043);
or U6856 (N_6856,N_5890,N_5664);
nand U6857 (N_6857,N_5511,N_5206);
or U6858 (N_6858,N_5553,N_5325);
xor U6859 (N_6859,N_5738,N_5244);
nand U6860 (N_6860,N_5758,N_5984);
xor U6861 (N_6861,N_5408,N_5258);
nand U6862 (N_6862,N_5698,N_5699);
xor U6863 (N_6863,N_5068,N_5073);
xnor U6864 (N_6864,N_5007,N_5440);
and U6865 (N_6865,N_5199,N_5042);
or U6866 (N_6866,N_5488,N_5622);
nand U6867 (N_6867,N_5953,N_5227);
nor U6868 (N_6868,N_5274,N_5942);
nor U6869 (N_6869,N_5464,N_5220);
and U6870 (N_6870,N_5377,N_5702);
xor U6871 (N_6871,N_5862,N_5379);
or U6872 (N_6872,N_5471,N_5388);
nand U6873 (N_6873,N_5537,N_5933);
nor U6874 (N_6874,N_5151,N_5114);
nor U6875 (N_6875,N_5088,N_5070);
nand U6876 (N_6876,N_5478,N_5339);
or U6877 (N_6877,N_5807,N_5383);
and U6878 (N_6878,N_5551,N_5693);
xnor U6879 (N_6879,N_5519,N_5050);
and U6880 (N_6880,N_5626,N_5875);
xor U6881 (N_6881,N_5972,N_5295);
and U6882 (N_6882,N_5221,N_5475);
and U6883 (N_6883,N_5246,N_5886);
nand U6884 (N_6884,N_5213,N_5300);
and U6885 (N_6885,N_5244,N_5737);
and U6886 (N_6886,N_5614,N_5208);
nand U6887 (N_6887,N_5311,N_5281);
nand U6888 (N_6888,N_5773,N_5116);
and U6889 (N_6889,N_5062,N_5392);
or U6890 (N_6890,N_5128,N_5498);
or U6891 (N_6891,N_5123,N_5201);
or U6892 (N_6892,N_5402,N_5654);
nand U6893 (N_6893,N_5156,N_5640);
xor U6894 (N_6894,N_5967,N_5038);
nor U6895 (N_6895,N_5449,N_5890);
and U6896 (N_6896,N_5885,N_5536);
nor U6897 (N_6897,N_5590,N_5625);
nor U6898 (N_6898,N_5147,N_5632);
or U6899 (N_6899,N_5733,N_5464);
or U6900 (N_6900,N_5778,N_5043);
or U6901 (N_6901,N_5964,N_5864);
or U6902 (N_6902,N_5100,N_5131);
or U6903 (N_6903,N_5214,N_5071);
or U6904 (N_6904,N_5785,N_5675);
and U6905 (N_6905,N_5988,N_5774);
and U6906 (N_6906,N_5903,N_5248);
and U6907 (N_6907,N_5288,N_5410);
and U6908 (N_6908,N_5801,N_5525);
or U6909 (N_6909,N_5040,N_5376);
and U6910 (N_6910,N_5631,N_5903);
or U6911 (N_6911,N_5494,N_5161);
or U6912 (N_6912,N_5286,N_5287);
and U6913 (N_6913,N_5807,N_5913);
or U6914 (N_6914,N_5377,N_5827);
nor U6915 (N_6915,N_5286,N_5542);
or U6916 (N_6916,N_5138,N_5765);
nand U6917 (N_6917,N_5625,N_5112);
nand U6918 (N_6918,N_5058,N_5572);
and U6919 (N_6919,N_5720,N_5631);
and U6920 (N_6920,N_5625,N_5039);
or U6921 (N_6921,N_5773,N_5034);
or U6922 (N_6922,N_5823,N_5746);
xnor U6923 (N_6923,N_5824,N_5994);
or U6924 (N_6924,N_5608,N_5632);
xnor U6925 (N_6925,N_5588,N_5429);
nand U6926 (N_6926,N_5646,N_5708);
or U6927 (N_6927,N_5890,N_5662);
and U6928 (N_6928,N_5464,N_5215);
nand U6929 (N_6929,N_5230,N_5516);
xnor U6930 (N_6930,N_5047,N_5111);
nor U6931 (N_6931,N_5766,N_5874);
and U6932 (N_6932,N_5970,N_5469);
or U6933 (N_6933,N_5595,N_5554);
xnor U6934 (N_6934,N_5844,N_5058);
xnor U6935 (N_6935,N_5180,N_5790);
nand U6936 (N_6936,N_5544,N_5256);
nor U6937 (N_6937,N_5778,N_5229);
or U6938 (N_6938,N_5011,N_5589);
and U6939 (N_6939,N_5824,N_5843);
or U6940 (N_6940,N_5929,N_5405);
and U6941 (N_6941,N_5245,N_5539);
and U6942 (N_6942,N_5726,N_5780);
nand U6943 (N_6943,N_5433,N_5711);
or U6944 (N_6944,N_5994,N_5606);
or U6945 (N_6945,N_5497,N_5922);
or U6946 (N_6946,N_5922,N_5729);
nor U6947 (N_6947,N_5486,N_5248);
or U6948 (N_6948,N_5369,N_5834);
nor U6949 (N_6949,N_5160,N_5788);
nand U6950 (N_6950,N_5041,N_5025);
nor U6951 (N_6951,N_5134,N_5766);
xnor U6952 (N_6952,N_5109,N_5323);
or U6953 (N_6953,N_5858,N_5576);
or U6954 (N_6954,N_5046,N_5303);
or U6955 (N_6955,N_5346,N_5239);
and U6956 (N_6956,N_5053,N_5307);
and U6957 (N_6957,N_5457,N_5659);
and U6958 (N_6958,N_5753,N_5810);
or U6959 (N_6959,N_5476,N_5671);
and U6960 (N_6960,N_5183,N_5243);
nand U6961 (N_6961,N_5076,N_5338);
and U6962 (N_6962,N_5848,N_5400);
or U6963 (N_6963,N_5680,N_5856);
nor U6964 (N_6964,N_5035,N_5723);
xnor U6965 (N_6965,N_5188,N_5844);
xnor U6966 (N_6966,N_5471,N_5249);
xor U6967 (N_6967,N_5234,N_5611);
nor U6968 (N_6968,N_5802,N_5102);
nand U6969 (N_6969,N_5541,N_5028);
xor U6970 (N_6970,N_5241,N_5773);
nor U6971 (N_6971,N_5915,N_5677);
and U6972 (N_6972,N_5398,N_5462);
nor U6973 (N_6973,N_5764,N_5623);
or U6974 (N_6974,N_5517,N_5863);
nand U6975 (N_6975,N_5008,N_5203);
or U6976 (N_6976,N_5676,N_5290);
xnor U6977 (N_6977,N_5603,N_5359);
and U6978 (N_6978,N_5851,N_5962);
and U6979 (N_6979,N_5576,N_5212);
nor U6980 (N_6980,N_5837,N_5090);
nor U6981 (N_6981,N_5229,N_5194);
nand U6982 (N_6982,N_5550,N_5983);
and U6983 (N_6983,N_5566,N_5422);
xor U6984 (N_6984,N_5393,N_5463);
nor U6985 (N_6985,N_5639,N_5575);
or U6986 (N_6986,N_5589,N_5493);
or U6987 (N_6987,N_5035,N_5576);
or U6988 (N_6988,N_5947,N_5842);
and U6989 (N_6989,N_5044,N_5394);
xnor U6990 (N_6990,N_5685,N_5430);
and U6991 (N_6991,N_5581,N_5752);
or U6992 (N_6992,N_5027,N_5353);
nor U6993 (N_6993,N_5168,N_5125);
or U6994 (N_6994,N_5963,N_5852);
xnor U6995 (N_6995,N_5776,N_5961);
nand U6996 (N_6996,N_5677,N_5536);
xor U6997 (N_6997,N_5053,N_5043);
and U6998 (N_6998,N_5452,N_5471);
nor U6999 (N_6999,N_5541,N_5819);
nor U7000 (N_7000,N_6530,N_6727);
or U7001 (N_7001,N_6301,N_6488);
nand U7002 (N_7002,N_6554,N_6533);
nor U7003 (N_7003,N_6775,N_6949);
xnor U7004 (N_7004,N_6563,N_6784);
nand U7005 (N_7005,N_6284,N_6306);
xor U7006 (N_7006,N_6996,N_6174);
xor U7007 (N_7007,N_6462,N_6670);
and U7008 (N_7008,N_6819,N_6092);
nor U7009 (N_7009,N_6211,N_6397);
or U7010 (N_7010,N_6409,N_6372);
xnor U7011 (N_7011,N_6641,N_6071);
and U7012 (N_7012,N_6149,N_6009);
or U7013 (N_7013,N_6401,N_6171);
nand U7014 (N_7014,N_6667,N_6357);
and U7015 (N_7015,N_6540,N_6853);
nand U7016 (N_7016,N_6236,N_6014);
nor U7017 (N_7017,N_6490,N_6651);
nand U7018 (N_7018,N_6606,N_6801);
nand U7019 (N_7019,N_6466,N_6732);
nand U7020 (N_7020,N_6035,N_6843);
and U7021 (N_7021,N_6820,N_6421);
nand U7022 (N_7022,N_6591,N_6779);
nor U7023 (N_7023,N_6386,N_6717);
or U7024 (N_7024,N_6756,N_6638);
xnor U7025 (N_7025,N_6525,N_6439);
nand U7026 (N_7026,N_6055,N_6322);
xor U7027 (N_7027,N_6643,N_6628);
and U7028 (N_7028,N_6391,N_6312);
nor U7029 (N_7029,N_6358,N_6511);
nor U7030 (N_7030,N_6550,N_6851);
nand U7031 (N_7031,N_6923,N_6152);
and U7032 (N_7032,N_6025,N_6362);
nand U7033 (N_7033,N_6690,N_6749);
nand U7034 (N_7034,N_6209,N_6581);
nand U7035 (N_7035,N_6895,N_6399);
xnor U7036 (N_7036,N_6430,N_6065);
xnor U7037 (N_7037,N_6745,N_6835);
or U7038 (N_7038,N_6267,N_6995);
and U7039 (N_7039,N_6791,N_6256);
nand U7040 (N_7040,N_6087,N_6221);
nand U7041 (N_7041,N_6882,N_6771);
xor U7042 (N_7042,N_6596,N_6645);
nand U7043 (N_7043,N_6451,N_6164);
nand U7044 (N_7044,N_6038,N_6860);
and U7045 (N_7045,N_6299,N_6766);
nand U7046 (N_7046,N_6828,N_6498);
nand U7047 (N_7047,N_6868,N_6004);
xnor U7048 (N_7048,N_6226,N_6751);
xnor U7049 (N_7049,N_6443,N_6750);
nor U7050 (N_7050,N_6273,N_6519);
xnor U7051 (N_7051,N_6185,N_6684);
and U7052 (N_7052,N_6176,N_6257);
or U7053 (N_7053,N_6547,N_6634);
nor U7054 (N_7054,N_6869,N_6531);
and U7055 (N_7055,N_6286,N_6011);
nor U7056 (N_7056,N_6348,N_6313);
nor U7057 (N_7057,N_6140,N_6197);
nand U7058 (N_7058,N_6944,N_6826);
and U7059 (N_7059,N_6818,N_6405);
nand U7060 (N_7060,N_6376,N_6446);
nor U7061 (N_7061,N_6161,N_6030);
or U7062 (N_7062,N_6447,N_6798);
nor U7063 (N_7063,N_6107,N_6415);
and U7064 (N_7064,N_6241,N_6005);
or U7065 (N_7065,N_6668,N_6746);
xor U7066 (N_7066,N_6237,N_6700);
nand U7067 (N_7067,N_6911,N_6761);
nor U7068 (N_7068,N_6617,N_6821);
and U7069 (N_7069,N_6551,N_6037);
xor U7070 (N_7070,N_6184,N_6253);
nand U7071 (N_7071,N_6747,N_6235);
xor U7072 (N_7072,N_6469,N_6876);
nor U7073 (N_7073,N_6827,N_6106);
and U7074 (N_7074,N_6958,N_6546);
nor U7075 (N_7075,N_6935,N_6527);
and U7076 (N_7076,N_6537,N_6752);
xor U7077 (N_7077,N_6767,N_6514);
nand U7078 (N_7078,N_6859,N_6977);
and U7079 (N_7079,N_6001,N_6637);
and U7080 (N_7080,N_6042,N_6815);
and U7081 (N_7081,N_6223,N_6658);
or U7082 (N_7082,N_6941,N_6100);
and U7083 (N_7083,N_6134,N_6111);
nand U7084 (N_7084,N_6742,N_6532);
xnor U7085 (N_7085,N_6189,N_6660);
nor U7086 (N_7086,N_6763,N_6353);
nand U7087 (N_7087,N_6325,N_6769);
and U7088 (N_7088,N_6308,N_6806);
and U7089 (N_7089,N_6109,N_6057);
nand U7090 (N_7090,N_6889,N_6683);
nand U7091 (N_7091,N_6167,N_6865);
or U7092 (N_7092,N_6458,N_6148);
nand U7093 (N_7093,N_6179,N_6154);
or U7094 (N_7094,N_6794,N_6852);
nor U7095 (N_7095,N_6957,N_6328);
or U7096 (N_7096,N_6604,N_6493);
or U7097 (N_7097,N_6268,N_6847);
nand U7098 (N_7098,N_6654,N_6385);
xnor U7099 (N_7099,N_6034,N_6981);
and U7100 (N_7100,N_6233,N_6564);
and U7101 (N_7101,N_6665,N_6925);
nand U7102 (N_7102,N_6311,N_6371);
nand U7103 (N_7103,N_6561,N_6460);
or U7104 (N_7104,N_6661,N_6411);
nor U7105 (N_7105,N_6496,N_6455);
and U7106 (N_7106,N_6983,N_6433);
xor U7107 (N_7107,N_6390,N_6129);
or U7108 (N_7108,N_6016,N_6196);
xnor U7109 (N_7109,N_6465,N_6762);
and U7110 (N_7110,N_6934,N_6612);
nand U7111 (N_7111,N_6029,N_6543);
xor U7112 (N_7112,N_6445,N_6053);
xor U7113 (N_7113,N_6679,N_6225);
and U7114 (N_7114,N_6010,N_6568);
nand U7115 (N_7115,N_6374,N_6516);
and U7116 (N_7116,N_6017,N_6317);
nor U7117 (N_7117,N_6698,N_6248);
nand U7118 (N_7118,N_6373,N_6126);
or U7119 (N_7119,N_6359,N_6146);
and U7120 (N_7120,N_6259,N_6985);
and U7121 (N_7121,N_6406,N_6553);
xnor U7122 (N_7122,N_6410,N_6491);
nor U7123 (N_7123,N_6922,N_6292);
and U7124 (N_7124,N_6020,N_6930);
xor U7125 (N_7125,N_6015,N_6989);
and U7126 (N_7126,N_6040,N_6250);
or U7127 (N_7127,N_6846,N_6157);
nor U7128 (N_7128,N_6125,N_6902);
and U7129 (N_7129,N_6862,N_6370);
xnor U7130 (N_7130,N_6836,N_6249);
nand U7131 (N_7131,N_6731,N_6091);
nor U7132 (N_7132,N_6730,N_6408);
or U7133 (N_7133,N_6621,N_6105);
nand U7134 (N_7134,N_6816,N_6694);
nor U7135 (N_7135,N_6890,N_6168);
and U7136 (N_7136,N_6444,N_6610);
or U7137 (N_7137,N_6150,N_6291);
xnor U7138 (N_7138,N_6090,N_6018);
nor U7139 (N_7139,N_6441,N_6201);
and U7140 (N_7140,N_6597,N_6897);
and U7141 (N_7141,N_6394,N_6419);
and U7142 (N_7142,N_6512,N_6266);
xor U7143 (N_7143,N_6175,N_6672);
xnor U7144 (N_7144,N_6518,N_6337);
or U7145 (N_7145,N_6738,N_6630);
nor U7146 (N_7146,N_6000,N_6669);
nand U7147 (N_7147,N_6973,N_6601);
xnor U7148 (N_7148,N_6243,N_6497);
nor U7149 (N_7149,N_6510,N_6432);
xnor U7150 (N_7150,N_6471,N_6422);
and U7151 (N_7151,N_6287,N_6653);
xnor U7152 (N_7152,N_6191,N_6802);
or U7153 (N_7153,N_6829,N_6160);
nand U7154 (N_7154,N_6319,N_6577);
nand U7155 (N_7155,N_6692,N_6470);
nand U7156 (N_7156,N_6813,N_6127);
or U7157 (N_7157,N_6954,N_6968);
and U7158 (N_7158,N_6593,N_6208);
nor U7159 (N_7159,N_6704,N_6842);
and U7160 (N_7160,N_6137,N_6324);
nor U7161 (N_7161,N_6217,N_6457);
and U7162 (N_7162,N_6162,N_6392);
and U7163 (N_7163,N_6461,N_6307);
nand U7164 (N_7164,N_6420,N_6494);
nand U7165 (N_7165,N_6896,N_6887);
xnor U7166 (N_7166,N_6332,N_6521);
or U7167 (N_7167,N_6875,N_6567);
xnor U7168 (N_7168,N_6986,N_6541);
and U7169 (N_7169,N_6863,N_6294);
or U7170 (N_7170,N_6964,N_6356);
and U7171 (N_7171,N_6327,N_6335);
xnor U7172 (N_7172,N_6585,N_6783);
or U7173 (N_7173,N_6913,N_6407);
nand U7174 (N_7174,N_6528,N_6759);
and U7175 (N_7175,N_6900,N_6023);
nand U7176 (N_7176,N_6620,N_6073);
or U7177 (N_7177,N_6720,N_6382);
xnor U7178 (N_7178,N_6123,N_6500);
and U7179 (N_7179,N_6753,N_6713);
nand U7180 (N_7180,N_6442,N_6387);
xor U7181 (N_7181,N_6579,N_6060);
or U7182 (N_7182,N_6832,N_6970);
nand U7183 (N_7183,N_6603,N_6426);
nand U7184 (N_7184,N_6288,N_6793);
xor U7185 (N_7185,N_6198,N_6960);
nor U7186 (N_7186,N_6141,N_6706);
nand U7187 (N_7187,N_6377,N_6424);
nor U7188 (N_7188,N_6515,N_6027);
or U7189 (N_7189,N_6962,N_6271);
and U7190 (N_7190,N_6166,N_6790);
xnor U7191 (N_7191,N_6276,N_6702);
nor U7192 (N_7192,N_6234,N_6772);
and U7193 (N_7193,N_6290,N_6467);
and U7194 (N_7194,N_6403,N_6228);
and U7195 (N_7195,N_6594,N_6691);
or U7196 (N_7196,N_6350,N_6979);
or U7197 (N_7197,N_6238,N_6714);
nand U7198 (N_7198,N_6991,N_6939);
and U7199 (N_7199,N_6582,N_6788);
nand U7200 (N_7200,N_6874,N_6245);
xnor U7201 (N_7201,N_6576,N_6272);
or U7202 (N_7202,N_6735,N_6108);
xor U7203 (N_7203,N_6590,N_6118);
xor U7204 (N_7204,N_6078,N_6880);
or U7205 (N_7205,N_6365,N_6549);
nand U7206 (N_7206,N_6240,N_6220);
nand U7207 (N_7207,N_6247,N_6026);
xor U7208 (N_7208,N_6048,N_6845);
xor U7209 (N_7209,N_6041,N_6782);
and U7210 (N_7210,N_6069,N_6557);
and U7211 (N_7211,N_6320,N_6931);
nand U7212 (N_7212,N_6739,N_6797);
and U7213 (N_7213,N_6854,N_6440);
and U7214 (N_7214,N_6507,N_6427);
xor U7215 (N_7215,N_6264,N_6659);
nand U7216 (N_7216,N_6338,N_6773);
nor U7217 (N_7217,N_6429,N_6003);
and U7218 (N_7218,N_6381,N_6921);
nor U7219 (N_7219,N_6652,N_6810);
nor U7220 (N_7220,N_6054,N_6602);
xnor U7221 (N_7221,N_6624,N_6449);
xor U7222 (N_7222,N_6589,N_6997);
nor U7223 (N_7223,N_6032,N_6165);
xor U7224 (N_7224,N_6074,N_6770);
and U7225 (N_7225,N_6050,N_6033);
xnor U7226 (N_7226,N_6346,N_6777);
nor U7227 (N_7227,N_6710,N_6536);
nand U7228 (N_7228,N_6644,N_6463);
nor U7229 (N_7229,N_6281,N_6688);
xnor U7230 (N_7230,N_6656,N_6663);
nand U7231 (N_7231,N_6905,N_6898);
xor U7232 (N_7232,N_6805,N_6082);
nand U7233 (N_7233,N_6578,N_6482);
nor U7234 (N_7234,N_6574,N_6119);
xor U7235 (N_7235,N_6275,N_6718);
or U7236 (N_7236,N_6992,N_6066);
nand U7237 (N_7237,N_6378,N_6438);
nor U7238 (N_7238,N_6844,N_6539);
xnor U7239 (N_7239,N_6450,N_6064);
and U7240 (N_7240,N_6883,N_6354);
and U7241 (N_7241,N_6051,N_6366);
nand U7242 (N_7242,N_6384,N_6110);
nor U7243 (N_7243,N_6193,N_6113);
or U7244 (N_7244,N_6204,N_6837);
nor U7245 (N_7245,N_6503,N_6400);
xor U7246 (N_7246,N_6423,N_6947);
nand U7247 (N_7247,N_6195,N_6219);
and U7248 (N_7248,N_6133,N_6636);
nand U7249 (N_7249,N_6468,N_6833);
nor U7250 (N_7250,N_6831,N_6120);
and U7251 (N_7251,N_6560,N_6310);
and U7252 (N_7252,N_6840,N_6187);
xor U7253 (N_7253,N_6881,N_6674);
nand U7254 (N_7254,N_6849,N_6389);
or U7255 (N_7255,N_6402,N_6413);
and U7256 (N_7256,N_6484,N_6347);
nor U7257 (N_7257,N_6128,N_6916);
nor U7258 (N_7258,N_6936,N_6618);
xnor U7259 (N_7259,N_6177,N_6956);
or U7260 (N_7260,N_6729,N_6024);
nand U7261 (N_7261,N_6850,N_6583);
and U7262 (N_7262,N_6888,N_6625);
nor U7263 (N_7263,N_6722,N_6435);
nand U7264 (N_7264,N_6339,N_6230);
xor U7265 (N_7265,N_6089,N_6203);
nor U7266 (N_7266,N_6116,N_6919);
or U7267 (N_7267,N_6300,N_6580);
or U7268 (N_7268,N_6676,N_6908);
nand U7269 (N_7269,N_6703,N_6117);
or U7270 (N_7270,N_6914,N_6464);
and U7271 (N_7271,N_6183,N_6019);
nand U7272 (N_7272,N_6937,N_6489);
nor U7273 (N_7273,N_6523,N_6210);
or U7274 (N_7274,N_6565,N_6943);
xnor U7275 (N_7275,N_6792,N_6428);
xnor U7276 (N_7276,N_6719,N_6901);
nand U7277 (N_7277,N_6122,N_6473);
nor U7278 (N_7278,N_6093,N_6899);
or U7279 (N_7279,N_6232,N_6448);
or U7280 (N_7280,N_6613,N_6006);
xor U7281 (N_7281,N_6942,N_6072);
nor U7282 (N_7282,N_6666,N_6112);
nor U7283 (N_7283,N_6315,N_6795);
xnor U7284 (N_7284,N_6912,N_6733);
xor U7285 (N_7285,N_6926,N_6906);
xor U7286 (N_7286,N_6715,N_6095);
nor U7287 (N_7287,N_6619,N_6969);
or U7288 (N_7288,N_6861,N_6258);
nor U7289 (N_7289,N_6920,N_6058);
nand U7290 (N_7290,N_6084,N_6336);
and U7291 (N_7291,N_6608,N_6155);
xor U7292 (N_7292,N_6039,N_6701);
nand U7293 (N_7293,N_6251,N_6139);
and U7294 (N_7294,N_6115,N_6664);
and U7295 (N_7295,N_6974,N_6340);
nand U7296 (N_7296,N_6067,N_6627);
and U7297 (N_7297,N_6326,N_6478);
nand U7298 (N_7298,N_6823,N_6224);
nor U7299 (N_7299,N_6002,N_6544);
or U7300 (N_7300,N_6548,N_6136);
nor U7301 (N_7301,N_6605,N_6008);
nand U7302 (N_7302,N_6909,N_6562);
and U7303 (N_7303,N_6043,N_6972);
nor U7304 (N_7304,N_6437,N_6364);
xnor U7305 (N_7305,N_6333,N_6526);
nor U7306 (N_7306,N_6787,N_6099);
nand U7307 (N_7307,N_6098,N_6296);
and U7308 (N_7308,N_6633,N_6980);
or U7309 (N_7309,N_6953,N_6088);
xor U7310 (N_7310,N_6323,N_6566);
or U7311 (N_7311,N_6675,N_6163);
xor U7312 (N_7312,N_6556,N_6904);
nor U7313 (N_7313,N_6007,N_6158);
or U7314 (N_7314,N_6363,N_6607);
and U7315 (N_7315,N_6431,N_6649);
nor U7316 (N_7316,N_6262,N_6884);
xnor U7317 (N_7317,N_6907,N_6061);
and U7318 (N_7318,N_6959,N_6812);
nand U7319 (N_7319,N_6927,N_6205);
or U7320 (N_7320,N_6452,N_6830);
nor U7321 (N_7321,N_6246,N_6505);
xor U7322 (N_7322,N_6768,N_6342);
xor U7323 (N_7323,N_6864,N_6477);
nor U7324 (N_7324,N_6282,N_6255);
xnor U7325 (N_7325,N_6534,N_6086);
nand U7326 (N_7326,N_6044,N_6056);
xor U7327 (N_7327,N_6774,N_6611);
nand U7328 (N_7328,N_6309,N_6685);
and U7329 (N_7329,N_6062,N_6206);
and U7330 (N_7330,N_6623,N_6552);
and U7331 (N_7331,N_6472,N_6796);
or U7332 (N_7332,N_6181,N_6212);
nand U7333 (N_7333,N_6022,N_6975);
nand U7334 (N_7334,N_6341,N_6501);
nand U7335 (N_7335,N_6144,N_6261);
or U7336 (N_7336,N_6910,N_6696);
xor U7337 (N_7337,N_6080,N_6270);
or U7338 (N_7338,N_6021,N_6573);
and U7339 (N_7339,N_6383,N_6814);
xor U7340 (N_7340,N_6475,N_6786);
nand U7341 (N_7341,N_6699,N_6194);
or U7342 (N_7342,N_6724,N_6571);
nor U7343 (N_7343,N_6781,N_6933);
and U7344 (N_7344,N_6131,N_6778);
and U7345 (N_7345,N_6269,N_6740);
xnor U7346 (N_7346,N_6535,N_6159);
or U7347 (N_7347,N_6677,N_6231);
or U7348 (N_7348,N_6263,N_6858);
nand U7349 (N_7349,N_6575,N_6207);
and U7350 (N_7350,N_6114,N_6213);
or U7351 (N_7351,N_6555,N_6479);
or U7352 (N_7352,N_6298,N_6329);
nor U7353 (N_7353,N_6824,N_6031);
nor U7354 (N_7354,N_6609,N_6485);
nand U7355 (N_7355,N_6036,N_6277);
and U7356 (N_7356,N_6481,N_6799);
or U7357 (N_7357,N_6877,N_6678);
nor U7358 (N_7358,N_6101,N_6130);
xnor U7359 (N_7359,N_6946,N_6712);
or U7360 (N_7360,N_6388,N_6542);
nor U7361 (N_7361,N_6595,N_6151);
xor U7362 (N_7362,N_6345,N_6707);
or U7363 (N_7363,N_6873,N_6436);
nor U7364 (N_7364,N_6616,N_6695);
or U7365 (N_7365,N_6013,N_6632);
nand U7366 (N_7366,N_6121,N_6520);
nor U7367 (N_7367,N_6776,N_6758);
or U7368 (N_7368,N_6894,N_6950);
and U7369 (N_7369,N_6351,N_6629);
nand U7370 (N_7370,N_6289,N_6808);
or U7371 (N_7371,N_6697,N_6999);
or U7372 (N_7372,N_6716,N_6517);
nor U7373 (N_7373,N_6838,N_6807);
nand U7374 (N_7374,N_6955,N_6425);
and U7375 (N_7375,N_6417,N_6891);
and U7376 (N_7376,N_6360,N_6689);
or U7377 (N_7377,N_6081,N_6570);
and U7378 (N_7378,N_6903,N_6254);
xor U7379 (N_7379,N_6395,N_6124);
nand U7380 (N_7380,N_6104,N_6822);
xor U7381 (N_7381,N_6499,N_6487);
or U7382 (N_7382,N_6334,N_6924);
xnor U7383 (N_7383,N_6486,N_6988);
nor U7384 (N_7384,N_6635,N_6693);
and U7385 (N_7385,N_6648,N_6283);
nor U7386 (N_7386,N_6834,N_6361);
xor U7387 (N_7387,N_6285,N_6222);
or U7388 (N_7388,N_6097,N_6734);
and U7389 (N_7389,N_6103,N_6379);
and U7390 (N_7390,N_6138,N_6079);
nor U7391 (N_7391,N_6917,N_6524);
and U7392 (N_7392,N_6757,N_6047);
xnor U7393 (N_7393,N_6229,N_6893);
xor U7394 (N_7394,N_6600,N_6588);
xnor U7395 (N_7395,N_6711,N_6687);
and U7396 (N_7396,N_6083,N_6012);
or U7397 (N_7397,N_6982,N_6723);
nand U7398 (N_7398,N_6709,N_6841);
and U7399 (N_7399,N_6369,N_6153);
and U7400 (N_7400,N_6173,N_6330);
nand U7401 (N_7401,N_6456,N_6199);
and U7402 (N_7402,N_6726,N_6755);
xor U7403 (N_7403,N_6599,N_6352);
nand U7404 (N_7404,N_6380,N_6316);
and U7405 (N_7405,N_6416,N_6476);
nand U7406 (N_7406,N_6848,N_6045);
nor U7407 (N_7407,N_6509,N_6785);
nor U7408 (N_7408,N_6764,N_6367);
nand U7409 (N_7409,N_6180,N_6626);
nor U7410 (N_7410,N_6070,N_6765);
xor U7411 (N_7411,N_6147,N_6961);
xor U7412 (N_7412,N_6538,N_6945);
and U7413 (N_7413,N_6736,N_6412);
xor U7414 (N_7414,N_6303,N_6800);
or U7415 (N_7415,N_6615,N_6454);
xor U7416 (N_7416,N_6855,N_6102);
nand U7417 (N_7417,N_6522,N_6886);
or U7418 (N_7418,N_6655,N_6495);
nor U7419 (N_7419,N_6856,N_6640);
nand U7420 (N_7420,N_6063,N_6046);
nor U7421 (N_7421,N_6971,N_6948);
nand U7422 (N_7422,N_6214,N_6789);
and U7423 (N_7423,N_6186,N_6178);
or U7424 (N_7424,N_6631,N_6169);
nor U7425 (N_7425,N_6639,N_6987);
nand U7426 (N_7426,N_6508,N_6990);
and U7427 (N_7427,N_6614,N_6872);
xnor U7428 (N_7428,N_6867,N_6349);
and U7429 (N_7429,N_6052,N_6239);
and U7430 (N_7430,N_6725,N_6647);
xor U7431 (N_7431,N_6192,N_6839);
xnor U7432 (N_7432,N_6393,N_6809);
and U7433 (N_7433,N_6156,N_6915);
or U7434 (N_7434,N_6059,N_6938);
and U7435 (N_7435,N_6295,N_6344);
and U7436 (N_7436,N_6592,N_6068);
and U7437 (N_7437,N_6572,N_6871);
xnor U7438 (N_7438,N_6728,N_6355);
and U7439 (N_7439,N_6279,N_6242);
nand U7440 (N_7440,N_6780,N_6825);
or U7441 (N_7441,N_6878,N_6502);
xor U7442 (N_7442,N_6145,N_6049);
xnor U7443 (N_7443,N_6622,N_6077);
nand U7444 (N_7444,N_6218,N_6993);
and U7445 (N_7445,N_6984,N_6598);
nor U7446 (N_7446,N_6857,N_6705);
xnor U7447 (N_7447,N_6331,N_6398);
nor U7448 (N_7448,N_6686,N_6318);
xnor U7449 (N_7449,N_6545,N_6744);
xor U7450 (N_7450,N_6459,N_6650);
nand U7451 (N_7451,N_6513,N_6929);
and U7452 (N_7452,N_6075,N_6483);
nand U7453 (N_7453,N_6280,N_6142);
and U7454 (N_7454,N_6314,N_6803);
or U7455 (N_7455,N_6673,N_6343);
nor U7456 (N_7456,N_6321,N_6396);
or U7457 (N_7457,N_6094,N_6304);
and U7458 (N_7458,N_6892,N_6879);
nor U7459 (N_7459,N_6418,N_6368);
nor U7460 (N_7460,N_6584,N_6967);
or U7461 (N_7461,N_6952,N_6434);
nor U7462 (N_7462,N_6998,N_6216);
and U7463 (N_7463,N_6741,N_6265);
xnor U7464 (N_7464,N_6642,N_6492);
xor U7465 (N_7465,N_6681,N_6743);
nor U7466 (N_7466,N_6252,N_6737);
nand U7467 (N_7467,N_6721,N_6760);
nor U7468 (N_7468,N_6227,N_6804);
xor U7469 (N_7469,N_6586,N_6940);
or U7470 (N_7470,N_6885,N_6135);
or U7471 (N_7471,N_6866,N_6559);
nand U7472 (N_7472,N_6293,N_6480);
nor U7473 (N_7473,N_6928,N_6932);
xor U7474 (N_7474,N_6646,N_6708);
and U7475 (N_7475,N_6375,N_6188);
and U7476 (N_7476,N_6202,N_6994);
nor U7477 (N_7477,N_6200,N_6657);
or U7478 (N_7478,N_6143,N_6453);
nor U7479 (N_7479,N_6474,N_6172);
nor U7480 (N_7480,N_6132,N_6085);
and U7481 (N_7481,N_6244,N_6404);
nand U7482 (N_7482,N_6966,N_6951);
nand U7483 (N_7483,N_6076,N_6918);
or U7484 (N_7484,N_6028,N_6754);
xnor U7485 (N_7485,N_6817,N_6297);
xnor U7486 (N_7486,N_6260,N_6963);
nor U7487 (N_7487,N_6870,N_6569);
and U7488 (N_7488,N_6504,N_6274);
or U7489 (N_7489,N_6587,N_6414);
or U7490 (N_7490,N_6978,N_6965);
nor U7491 (N_7491,N_6558,N_6305);
and U7492 (N_7492,N_6976,N_6302);
nor U7493 (N_7493,N_6680,N_6190);
xor U7494 (N_7494,N_6529,N_6748);
nor U7495 (N_7495,N_6170,N_6682);
and U7496 (N_7496,N_6671,N_6182);
nand U7497 (N_7497,N_6215,N_6811);
nor U7498 (N_7498,N_6662,N_6278);
nand U7499 (N_7499,N_6506,N_6096);
xor U7500 (N_7500,N_6656,N_6056);
or U7501 (N_7501,N_6069,N_6853);
nor U7502 (N_7502,N_6249,N_6181);
nand U7503 (N_7503,N_6347,N_6556);
nand U7504 (N_7504,N_6567,N_6134);
or U7505 (N_7505,N_6024,N_6572);
or U7506 (N_7506,N_6398,N_6505);
or U7507 (N_7507,N_6040,N_6289);
nor U7508 (N_7508,N_6649,N_6499);
xnor U7509 (N_7509,N_6355,N_6920);
nor U7510 (N_7510,N_6656,N_6640);
or U7511 (N_7511,N_6435,N_6286);
and U7512 (N_7512,N_6554,N_6999);
and U7513 (N_7513,N_6909,N_6927);
xor U7514 (N_7514,N_6975,N_6221);
nor U7515 (N_7515,N_6794,N_6562);
nor U7516 (N_7516,N_6238,N_6686);
or U7517 (N_7517,N_6118,N_6827);
or U7518 (N_7518,N_6696,N_6323);
xor U7519 (N_7519,N_6218,N_6158);
or U7520 (N_7520,N_6471,N_6160);
xor U7521 (N_7521,N_6952,N_6798);
xor U7522 (N_7522,N_6126,N_6664);
xor U7523 (N_7523,N_6817,N_6247);
or U7524 (N_7524,N_6848,N_6761);
and U7525 (N_7525,N_6423,N_6819);
xnor U7526 (N_7526,N_6668,N_6245);
nand U7527 (N_7527,N_6980,N_6381);
nor U7528 (N_7528,N_6153,N_6107);
or U7529 (N_7529,N_6300,N_6583);
or U7530 (N_7530,N_6362,N_6835);
nor U7531 (N_7531,N_6434,N_6933);
nor U7532 (N_7532,N_6763,N_6351);
nand U7533 (N_7533,N_6770,N_6183);
or U7534 (N_7534,N_6874,N_6437);
and U7535 (N_7535,N_6066,N_6253);
nand U7536 (N_7536,N_6464,N_6904);
xnor U7537 (N_7537,N_6821,N_6775);
nor U7538 (N_7538,N_6705,N_6727);
or U7539 (N_7539,N_6321,N_6901);
xor U7540 (N_7540,N_6226,N_6181);
and U7541 (N_7541,N_6534,N_6245);
and U7542 (N_7542,N_6618,N_6180);
nor U7543 (N_7543,N_6693,N_6762);
xnor U7544 (N_7544,N_6375,N_6784);
xor U7545 (N_7545,N_6348,N_6227);
and U7546 (N_7546,N_6073,N_6565);
nand U7547 (N_7547,N_6631,N_6698);
and U7548 (N_7548,N_6661,N_6590);
nand U7549 (N_7549,N_6813,N_6093);
or U7550 (N_7550,N_6384,N_6273);
xor U7551 (N_7551,N_6400,N_6903);
xor U7552 (N_7552,N_6643,N_6529);
nand U7553 (N_7553,N_6769,N_6632);
nor U7554 (N_7554,N_6977,N_6905);
nand U7555 (N_7555,N_6964,N_6549);
xnor U7556 (N_7556,N_6727,N_6359);
or U7557 (N_7557,N_6091,N_6566);
nand U7558 (N_7558,N_6782,N_6209);
nand U7559 (N_7559,N_6593,N_6698);
or U7560 (N_7560,N_6086,N_6550);
nand U7561 (N_7561,N_6935,N_6565);
or U7562 (N_7562,N_6420,N_6383);
nand U7563 (N_7563,N_6116,N_6334);
nand U7564 (N_7564,N_6460,N_6489);
or U7565 (N_7565,N_6540,N_6708);
nor U7566 (N_7566,N_6733,N_6075);
or U7567 (N_7567,N_6689,N_6865);
nand U7568 (N_7568,N_6122,N_6070);
xor U7569 (N_7569,N_6619,N_6578);
and U7570 (N_7570,N_6183,N_6200);
nand U7571 (N_7571,N_6255,N_6378);
nor U7572 (N_7572,N_6016,N_6480);
xor U7573 (N_7573,N_6022,N_6856);
and U7574 (N_7574,N_6716,N_6004);
nor U7575 (N_7575,N_6596,N_6727);
or U7576 (N_7576,N_6031,N_6272);
nor U7577 (N_7577,N_6649,N_6335);
nor U7578 (N_7578,N_6512,N_6677);
or U7579 (N_7579,N_6354,N_6100);
and U7580 (N_7580,N_6065,N_6746);
nand U7581 (N_7581,N_6055,N_6141);
and U7582 (N_7582,N_6505,N_6676);
or U7583 (N_7583,N_6754,N_6095);
nand U7584 (N_7584,N_6936,N_6763);
xnor U7585 (N_7585,N_6265,N_6026);
xnor U7586 (N_7586,N_6903,N_6029);
xor U7587 (N_7587,N_6152,N_6957);
or U7588 (N_7588,N_6604,N_6077);
xor U7589 (N_7589,N_6265,N_6422);
nand U7590 (N_7590,N_6652,N_6231);
xnor U7591 (N_7591,N_6115,N_6218);
or U7592 (N_7592,N_6753,N_6577);
nor U7593 (N_7593,N_6866,N_6091);
or U7594 (N_7594,N_6428,N_6326);
nor U7595 (N_7595,N_6996,N_6714);
nand U7596 (N_7596,N_6123,N_6399);
or U7597 (N_7597,N_6750,N_6700);
and U7598 (N_7598,N_6399,N_6289);
nor U7599 (N_7599,N_6054,N_6381);
or U7600 (N_7600,N_6443,N_6128);
and U7601 (N_7601,N_6720,N_6019);
xor U7602 (N_7602,N_6229,N_6829);
nor U7603 (N_7603,N_6283,N_6315);
nor U7604 (N_7604,N_6464,N_6937);
and U7605 (N_7605,N_6925,N_6692);
xor U7606 (N_7606,N_6149,N_6255);
xor U7607 (N_7607,N_6960,N_6941);
and U7608 (N_7608,N_6193,N_6620);
xnor U7609 (N_7609,N_6515,N_6625);
xor U7610 (N_7610,N_6591,N_6058);
or U7611 (N_7611,N_6261,N_6085);
nand U7612 (N_7612,N_6569,N_6446);
and U7613 (N_7613,N_6033,N_6093);
nor U7614 (N_7614,N_6489,N_6181);
and U7615 (N_7615,N_6863,N_6566);
or U7616 (N_7616,N_6522,N_6597);
nand U7617 (N_7617,N_6180,N_6883);
or U7618 (N_7618,N_6119,N_6756);
and U7619 (N_7619,N_6313,N_6281);
nand U7620 (N_7620,N_6773,N_6385);
nor U7621 (N_7621,N_6590,N_6353);
nor U7622 (N_7622,N_6500,N_6184);
or U7623 (N_7623,N_6131,N_6047);
nor U7624 (N_7624,N_6064,N_6665);
nor U7625 (N_7625,N_6210,N_6067);
or U7626 (N_7626,N_6757,N_6056);
xnor U7627 (N_7627,N_6922,N_6789);
nand U7628 (N_7628,N_6072,N_6757);
nand U7629 (N_7629,N_6345,N_6645);
or U7630 (N_7630,N_6764,N_6607);
or U7631 (N_7631,N_6957,N_6870);
and U7632 (N_7632,N_6677,N_6865);
nand U7633 (N_7633,N_6880,N_6301);
and U7634 (N_7634,N_6849,N_6494);
and U7635 (N_7635,N_6272,N_6510);
or U7636 (N_7636,N_6447,N_6276);
nor U7637 (N_7637,N_6513,N_6760);
xor U7638 (N_7638,N_6348,N_6431);
or U7639 (N_7639,N_6468,N_6665);
nand U7640 (N_7640,N_6359,N_6317);
or U7641 (N_7641,N_6720,N_6783);
or U7642 (N_7642,N_6543,N_6736);
nand U7643 (N_7643,N_6755,N_6215);
and U7644 (N_7644,N_6319,N_6404);
and U7645 (N_7645,N_6214,N_6799);
and U7646 (N_7646,N_6030,N_6104);
xor U7647 (N_7647,N_6350,N_6478);
xnor U7648 (N_7648,N_6260,N_6482);
xnor U7649 (N_7649,N_6954,N_6896);
nand U7650 (N_7650,N_6083,N_6454);
nor U7651 (N_7651,N_6497,N_6038);
and U7652 (N_7652,N_6360,N_6929);
xor U7653 (N_7653,N_6046,N_6253);
nor U7654 (N_7654,N_6641,N_6737);
or U7655 (N_7655,N_6979,N_6091);
or U7656 (N_7656,N_6825,N_6627);
and U7657 (N_7657,N_6263,N_6200);
nand U7658 (N_7658,N_6023,N_6370);
and U7659 (N_7659,N_6400,N_6218);
nor U7660 (N_7660,N_6998,N_6711);
nand U7661 (N_7661,N_6433,N_6883);
xnor U7662 (N_7662,N_6550,N_6753);
nor U7663 (N_7663,N_6122,N_6630);
xor U7664 (N_7664,N_6309,N_6966);
nand U7665 (N_7665,N_6872,N_6127);
xor U7666 (N_7666,N_6413,N_6190);
or U7667 (N_7667,N_6447,N_6595);
and U7668 (N_7668,N_6894,N_6031);
nand U7669 (N_7669,N_6190,N_6063);
nand U7670 (N_7670,N_6095,N_6659);
nand U7671 (N_7671,N_6592,N_6968);
xor U7672 (N_7672,N_6605,N_6123);
nand U7673 (N_7673,N_6124,N_6821);
nand U7674 (N_7674,N_6869,N_6999);
or U7675 (N_7675,N_6479,N_6729);
nor U7676 (N_7676,N_6487,N_6948);
and U7677 (N_7677,N_6941,N_6704);
nand U7678 (N_7678,N_6861,N_6725);
and U7679 (N_7679,N_6661,N_6842);
nor U7680 (N_7680,N_6595,N_6981);
xnor U7681 (N_7681,N_6737,N_6721);
and U7682 (N_7682,N_6269,N_6306);
xnor U7683 (N_7683,N_6613,N_6940);
nand U7684 (N_7684,N_6541,N_6954);
and U7685 (N_7685,N_6318,N_6743);
and U7686 (N_7686,N_6205,N_6545);
and U7687 (N_7687,N_6772,N_6595);
xor U7688 (N_7688,N_6538,N_6255);
or U7689 (N_7689,N_6093,N_6219);
xnor U7690 (N_7690,N_6678,N_6030);
and U7691 (N_7691,N_6644,N_6243);
and U7692 (N_7692,N_6461,N_6201);
nor U7693 (N_7693,N_6374,N_6187);
xor U7694 (N_7694,N_6096,N_6806);
or U7695 (N_7695,N_6251,N_6765);
nand U7696 (N_7696,N_6752,N_6009);
and U7697 (N_7697,N_6228,N_6108);
nor U7698 (N_7698,N_6914,N_6170);
xor U7699 (N_7699,N_6303,N_6690);
nand U7700 (N_7700,N_6456,N_6684);
xor U7701 (N_7701,N_6876,N_6785);
and U7702 (N_7702,N_6451,N_6778);
nor U7703 (N_7703,N_6468,N_6692);
xor U7704 (N_7704,N_6760,N_6686);
nand U7705 (N_7705,N_6549,N_6401);
nand U7706 (N_7706,N_6705,N_6799);
nand U7707 (N_7707,N_6885,N_6578);
or U7708 (N_7708,N_6972,N_6732);
nand U7709 (N_7709,N_6199,N_6582);
or U7710 (N_7710,N_6119,N_6791);
xor U7711 (N_7711,N_6738,N_6476);
nor U7712 (N_7712,N_6743,N_6190);
and U7713 (N_7713,N_6439,N_6841);
xnor U7714 (N_7714,N_6604,N_6244);
nand U7715 (N_7715,N_6660,N_6540);
nand U7716 (N_7716,N_6420,N_6714);
xor U7717 (N_7717,N_6035,N_6257);
or U7718 (N_7718,N_6450,N_6292);
nor U7719 (N_7719,N_6076,N_6472);
or U7720 (N_7720,N_6154,N_6425);
xnor U7721 (N_7721,N_6498,N_6908);
and U7722 (N_7722,N_6765,N_6093);
and U7723 (N_7723,N_6054,N_6798);
and U7724 (N_7724,N_6382,N_6060);
nand U7725 (N_7725,N_6209,N_6960);
and U7726 (N_7726,N_6651,N_6944);
nor U7727 (N_7727,N_6163,N_6232);
or U7728 (N_7728,N_6717,N_6918);
and U7729 (N_7729,N_6580,N_6152);
nand U7730 (N_7730,N_6375,N_6540);
nand U7731 (N_7731,N_6334,N_6675);
and U7732 (N_7732,N_6911,N_6415);
or U7733 (N_7733,N_6597,N_6466);
and U7734 (N_7734,N_6208,N_6631);
nor U7735 (N_7735,N_6779,N_6706);
or U7736 (N_7736,N_6911,N_6201);
and U7737 (N_7737,N_6144,N_6508);
or U7738 (N_7738,N_6653,N_6849);
and U7739 (N_7739,N_6839,N_6065);
or U7740 (N_7740,N_6529,N_6407);
and U7741 (N_7741,N_6547,N_6794);
and U7742 (N_7742,N_6940,N_6281);
nor U7743 (N_7743,N_6726,N_6224);
xnor U7744 (N_7744,N_6786,N_6820);
and U7745 (N_7745,N_6788,N_6362);
xor U7746 (N_7746,N_6627,N_6508);
and U7747 (N_7747,N_6807,N_6967);
nand U7748 (N_7748,N_6911,N_6467);
and U7749 (N_7749,N_6880,N_6628);
xor U7750 (N_7750,N_6780,N_6897);
and U7751 (N_7751,N_6952,N_6961);
nand U7752 (N_7752,N_6829,N_6063);
nand U7753 (N_7753,N_6188,N_6292);
and U7754 (N_7754,N_6647,N_6993);
nor U7755 (N_7755,N_6133,N_6533);
xnor U7756 (N_7756,N_6543,N_6970);
xor U7757 (N_7757,N_6916,N_6210);
and U7758 (N_7758,N_6217,N_6705);
xor U7759 (N_7759,N_6843,N_6529);
nor U7760 (N_7760,N_6741,N_6554);
and U7761 (N_7761,N_6080,N_6332);
and U7762 (N_7762,N_6454,N_6909);
nand U7763 (N_7763,N_6451,N_6805);
nand U7764 (N_7764,N_6242,N_6469);
or U7765 (N_7765,N_6105,N_6908);
nand U7766 (N_7766,N_6307,N_6581);
and U7767 (N_7767,N_6200,N_6346);
and U7768 (N_7768,N_6728,N_6481);
nand U7769 (N_7769,N_6888,N_6938);
xor U7770 (N_7770,N_6353,N_6829);
or U7771 (N_7771,N_6608,N_6499);
or U7772 (N_7772,N_6301,N_6879);
nor U7773 (N_7773,N_6850,N_6141);
nor U7774 (N_7774,N_6760,N_6802);
nand U7775 (N_7775,N_6926,N_6429);
or U7776 (N_7776,N_6508,N_6129);
xnor U7777 (N_7777,N_6922,N_6531);
and U7778 (N_7778,N_6861,N_6182);
or U7779 (N_7779,N_6126,N_6572);
nor U7780 (N_7780,N_6525,N_6064);
xor U7781 (N_7781,N_6177,N_6073);
nand U7782 (N_7782,N_6094,N_6312);
xnor U7783 (N_7783,N_6177,N_6329);
nand U7784 (N_7784,N_6857,N_6720);
or U7785 (N_7785,N_6214,N_6515);
xnor U7786 (N_7786,N_6212,N_6950);
or U7787 (N_7787,N_6253,N_6192);
nand U7788 (N_7788,N_6249,N_6325);
nor U7789 (N_7789,N_6057,N_6159);
nand U7790 (N_7790,N_6256,N_6709);
nor U7791 (N_7791,N_6617,N_6851);
and U7792 (N_7792,N_6408,N_6673);
or U7793 (N_7793,N_6254,N_6767);
and U7794 (N_7794,N_6373,N_6259);
xnor U7795 (N_7795,N_6007,N_6769);
nand U7796 (N_7796,N_6346,N_6427);
and U7797 (N_7797,N_6170,N_6184);
xor U7798 (N_7798,N_6730,N_6745);
nand U7799 (N_7799,N_6953,N_6434);
xnor U7800 (N_7800,N_6975,N_6408);
or U7801 (N_7801,N_6970,N_6536);
and U7802 (N_7802,N_6407,N_6265);
nand U7803 (N_7803,N_6475,N_6605);
nor U7804 (N_7804,N_6405,N_6585);
nand U7805 (N_7805,N_6387,N_6342);
nor U7806 (N_7806,N_6224,N_6294);
nor U7807 (N_7807,N_6264,N_6306);
xnor U7808 (N_7808,N_6021,N_6862);
or U7809 (N_7809,N_6104,N_6760);
nand U7810 (N_7810,N_6503,N_6080);
xnor U7811 (N_7811,N_6235,N_6769);
nand U7812 (N_7812,N_6286,N_6053);
nand U7813 (N_7813,N_6557,N_6434);
or U7814 (N_7814,N_6566,N_6656);
xnor U7815 (N_7815,N_6529,N_6640);
nand U7816 (N_7816,N_6299,N_6192);
and U7817 (N_7817,N_6309,N_6841);
xor U7818 (N_7818,N_6219,N_6847);
xor U7819 (N_7819,N_6953,N_6780);
or U7820 (N_7820,N_6344,N_6634);
xnor U7821 (N_7821,N_6088,N_6452);
xor U7822 (N_7822,N_6714,N_6018);
nor U7823 (N_7823,N_6857,N_6641);
nor U7824 (N_7824,N_6796,N_6536);
and U7825 (N_7825,N_6641,N_6939);
nor U7826 (N_7826,N_6109,N_6712);
nand U7827 (N_7827,N_6142,N_6216);
or U7828 (N_7828,N_6979,N_6189);
or U7829 (N_7829,N_6346,N_6326);
xor U7830 (N_7830,N_6943,N_6040);
or U7831 (N_7831,N_6261,N_6200);
and U7832 (N_7832,N_6078,N_6817);
or U7833 (N_7833,N_6433,N_6387);
xor U7834 (N_7834,N_6625,N_6783);
nand U7835 (N_7835,N_6130,N_6630);
xor U7836 (N_7836,N_6826,N_6276);
xnor U7837 (N_7837,N_6072,N_6587);
and U7838 (N_7838,N_6288,N_6955);
nand U7839 (N_7839,N_6824,N_6977);
xor U7840 (N_7840,N_6801,N_6177);
and U7841 (N_7841,N_6031,N_6721);
nor U7842 (N_7842,N_6612,N_6357);
xnor U7843 (N_7843,N_6381,N_6490);
or U7844 (N_7844,N_6799,N_6741);
nand U7845 (N_7845,N_6509,N_6056);
and U7846 (N_7846,N_6301,N_6583);
or U7847 (N_7847,N_6227,N_6354);
nor U7848 (N_7848,N_6318,N_6150);
nand U7849 (N_7849,N_6708,N_6547);
nor U7850 (N_7850,N_6558,N_6449);
nor U7851 (N_7851,N_6570,N_6401);
nand U7852 (N_7852,N_6086,N_6448);
nor U7853 (N_7853,N_6949,N_6791);
and U7854 (N_7854,N_6834,N_6856);
nand U7855 (N_7855,N_6692,N_6660);
nand U7856 (N_7856,N_6940,N_6178);
nand U7857 (N_7857,N_6500,N_6363);
nand U7858 (N_7858,N_6400,N_6461);
xor U7859 (N_7859,N_6642,N_6753);
nor U7860 (N_7860,N_6062,N_6667);
nor U7861 (N_7861,N_6806,N_6159);
or U7862 (N_7862,N_6077,N_6413);
nor U7863 (N_7863,N_6829,N_6997);
and U7864 (N_7864,N_6327,N_6299);
or U7865 (N_7865,N_6907,N_6073);
or U7866 (N_7866,N_6872,N_6992);
nor U7867 (N_7867,N_6243,N_6226);
and U7868 (N_7868,N_6672,N_6324);
and U7869 (N_7869,N_6034,N_6974);
nand U7870 (N_7870,N_6985,N_6780);
nand U7871 (N_7871,N_6494,N_6691);
nand U7872 (N_7872,N_6414,N_6306);
xor U7873 (N_7873,N_6449,N_6222);
xor U7874 (N_7874,N_6903,N_6813);
and U7875 (N_7875,N_6016,N_6746);
and U7876 (N_7876,N_6695,N_6460);
and U7877 (N_7877,N_6038,N_6293);
nor U7878 (N_7878,N_6171,N_6509);
nand U7879 (N_7879,N_6035,N_6100);
and U7880 (N_7880,N_6558,N_6092);
or U7881 (N_7881,N_6263,N_6434);
nor U7882 (N_7882,N_6695,N_6192);
or U7883 (N_7883,N_6874,N_6361);
or U7884 (N_7884,N_6061,N_6868);
or U7885 (N_7885,N_6077,N_6621);
or U7886 (N_7886,N_6512,N_6819);
nand U7887 (N_7887,N_6950,N_6588);
and U7888 (N_7888,N_6647,N_6399);
and U7889 (N_7889,N_6313,N_6264);
and U7890 (N_7890,N_6993,N_6076);
nor U7891 (N_7891,N_6341,N_6743);
or U7892 (N_7892,N_6111,N_6321);
or U7893 (N_7893,N_6639,N_6955);
nand U7894 (N_7894,N_6665,N_6415);
xor U7895 (N_7895,N_6849,N_6085);
nand U7896 (N_7896,N_6472,N_6337);
and U7897 (N_7897,N_6466,N_6206);
xor U7898 (N_7898,N_6202,N_6739);
xor U7899 (N_7899,N_6821,N_6731);
or U7900 (N_7900,N_6835,N_6144);
nand U7901 (N_7901,N_6048,N_6628);
xor U7902 (N_7902,N_6261,N_6544);
nor U7903 (N_7903,N_6674,N_6613);
nor U7904 (N_7904,N_6172,N_6280);
and U7905 (N_7905,N_6806,N_6420);
nor U7906 (N_7906,N_6287,N_6939);
and U7907 (N_7907,N_6489,N_6991);
nor U7908 (N_7908,N_6718,N_6327);
xnor U7909 (N_7909,N_6383,N_6412);
xor U7910 (N_7910,N_6738,N_6554);
xnor U7911 (N_7911,N_6137,N_6599);
xor U7912 (N_7912,N_6843,N_6261);
nand U7913 (N_7913,N_6902,N_6801);
or U7914 (N_7914,N_6363,N_6437);
nand U7915 (N_7915,N_6197,N_6033);
and U7916 (N_7916,N_6372,N_6724);
nand U7917 (N_7917,N_6716,N_6302);
nor U7918 (N_7918,N_6359,N_6010);
or U7919 (N_7919,N_6858,N_6673);
and U7920 (N_7920,N_6260,N_6033);
and U7921 (N_7921,N_6822,N_6406);
or U7922 (N_7922,N_6224,N_6001);
xor U7923 (N_7923,N_6818,N_6992);
nor U7924 (N_7924,N_6513,N_6526);
nor U7925 (N_7925,N_6980,N_6300);
xor U7926 (N_7926,N_6329,N_6708);
and U7927 (N_7927,N_6115,N_6506);
xnor U7928 (N_7928,N_6175,N_6124);
nor U7929 (N_7929,N_6262,N_6879);
nand U7930 (N_7930,N_6641,N_6153);
nand U7931 (N_7931,N_6387,N_6525);
or U7932 (N_7932,N_6061,N_6347);
and U7933 (N_7933,N_6267,N_6907);
nand U7934 (N_7934,N_6142,N_6447);
or U7935 (N_7935,N_6287,N_6273);
nor U7936 (N_7936,N_6729,N_6623);
and U7937 (N_7937,N_6683,N_6874);
nor U7938 (N_7938,N_6478,N_6158);
xnor U7939 (N_7939,N_6879,N_6198);
nor U7940 (N_7940,N_6663,N_6754);
nor U7941 (N_7941,N_6321,N_6821);
and U7942 (N_7942,N_6995,N_6154);
or U7943 (N_7943,N_6860,N_6691);
or U7944 (N_7944,N_6006,N_6040);
or U7945 (N_7945,N_6380,N_6783);
xnor U7946 (N_7946,N_6131,N_6152);
xnor U7947 (N_7947,N_6982,N_6618);
and U7948 (N_7948,N_6488,N_6854);
nand U7949 (N_7949,N_6898,N_6999);
nor U7950 (N_7950,N_6073,N_6354);
nor U7951 (N_7951,N_6625,N_6947);
xor U7952 (N_7952,N_6017,N_6819);
and U7953 (N_7953,N_6021,N_6344);
nor U7954 (N_7954,N_6105,N_6969);
nor U7955 (N_7955,N_6217,N_6927);
or U7956 (N_7956,N_6791,N_6087);
nor U7957 (N_7957,N_6586,N_6450);
or U7958 (N_7958,N_6547,N_6121);
xnor U7959 (N_7959,N_6968,N_6366);
or U7960 (N_7960,N_6067,N_6892);
and U7961 (N_7961,N_6496,N_6928);
and U7962 (N_7962,N_6437,N_6234);
and U7963 (N_7963,N_6303,N_6182);
and U7964 (N_7964,N_6621,N_6950);
nor U7965 (N_7965,N_6743,N_6303);
and U7966 (N_7966,N_6136,N_6153);
or U7967 (N_7967,N_6721,N_6882);
xnor U7968 (N_7968,N_6924,N_6399);
xnor U7969 (N_7969,N_6306,N_6165);
or U7970 (N_7970,N_6870,N_6382);
xor U7971 (N_7971,N_6086,N_6546);
or U7972 (N_7972,N_6062,N_6973);
xnor U7973 (N_7973,N_6391,N_6749);
xnor U7974 (N_7974,N_6888,N_6972);
nor U7975 (N_7975,N_6908,N_6897);
and U7976 (N_7976,N_6617,N_6838);
or U7977 (N_7977,N_6599,N_6942);
nor U7978 (N_7978,N_6743,N_6678);
nor U7979 (N_7979,N_6082,N_6702);
nand U7980 (N_7980,N_6786,N_6745);
xor U7981 (N_7981,N_6074,N_6071);
nor U7982 (N_7982,N_6071,N_6065);
and U7983 (N_7983,N_6677,N_6838);
xnor U7984 (N_7984,N_6554,N_6868);
or U7985 (N_7985,N_6397,N_6881);
and U7986 (N_7986,N_6569,N_6055);
nand U7987 (N_7987,N_6979,N_6899);
and U7988 (N_7988,N_6626,N_6582);
nand U7989 (N_7989,N_6833,N_6634);
or U7990 (N_7990,N_6017,N_6272);
nand U7991 (N_7991,N_6275,N_6663);
or U7992 (N_7992,N_6562,N_6657);
xnor U7993 (N_7993,N_6157,N_6908);
xnor U7994 (N_7994,N_6034,N_6823);
nand U7995 (N_7995,N_6966,N_6458);
and U7996 (N_7996,N_6871,N_6420);
and U7997 (N_7997,N_6445,N_6594);
xnor U7998 (N_7998,N_6611,N_6607);
nand U7999 (N_7999,N_6518,N_6081);
or U8000 (N_8000,N_7313,N_7325);
xor U8001 (N_8001,N_7948,N_7234);
nor U8002 (N_8002,N_7595,N_7020);
nand U8003 (N_8003,N_7152,N_7400);
nand U8004 (N_8004,N_7332,N_7495);
xnor U8005 (N_8005,N_7968,N_7704);
nor U8006 (N_8006,N_7046,N_7115);
nor U8007 (N_8007,N_7854,N_7838);
and U8008 (N_8008,N_7190,N_7006);
and U8009 (N_8009,N_7914,N_7412);
nor U8010 (N_8010,N_7677,N_7493);
nor U8011 (N_8011,N_7244,N_7870);
and U8012 (N_8012,N_7195,N_7167);
and U8013 (N_8013,N_7377,N_7408);
and U8014 (N_8014,N_7370,N_7524);
xnor U8015 (N_8015,N_7305,N_7077);
and U8016 (N_8016,N_7315,N_7140);
or U8017 (N_8017,N_7731,N_7442);
nand U8018 (N_8018,N_7534,N_7038);
xor U8019 (N_8019,N_7229,N_7398);
and U8020 (N_8020,N_7894,N_7798);
xor U8021 (N_8021,N_7269,N_7245);
nor U8022 (N_8022,N_7597,N_7171);
xor U8023 (N_8023,N_7317,N_7754);
or U8024 (N_8024,N_7910,N_7949);
or U8025 (N_8025,N_7753,N_7456);
or U8026 (N_8026,N_7516,N_7438);
nor U8027 (N_8027,N_7337,N_7354);
nand U8028 (N_8028,N_7248,N_7514);
nand U8029 (N_8029,N_7805,N_7686);
nand U8030 (N_8030,N_7471,N_7458);
or U8031 (N_8031,N_7070,N_7581);
xor U8032 (N_8032,N_7013,N_7876);
xor U8033 (N_8033,N_7735,N_7364);
nand U8034 (N_8034,N_7341,N_7027);
nor U8035 (N_8035,N_7542,N_7537);
xnor U8036 (N_8036,N_7003,N_7764);
or U8037 (N_8037,N_7952,N_7128);
nor U8038 (N_8038,N_7904,N_7201);
nand U8039 (N_8039,N_7703,N_7921);
nand U8040 (N_8040,N_7622,N_7053);
nand U8041 (N_8041,N_7843,N_7559);
xor U8042 (N_8042,N_7963,N_7821);
xnor U8043 (N_8043,N_7088,N_7886);
and U8044 (N_8044,N_7182,N_7634);
and U8045 (N_8045,N_7819,N_7574);
xor U8046 (N_8046,N_7085,N_7688);
or U8047 (N_8047,N_7453,N_7959);
xor U8048 (N_8048,N_7209,N_7746);
nand U8049 (N_8049,N_7800,N_7094);
and U8050 (N_8050,N_7065,N_7306);
or U8051 (N_8051,N_7916,N_7226);
or U8052 (N_8052,N_7454,N_7874);
or U8053 (N_8053,N_7426,N_7506);
and U8054 (N_8054,N_7625,N_7186);
and U8055 (N_8055,N_7452,N_7745);
nor U8056 (N_8056,N_7270,N_7416);
or U8057 (N_8057,N_7931,N_7722);
nor U8058 (N_8058,N_7814,N_7668);
nand U8059 (N_8059,N_7199,N_7486);
or U8060 (N_8060,N_7738,N_7338);
and U8061 (N_8061,N_7799,N_7518);
nand U8062 (N_8062,N_7974,N_7335);
nor U8063 (N_8063,N_7969,N_7715);
or U8064 (N_8064,N_7002,N_7233);
nand U8065 (N_8065,N_7767,N_7449);
or U8066 (N_8066,N_7241,N_7250);
nor U8067 (N_8067,N_7355,N_7051);
nand U8068 (N_8068,N_7276,N_7385);
nor U8069 (N_8069,N_7889,N_7784);
nand U8070 (N_8070,N_7112,N_7267);
nor U8071 (N_8071,N_7797,N_7845);
nand U8072 (N_8072,N_7594,N_7697);
or U8073 (N_8073,N_7009,N_7905);
and U8074 (N_8074,N_7425,N_7836);
xor U8075 (N_8075,N_7627,N_7258);
xnor U8076 (N_8076,N_7601,N_7073);
nor U8077 (N_8077,N_7175,N_7732);
nor U8078 (N_8078,N_7379,N_7494);
nor U8079 (N_8079,N_7928,N_7345);
xor U8080 (N_8080,N_7380,N_7392);
nand U8081 (N_8081,N_7823,N_7173);
and U8082 (N_8082,N_7641,N_7624);
nand U8083 (N_8083,N_7915,N_7168);
nor U8084 (N_8084,N_7110,N_7163);
nand U8085 (N_8085,N_7585,N_7455);
or U8086 (N_8086,N_7960,N_7221);
xnor U8087 (N_8087,N_7118,N_7719);
nor U8088 (N_8088,N_7272,N_7129);
nand U8089 (N_8089,N_7620,N_7706);
xor U8090 (N_8090,N_7042,N_7950);
xnor U8091 (N_8091,N_7919,N_7447);
and U8092 (N_8092,N_7582,N_7146);
or U8093 (N_8093,N_7045,N_7639);
xnor U8094 (N_8094,N_7057,N_7104);
nand U8095 (N_8095,N_7353,N_7564);
nand U8096 (N_8096,N_7406,N_7975);
xor U8097 (N_8097,N_7461,N_7145);
xnor U8098 (N_8098,N_7572,N_7161);
nor U8099 (N_8099,N_7419,N_7551);
nand U8100 (N_8100,N_7228,N_7888);
and U8101 (N_8101,N_7763,N_7293);
xnor U8102 (N_8102,N_7203,N_7737);
or U8103 (N_8103,N_7039,N_7774);
nand U8104 (N_8104,N_7060,N_7211);
xor U8105 (N_8105,N_7890,N_7154);
or U8106 (N_8106,N_7159,N_7972);
nand U8107 (N_8107,N_7047,N_7691);
nor U8108 (N_8108,N_7074,N_7899);
xnor U8109 (N_8109,N_7106,N_7547);
and U8110 (N_8110,N_7566,N_7718);
and U8111 (N_8111,N_7290,N_7980);
nor U8112 (N_8112,N_7391,N_7658);
nand U8113 (N_8113,N_7583,N_7119);
nand U8114 (N_8114,N_7635,N_7956);
nor U8115 (N_8115,N_7608,N_7422);
or U8116 (N_8116,N_7428,N_7897);
nand U8117 (N_8117,N_7288,N_7664);
nand U8118 (N_8118,N_7067,N_7028);
nand U8119 (N_8119,N_7089,N_7786);
xor U8120 (N_8120,N_7298,N_7589);
or U8121 (N_8121,N_7103,N_7708);
and U8122 (N_8122,N_7696,N_7123);
xnor U8123 (N_8123,N_7436,N_7661);
xor U8124 (N_8124,N_7176,N_7810);
or U8125 (N_8125,N_7184,N_7479);
and U8126 (N_8126,N_7212,N_7144);
and U8127 (N_8127,N_7394,N_7296);
nor U8128 (N_8128,N_7314,N_7008);
nand U8129 (N_8129,N_7382,N_7435);
and U8130 (N_8130,N_7695,N_7091);
nor U8131 (N_8131,N_7979,N_7177);
nand U8132 (N_8132,N_7565,N_7496);
xnor U8133 (N_8133,N_7670,N_7302);
nand U8134 (N_8134,N_7049,N_7026);
nand U8135 (N_8135,N_7557,N_7985);
and U8136 (N_8136,N_7265,N_7474);
xnor U8137 (N_8137,N_7059,N_7035);
nand U8138 (N_8138,N_7917,N_7730);
xor U8139 (N_8139,N_7157,N_7183);
and U8140 (N_8140,N_7384,N_7812);
or U8141 (N_8141,N_7365,N_7993);
or U8142 (N_8142,N_7510,N_7022);
nand U8143 (N_8143,N_7623,N_7371);
nand U8144 (N_8144,N_7934,N_7102);
nor U8145 (N_8145,N_7587,N_7082);
and U8146 (N_8146,N_7194,N_7793);
nand U8147 (N_8147,N_7411,N_7644);
nand U8148 (N_8148,N_7071,N_7857);
or U8149 (N_8149,N_7803,N_7882);
xnor U8150 (N_8150,N_7809,N_7504);
xor U8151 (N_8151,N_7673,N_7726);
nor U8152 (N_8152,N_7947,N_7604);
nor U8153 (N_8153,N_7366,N_7853);
or U8154 (N_8154,N_7871,N_7257);
xor U8155 (N_8155,N_7232,N_7900);
and U8156 (N_8156,N_7259,N_7058);
xor U8157 (N_8157,N_7023,N_7395);
or U8158 (N_8158,N_7909,N_7877);
xnor U8159 (N_8159,N_7707,N_7043);
xnor U8160 (N_8160,N_7817,N_7283);
or U8161 (N_8161,N_7381,N_7142);
and U8162 (N_8162,N_7470,N_7503);
nor U8163 (N_8163,N_7036,N_7858);
nor U8164 (N_8164,N_7961,N_7410);
nand U8165 (N_8165,N_7811,N_7260);
xor U8166 (N_8166,N_7390,N_7598);
nand U8167 (N_8167,N_7989,N_7373);
nor U8168 (N_8168,N_7090,N_7613);
nor U8169 (N_8169,N_7775,N_7881);
nor U8170 (N_8170,N_7356,N_7433);
or U8171 (N_8171,N_7308,N_7614);
or U8172 (N_8172,N_7117,N_7951);
nor U8173 (N_8173,N_7662,N_7507);
nand U8174 (N_8174,N_7001,N_7367);
nor U8175 (N_8175,N_7723,N_7463);
nor U8176 (N_8176,N_7702,N_7297);
nor U8177 (N_8177,N_7586,N_7740);
or U8178 (N_8178,N_7443,N_7711);
xnor U8179 (N_8179,N_7652,N_7728);
nor U8180 (N_8180,N_7781,N_7213);
or U8181 (N_8181,N_7124,N_7602);
nand U8182 (N_8182,N_7649,N_7206);
nand U8183 (N_8183,N_7663,N_7519);
and U8184 (N_8184,N_7698,N_7512);
nor U8185 (N_8185,N_7590,N_7864);
nand U8186 (N_8186,N_7359,N_7252);
or U8187 (N_8187,N_7374,N_7467);
nor U8188 (N_8188,N_7116,N_7238);
and U8189 (N_8189,N_7230,N_7713);
and U8190 (N_8190,N_7300,N_7879);
or U8191 (N_8191,N_7240,N_7760);
nor U8192 (N_8192,N_7350,N_7417);
nand U8193 (N_8193,N_7434,N_7923);
or U8194 (N_8194,N_7351,N_7908);
nor U8195 (N_8195,N_7683,N_7527);
and U8196 (N_8196,N_7149,N_7827);
xnor U8197 (N_8197,N_7901,N_7619);
xor U8198 (N_8198,N_7048,N_7941);
nand U8199 (N_8199,N_7606,N_7466);
xnor U8200 (N_8200,N_7592,N_7848);
nor U8201 (N_8201,N_7347,N_7808);
xor U8202 (N_8202,N_7762,N_7076);
nand U8203 (N_8203,N_7450,N_7513);
and U8204 (N_8204,N_7561,N_7277);
xor U8205 (N_8205,N_7891,N_7185);
xnor U8206 (N_8206,N_7137,N_7062);
nor U8207 (N_8207,N_7488,N_7717);
xnor U8208 (N_8208,N_7200,N_7958);
nor U8209 (N_8209,N_7852,N_7813);
nand U8210 (N_8210,N_7135,N_7539);
xnor U8211 (N_8211,N_7727,N_7247);
nand U8212 (N_8212,N_7840,N_7650);
xnor U8213 (N_8213,N_7536,N_7205);
xor U8214 (N_8214,N_7399,N_7892);
or U8215 (N_8215,N_7567,N_7878);
and U8216 (N_8216,N_7694,N_7299);
xnor U8217 (N_8217,N_7019,N_7268);
nor U8218 (N_8218,N_7286,N_7440);
xor U8219 (N_8219,N_7284,N_7339);
nor U8220 (N_8220,N_7148,N_7679);
nand U8221 (N_8221,N_7424,N_7386);
xor U8222 (N_8222,N_7114,N_7285);
or U8223 (N_8223,N_7884,N_7204);
nor U8224 (N_8224,N_7402,N_7121);
or U8225 (N_8225,N_7464,N_7349);
nand U8226 (N_8226,N_7875,N_7301);
and U8227 (N_8227,N_7362,N_7388);
or U8228 (N_8228,N_7943,N_7749);
nor U8229 (N_8229,N_7136,N_7012);
or U8230 (N_8230,N_7543,N_7389);
nand U8231 (N_8231,N_7033,N_7162);
xor U8232 (N_8232,N_7180,N_7954);
or U8233 (N_8233,N_7570,N_7938);
nand U8234 (N_8234,N_7092,N_7788);
nor U8235 (N_8235,N_7842,N_7787);
nor U8236 (N_8236,N_7465,N_7500);
xor U8237 (N_8237,N_7521,N_7423);
nor U8238 (N_8238,N_7225,N_7801);
nand U8239 (N_8239,N_7334,N_7846);
nor U8240 (N_8240,N_7319,N_7841);
nand U8241 (N_8241,N_7682,N_7397);
nand U8242 (N_8242,N_7758,N_7946);
nor U8243 (N_8243,N_7692,N_7967);
or U8244 (N_8244,N_7593,N_7346);
nor U8245 (N_8245,N_7083,N_7188);
xnor U8246 (N_8246,N_7295,N_7271);
nor U8247 (N_8247,N_7633,N_7418);
nand U8248 (N_8248,N_7475,N_7040);
nand U8249 (N_8249,N_7755,N_7747);
or U8250 (N_8250,N_7554,N_7477);
nor U8251 (N_8251,N_7665,N_7109);
nand U8252 (N_8252,N_7957,N_7025);
and U8253 (N_8253,N_7672,N_7765);
and U8254 (N_8254,N_7869,N_7898);
and U8255 (N_8255,N_7930,N_7321);
nor U8256 (N_8256,N_7712,N_7548);
nor U8257 (N_8257,N_7637,N_7887);
xnor U8258 (N_8258,N_7393,N_7829);
or U8259 (N_8259,N_7978,N_7820);
and U8260 (N_8260,N_7480,N_7169);
xnor U8261 (N_8261,N_7666,N_7156);
nand U8262 (N_8262,N_7669,N_7802);
nand U8263 (N_8263,N_7657,N_7626);
xor U8264 (N_8264,N_7187,N_7535);
nand U8265 (N_8265,N_7029,N_7063);
or U8266 (N_8266,N_7655,N_7056);
and U8267 (N_8267,N_7970,N_7924);
or U8268 (N_8268,N_7942,N_7520);
nor U8269 (N_8269,N_7231,N_7143);
nor U8270 (N_8270,N_7588,N_7403);
nand U8271 (N_8271,N_7933,N_7860);
nor U8272 (N_8272,N_7138,N_7981);
xnor U8273 (N_8273,N_7511,N_7153);
and U8274 (N_8274,N_7632,N_7310);
and U8275 (N_8275,N_7255,N_7214);
xnor U8276 (N_8276,N_7739,N_7172);
and U8277 (N_8277,N_7578,N_7444);
nor U8278 (N_8278,N_7401,N_7533);
or U8279 (N_8279,N_7752,N_7275);
or U8280 (N_8280,N_7080,N_7709);
and U8281 (N_8281,N_7150,N_7484);
nand U8282 (N_8282,N_7913,N_7273);
nor U8283 (N_8283,N_7883,N_7376);
nor U8284 (N_8284,N_7105,N_7856);
xor U8285 (N_8285,N_7030,N_7031);
nor U8286 (N_8286,N_7906,N_7108);
or U8287 (N_8287,N_7789,N_7243);
nand U8288 (N_8288,N_7432,N_7575);
nand U8289 (N_8289,N_7427,N_7125);
and U8290 (N_8290,N_7645,N_7994);
nor U8291 (N_8291,N_7266,N_7217);
and U8292 (N_8292,N_7676,N_7193);
xor U8293 (N_8293,N_7358,N_7107);
xor U8294 (N_8294,N_7352,N_7441);
or U8295 (N_8295,N_7568,N_7000);
xor U8296 (N_8296,N_7281,N_7660);
or U8297 (N_8297,N_7911,N_7806);
and U8298 (N_8298,N_7100,N_7822);
and U8299 (N_8299,N_7126,N_7404);
or U8300 (N_8300,N_7360,N_7544);
xor U8301 (N_8301,N_7368,N_7330);
xor U8302 (N_8302,N_7873,N_7868);
xor U8303 (N_8303,N_7131,N_7609);
nor U8304 (N_8304,N_7196,N_7218);
xnor U8305 (N_8305,N_7378,N_7807);
and U8306 (N_8306,N_7556,N_7055);
or U8307 (N_8307,N_7849,N_7348);
nor U8308 (N_8308,N_7280,N_7113);
and U8309 (N_8309,N_7847,N_7546);
or U8310 (N_8310,N_7724,N_7940);
and U8311 (N_8311,N_7725,N_7998);
nor U8312 (N_8312,N_7859,N_7253);
or U8313 (N_8313,N_7816,N_7502);
and U8314 (N_8314,N_7584,N_7499);
and U8315 (N_8315,N_7839,N_7178);
nor U8316 (N_8316,N_7224,N_7476);
xnor U8317 (N_8317,N_7618,N_7850);
nor U8318 (N_8318,N_7487,N_7832);
xor U8319 (N_8319,N_7361,N_7988);
xnor U8320 (N_8320,N_7796,N_7430);
and U8321 (N_8321,N_7050,N_7015);
and U8322 (N_8322,N_7208,N_7790);
and U8323 (N_8323,N_7084,N_7538);
nor U8324 (N_8324,N_7830,N_7643);
xnor U8325 (N_8325,N_7174,N_7294);
and U8326 (N_8326,N_7079,N_7987);
nand U8327 (N_8327,N_7099,N_7638);
nor U8328 (N_8328,N_7835,N_7550);
nor U8329 (N_8329,N_7197,N_7929);
xor U8330 (N_8330,N_7647,N_7734);
and U8331 (N_8331,N_7563,N_7215);
or U8332 (N_8332,N_7120,N_7654);
or U8333 (N_8333,N_7387,N_7750);
and U8334 (N_8334,N_7237,N_7701);
and U8335 (N_8335,N_7437,N_7515);
nand U8336 (N_8336,N_7497,N_7700);
and U8337 (N_8337,N_7498,N_7041);
and U8338 (N_8338,N_7414,N_7421);
and U8339 (N_8339,N_7101,N_7855);
nand U8340 (N_8340,N_7192,N_7469);
xnor U8341 (N_8341,N_7485,N_7603);
or U8342 (N_8342,N_7420,N_7307);
and U8343 (N_8343,N_7405,N_7945);
xor U8344 (N_8344,N_7251,N_7044);
and U8345 (N_8345,N_7674,N_7893);
or U8346 (N_8346,N_7292,N_7766);
nor U8347 (N_8347,N_7522,N_7457);
and U8348 (N_8348,N_7236,N_7944);
and U8349 (N_8349,N_7459,N_7505);
or U8350 (N_8350,N_7489,N_7605);
nand U8351 (N_8351,N_7792,N_7483);
xor U8352 (N_8352,N_7525,N_7151);
or U8353 (N_8353,N_7014,N_7780);
or U8354 (N_8354,N_7482,N_7865);
and U8355 (N_8355,N_7478,N_7577);
nand U8356 (N_8356,N_7834,N_7078);
xor U8357 (N_8357,N_7309,N_7553);
or U8358 (N_8358,N_7097,N_7689);
and U8359 (N_8359,N_7531,N_7617);
nand U8360 (N_8360,N_7680,N_7363);
or U8361 (N_8361,N_7468,N_7096);
or U8362 (N_8362,N_7034,N_7628);
nor U8363 (N_8363,N_7329,N_7235);
nor U8364 (N_8364,N_7165,N_7278);
nor U8365 (N_8365,N_7344,N_7439);
nor U8366 (N_8366,N_7571,N_7075);
nor U8367 (N_8367,N_7254,N_7962);
nor U8368 (N_8368,N_7687,N_7220);
nor U8369 (N_8369,N_7227,N_7133);
and U8370 (N_8370,N_7021,N_7610);
or U8371 (N_8371,N_7815,N_7971);
or U8372 (N_8372,N_7261,N_7331);
xor U8373 (N_8373,N_7920,N_7636);
or U8374 (N_8374,N_7242,N_7409);
xnor U8375 (N_8375,N_7999,N_7445);
or U8376 (N_8376,N_7492,N_7462);
nand U8377 (N_8377,N_7052,N_7785);
and U8378 (N_8378,N_7287,N_7937);
xnor U8379 (N_8379,N_7383,N_7705);
or U8380 (N_8380,N_7164,N_7326);
nor U8381 (N_8381,N_7656,N_7407);
xor U8382 (N_8382,N_7446,N_7005);
or U8383 (N_8383,N_7776,N_7895);
or U8384 (N_8384,N_7291,N_7828);
nand U8385 (N_8385,N_7246,N_7132);
nand U8386 (N_8386,N_7179,N_7139);
nand U8387 (N_8387,N_7714,N_7939);
or U8388 (N_8388,N_7327,N_7616);
nand U8389 (N_8389,N_7659,N_7451);
or U8390 (N_8390,N_7086,N_7851);
and U8391 (N_8391,N_7902,N_7130);
and U8392 (N_8392,N_7202,N_7262);
or U8393 (N_8393,N_7837,N_7098);
nand U8394 (N_8394,N_7303,N_7460);
nor U8395 (N_8395,N_7526,N_7342);
nand U8396 (N_8396,N_7501,N_7791);
and U8397 (N_8397,N_7751,N_7508);
or U8398 (N_8398,N_7768,N_7032);
nor U8399 (N_8399,N_7181,N_7862);
or U8400 (N_8400,N_7198,N_7491);
xor U8401 (N_8401,N_7642,N_7016);
nor U8402 (N_8402,N_7579,N_7448);
and U8403 (N_8403,N_7885,N_7991);
nand U8404 (N_8404,N_7095,N_7742);
nand U8405 (N_8405,N_7087,N_7757);
xnor U8406 (N_8406,N_7648,N_7037);
xor U8407 (N_8407,N_7710,N_7576);
and U8408 (N_8408,N_7007,N_7322);
and U8409 (N_8409,N_7804,N_7861);
nand U8410 (N_8410,N_7778,N_7863);
nand U8411 (N_8411,N_7413,N_7986);
or U8412 (N_8412,N_7372,N_7264);
nand U8413 (N_8413,N_7064,N_7068);
nand U8414 (N_8414,N_7573,N_7328);
nand U8415 (N_8415,N_7170,N_7922);
nor U8416 (N_8416,N_7134,N_7160);
nand U8417 (N_8417,N_7473,N_7671);
and U8418 (N_8418,N_7141,N_7562);
nand U8419 (N_8419,N_7795,N_7429);
or U8420 (N_8420,N_7396,N_7982);
and U8421 (N_8421,N_7782,N_7646);
nand U8422 (N_8422,N_7011,N_7651);
or U8423 (N_8423,N_7530,N_7684);
nor U8424 (N_8424,N_7611,N_7207);
or U8425 (N_8425,N_7263,N_7777);
nand U8426 (N_8426,N_7481,N_7772);
nor U8427 (N_8427,N_7997,N_7066);
nand U8428 (N_8428,N_7685,N_7552);
nor U8429 (N_8429,N_7111,N_7984);
nand U8430 (N_8430,N_7336,N_7312);
nor U8431 (N_8431,N_7155,N_7333);
xnor U8432 (N_8432,N_7729,N_7517);
xor U8433 (N_8433,N_7761,N_7748);
nand U8434 (N_8434,N_7690,N_7743);
nor U8435 (N_8435,N_7311,N_7010);
nand U8436 (N_8436,N_7681,N_7976);
nand U8437 (N_8437,N_7054,N_7239);
or U8438 (N_8438,N_7093,N_7736);
nand U8439 (N_8439,N_7289,N_7081);
nand U8440 (N_8440,N_7918,N_7783);
and U8441 (N_8441,N_7631,N_7532);
and U8442 (N_8442,N_7973,N_7675);
and U8443 (N_8443,N_7640,N_7318);
nand U8444 (N_8444,N_7779,N_7490);
nor U8445 (N_8445,N_7794,N_7744);
and U8446 (N_8446,N_7569,N_7955);
nand U8447 (N_8447,N_7279,N_7759);
xor U8448 (N_8448,N_7061,N_7896);
nand U8449 (N_8449,N_7953,N_7558);
xnor U8450 (N_8450,N_7216,N_7549);
and U8451 (N_8451,N_7990,N_7615);
or U8452 (N_8452,N_7580,N_7867);
xor U8453 (N_8453,N_7831,N_7596);
nor U8454 (N_8454,N_7964,N_7667);
and U8455 (N_8455,N_7166,N_7523);
and U8456 (N_8456,N_7357,N_7528);
xor U8457 (N_8457,N_7983,N_7833);
nand U8458 (N_8458,N_7189,N_7699);
xnor U8459 (N_8459,N_7127,N_7769);
and U8460 (N_8460,N_7369,N_7210);
and U8461 (N_8461,N_7599,N_7018);
or U8462 (N_8462,N_7600,N_7158);
and U8463 (N_8463,N_7720,N_7223);
or U8464 (N_8464,N_7716,N_7324);
nor U8465 (N_8465,N_7653,N_7741);
xor U8466 (N_8466,N_7509,N_7995);
nand U8467 (N_8467,N_7545,N_7721);
and U8468 (N_8468,N_7282,N_7147);
and U8469 (N_8469,N_7880,N_7541);
or U8470 (N_8470,N_7907,N_7977);
or U8471 (N_8471,N_7472,N_7017);
nor U8472 (N_8472,N_7004,N_7274);
nor U8473 (N_8473,N_7912,N_7323);
nor U8474 (N_8474,N_7826,N_7122);
or U8475 (N_8475,N_7927,N_7965);
and U8476 (N_8476,N_7770,N_7316);
and U8477 (N_8477,N_7996,N_7560);
or U8478 (N_8478,N_7304,N_7024);
xor U8479 (N_8479,N_7678,N_7555);
nor U8480 (N_8480,N_7936,N_7925);
nand U8481 (N_8481,N_7824,N_7693);
nor U8482 (N_8482,N_7249,N_7219);
and U8483 (N_8483,N_7866,N_7072);
nor U8484 (N_8484,N_7773,N_7733);
or U8485 (N_8485,N_7069,N_7612);
nand U8486 (N_8486,N_7191,N_7926);
xor U8487 (N_8487,N_7591,N_7935);
and U8488 (N_8488,N_7903,N_7415);
xnor U8489 (N_8489,N_7431,N_7825);
and U8490 (N_8490,N_7320,N_7540);
or U8491 (N_8491,N_7621,N_7844);
xor U8492 (N_8492,N_7992,N_7375);
nand U8493 (N_8493,N_7756,N_7818);
xor U8494 (N_8494,N_7932,N_7629);
or U8495 (N_8495,N_7630,N_7340);
xor U8496 (N_8496,N_7256,N_7343);
or U8497 (N_8497,N_7607,N_7966);
nor U8498 (N_8498,N_7771,N_7222);
nor U8499 (N_8499,N_7529,N_7872);
xnor U8500 (N_8500,N_7501,N_7460);
xor U8501 (N_8501,N_7324,N_7818);
or U8502 (N_8502,N_7795,N_7837);
xnor U8503 (N_8503,N_7848,N_7750);
and U8504 (N_8504,N_7419,N_7783);
xor U8505 (N_8505,N_7566,N_7558);
xor U8506 (N_8506,N_7795,N_7117);
nand U8507 (N_8507,N_7450,N_7317);
nand U8508 (N_8508,N_7111,N_7083);
or U8509 (N_8509,N_7988,N_7840);
nor U8510 (N_8510,N_7158,N_7457);
xnor U8511 (N_8511,N_7123,N_7266);
xnor U8512 (N_8512,N_7902,N_7400);
nand U8513 (N_8513,N_7925,N_7502);
xnor U8514 (N_8514,N_7835,N_7331);
nand U8515 (N_8515,N_7276,N_7240);
nor U8516 (N_8516,N_7847,N_7407);
and U8517 (N_8517,N_7701,N_7594);
xnor U8518 (N_8518,N_7507,N_7247);
or U8519 (N_8519,N_7686,N_7582);
nor U8520 (N_8520,N_7154,N_7391);
nand U8521 (N_8521,N_7358,N_7509);
nand U8522 (N_8522,N_7968,N_7973);
xor U8523 (N_8523,N_7481,N_7638);
or U8524 (N_8524,N_7939,N_7444);
nor U8525 (N_8525,N_7078,N_7404);
and U8526 (N_8526,N_7840,N_7597);
xnor U8527 (N_8527,N_7865,N_7750);
and U8528 (N_8528,N_7939,N_7960);
nand U8529 (N_8529,N_7447,N_7994);
or U8530 (N_8530,N_7155,N_7291);
xor U8531 (N_8531,N_7089,N_7612);
nor U8532 (N_8532,N_7497,N_7817);
nor U8533 (N_8533,N_7874,N_7619);
and U8534 (N_8534,N_7378,N_7012);
and U8535 (N_8535,N_7775,N_7056);
or U8536 (N_8536,N_7242,N_7365);
or U8537 (N_8537,N_7589,N_7577);
nor U8538 (N_8538,N_7053,N_7170);
and U8539 (N_8539,N_7569,N_7564);
nand U8540 (N_8540,N_7019,N_7904);
nand U8541 (N_8541,N_7358,N_7013);
nand U8542 (N_8542,N_7650,N_7015);
xnor U8543 (N_8543,N_7256,N_7980);
nor U8544 (N_8544,N_7704,N_7180);
xnor U8545 (N_8545,N_7029,N_7128);
or U8546 (N_8546,N_7545,N_7419);
or U8547 (N_8547,N_7509,N_7066);
and U8548 (N_8548,N_7754,N_7370);
nand U8549 (N_8549,N_7900,N_7649);
or U8550 (N_8550,N_7707,N_7188);
and U8551 (N_8551,N_7805,N_7597);
nand U8552 (N_8552,N_7217,N_7825);
or U8553 (N_8553,N_7405,N_7542);
xor U8554 (N_8554,N_7863,N_7209);
and U8555 (N_8555,N_7623,N_7979);
nand U8556 (N_8556,N_7451,N_7384);
xor U8557 (N_8557,N_7120,N_7376);
xnor U8558 (N_8558,N_7100,N_7970);
xnor U8559 (N_8559,N_7776,N_7546);
xnor U8560 (N_8560,N_7955,N_7521);
nand U8561 (N_8561,N_7181,N_7821);
xor U8562 (N_8562,N_7679,N_7604);
nand U8563 (N_8563,N_7946,N_7146);
xor U8564 (N_8564,N_7269,N_7180);
xnor U8565 (N_8565,N_7404,N_7249);
nand U8566 (N_8566,N_7703,N_7431);
or U8567 (N_8567,N_7770,N_7689);
and U8568 (N_8568,N_7622,N_7690);
and U8569 (N_8569,N_7683,N_7649);
nand U8570 (N_8570,N_7315,N_7318);
xnor U8571 (N_8571,N_7606,N_7460);
or U8572 (N_8572,N_7486,N_7755);
xor U8573 (N_8573,N_7694,N_7202);
or U8574 (N_8574,N_7290,N_7282);
nor U8575 (N_8575,N_7669,N_7038);
nand U8576 (N_8576,N_7657,N_7123);
nand U8577 (N_8577,N_7580,N_7221);
nand U8578 (N_8578,N_7115,N_7174);
or U8579 (N_8579,N_7216,N_7587);
xnor U8580 (N_8580,N_7681,N_7634);
or U8581 (N_8581,N_7719,N_7538);
or U8582 (N_8582,N_7127,N_7613);
or U8583 (N_8583,N_7447,N_7661);
or U8584 (N_8584,N_7567,N_7353);
and U8585 (N_8585,N_7856,N_7149);
nand U8586 (N_8586,N_7337,N_7241);
xor U8587 (N_8587,N_7583,N_7528);
or U8588 (N_8588,N_7867,N_7705);
or U8589 (N_8589,N_7638,N_7696);
nand U8590 (N_8590,N_7787,N_7798);
and U8591 (N_8591,N_7090,N_7440);
nand U8592 (N_8592,N_7505,N_7432);
or U8593 (N_8593,N_7145,N_7620);
nand U8594 (N_8594,N_7724,N_7115);
and U8595 (N_8595,N_7626,N_7865);
and U8596 (N_8596,N_7801,N_7697);
nor U8597 (N_8597,N_7531,N_7209);
or U8598 (N_8598,N_7835,N_7392);
nor U8599 (N_8599,N_7508,N_7637);
xnor U8600 (N_8600,N_7462,N_7898);
or U8601 (N_8601,N_7849,N_7323);
nand U8602 (N_8602,N_7910,N_7941);
nand U8603 (N_8603,N_7600,N_7292);
or U8604 (N_8604,N_7359,N_7413);
and U8605 (N_8605,N_7419,N_7520);
nor U8606 (N_8606,N_7287,N_7404);
xnor U8607 (N_8607,N_7550,N_7538);
or U8608 (N_8608,N_7256,N_7670);
and U8609 (N_8609,N_7889,N_7227);
or U8610 (N_8610,N_7794,N_7532);
nand U8611 (N_8611,N_7162,N_7836);
xnor U8612 (N_8612,N_7580,N_7885);
or U8613 (N_8613,N_7084,N_7316);
nand U8614 (N_8614,N_7299,N_7972);
nand U8615 (N_8615,N_7443,N_7108);
and U8616 (N_8616,N_7816,N_7443);
and U8617 (N_8617,N_7528,N_7750);
or U8618 (N_8618,N_7282,N_7998);
and U8619 (N_8619,N_7144,N_7063);
and U8620 (N_8620,N_7371,N_7127);
xor U8621 (N_8621,N_7620,N_7994);
and U8622 (N_8622,N_7056,N_7836);
nand U8623 (N_8623,N_7596,N_7682);
nor U8624 (N_8624,N_7330,N_7385);
xnor U8625 (N_8625,N_7653,N_7397);
or U8626 (N_8626,N_7352,N_7791);
and U8627 (N_8627,N_7632,N_7045);
xnor U8628 (N_8628,N_7934,N_7993);
nor U8629 (N_8629,N_7375,N_7352);
and U8630 (N_8630,N_7794,N_7665);
nor U8631 (N_8631,N_7547,N_7415);
xor U8632 (N_8632,N_7732,N_7751);
nor U8633 (N_8633,N_7900,N_7277);
xnor U8634 (N_8634,N_7404,N_7181);
nor U8635 (N_8635,N_7878,N_7176);
xnor U8636 (N_8636,N_7828,N_7152);
nor U8637 (N_8637,N_7846,N_7776);
xor U8638 (N_8638,N_7789,N_7445);
or U8639 (N_8639,N_7626,N_7110);
or U8640 (N_8640,N_7152,N_7629);
nand U8641 (N_8641,N_7311,N_7264);
nor U8642 (N_8642,N_7712,N_7184);
nor U8643 (N_8643,N_7529,N_7010);
nand U8644 (N_8644,N_7343,N_7372);
xnor U8645 (N_8645,N_7310,N_7140);
nor U8646 (N_8646,N_7954,N_7541);
nand U8647 (N_8647,N_7520,N_7704);
or U8648 (N_8648,N_7934,N_7888);
and U8649 (N_8649,N_7562,N_7026);
xor U8650 (N_8650,N_7313,N_7108);
nor U8651 (N_8651,N_7163,N_7622);
or U8652 (N_8652,N_7130,N_7675);
nor U8653 (N_8653,N_7274,N_7183);
and U8654 (N_8654,N_7621,N_7208);
xor U8655 (N_8655,N_7583,N_7974);
nand U8656 (N_8656,N_7484,N_7180);
nor U8657 (N_8657,N_7827,N_7456);
and U8658 (N_8658,N_7346,N_7952);
or U8659 (N_8659,N_7696,N_7352);
nor U8660 (N_8660,N_7799,N_7648);
or U8661 (N_8661,N_7915,N_7418);
nand U8662 (N_8662,N_7900,N_7613);
xor U8663 (N_8663,N_7358,N_7526);
nand U8664 (N_8664,N_7168,N_7878);
or U8665 (N_8665,N_7922,N_7783);
xnor U8666 (N_8666,N_7816,N_7984);
or U8667 (N_8667,N_7573,N_7667);
xor U8668 (N_8668,N_7617,N_7169);
nor U8669 (N_8669,N_7062,N_7566);
or U8670 (N_8670,N_7313,N_7163);
xor U8671 (N_8671,N_7776,N_7544);
nor U8672 (N_8672,N_7352,N_7914);
or U8673 (N_8673,N_7703,N_7865);
nand U8674 (N_8674,N_7879,N_7031);
nand U8675 (N_8675,N_7487,N_7798);
nand U8676 (N_8676,N_7697,N_7640);
nand U8677 (N_8677,N_7001,N_7672);
xnor U8678 (N_8678,N_7435,N_7626);
and U8679 (N_8679,N_7908,N_7909);
or U8680 (N_8680,N_7238,N_7244);
and U8681 (N_8681,N_7841,N_7152);
xnor U8682 (N_8682,N_7717,N_7048);
nand U8683 (N_8683,N_7992,N_7956);
xnor U8684 (N_8684,N_7364,N_7581);
nand U8685 (N_8685,N_7634,N_7373);
nand U8686 (N_8686,N_7692,N_7784);
nand U8687 (N_8687,N_7407,N_7618);
xnor U8688 (N_8688,N_7259,N_7638);
and U8689 (N_8689,N_7182,N_7824);
nand U8690 (N_8690,N_7957,N_7509);
and U8691 (N_8691,N_7381,N_7203);
xnor U8692 (N_8692,N_7490,N_7397);
nor U8693 (N_8693,N_7453,N_7491);
nand U8694 (N_8694,N_7985,N_7755);
xnor U8695 (N_8695,N_7924,N_7285);
or U8696 (N_8696,N_7594,N_7615);
nand U8697 (N_8697,N_7319,N_7105);
nor U8698 (N_8698,N_7461,N_7921);
nor U8699 (N_8699,N_7574,N_7552);
nor U8700 (N_8700,N_7281,N_7341);
nand U8701 (N_8701,N_7038,N_7784);
and U8702 (N_8702,N_7280,N_7310);
and U8703 (N_8703,N_7465,N_7573);
or U8704 (N_8704,N_7335,N_7698);
nor U8705 (N_8705,N_7538,N_7385);
xor U8706 (N_8706,N_7400,N_7654);
and U8707 (N_8707,N_7112,N_7188);
nand U8708 (N_8708,N_7017,N_7683);
nor U8709 (N_8709,N_7281,N_7616);
and U8710 (N_8710,N_7544,N_7689);
nor U8711 (N_8711,N_7735,N_7659);
nor U8712 (N_8712,N_7374,N_7732);
nor U8713 (N_8713,N_7313,N_7282);
xnor U8714 (N_8714,N_7523,N_7384);
or U8715 (N_8715,N_7804,N_7867);
nor U8716 (N_8716,N_7915,N_7264);
nand U8717 (N_8717,N_7048,N_7568);
and U8718 (N_8718,N_7610,N_7801);
or U8719 (N_8719,N_7323,N_7350);
and U8720 (N_8720,N_7445,N_7365);
nor U8721 (N_8721,N_7115,N_7336);
nor U8722 (N_8722,N_7368,N_7060);
xnor U8723 (N_8723,N_7186,N_7583);
or U8724 (N_8724,N_7299,N_7425);
nor U8725 (N_8725,N_7634,N_7124);
nor U8726 (N_8726,N_7067,N_7018);
and U8727 (N_8727,N_7019,N_7646);
nor U8728 (N_8728,N_7472,N_7324);
nand U8729 (N_8729,N_7662,N_7438);
xnor U8730 (N_8730,N_7881,N_7921);
nor U8731 (N_8731,N_7246,N_7520);
nor U8732 (N_8732,N_7889,N_7336);
or U8733 (N_8733,N_7766,N_7885);
or U8734 (N_8734,N_7212,N_7270);
or U8735 (N_8735,N_7357,N_7813);
nand U8736 (N_8736,N_7727,N_7781);
nor U8737 (N_8737,N_7672,N_7044);
and U8738 (N_8738,N_7313,N_7863);
or U8739 (N_8739,N_7428,N_7437);
nor U8740 (N_8740,N_7326,N_7308);
xnor U8741 (N_8741,N_7418,N_7801);
or U8742 (N_8742,N_7865,N_7485);
nand U8743 (N_8743,N_7428,N_7523);
nor U8744 (N_8744,N_7305,N_7405);
or U8745 (N_8745,N_7466,N_7400);
nand U8746 (N_8746,N_7619,N_7764);
or U8747 (N_8747,N_7886,N_7853);
xnor U8748 (N_8748,N_7502,N_7376);
nor U8749 (N_8749,N_7387,N_7258);
or U8750 (N_8750,N_7128,N_7501);
nand U8751 (N_8751,N_7546,N_7650);
or U8752 (N_8752,N_7653,N_7717);
xor U8753 (N_8753,N_7041,N_7485);
or U8754 (N_8754,N_7063,N_7211);
xnor U8755 (N_8755,N_7189,N_7128);
nand U8756 (N_8756,N_7571,N_7343);
xnor U8757 (N_8757,N_7713,N_7574);
xor U8758 (N_8758,N_7003,N_7448);
xor U8759 (N_8759,N_7445,N_7582);
and U8760 (N_8760,N_7420,N_7143);
xnor U8761 (N_8761,N_7525,N_7232);
or U8762 (N_8762,N_7477,N_7108);
nor U8763 (N_8763,N_7959,N_7688);
nor U8764 (N_8764,N_7899,N_7415);
xor U8765 (N_8765,N_7442,N_7046);
nor U8766 (N_8766,N_7392,N_7432);
nor U8767 (N_8767,N_7025,N_7094);
nor U8768 (N_8768,N_7689,N_7688);
or U8769 (N_8769,N_7446,N_7673);
and U8770 (N_8770,N_7155,N_7825);
or U8771 (N_8771,N_7633,N_7803);
nor U8772 (N_8772,N_7763,N_7927);
or U8773 (N_8773,N_7529,N_7265);
nor U8774 (N_8774,N_7053,N_7832);
nor U8775 (N_8775,N_7886,N_7239);
nand U8776 (N_8776,N_7442,N_7402);
nand U8777 (N_8777,N_7173,N_7146);
nand U8778 (N_8778,N_7507,N_7080);
nor U8779 (N_8779,N_7215,N_7526);
nor U8780 (N_8780,N_7016,N_7540);
nor U8781 (N_8781,N_7993,N_7463);
or U8782 (N_8782,N_7071,N_7970);
nand U8783 (N_8783,N_7769,N_7748);
nor U8784 (N_8784,N_7583,N_7918);
xor U8785 (N_8785,N_7169,N_7592);
nor U8786 (N_8786,N_7849,N_7547);
and U8787 (N_8787,N_7821,N_7071);
nand U8788 (N_8788,N_7054,N_7594);
and U8789 (N_8789,N_7017,N_7529);
nor U8790 (N_8790,N_7991,N_7316);
and U8791 (N_8791,N_7306,N_7950);
xnor U8792 (N_8792,N_7623,N_7661);
and U8793 (N_8793,N_7826,N_7302);
or U8794 (N_8794,N_7969,N_7424);
xnor U8795 (N_8795,N_7996,N_7746);
nor U8796 (N_8796,N_7901,N_7351);
nand U8797 (N_8797,N_7247,N_7229);
xor U8798 (N_8798,N_7188,N_7682);
or U8799 (N_8799,N_7079,N_7140);
or U8800 (N_8800,N_7811,N_7589);
xnor U8801 (N_8801,N_7924,N_7726);
xor U8802 (N_8802,N_7777,N_7500);
nand U8803 (N_8803,N_7851,N_7528);
and U8804 (N_8804,N_7827,N_7782);
xor U8805 (N_8805,N_7988,N_7781);
and U8806 (N_8806,N_7807,N_7465);
and U8807 (N_8807,N_7922,N_7060);
xor U8808 (N_8808,N_7767,N_7315);
and U8809 (N_8809,N_7596,N_7311);
xnor U8810 (N_8810,N_7564,N_7222);
nand U8811 (N_8811,N_7250,N_7621);
nor U8812 (N_8812,N_7855,N_7302);
and U8813 (N_8813,N_7773,N_7637);
nor U8814 (N_8814,N_7294,N_7433);
nor U8815 (N_8815,N_7154,N_7012);
nor U8816 (N_8816,N_7695,N_7792);
nand U8817 (N_8817,N_7986,N_7257);
nor U8818 (N_8818,N_7882,N_7861);
xnor U8819 (N_8819,N_7913,N_7686);
nor U8820 (N_8820,N_7338,N_7848);
and U8821 (N_8821,N_7445,N_7844);
or U8822 (N_8822,N_7315,N_7184);
and U8823 (N_8823,N_7287,N_7437);
and U8824 (N_8824,N_7211,N_7516);
and U8825 (N_8825,N_7039,N_7131);
or U8826 (N_8826,N_7919,N_7772);
or U8827 (N_8827,N_7038,N_7284);
xnor U8828 (N_8828,N_7949,N_7948);
nor U8829 (N_8829,N_7360,N_7178);
nor U8830 (N_8830,N_7955,N_7812);
and U8831 (N_8831,N_7119,N_7095);
nor U8832 (N_8832,N_7131,N_7525);
nand U8833 (N_8833,N_7481,N_7751);
xor U8834 (N_8834,N_7301,N_7682);
nor U8835 (N_8835,N_7284,N_7041);
nand U8836 (N_8836,N_7398,N_7976);
xnor U8837 (N_8837,N_7861,N_7850);
nand U8838 (N_8838,N_7546,N_7596);
nor U8839 (N_8839,N_7409,N_7349);
and U8840 (N_8840,N_7226,N_7293);
nand U8841 (N_8841,N_7939,N_7926);
nor U8842 (N_8842,N_7571,N_7111);
xnor U8843 (N_8843,N_7150,N_7659);
or U8844 (N_8844,N_7577,N_7551);
or U8845 (N_8845,N_7035,N_7763);
nand U8846 (N_8846,N_7919,N_7412);
nand U8847 (N_8847,N_7505,N_7974);
and U8848 (N_8848,N_7868,N_7445);
xnor U8849 (N_8849,N_7280,N_7472);
nor U8850 (N_8850,N_7814,N_7290);
nor U8851 (N_8851,N_7930,N_7842);
nand U8852 (N_8852,N_7741,N_7237);
xnor U8853 (N_8853,N_7945,N_7713);
or U8854 (N_8854,N_7649,N_7748);
xnor U8855 (N_8855,N_7977,N_7261);
xor U8856 (N_8856,N_7426,N_7636);
nand U8857 (N_8857,N_7409,N_7715);
nand U8858 (N_8858,N_7555,N_7472);
nand U8859 (N_8859,N_7808,N_7981);
and U8860 (N_8860,N_7173,N_7495);
xor U8861 (N_8861,N_7115,N_7280);
xor U8862 (N_8862,N_7339,N_7081);
xnor U8863 (N_8863,N_7917,N_7906);
nand U8864 (N_8864,N_7856,N_7075);
nand U8865 (N_8865,N_7508,N_7633);
and U8866 (N_8866,N_7664,N_7387);
or U8867 (N_8867,N_7211,N_7257);
nand U8868 (N_8868,N_7963,N_7083);
and U8869 (N_8869,N_7638,N_7036);
xor U8870 (N_8870,N_7097,N_7073);
and U8871 (N_8871,N_7047,N_7222);
and U8872 (N_8872,N_7225,N_7014);
or U8873 (N_8873,N_7244,N_7336);
and U8874 (N_8874,N_7933,N_7791);
nand U8875 (N_8875,N_7027,N_7552);
and U8876 (N_8876,N_7160,N_7741);
nand U8877 (N_8877,N_7305,N_7611);
nand U8878 (N_8878,N_7732,N_7087);
xnor U8879 (N_8879,N_7884,N_7642);
or U8880 (N_8880,N_7159,N_7399);
xor U8881 (N_8881,N_7375,N_7850);
xnor U8882 (N_8882,N_7882,N_7237);
and U8883 (N_8883,N_7457,N_7252);
or U8884 (N_8884,N_7195,N_7353);
nand U8885 (N_8885,N_7197,N_7467);
xor U8886 (N_8886,N_7909,N_7491);
nor U8887 (N_8887,N_7540,N_7463);
and U8888 (N_8888,N_7443,N_7461);
and U8889 (N_8889,N_7037,N_7303);
nor U8890 (N_8890,N_7937,N_7794);
nor U8891 (N_8891,N_7005,N_7277);
nor U8892 (N_8892,N_7746,N_7138);
nor U8893 (N_8893,N_7089,N_7866);
nand U8894 (N_8894,N_7603,N_7913);
nor U8895 (N_8895,N_7799,N_7668);
nand U8896 (N_8896,N_7256,N_7940);
xnor U8897 (N_8897,N_7303,N_7892);
xnor U8898 (N_8898,N_7620,N_7290);
nor U8899 (N_8899,N_7703,N_7808);
nor U8900 (N_8900,N_7703,N_7237);
or U8901 (N_8901,N_7305,N_7357);
and U8902 (N_8902,N_7359,N_7831);
and U8903 (N_8903,N_7660,N_7143);
nor U8904 (N_8904,N_7952,N_7320);
nand U8905 (N_8905,N_7921,N_7653);
or U8906 (N_8906,N_7349,N_7519);
nor U8907 (N_8907,N_7349,N_7437);
or U8908 (N_8908,N_7576,N_7080);
or U8909 (N_8909,N_7611,N_7998);
nand U8910 (N_8910,N_7088,N_7670);
xnor U8911 (N_8911,N_7631,N_7297);
nand U8912 (N_8912,N_7455,N_7592);
nor U8913 (N_8913,N_7308,N_7957);
nor U8914 (N_8914,N_7874,N_7847);
nor U8915 (N_8915,N_7903,N_7554);
and U8916 (N_8916,N_7946,N_7524);
or U8917 (N_8917,N_7698,N_7184);
or U8918 (N_8918,N_7924,N_7006);
nor U8919 (N_8919,N_7079,N_7292);
nand U8920 (N_8920,N_7688,N_7910);
or U8921 (N_8921,N_7450,N_7831);
and U8922 (N_8922,N_7979,N_7572);
nor U8923 (N_8923,N_7659,N_7879);
nor U8924 (N_8924,N_7359,N_7759);
nand U8925 (N_8925,N_7259,N_7082);
nand U8926 (N_8926,N_7377,N_7608);
and U8927 (N_8927,N_7375,N_7465);
or U8928 (N_8928,N_7802,N_7154);
and U8929 (N_8929,N_7956,N_7507);
and U8930 (N_8930,N_7311,N_7393);
and U8931 (N_8931,N_7195,N_7295);
nor U8932 (N_8932,N_7281,N_7975);
nand U8933 (N_8933,N_7935,N_7128);
nor U8934 (N_8934,N_7493,N_7442);
and U8935 (N_8935,N_7264,N_7459);
xnor U8936 (N_8936,N_7341,N_7514);
and U8937 (N_8937,N_7963,N_7304);
nand U8938 (N_8938,N_7151,N_7402);
nor U8939 (N_8939,N_7672,N_7974);
and U8940 (N_8940,N_7183,N_7105);
nand U8941 (N_8941,N_7968,N_7080);
xnor U8942 (N_8942,N_7499,N_7692);
and U8943 (N_8943,N_7708,N_7402);
or U8944 (N_8944,N_7519,N_7723);
or U8945 (N_8945,N_7352,N_7403);
nand U8946 (N_8946,N_7378,N_7753);
nand U8947 (N_8947,N_7515,N_7983);
nor U8948 (N_8948,N_7529,N_7620);
or U8949 (N_8949,N_7468,N_7205);
or U8950 (N_8950,N_7046,N_7060);
or U8951 (N_8951,N_7401,N_7550);
nand U8952 (N_8952,N_7437,N_7247);
nor U8953 (N_8953,N_7124,N_7484);
xor U8954 (N_8954,N_7863,N_7753);
nand U8955 (N_8955,N_7546,N_7203);
or U8956 (N_8956,N_7368,N_7749);
xnor U8957 (N_8957,N_7000,N_7593);
xor U8958 (N_8958,N_7517,N_7858);
xor U8959 (N_8959,N_7417,N_7237);
xnor U8960 (N_8960,N_7592,N_7362);
nor U8961 (N_8961,N_7115,N_7519);
nor U8962 (N_8962,N_7315,N_7899);
xor U8963 (N_8963,N_7849,N_7554);
and U8964 (N_8964,N_7999,N_7663);
or U8965 (N_8965,N_7701,N_7498);
xor U8966 (N_8966,N_7253,N_7359);
nor U8967 (N_8967,N_7729,N_7659);
or U8968 (N_8968,N_7492,N_7387);
nand U8969 (N_8969,N_7388,N_7669);
or U8970 (N_8970,N_7166,N_7096);
xor U8971 (N_8971,N_7822,N_7402);
nor U8972 (N_8972,N_7967,N_7884);
nand U8973 (N_8973,N_7463,N_7188);
and U8974 (N_8974,N_7732,N_7848);
xnor U8975 (N_8975,N_7574,N_7160);
and U8976 (N_8976,N_7850,N_7780);
nor U8977 (N_8977,N_7622,N_7140);
xnor U8978 (N_8978,N_7408,N_7844);
nor U8979 (N_8979,N_7333,N_7343);
xor U8980 (N_8980,N_7767,N_7492);
and U8981 (N_8981,N_7259,N_7888);
and U8982 (N_8982,N_7671,N_7672);
nand U8983 (N_8983,N_7735,N_7533);
or U8984 (N_8984,N_7003,N_7627);
xor U8985 (N_8985,N_7208,N_7091);
or U8986 (N_8986,N_7303,N_7017);
xor U8987 (N_8987,N_7859,N_7411);
nand U8988 (N_8988,N_7694,N_7562);
nand U8989 (N_8989,N_7962,N_7039);
xor U8990 (N_8990,N_7943,N_7289);
or U8991 (N_8991,N_7115,N_7866);
xnor U8992 (N_8992,N_7341,N_7605);
or U8993 (N_8993,N_7402,N_7203);
and U8994 (N_8994,N_7203,N_7732);
xnor U8995 (N_8995,N_7230,N_7762);
nand U8996 (N_8996,N_7912,N_7296);
xor U8997 (N_8997,N_7514,N_7405);
and U8998 (N_8998,N_7970,N_7948);
nor U8999 (N_8999,N_7009,N_7773);
xnor U9000 (N_9000,N_8288,N_8290);
nand U9001 (N_9001,N_8164,N_8285);
or U9002 (N_9002,N_8108,N_8435);
and U9003 (N_9003,N_8217,N_8909);
and U9004 (N_9004,N_8201,N_8843);
or U9005 (N_9005,N_8536,N_8558);
and U9006 (N_9006,N_8944,N_8351);
nand U9007 (N_9007,N_8865,N_8762);
nand U9008 (N_9008,N_8325,N_8141);
or U9009 (N_9009,N_8896,N_8229);
or U9010 (N_9010,N_8583,N_8265);
and U9011 (N_9011,N_8375,N_8993);
xnor U9012 (N_9012,N_8406,N_8342);
nand U9013 (N_9013,N_8639,N_8304);
nand U9014 (N_9014,N_8115,N_8739);
nor U9015 (N_9015,N_8580,N_8082);
nand U9016 (N_9016,N_8198,N_8291);
and U9017 (N_9017,N_8356,N_8619);
nand U9018 (N_9018,N_8233,N_8034);
nor U9019 (N_9019,N_8565,N_8885);
or U9020 (N_9020,N_8972,N_8617);
or U9021 (N_9021,N_8299,N_8818);
nor U9022 (N_9022,N_8344,N_8743);
or U9023 (N_9023,N_8939,N_8677);
nor U9024 (N_9024,N_8365,N_8220);
and U9025 (N_9025,N_8432,N_8471);
or U9026 (N_9026,N_8576,N_8110);
nand U9027 (N_9027,N_8995,N_8402);
or U9028 (N_9028,N_8457,N_8231);
xor U9029 (N_9029,N_8815,N_8609);
or U9030 (N_9030,N_8292,N_8400);
or U9031 (N_9031,N_8200,N_8641);
nand U9032 (N_9032,N_8712,N_8856);
or U9033 (N_9033,N_8537,N_8538);
nand U9034 (N_9034,N_8685,N_8530);
nand U9035 (N_9035,N_8914,N_8343);
nand U9036 (N_9036,N_8690,N_8149);
nand U9037 (N_9037,N_8611,N_8479);
xnor U9038 (N_9038,N_8173,N_8938);
nor U9039 (N_9039,N_8066,N_8785);
nand U9040 (N_9040,N_8635,N_8737);
or U9041 (N_9041,N_8973,N_8429);
and U9042 (N_9042,N_8262,N_8236);
xor U9043 (N_9043,N_8545,N_8563);
and U9044 (N_9044,N_8323,N_8372);
nand U9045 (N_9045,N_8509,N_8297);
and U9046 (N_9046,N_8513,N_8741);
and U9047 (N_9047,N_8651,N_8336);
nor U9048 (N_9048,N_8936,N_8780);
xor U9049 (N_9049,N_8599,N_8753);
and U9050 (N_9050,N_8086,N_8531);
or U9051 (N_9051,N_8003,N_8393);
and U9052 (N_9052,N_8459,N_8966);
xor U9053 (N_9053,N_8187,N_8933);
or U9054 (N_9054,N_8355,N_8757);
nand U9055 (N_9055,N_8409,N_8898);
nor U9056 (N_9056,N_8455,N_8915);
nor U9057 (N_9057,N_8584,N_8386);
and U9058 (N_9058,N_8508,N_8042);
or U9059 (N_9059,N_8259,N_8610);
xnor U9060 (N_9060,N_8771,N_8642);
or U9061 (N_9061,N_8997,N_8729);
xor U9062 (N_9062,N_8602,N_8812);
or U9063 (N_9063,N_8495,N_8489);
nand U9064 (N_9064,N_8860,N_8855);
xnor U9065 (N_9065,N_8051,N_8965);
nand U9066 (N_9066,N_8632,N_8474);
nand U9067 (N_9067,N_8458,N_8060);
xnor U9068 (N_9068,N_8048,N_8614);
xnor U9069 (N_9069,N_8983,N_8722);
or U9070 (N_9070,N_8691,N_8601);
or U9071 (N_9071,N_8329,N_8660);
and U9072 (N_9072,N_8674,N_8624);
nand U9073 (N_9073,N_8745,N_8572);
nor U9074 (N_9074,N_8512,N_8100);
nand U9075 (N_9075,N_8013,N_8475);
nor U9076 (N_9076,N_8961,N_8267);
nand U9077 (N_9077,N_8181,N_8831);
or U9078 (N_9078,N_8647,N_8129);
nor U9079 (N_9079,N_8925,N_8077);
nand U9080 (N_9080,N_8974,N_8184);
or U9081 (N_9081,N_8932,N_8261);
nor U9082 (N_9082,N_8754,N_8358);
or U9083 (N_9083,N_8162,N_8283);
xnor U9084 (N_9084,N_8247,N_8571);
nand U9085 (N_9085,N_8850,N_8018);
nand U9086 (N_9086,N_8946,N_8121);
and U9087 (N_9087,N_8269,N_8466);
nor U9088 (N_9088,N_8353,N_8485);
and U9089 (N_9089,N_8152,N_8874);
xor U9090 (N_9090,N_8561,N_8151);
xnor U9091 (N_9091,N_8190,N_8582);
nand U9092 (N_9092,N_8235,N_8258);
nand U9093 (N_9093,N_8085,N_8234);
or U9094 (N_9094,N_8649,N_8067);
nand U9095 (N_9095,N_8721,N_8410);
nand U9096 (N_9096,N_8011,N_8643);
xor U9097 (N_9097,N_8431,N_8954);
xor U9098 (N_9098,N_8315,N_8543);
nor U9099 (N_9099,N_8811,N_8695);
nor U9100 (N_9100,N_8046,N_8989);
xor U9101 (N_9101,N_8652,N_8775);
or U9102 (N_9102,N_8532,N_8055);
nand U9103 (N_9103,N_8730,N_8628);
and U9104 (N_9104,N_8109,N_8027);
or U9105 (N_9105,N_8442,N_8986);
nor U9106 (N_9106,N_8472,N_8560);
nor U9107 (N_9107,N_8196,N_8090);
nor U9108 (N_9108,N_8706,N_8581);
and U9109 (N_9109,N_8056,N_8021);
or U9110 (N_9110,N_8408,N_8862);
xor U9111 (N_9111,N_8907,N_8819);
xnor U9112 (N_9112,N_8963,N_8123);
xor U9113 (N_9113,N_8985,N_8370);
and U9114 (N_9114,N_8881,N_8371);
nand U9115 (N_9115,N_8703,N_8126);
nand U9116 (N_9116,N_8585,N_8145);
and U9117 (N_9117,N_8125,N_8140);
xor U9118 (N_9118,N_8595,N_8394);
xor U9119 (N_9119,N_8878,N_8089);
or U9120 (N_9120,N_8945,N_8096);
nand U9121 (N_9121,N_8764,N_8675);
xor U9122 (N_9122,N_8491,N_8071);
xor U9123 (N_9123,N_8988,N_8636);
and U9124 (N_9124,N_8822,N_8147);
and U9125 (N_9125,N_8070,N_8788);
or U9126 (N_9126,N_8888,N_8622);
xnor U9127 (N_9127,N_8063,N_8990);
xor U9128 (N_9128,N_8700,N_8923);
or U9129 (N_9129,N_8903,N_8734);
xnor U9130 (N_9130,N_8931,N_8367);
nor U9131 (N_9131,N_8176,N_8807);
and U9132 (N_9132,N_8303,N_8648);
nor U9133 (N_9133,N_8423,N_8310);
and U9134 (N_9134,N_8248,N_8994);
or U9135 (N_9135,N_8237,N_8550);
and U9136 (N_9136,N_8593,N_8638);
or U9137 (N_9137,N_8270,N_8287);
xnor U9138 (N_9138,N_8332,N_8701);
nor U9139 (N_9139,N_8710,N_8156);
xnor U9140 (N_9140,N_8801,N_8163);
or U9141 (N_9141,N_8094,N_8964);
nand U9142 (N_9142,N_8767,N_8518);
and U9143 (N_9143,N_8520,N_8752);
and U9144 (N_9144,N_8028,N_8135);
xnor U9145 (N_9145,N_8943,N_8481);
nand U9146 (N_9146,N_8037,N_8742);
nor U9147 (N_9147,N_8437,N_8180);
xor U9148 (N_9148,N_8846,N_8553);
or U9149 (N_9149,N_8864,N_8918);
xnor U9150 (N_9150,N_8068,N_8792);
or U9151 (N_9151,N_8340,N_8655);
nand U9152 (N_9152,N_8047,N_8033);
or U9153 (N_9153,N_8894,N_8454);
or U9154 (N_9154,N_8620,N_8319);
nor U9155 (N_9155,N_8260,N_8482);
nand U9156 (N_9156,N_8391,N_8249);
and U9157 (N_9157,N_8820,N_8646);
or U9158 (N_9158,N_8924,N_8694);
and U9159 (N_9159,N_8806,N_8373);
nand U9160 (N_9160,N_8656,N_8146);
xor U9161 (N_9161,N_8362,N_8523);
xnor U9162 (N_9162,N_8460,N_8566);
xor U9163 (N_9163,N_8369,N_8004);
and U9164 (N_9164,N_8879,N_8746);
xor U9165 (N_9165,N_8594,N_8257);
and U9166 (N_9166,N_8240,N_8616);
and U9167 (N_9167,N_8511,N_8547);
xor U9168 (N_9168,N_8687,N_8733);
and U9169 (N_9169,N_8670,N_8078);
nand U9170 (N_9170,N_8010,N_8144);
xor U9171 (N_9171,N_8836,N_8505);
and U9172 (N_9172,N_8421,N_8389);
nor U9173 (N_9173,N_8464,N_8031);
and U9174 (N_9174,N_8814,N_8625);
and U9175 (N_9175,N_8496,N_8663);
and U9176 (N_9176,N_8662,N_8219);
nor U9177 (N_9177,N_8134,N_8405);
nor U9178 (N_9178,N_8615,N_8606);
xnor U9179 (N_9179,N_8483,N_8574);
nor U9180 (N_9180,N_8699,N_8919);
or U9181 (N_9181,N_8917,N_8054);
and U9182 (N_9182,N_8922,N_8256);
nand U9183 (N_9183,N_8837,N_8415);
nor U9184 (N_9184,N_8608,N_8449);
nor U9185 (N_9185,N_8779,N_8349);
or U9186 (N_9186,N_8838,N_8264);
and U9187 (N_9187,N_8724,N_8193);
nor U9188 (N_9188,N_8058,N_8631);
nand U9189 (N_9189,N_8603,N_8927);
and U9190 (N_9190,N_8320,N_8782);
xor U9191 (N_9191,N_8441,N_8492);
xor U9192 (N_9192,N_8440,N_8012);
nand U9193 (N_9193,N_8910,N_8740);
or U9194 (N_9194,N_8470,N_8216);
or U9195 (N_9195,N_8809,N_8207);
xnor U9196 (N_9196,N_8322,N_8667);
nor U9197 (N_9197,N_8890,N_8128);
or U9198 (N_9198,N_8852,N_8555);
nand U9199 (N_9199,N_8168,N_8242);
and U9200 (N_9200,N_8473,N_8787);
or U9201 (N_9201,N_8678,N_8784);
and U9202 (N_9202,N_8334,N_8588);
nor U9203 (N_9203,N_8398,N_8659);
or U9204 (N_9204,N_8681,N_8253);
nor U9205 (N_9205,N_8817,N_8870);
or U9206 (N_9206,N_8118,N_8790);
nand U9207 (N_9207,N_8213,N_8490);
and U9208 (N_9208,N_8825,N_8793);
xor U9209 (N_9209,N_8516,N_8720);
nand U9210 (N_9210,N_8789,N_8113);
and U9211 (N_9211,N_8225,N_8266);
xnor U9212 (N_9212,N_8866,N_8453);
xnor U9213 (N_9213,N_8950,N_8503);
or U9214 (N_9214,N_8218,N_8967);
or U9215 (N_9215,N_8243,N_8998);
nor U9216 (N_9216,N_8666,N_8337);
nor U9217 (N_9217,N_8254,N_8766);
nand U9218 (N_9218,N_8810,N_8169);
nand U9219 (N_9219,N_8597,N_8851);
nand U9220 (N_9220,N_8707,N_8877);
and U9221 (N_9221,N_8981,N_8901);
nand U9222 (N_9222,N_8697,N_8321);
and U9223 (N_9223,N_8174,N_8478);
and U9224 (N_9224,N_8080,N_8893);
xnor U9225 (N_9225,N_8867,N_8952);
nand U9226 (N_9226,N_8761,N_8183);
nor U9227 (N_9227,N_8501,N_8692);
or U9228 (N_9228,N_8105,N_8317);
xor U9229 (N_9229,N_8556,N_8025);
and U9230 (N_9230,N_8913,N_8926);
and U9231 (N_9231,N_8452,N_8827);
or U9232 (N_9232,N_8668,N_8330);
or U9233 (N_9233,N_8143,N_8157);
nand U9234 (N_9234,N_8960,N_8544);
or U9235 (N_9235,N_8395,N_8984);
and U9236 (N_9236,N_8506,N_8305);
nand U9237 (N_9237,N_8569,N_8368);
nor U9238 (N_9238,N_8600,N_8061);
or U9239 (N_9239,N_8630,N_8079);
or U9240 (N_9240,N_8212,N_8274);
nand U9241 (N_9241,N_8686,N_8192);
xnor U9242 (N_9242,N_8634,N_8527);
or U9243 (N_9243,N_8828,N_8804);
nor U9244 (N_9244,N_8891,N_8221);
and U9245 (N_9245,N_8476,N_8982);
nand U9246 (N_9246,N_8194,N_8084);
and U9247 (N_9247,N_8255,N_8127);
or U9248 (N_9248,N_8185,N_8921);
or U9249 (N_9249,N_8736,N_8562);
and U9250 (N_9250,N_8308,N_8397);
xnor U9251 (N_9251,N_8314,N_8959);
nor U9252 (N_9252,N_8549,N_8436);
xor U9253 (N_9253,N_8887,N_8499);
or U9254 (N_9254,N_8107,N_8049);
or U9255 (N_9255,N_8979,N_8956);
and U9256 (N_9256,N_8644,N_8542);
and U9257 (N_9257,N_8968,N_8222);
nand U9258 (N_9258,N_8940,N_8839);
nand U9259 (N_9259,N_8425,N_8131);
or U9260 (N_9260,N_8570,N_8920);
nand U9261 (N_9261,N_8645,N_8403);
or U9262 (N_9262,N_8680,N_8117);
and U9263 (N_9263,N_8382,N_8101);
nand U9264 (N_9264,N_8709,N_8484);
and U9265 (N_9265,N_8136,N_8504);
xnor U9266 (N_9266,N_8407,N_8103);
or U9267 (N_9267,N_8525,N_8847);
and U9268 (N_9268,N_8904,N_8230);
or U9269 (N_9269,N_8433,N_8906);
and U9270 (N_9270,N_8087,N_8769);
or U9271 (N_9271,N_8705,N_8726);
xnor U9272 (N_9272,N_8102,N_8744);
nor U9273 (N_9273,N_8684,N_8497);
nand U9274 (N_9274,N_8281,N_8975);
nor U9275 (N_9275,N_8738,N_8211);
and U9276 (N_9276,N_8586,N_8309);
xnor U9277 (N_9277,N_8227,N_8298);
nor U9278 (N_9278,N_8612,N_8477);
and U9279 (N_9279,N_8480,N_8462);
and U9280 (N_9280,N_8682,N_8696);
and U9281 (N_9281,N_8142,N_8179);
nand U9282 (N_9282,N_8872,N_8596);
nor U9283 (N_9283,N_8426,N_8731);
xnor U9284 (N_9284,N_8533,N_8448);
nand U9285 (N_9285,N_8081,N_8347);
and U9286 (N_9286,N_8199,N_8849);
xnor U9287 (N_9287,N_8669,N_8834);
nand U9288 (N_9288,N_8564,N_8702);
or U9289 (N_9289,N_8348,N_8942);
nand U9290 (N_9290,N_8384,N_8808);
nor U9291 (N_9291,N_8053,N_8665);
xnor U9292 (N_9292,N_8568,N_8607);
or U9293 (N_9293,N_8106,N_8991);
xnor U9294 (N_9294,N_8419,N_8271);
or U9295 (N_9295,N_8158,N_8579);
nor U9296 (N_9296,N_8364,N_8770);
nand U9297 (N_9297,N_8098,N_8188);
nor U9298 (N_9298,N_8114,N_8725);
xnor U9299 (N_9299,N_8951,N_8122);
nand U9300 (N_9300,N_8573,N_8275);
nand U9301 (N_9301,N_8392,N_8273);
xor U9302 (N_9302,N_8708,N_8293);
xnor U9303 (N_9303,N_8786,N_8428);
xor U9304 (N_9304,N_8420,N_8195);
and U9305 (N_9305,N_8575,N_8816);
nor U9306 (N_9306,N_8328,N_8418);
nor U9307 (N_9307,N_8023,N_8014);
xor U9308 (N_9308,N_8949,N_8451);
nand U9309 (N_9309,N_8171,N_8640);
xor U9310 (N_9310,N_8953,N_8165);
nor U9311 (N_9311,N_8388,N_8493);
or U9312 (N_9312,N_8244,N_8899);
nand U9313 (N_9313,N_8434,N_8999);
nor U9314 (N_9314,N_8302,N_8772);
nand U9315 (N_9315,N_8930,N_8517);
nand U9316 (N_9316,N_8166,N_8908);
or U9317 (N_9317,N_8657,N_8911);
nand U9318 (N_9318,N_8150,N_8510);
and U9319 (N_9319,N_8521,N_8854);
nor U9320 (N_9320,N_8627,N_8280);
xor U9321 (N_9321,N_8411,N_8704);
nand U9322 (N_9322,N_8387,N_8250);
or U9323 (N_9323,N_8414,N_8800);
or U9324 (N_9324,N_8030,N_8205);
or U9325 (N_9325,N_8005,N_8794);
nand U9326 (N_9326,N_8673,N_8783);
nor U9327 (N_9327,N_8519,N_8272);
or U9328 (N_9328,N_8781,N_8826);
nor U9329 (N_9329,N_8498,N_8876);
nand U9330 (N_9330,N_8245,N_8016);
and U9331 (N_9331,N_8935,N_8316);
xnor U9332 (N_9332,N_8842,N_8252);
and U9333 (N_9333,N_8755,N_8399);
nand U9334 (N_9334,N_8357,N_8238);
xor U9335 (N_9335,N_8312,N_8036);
and U9336 (N_9336,N_8886,N_8282);
and U9337 (N_9337,N_8500,N_8246);
nand U9338 (N_9338,N_8172,N_8980);
nand U9339 (N_9339,N_8001,N_8535);
and U9340 (N_9340,N_8534,N_8689);
and U9341 (N_9341,N_8331,N_8072);
nor U9342 (N_9342,N_8824,N_8621);
nor U9343 (N_9343,N_8868,N_8024);
or U9344 (N_9344,N_8773,N_8017);
or U9345 (N_9345,N_8883,N_8139);
nor U9346 (N_9346,N_8776,N_8578);
nand U9347 (N_9347,N_8654,N_8381);
and U9348 (N_9348,N_8463,N_8735);
xnor U9349 (N_9349,N_8514,N_8112);
nand U9350 (N_9350,N_8859,N_8747);
nand U9351 (N_9351,N_8884,N_8941);
nor U9352 (N_9352,N_8326,N_8486);
xor U9353 (N_9353,N_8020,N_8823);
or U9354 (N_9354,N_8294,N_8969);
or U9355 (N_9355,N_8132,N_8360);
xnor U9356 (N_9356,N_8714,N_8301);
nand U9357 (N_9357,N_8374,N_8937);
and U9358 (N_9358,N_8661,N_8774);
nand U9359 (N_9359,N_8955,N_8413);
xnor U9360 (N_9360,N_8300,N_8494);
nor U9361 (N_9361,N_8718,N_8443);
or U9362 (N_9362,N_8279,N_8797);
or U9363 (N_9363,N_8401,N_8352);
nor U9364 (N_9364,N_8803,N_8992);
and U9365 (N_9365,N_8613,N_8591);
or U9366 (N_9366,N_8366,N_8507);
nor U9367 (N_9367,N_8186,N_8763);
or U9368 (N_9368,N_8833,N_8522);
xnor U9369 (N_9369,N_8191,N_8947);
and U9370 (N_9370,N_8658,N_8557);
xnor U9371 (N_9371,N_8756,N_8698);
and U9372 (N_9372,N_8045,N_8768);
and U9373 (N_9373,N_8526,N_8875);
nand U9374 (N_9374,N_8160,N_8044);
or U9375 (N_9375,N_8528,N_8664);
nor U9376 (N_9376,N_8223,N_8805);
nor U9377 (N_9377,N_8209,N_8439);
and U9378 (N_9378,N_8604,N_8170);
or U9379 (N_9379,N_8052,N_8618);
or U9380 (N_9380,N_8154,N_8524);
or U9381 (N_9381,N_8099,N_8765);
or U9382 (N_9382,N_8559,N_8026);
or U9383 (N_9383,N_8313,N_8263);
nor U9384 (N_9384,N_8093,N_8111);
xnor U9385 (N_9385,N_8853,N_8465);
nor U9386 (N_9386,N_8653,N_8376);
xnor U9387 (N_9387,N_8307,N_8296);
or U9388 (N_9388,N_8540,N_8385);
nand U9389 (N_9389,N_8889,N_8929);
or U9390 (N_9390,N_8857,N_8679);
or U9391 (N_9391,N_8840,N_8155);
nor U9392 (N_9392,N_8124,N_8717);
nand U9393 (N_9393,N_8934,N_8487);
and U9394 (N_9394,N_8554,N_8324);
or U9395 (N_9395,N_8361,N_8948);
nor U9396 (N_9396,N_8069,N_8359);
xnor U9397 (N_9397,N_8777,N_8728);
nand U9398 (N_9398,N_8206,N_8749);
xor U9399 (N_9399,N_8363,N_8333);
and U9400 (N_9400,N_8153,N_8683);
nor U9401 (N_9401,N_8897,N_8339);
nor U9402 (N_9402,N_8715,N_8215);
nand U9403 (N_9403,N_8795,N_8905);
xor U9404 (N_9404,N_8590,N_8417);
or U9405 (N_9405,N_8383,N_8204);
nand U9406 (N_9406,N_8039,N_8928);
and U9407 (N_9407,N_8895,N_8083);
xor U9408 (N_9408,N_8120,N_8041);
nand U9409 (N_9409,N_8727,N_8064);
xnor U9410 (N_9410,N_8541,N_8006);
or U9411 (N_9411,N_8446,N_8845);
xor U9412 (N_9412,N_8002,N_8882);
and U9413 (N_9413,N_8830,N_8488);
nor U9414 (N_9414,N_8197,N_8019);
xnor U9415 (N_9415,N_8378,N_8427);
nand U9416 (N_9416,N_8650,N_8159);
xnor U9417 (N_9417,N_8987,N_8858);
nor U9418 (N_9418,N_8829,N_8529);
nand U9419 (N_9419,N_8567,N_8623);
or U9420 (N_9420,N_8880,N_8203);
and U9421 (N_9421,N_8444,N_8548);
nand U9422 (N_9422,N_8354,N_8438);
nand U9423 (N_9423,N_8210,N_8032);
and U9424 (N_9424,N_8732,N_8295);
nand U9425 (N_9425,N_8059,N_8073);
and U9426 (N_9426,N_8871,N_8587);
or U9427 (N_9427,N_8672,N_8813);
or U9428 (N_9428,N_8916,N_8751);
xnor U9429 (N_9429,N_8748,N_8416);
or U9430 (N_9430,N_8009,N_8284);
nand U9431 (N_9431,N_8902,N_8821);
or U9432 (N_9432,N_8430,N_8133);
or U9433 (N_9433,N_8130,N_8097);
and U9434 (N_9434,N_8461,N_8390);
nand U9435 (N_9435,N_8057,N_8379);
nand U9436 (N_9436,N_8633,N_8957);
nand U9437 (N_9437,N_8637,N_8268);
and U9438 (N_9438,N_8469,N_8232);
and U9439 (N_9439,N_8050,N_8177);
xor U9440 (N_9440,N_8043,N_8182);
xor U9441 (N_9441,N_8716,N_8841);
or U9442 (N_9442,N_8977,N_8598);
nor U9443 (N_9443,N_8798,N_8104);
and U9444 (N_9444,N_8456,N_8075);
nand U9445 (N_9445,N_8278,N_8116);
nand U9446 (N_9446,N_8338,N_8062);
or U9447 (N_9447,N_8277,N_8346);
or U9448 (N_9448,N_8241,N_8863);
nand U9449 (N_9449,N_8424,N_8467);
xor U9450 (N_9450,N_8178,N_8228);
xnor U9451 (N_9451,N_8750,N_8760);
xnor U9452 (N_9452,N_8022,N_8844);
and U9453 (N_9453,N_8873,N_8445);
and U9454 (N_9454,N_8791,N_8552);
and U9455 (N_9455,N_8958,N_8869);
nor U9456 (N_9456,N_8074,N_8008);
nand U9457 (N_9457,N_8286,N_8971);
and U9458 (N_9458,N_8306,N_8092);
nand U9459 (N_9459,N_8239,N_8693);
or U9460 (N_9460,N_8311,N_8137);
and U9461 (N_9461,N_8088,N_8861);
nor U9462 (N_9462,N_8515,N_8778);
or U9463 (N_9463,N_8119,N_8832);
nor U9464 (N_9464,N_8345,N_8007);
xor U9465 (N_9465,N_8189,N_8450);
nand U9466 (N_9466,N_8015,N_8161);
nor U9467 (N_9467,N_8976,N_8577);
xor U9468 (N_9468,N_8626,N_8076);
or U9469 (N_9469,N_8327,N_8551);
or U9470 (N_9470,N_8035,N_8711);
xor U9471 (N_9471,N_8167,N_8759);
nand U9472 (N_9472,N_8996,N_8202);
and U9473 (N_9473,N_8539,N_8912);
and U9474 (N_9474,N_8396,N_8038);
nor U9475 (N_9475,N_8629,N_8289);
or U9476 (N_9476,N_8799,N_8341);
nor U9477 (N_9477,N_8029,N_8723);
nand U9478 (N_9478,N_8040,N_8589);
nand U9479 (N_9479,N_8719,N_8900);
nand U9480 (N_9480,N_8978,N_8175);
and U9481 (N_9481,N_8970,N_8251);
xnor U9482 (N_9482,N_8276,N_8412);
and U9483 (N_9483,N_8713,N_8148);
xor U9484 (N_9484,N_8335,N_8802);
nand U9485 (N_9485,N_8138,N_8605);
or U9486 (N_9486,N_8892,N_8848);
nand U9487 (N_9487,N_8091,N_8065);
xor U9488 (N_9488,N_8404,N_8226);
nor U9489 (N_9489,N_8468,N_8208);
and U9490 (N_9490,N_8224,N_8592);
or U9491 (N_9491,N_8350,N_8546);
nor U9492 (N_9492,N_8796,N_8758);
and U9493 (N_9493,N_8422,N_8214);
or U9494 (N_9494,N_8000,N_8688);
and U9495 (N_9495,N_8447,N_8095);
and U9496 (N_9496,N_8676,N_8962);
xnor U9497 (N_9497,N_8380,N_8671);
or U9498 (N_9498,N_8377,N_8502);
xor U9499 (N_9499,N_8318,N_8835);
nor U9500 (N_9500,N_8435,N_8843);
xor U9501 (N_9501,N_8826,N_8708);
xor U9502 (N_9502,N_8843,N_8135);
nand U9503 (N_9503,N_8118,N_8094);
nand U9504 (N_9504,N_8138,N_8641);
nand U9505 (N_9505,N_8775,N_8736);
and U9506 (N_9506,N_8684,N_8624);
xor U9507 (N_9507,N_8110,N_8406);
nand U9508 (N_9508,N_8678,N_8188);
or U9509 (N_9509,N_8841,N_8646);
or U9510 (N_9510,N_8800,N_8131);
nand U9511 (N_9511,N_8381,N_8846);
or U9512 (N_9512,N_8963,N_8953);
xnor U9513 (N_9513,N_8985,N_8426);
and U9514 (N_9514,N_8323,N_8145);
xnor U9515 (N_9515,N_8206,N_8149);
or U9516 (N_9516,N_8402,N_8828);
nor U9517 (N_9517,N_8371,N_8319);
nand U9518 (N_9518,N_8912,N_8952);
or U9519 (N_9519,N_8520,N_8775);
or U9520 (N_9520,N_8927,N_8651);
xor U9521 (N_9521,N_8067,N_8579);
or U9522 (N_9522,N_8988,N_8845);
nor U9523 (N_9523,N_8166,N_8701);
and U9524 (N_9524,N_8476,N_8252);
nand U9525 (N_9525,N_8444,N_8261);
and U9526 (N_9526,N_8395,N_8564);
and U9527 (N_9527,N_8102,N_8733);
nor U9528 (N_9528,N_8352,N_8415);
nor U9529 (N_9529,N_8551,N_8333);
or U9530 (N_9530,N_8727,N_8673);
and U9531 (N_9531,N_8972,N_8895);
and U9532 (N_9532,N_8557,N_8588);
or U9533 (N_9533,N_8133,N_8232);
or U9534 (N_9534,N_8388,N_8948);
or U9535 (N_9535,N_8540,N_8055);
or U9536 (N_9536,N_8375,N_8076);
and U9537 (N_9537,N_8432,N_8842);
nand U9538 (N_9538,N_8792,N_8392);
nor U9539 (N_9539,N_8798,N_8431);
xnor U9540 (N_9540,N_8030,N_8973);
xnor U9541 (N_9541,N_8614,N_8381);
nand U9542 (N_9542,N_8418,N_8719);
or U9543 (N_9543,N_8447,N_8479);
xnor U9544 (N_9544,N_8437,N_8458);
xnor U9545 (N_9545,N_8083,N_8116);
and U9546 (N_9546,N_8494,N_8617);
and U9547 (N_9547,N_8705,N_8575);
nor U9548 (N_9548,N_8772,N_8401);
xor U9549 (N_9549,N_8321,N_8766);
nor U9550 (N_9550,N_8896,N_8336);
or U9551 (N_9551,N_8166,N_8772);
nand U9552 (N_9552,N_8574,N_8119);
nand U9553 (N_9553,N_8082,N_8609);
and U9554 (N_9554,N_8123,N_8441);
nand U9555 (N_9555,N_8222,N_8820);
xor U9556 (N_9556,N_8396,N_8656);
nand U9557 (N_9557,N_8615,N_8809);
and U9558 (N_9558,N_8381,N_8865);
nor U9559 (N_9559,N_8741,N_8119);
nor U9560 (N_9560,N_8428,N_8654);
or U9561 (N_9561,N_8364,N_8411);
and U9562 (N_9562,N_8748,N_8292);
nor U9563 (N_9563,N_8654,N_8502);
xor U9564 (N_9564,N_8292,N_8641);
xnor U9565 (N_9565,N_8491,N_8542);
nor U9566 (N_9566,N_8603,N_8013);
and U9567 (N_9567,N_8434,N_8443);
xnor U9568 (N_9568,N_8382,N_8193);
xor U9569 (N_9569,N_8931,N_8409);
xor U9570 (N_9570,N_8218,N_8579);
or U9571 (N_9571,N_8390,N_8268);
xnor U9572 (N_9572,N_8416,N_8443);
nor U9573 (N_9573,N_8984,N_8527);
nand U9574 (N_9574,N_8476,N_8653);
nand U9575 (N_9575,N_8075,N_8952);
nor U9576 (N_9576,N_8988,N_8794);
nor U9577 (N_9577,N_8957,N_8732);
xor U9578 (N_9578,N_8010,N_8280);
nor U9579 (N_9579,N_8911,N_8908);
nor U9580 (N_9580,N_8941,N_8509);
nor U9581 (N_9581,N_8972,N_8399);
or U9582 (N_9582,N_8658,N_8259);
nand U9583 (N_9583,N_8748,N_8013);
nand U9584 (N_9584,N_8297,N_8789);
nor U9585 (N_9585,N_8264,N_8212);
and U9586 (N_9586,N_8834,N_8858);
or U9587 (N_9587,N_8288,N_8001);
and U9588 (N_9588,N_8233,N_8933);
nand U9589 (N_9589,N_8920,N_8045);
nand U9590 (N_9590,N_8301,N_8473);
and U9591 (N_9591,N_8517,N_8059);
or U9592 (N_9592,N_8172,N_8418);
xor U9593 (N_9593,N_8682,N_8813);
and U9594 (N_9594,N_8713,N_8974);
nand U9595 (N_9595,N_8232,N_8513);
or U9596 (N_9596,N_8498,N_8274);
nand U9597 (N_9597,N_8631,N_8704);
and U9598 (N_9598,N_8781,N_8074);
nor U9599 (N_9599,N_8144,N_8613);
xnor U9600 (N_9600,N_8451,N_8054);
nand U9601 (N_9601,N_8514,N_8380);
or U9602 (N_9602,N_8236,N_8917);
nand U9603 (N_9603,N_8546,N_8129);
and U9604 (N_9604,N_8984,N_8575);
nor U9605 (N_9605,N_8905,N_8951);
nand U9606 (N_9606,N_8991,N_8555);
and U9607 (N_9607,N_8870,N_8463);
nor U9608 (N_9608,N_8616,N_8269);
xor U9609 (N_9609,N_8213,N_8296);
and U9610 (N_9610,N_8239,N_8343);
nand U9611 (N_9611,N_8126,N_8651);
or U9612 (N_9612,N_8535,N_8510);
or U9613 (N_9613,N_8993,N_8230);
and U9614 (N_9614,N_8923,N_8030);
nor U9615 (N_9615,N_8025,N_8283);
xor U9616 (N_9616,N_8529,N_8454);
and U9617 (N_9617,N_8660,N_8471);
nand U9618 (N_9618,N_8581,N_8441);
or U9619 (N_9619,N_8466,N_8260);
and U9620 (N_9620,N_8044,N_8668);
and U9621 (N_9621,N_8177,N_8185);
nand U9622 (N_9622,N_8941,N_8176);
or U9623 (N_9623,N_8454,N_8482);
nor U9624 (N_9624,N_8533,N_8949);
nor U9625 (N_9625,N_8975,N_8233);
or U9626 (N_9626,N_8646,N_8980);
and U9627 (N_9627,N_8890,N_8662);
and U9628 (N_9628,N_8141,N_8386);
or U9629 (N_9629,N_8621,N_8160);
or U9630 (N_9630,N_8771,N_8824);
or U9631 (N_9631,N_8521,N_8186);
xor U9632 (N_9632,N_8920,N_8701);
xor U9633 (N_9633,N_8714,N_8663);
xnor U9634 (N_9634,N_8207,N_8887);
and U9635 (N_9635,N_8286,N_8588);
nand U9636 (N_9636,N_8650,N_8651);
or U9637 (N_9637,N_8101,N_8408);
and U9638 (N_9638,N_8974,N_8139);
nor U9639 (N_9639,N_8163,N_8717);
nor U9640 (N_9640,N_8988,N_8762);
xnor U9641 (N_9641,N_8356,N_8248);
or U9642 (N_9642,N_8572,N_8095);
nor U9643 (N_9643,N_8047,N_8170);
and U9644 (N_9644,N_8300,N_8056);
nand U9645 (N_9645,N_8142,N_8201);
nand U9646 (N_9646,N_8209,N_8279);
and U9647 (N_9647,N_8243,N_8958);
and U9648 (N_9648,N_8809,N_8790);
or U9649 (N_9649,N_8139,N_8575);
xor U9650 (N_9650,N_8209,N_8740);
and U9651 (N_9651,N_8755,N_8356);
nand U9652 (N_9652,N_8071,N_8322);
or U9653 (N_9653,N_8888,N_8871);
and U9654 (N_9654,N_8106,N_8658);
and U9655 (N_9655,N_8883,N_8159);
nor U9656 (N_9656,N_8438,N_8623);
nand U9657 (N_9657,N_8872,N_8861);
nor U9658 (N_9658,N_8868,N_8598);
nor U9659 (N_9659,N_8147,N_8166);
nor U9660 (N_9660,N_8091,N_8329);
nor U9661 (N_9661,N_8260,N_8404);
or U9662 (N_9662,N_8254,N_8181);
nor U9663 (N_9663,N_8282,N_8099);
nor U9664 (N_9664,N_8842,N_8117);
and U9665 (N_9665,N_8929,N_8986);
xor U9666 (N_9666,N_8855,N_8212);
and U9667 (N_9667,N_8224,N_8949);
xor U9668 (N_9668,N_8712,N_8748);
or U9669 (N_9669,N_8257,N_8958);
and U9670 (N_9670,N_8825,N_8335);
xor U9671 (N_9671,N_8163,N_8273);
nand U9672 (N_9672,N_8818,N_8943);
and U9673 (N_9673,N_8980,N_8693);
nand U9674 (N_9674,N_8645,N_8412);
nand U9675 (N_9675,N_8316,N_8267);
nor U9676 (N_9676,N_8268,N_8479);
and U9677 (N_9677,N_8618,N_8026);
xnor U9678 (N_9678,N_8327,N_8337);
and U9679 (N_9679,N_8383,N_8927);
xnor U9680 (N_9680,N_8459,N_8329);
nor U9681 (N_9681,N_8526,N_8356);
and U9682 (N_9682,N_8359,N_8177);
or U9683 (N_9683,N_8023,N_8525);
nand U9684 (N_9684,N_8488,N_8903);
nor U9685 (N_9685,N_8967,N_8002);
and U9686 (N_9686,N_8255,N_8215);
nand U9687 (N_9687,N_8323,N_8120);
or U9688 (N_9688,N_8280,N_8611);
xor U9689 (N_9689,N_8199,N_8380);
or U9690 (N_9690,N_8870,N_8763);
and U9691 (N_9691,N_8393,N_8043);
nor U9692 (N_9692,N_8021,N_8243);
and U9693 (N_9693,N_8413,N_8672);
nand U9694 (N_9694,N_8813,N_8636);
and U9695 (N_9695,N_8343,N_8895);
nand U9696 (N_9696,N_8156,N_8268);
xor U9697 (N_9697,N_8022,N_8282);
or U9698 (N_9698,N_8581,N_8096);
xnor U9699 (N_9699,N_8136,N_8509);
or U9700 (N_9700,N_8852,N_8580);
or U9701 (N_9701,N_8307,N_8253);
nand U9702 (N_9702,N_8304,N_8382);
nor U9703 (N_9703,N_8147,N_8003);
xor U9704 (N_9704,N_8678,N_8479);
nand U9705 (N_9705,N_8764,N_8514);
and U9706 (N_9706,N_8400,N_8135);
and U9707 (N_9707,N_8376,N_8749);
and U9708 (N_9708,N_8709,N_8864);
or U9709 (N_9709,N_8796,N_8908);
nand U9710 (N_9710,N_8260,N_8081);
or U9711 (N_9711,N_8048,N_8650);
nor U9712 (N_9712,N_8450,N_8826);
xor U9713 (N_9713,N_8083,N_8194);
nand U9714 (N_9714,N_8743,N_8873);
xnor U9715 (N_9715,N_8548,N_8541);
xnor U9716 (N_9716,N_8590,N_8431);
xnor U9717 (N_9717,N_8440,N_8656);
nor U9718 (N_9718,N_8153,N_8986);
and U9719 (N_9719,N_8609,N_8971);
and U9720 (N_9720,N_8727,N_8509);
nor U9721 (N_9721,N_8244,N_8401);
xor U9722 (N_9722,N_8611,N_8261);
xor U9723 (N_9723,N_8193,N_8218);
nor U9724 (N_9724,N_8484,N_8168);
xnor U9725 (N_9725,N_8558,N_8273);
or U9726 (N_9726,N_8996,N_8892);
xnor U9727 (N_9727,N_8412,N_8246);
and U9728 (N_9728,N_8197,N_8205);
nor U9729 (N_9729,N_8486,N_8851);
nand U9730 (N_9730,N_8448,N_8597);
xor U9731 (N_9731,N_8483,N_8803);
or U9732 (N_9732,N_8754,N_8345);
nor U9733 (N_9733,N_8993,N_8579);
xor U9734 (N_9734,N_8325,N_8226);
nor U9735 (N_9735,N_8659,N_8055);
xnor U9736 (N_9736,N_8729,N_8736);
nor U9737 (N_9737,N_8369,N_8048);
nor U9738 (N_9738,N_8346,N_8474);
xnor U9739 (N_9739,N_8838,N_8030);
nand U9740 (N_9740,N_8779,N_8213);
xnor U9741 (N_9741,N_8963,N_8654);
nand U9742 (N_9742,N_8661,N_8509);
nor U9743 (N_9743,N_8270,N_8505);
nand U9744 (N_9744,N_8897,N_8079);
nand U9745 (N_9745,N_8923,N_8278);
xor U9746 (N_9746,N_8904,N_8475);
nand U9747 (N_9747,N_8771,N_8474);
or U9748 (N_9748,N_8038,N_8782);
nand U9749 (N_9749,N_8600,N_8324);
or U9750 (N_9750,N_8591,N_8024);
or U9751 (N_9751,N_8073,N_8524);
and U9752 (N_9752,N_8959,N_8847);
or U9753 (N_9753,N_8374,N_8807);
xnor U9754 (N_9754,N_8783,N_8353);
nor U9755 (N_9755,N_8997,N_8880);
nor U9756 (N_9756,N_8497,N_8460);
and U9757 (N_9757,N_8148,N_8982);
or U9758 (N_9758,N_8906,N_8443);
nand U9759 (N_9759,N_8239,N_8649);
nor U9760 (N_9760,N_8957,N_8300);
or U9761 (N_9761,N_8460,N_8580);
nand U9762 (N_9762,N_8261,N_8377);
and U9763 (N_9763,N_8241,N_8227);
and U9764 (N_9764,N_8515,N_8024);
and U9765 (N_9765,N_8330,N_8447);
or U9766 (N_9766,N_8006,N_8055);
or U9767 (N_9767,N_8418,N_8377);
nor U9768 (N_9768,N_8186,N_8452);
nor U9769 (N_9769,N_8611,N_8073);
nand U9770 (N_9770,N_8046,N_8283);
xor U9771 (N_9771,N_8844,N_8093);
xnor U9772 (N_9772,N_8616,N_8709);
nand U9773 (N_9773,N_8396,N_8584);
and U9774 (N_9774,N_8810,N_8301);
or U9775 (N_9775,N_8919,N_8856);
xnor U9776 (N_9776,N_8588,N_8198);
nor U9777 (N_9777,N_8282,N_8911);
nor U9778 (N_9778,N_8022,N_8784);
or U9779 (N_9779,N_8224,N_8058);
or U9780 (N_9780,N_8136,N_8303);
or U9781 (N_9781,N_8533,N_8391);
nor U9782 (N_9782,N_8094,N_8219);
and U9783 (N_9783,N_8647,N_8140);
or U9784 (N_9784,N_8776,N_8823);
and U9785 (N_9785,N_8564,N_8009);
nor U9786 (N_9786,N_8333,N_8538);
or U9787 (N_9787,N_8361,N_8016);
nor U9788 (N_9788,N_8710,N_8429);
nor U9789 (N_9789,N_8216,N_8160);
nor U9790 (N_9790,N_8433,N_8353);
and U9791 (N_9791,N_8769,N_8978);
xnor U9792 (N_9792,N_8616,N_8546);
nand U9793 (N_9793,N_8295,N_8408);
xor U9794 (N_9794,N_8919,N_8692);
nor U9795 (N_9795,N_8058,N_8968);
nand U9796 (N_9796,N_8796,N_8381);
nor U9797 (N_9797,N_8404,N_8281);
nand U9798 (N_9798,N_8504,N_8800);
xnor U9799 (N_9799,N_8785,N_8675);
and U9800 (N_9800,N_8307,N_8676);
or U9801 (N_9801,N_8457,N_8503);
xor U9802 (N_9802,N_8240,N_8062);
nor U9803 (N_9803,N_8434,N_8480);
nor U9804 (N_9804,N_8405,N_8308);
and U9805 (N_9805,N_8826,N_8640);
and U9806 (N_9806,N_8483,N_8179);
or U9807 (N_9807,N_8597,N_8864);
xnor U9808 (N_9808,N_8911,N_8225);
xor U9809 (N_9809,N_8686,N_8401);
or U9810 (N_9810,N_8788,N_8434);
and U9811 (N_9811,N_8486,N_8639);
nand U9812 (N_9812,N_8111,N_8937);
nand U9813 (N_9813,N_8494,N_8629);
and U9814 (N_9814,N_8479,N_8590);
or U9815 (N_9815,N_8001,N_8689);
xor U9816 (N_9816,N_8350,N_8501);
nand U9817 (N_9817,N_8752,N_8603);
or U9818 (N_9818,N_8762,N_8741);
and U9819 (N_9819,N_8979,N_8269);
nor U9820 (N_9820,N_8836,N_8952);
nor U9821 (N_9821,N_8957,N_8842);
or U9822 (N_9822,N_8258,N_8103);
nand U9823 (N_9823,N_8362,N_8757);
xnor U9824 (N_9824,N_8101,N_8437);
or U9825 (N_9825,N_8038,N_8355);
and U9826 (N_9826,N_8621,N_8531);
xnor U9827 (N_9827,N_8725,N_8200);
or U9828 (N_9828,N_8350,N_8379);
nor U9829 (N_9829,N_8741,N_8093);
xor U9830 (N_9830,N_8260,N_8780);
xnor U9831 (N_9831,N_8053,N_8692);
nand U9832 (N_9832,N_8760,N_8471);
nand U9833 (N_9833,N_8589,N_8183);
or U9834 (N_9834,N_8807,N_8227);
nor U9835 (N_9835,N_8757,N_8950);
nand U9836 (N_9836,N_8863,N_8685);
or U9837 (N_9837,N_8492,N_8522);
and U9838 (N_9838,N_8511,N_8952);
or U9839 (N_9839,N_8760,N_8266);
xnor U9840 (N_9840,N_8601,N_8339);
or U9841 (N_9841,N_8313,N_8923);
or U9842 (N_9842,N_8512,N_8651);
xnor U9843 (N_9843,N_8089,N_8682);
or U9844 (N_9844,N_8674,N_8659);
nor U9845 (N_9845,N_8172,N_8699);
nor U9846 (N_9846,N_8034,N_8288);
and U9847 (N_9847,N_8468,N_8256);
nand U9848 (N_9848,N_8114,N_8238);
or U9849 (N_9849,N_8323,N_8621);
or U9850 (N_9850,N_8645,N_8366);
or U9851 (N_9851,N_8115,N_8187);
nor U9852 (N_9852,N_8701,N_8145);
or U9853 (N_9853,N_8918,N_8108);
and U9854 (N_9854,N_8231,N_8340);
nor U9855 (N_9855,N_8701,N_8536);
or U9856 (N_9856,N_8604,N_8369);
or U9857 (N_9857,N_8976,N_8736);
xnor U9858 (N_9858,N_8564,N_8467);
and U9859 (N_9859,N_8309,N_8658);
nand U9860 (N_9860,N_8739,N_8393);
and U9861 (N_9861,N_8578,N_8355);
or U9862 (N_9862,N_8951,N_8030);
nand U9863 (N_9863,N_8084,N_8639);
nor U9864 (N_9864,N_8534,N_8884);
nor U9865 (N_9865,N_8512,N_8932);
and U9866 (N_9866,N_8856,N_8129);
nor U9867 (N_9867,N_8209,N_8095);
nand U9868 (N_9868,N_8223,N_8561);
xnor U9869 (N_9869,N_8578,N_8158);
nor U9870 (N_9870,N_8598,N_8771);
nand U9871 (N_9871,N_8340,N_8511);
nand U9872 (N_9872,N_8005,N_8703);
nor U9873 (N_9873,N_8662,N_8350);
or U9874 (N_9874,N_8876,N_8379);
nand U9875 (N_9875,N_8725,N_8426);
and U9876 (N_9876,N_8838,N_8131);
nor U9877 (N_9877,N_8862,N_8582);
nor U9878 (N_9878,N_8646,N_8187);
or U9879 (N_9879,N_8418,N_8133);
nand U9880 (N_9880,N_8865,N_8283);
nor U9881 (N_9881,N_8604,N_8165);
nor U9882 (N_9882,N_8247,N_8980);
or U9883 (N_9883,N_8387,N_8996);
or U9884 (N_9884,N_8455,N_8985);
nand U9885 (N_9885,N_8795,N_8613);
or U9886 (N_9886,N_8621,N_8328);
and U9887 (N_9887,N_8922,N_8839);
and U9888 (N_9888,N_8638,N_8253);
nand U9889 (N_9889,N_8268,N_8975);
nor U9890 (N_9890,N_8034,N_8594);
nand U9891 (N_9891,N_8417,N_8146);
and U9892 (N_9892,N_8366,N_8260);
nand U9893 (N_9893,N_8172,N_8604);
xor U9894 (N_9894,N_8495,N_8692);
or U9895 (N_9895,N_8940,N_8256);
and U9896 (N_9896,N_8002,N_8720);
or U9897 (N_9897,N_8132,N_8700);
nand U9898 (N_9898,N_8090,N_8905);
nor U9899 (N_9899,N_8495,N_8367);
xor U9900 (N_9900,N_8398,N_8962);
or U9901 (N_9901,N_8713,N_8336);
and U9902 (N_9902,N_8599,N_8696);
nor U9903 (N_9903,N_8257,N_8575);
nand U9904 (N_9904,N_8788,N_8523);
and U9905 (N_9905,N_8415,N_8116);
nor U9906 (N_9906,N_8853,N_8511);
or U9907 (N_9907,N_8417,N_8686);
nand U9908 (N_9908,N_8347,N_8380);
nor U9909 (N_9909,N_8514,N_8555);
nand U9910 (N_9910,N_8690,N_8037);
xor U9911 (N_9911,N_8148,N_8651);
and U9912 (N_9912,N_8661,N_8457);
xnor U9913 (N_9913,N_8758,N_8169);
and U9914 (N_9914,N_8415,N_8335);
and U9915 (N_9915,N_8671,N_8261);
xor U9916 (N_9916,N_8652,N_8505);
xor U9917 (N_9917,N_8822,N_8763);
and U9918 (N_9918,N_8747,N_8093);
nand U9919 (N_9919,N_8948,N_8288);
nor U9920 (N_9920,N_8072,N_8816);
xor U9921 (N_9921,N_8723,N_8903);
or U9922 (N_9922,N_8852,N_8022);
and U9923 (N_9923,N_8695,N_8518);
nor U9924 (N_9924,N_8368,N_8907);
or U9925 (N_9925,N_8278,N_8105);
xor U9926 (N_9926,N_8376,N_8605);
xor U9927 (N_9927,N_8788,N_8511);
nand U9928 (N_9928,N_8198,N_8988);
nand U9929 (N_9929,N_8230,N_8253);
xnor U9930 (N_9930,N_8943,N_8246);
or U9931 (N_9931,N_8539,N_8527);
or U9932 (N_9932,N_8637,N_8779);
and U9933 (N_9933,N_8271,N_8547);
nand U9934 (N_9934,N_8074,N_8272);
nor U9935 (N_9935,N_8876,N_8740);
or U9936 (N_9936,N_8409,N_8139);
nor U9937 (N_9937,N_8266,N_8766);
or U9938 (N_9938,N_8602,N_8684);
and U9939 (N_9939,N_8369,N_8816);
nor U9940 (N_9940,N_8240,N_8780);
and U9941 (N_9941,N_8503,N_8720);
or U9942 (N_9942,N_8284,N_8781);
xor U9943 (N_9943,N_8045,N_8059);
or U9944 (N_9944,N_8745,N_8164);
nor U9945 (N_9945,N_8144,N_8320);
or U9946 (N_9946,N_8474,N_8511);
xnor U9947 (N_9947,N_8103,N_8625);
or U9948 (N_9948,N_8510,N_8652);
or U9949 (N_9949,N_8170,N_8394);
xnor U9950 (N_9950,N_8096,N_8510);
nor U9951 (N_9951,N_8630,N_8304);
xnor U9952 (N_9952,N_8736,N_8200);
or U9953 (N_9953,N_8189,N_8710);
xnor U9954 (N_9954,N_8515,N_8674);
nor U9955 (N_9955,N_8615,N_8588);
or U9956 (N_9956,N_8291,N_8972);
nand U9957 (N_9957,N_8405,N_8149);
nor U9958 (N_9958,N_8737,N_8118);
or U9959 (N_9959,N_8638,N_8194);
nor U9960 (N_9960,N_8714,N_8564);
or U9961 (N_9961,N_8832,N_8989);
nor U9962 (N_9962,N_8096,N_8641);
nand U9963 (N_9963,N_8457,N_8944);
or U9964 (N_9964,N_8525,N_8559);
nand U9965 (N_9965,N_8247,N_8487);
xor U9966 (N_9966,N_8854,N_8971);
nor U9967 (N_9967,N_8118,N_8107);
and U9968 (N_9968,N_8885,N_8477);
or U9969 (N_9969,N_8058,N_8434);
xnor U9970 (N_9970,N_8536,N_8073);
or U9971 (N_9971,N_8951,N_8986);
nand U9972 (N_9972,N_8120,N_8751);
and U9973 (N_9973,N_8185,N_8927);
and U9974 (N_9974,N_8281,N_8649);
nor U9975 (N_9975,N_8736,N_8766);
and U9976 (N_9976,N_8278,N_8864);
nor U9977 (N_9977,N_8854,N_8795);
or U9978 (N_9978,N_8137,N_8553);
nor U9979 (N_9979,N_8516,N_8840);
xor U9980 (N_9980,N_8191,N_8483);
or U9981 (N_9981,N_8443,N_8939);
nor U9982 (N_9982,N_8046,N_8275);
and U9983 (N_9983,N_8199,N_8585);
xor U9984 (N_9984,N_8981,N_8951);
nand U9985 (N_9985,N_8285,N_8137);
or U9986 (N_9986,N_8521,N_8082);
xnor U9987 (N_9987,N_8465,N_8154);
nand U9988 (N_9988,N_8286,N_8124);
nor U9989 (N_9989,N_8764,N_8507);
xnor U9990 (N_9990,N_8175,N_8511);
or U9991 (N_9991,N_8315,N_8895);
nand U9992 (N_9992,N_8478,N_8084);
and U9993 (N_9993,N_8407,N_8634);
nor U9994 (N_9994,N_8329,N_8549);
nand U9995 (N_9995,N_8902,N_8113);
or U9996 (N_9996,N_8951,N_8878);
and U9997 (N_9997,N_8130,N_8385);
nor U9998 (N_9998,N_8993,N_8735);
xor U9999 (N_9999,N_8794,N_8609);
xor U10000 (N_10000,N_9556,N_9466);
nand U10001 (N_10001,N_9634,N_9054);
nand U10002 (N_10002,N_9108,N_9195);
and U10003 (N_10003,N_9388,N_9975);
or U10004 (N_10004,N_9193,N_9589);
xor U10005 (N_10005,N_9212,N_9864);
and U10006 (N_10006,N_9962,N_9192);
xnor U10007 (N_10007,N_9246,N_9714);
nand U10008 (N_10008,N_9446,N_9127);
and U10009 (N_10009,N_9857,N_9028);
nor U10010 (N_10010,N_9264,N_9522);
nor U10011 (N_10011,N_9344,N_9262);
nand U10012 (N_10012,N_9009,N_9837);
nor U10013 (N_10013,N_9079,N_9667);
xnor U10014 (N_10014,N_9835,N_9162);
or U10015 (N_10015,N_9644,N_9257);
xor U10016 (N_10016,N_9378,N_9188);
xor U10017 (N_10017,N_9713,N_9819);
nor U10018 (N_10018,N_9218,N_9040);
xor U10019 (N_10019,N_9343,N_9968);
xnor U10020 (N_10020,N_9944,N_9880);
xor U10021 (N_10021,N_9992,N_9896);
or U10022 (N_10022,N_9694,N_9438);
and U10023 (N_10023,N_9507,N_9242);
and U10024 (N_10024,N_9220,N_9812);
nand U10025 (N_10025,N_9179,N_9704);
xor U10026 (N_10026,N_9329,N_9073);
xnor U10027 (N_10027,N_9672,N_9889);
or U10028 (N_10028,N_9940,N_9543);
nor U10029 (N_10029,N_9524,N_9987);
nor U10030 (N_10030,N_9364,N_9996);
xnor U10031 (N_10031,N_9965,N_9464);
xnor U10032 (N_10032,N_9610,N_9159);
xor U10033 (N_10033,N_9395,N_9414);
or U10034 (N_10034,N_9764,N_9389);
nand U10035 (N_10035,N_9984,N_9846);
and U10036 (N_10036,N_9983,N_9031);
nor U10037 (N_10037,N_9848,N_9902);
nor U10038 (N_10038,N_9790,N_9354);
xnor U10039 (N_10039,N_9788,N_9319);
nand U10040 (N_10040,N_9937,N_9461);
and U10041 (N_10041,N_9082,N_9025);
xnor U10042 (N_10042,N_9753,N_9649);
or U10043 (N_10043,N_9015,N_9850);
nor U10044 (N_10044,N_9055,N_9153);
xnor U10045 (N_10045,N_9725,N_9097);
and U10046 (N_10046,N_9290,N_9800);
or U10047 (N_10047,N_9733,N_9500);
and U10048 (N_10048,N_9805,N_9286);
nor U10049 (N_10049,N_9318,N_9576);
xor U10050 (N_10050,N_9105,N_9701);
and U10051 (N_10051,N_9460,N_9029);
or U10052 (N_10052,N_9299,N_9163);
xnor U10053 (N_10053,N_9831,N_9808);
nor U10054 (N_10054,N_9287,N_9165);
xnor U10055 (N_10055,N_9315,N_9597);
or U10056 (N_10056,N_9929,N_9310);
nor U10057 (N_10057,N_9912,N_9143);
xor U10058 (N_10058,N_9907,N_9309);
nor U10059 (N_10059,N_9488,N_9345);
and U10060 (N_10060,N_9666,N_9881);
nand U10061 (N_10061,N_9393,N_9527);
nor U10062 (N_10062,N_9718,N_9587);
nor U10063 (N_10063,N_9427,N_9605);
and U10064 (N_10064,N_9476,N_9600);
nand U10065 (N_10065,N_9441,N_9958);
or U10066 (N_10066,N_9209,N_9136);
nor U10067 (N_10067,N_9719,N_9140);
nand U10068 (N_10068,N_9633,N_9431);
nor U10069 (N_10069,N_9532,N_9386);
and U10070 (N_10070,N_9854,N_9664);
nor U10071 (N_10071,N_9780,N_9093);
and U10072 (N_10072,N_9871,N_9707);
nor U10073 (N_10073,N_9449,N_9551);
and U10074 (N_10074,N_9206,N_9530);
nor U10075 (N_10075,N_9722,N_9201);
xnor U10076 (N_10076,N_9828,N_9401);
xor U10077 (N_10077,N_9906,N_9976);
and U10078 (N_10078,N_9882,N_9170);
nor U10079 (N_10079,N_9064,N_9927);
nor U10080 (N_10080,N_9297,N_9643);
and U10081 (N_10081,N_9595,N_9408);
and U10082 (N_10082,N_9898,N_9771);
nand U10083 (N_10083,N_9624,N_9190);
and U10084 (N_10084,N_9801,N_9101);
xnor U10085 (N_10085,N_9394,N_9844);
or U10086 (N_10086,N_9475,N_9370);
or U10087 (N_10087,N_9196,N_9562);
nand U10088 (N_10088,N_9325,N_9341);
nor U10089 (N_10089,N_9544,N_9096);
nand U10090 (N_10090,N_9100,N_9281);
nor U10091 (N_10091,N_9497,N_9276);
and U10092 (N_10092,N_9300,N_9593);
nand U10093 (N_10093,N_9582,N_9558);
and U10094 (N_10094,N_9240,N_9385);
nor U10095 (N_10095,N_9570,N_9765);
nor U10096 (N_10096,N_9231,N_9747);
nand U10097 (N_10097,N_9072,N_9186);
nor U10098 (N_10098,N_9030,N_9526);
and U10099 (N_10099,N_9821,N_9550);
xor U10100 (N_10100,N_9826,N_9443);
nor U10101 (N_10101,N_9646,N_9489);
or U10102 (N_10102,N_9749,N_9629);
nor U10103 (N_10103,N_9618,N_9450);
and U10104 (N_10104,N_9061,N_9591);
xnor U10105 (N_10105,N_9226,N_9947);
nand U10106 (N_10106,N_9499,N_9151);
xnor U10107 (N_10107,N_9679,N_9545);
or U10108 (N_10108,N_9392,N_9365);
xnor U10109 (N_10109,N_9870,N_9567);
and U10110 (N_10110,N_9412,N_9843);
or U10111 (N_10111,N_9795,N_9862);
or U10112 (N_10112,N_9433,N_9743);
and U10113 (N_10113,N_9353,N_9791);
and U10114 (N_10114,N_9059,N_9440);
or U10115 (N_10115,N_9809,N_9782);
nor U10116 (N_10116,N_9807,N_9459);
and U10117 (N_10117,N_9684,N_9396);
or U10118 (N_10118,N_9210,N_9676);
nand U10119 (N_10119,N_9243,N_9458);
or U10120 (N_10120,N_9954,N_9038);
and U10121 (N_10121,N_9734,N_9516);
nor U10122 (N_10122,N_9278,N_9062);
nand U10123 (N_10123,N_9087,N_9052);
xnor U10124 (N_10124,N_9478,N_9171);
xor U10125 (N_10125,N_9227,N_9696);
nor U10126 (N_10126,N_9675,N_9298);
or U10127 (N_10127,N_9538,N_9372);
nand U10128 (N_10128,N_9083,N_9494);
nor U10129 (N_10129,N_9419,N_9729);
nor U10130 (N_10130,N_9953,N_9663);
nor U10131 (N_10131,N_9619,N_9482);
nor U10132 (N_10132,N_9448,N_9283);
or U10133 (N_10133,N_9363,N_9942);
nand U10134 (N_10134,N_9799,N_9737);
xnor U10135 (N_10135,N_9022,N_9811);
nand U10136 (N_10136,N_9293,N_9168);
and U10137 (N_10137,N_9893,N_9573);
and U10138 (N_10138,N_9360,N_9352);
xor U10139 (N_10139,N_9503,N_9081);
or U10140 (N_10140,N_9410,N_9739);
xnor U10141 (N_10141,N_9615,N_9540);
nor U10142 (N_10142,N_9307,N_9561);
and U10143 (N_10143,N_9012,N_9228);
nand U10144 (N_10144,N_9934,N_9537);
nand U10145 (N_10145,N_9091,N_9825);
or U10146 (N_10146,N_9838,N_9515);
and U10147 (N_10147,N_9781,N_9866);
nor U10148 (N_10148,N_9334,N_9185);
and U10149 (N_10149,N_9579,N_9580);
nor U10150 (N_10150,N_9049,N_9160);
and U10151 (N_10151,N_9452,N_9816);
and U10152 (N_10152,N_9581,N_9622);
xor U10153 (N_10153,N_9598,N_9122);
and U10154 (N_10154,N_9710,N_9036);
nor U10155 (N_10155,N_9088,N_9931);
nand U10156 (N_10156,N_9783,N_9203);
nor U10157 (N_10157,N_9956,N_9229);
or U10158 (N_10158,N_9111,N_9943);
or U10159 (N_10159,N_9736,N_9416);
and U10160 (N_10160,N_9470,N_9858);
xnor U10161 (N_10161,N_9523,N_9282);
nand U10162 (N_10162,N_9400,N_9071);
nand U10163 (N_10163,N_9237,N_9387);
nand U10164 (N_10164,N_9014,N_9042);
nor U10165 (N_10165,N_9640,N_9349);
xor U10166 (N_10166,N_9067,N_9258);
and U10167 (N_10167,N_9355,N_9121);
and U10168 (N_10168,N_9642,N_9603);
or U10169 (N_10169,N_9911,N_9280);
or U10170 (N_10170,N_9358,N_9511);
and U10171 (N_10171,N_9484,N_9144);
nand U10172 (N_10172,N_9407,N_9759);
nor U10173 (N_10173,N_9379,N_9892);
or U10174 (N_10174,N_9000,N_9625);
nor U10175 (N_10175,N_9614,N_9963);
nor U10176 (N_10176,N_9789,N_9648);
nor U10177 (N_10177,N_9322,N_9720);
or U10178 (N_10178,N_9207,N_9141);
nand U10179 (N_10179,N_9630,N_9018);
nand U10180 (N_10180,N_9045,N_9430);
xor U10181 (N_10181,N_9357,N_9462);
nand U10182 (N_10182,N_9342,N_9376);
or U10183 (N_10183,N_9685,N_9232);
and U10184 (N_10184,N_9048,N_9180);
xnor U10185 (N_10185,N_9620,N_9444);
nor U10186 (N_10186,N_9840,N_9474);
nand U10187 (N_10187,N_9382,N_9546);
nand U10188 (N_10188,N_9421,N_9697);
or U10189 (N_10189,N_9104,N_9842);
nor U10190 (N_10190,N_9745,N_9506);
nor U10191 (N_10191,N_9981,N_9536);
xor U10192 (N_10192,N_9690,N_9333);
nor U10193 (N_10193,N_9090,N_9779);
nor U10194 (N_10194,N_9999,N_9266);
and U10195 (N_10195,N_9026,N_9167);
and U10196 (N_10196,N_9909,N_9250);
nor U10197 (N_10197,N_9245,N_9123);
and U10198 (N_10198,N_9361,N_9712);
nand U10199 (N_10199,N_9873,N_9439);
or U10200 (N_10200,N_9883,N_9027);
nand U10201 (N_10201,N_9935,N_9017);
or U10202 (N_10202,N_9058,N_9606);
nor U10203 (N_10203,N_9994,N_9967);
and U10204 (N_10204,N_9888,N_9933);
nand U10205 (N_10205,N_9938,N_9867);
nor U10206 (N_10206,N_9949,N_9677);
xor U10207 (N_10207,N_9383,N_9485);
and U10208 (N_10208,N_9187,N_9554);
nand U10209 (N_10209,N_9741,N_9164);
nor U10210 (N_10210,N_9671,N_9773);
nand U10211 (N_10211,N_9886,N_9692);
and U10212 (N_10212,N_9374,N_9786);
or U10213 (N_10213,N_9897,N_9616);
nand U10214 (N_10214,N_9859,N_9295);
nand U10215 (N_10215,N_9323,N_9599);
nor U10216 (N_10216,N_9590,N_9356);
xor U10217 (N_10217,N_9752,N_9763);
nor U10218 (N_10218,N_9723,N_9256);
xnor U10219 (N_10219,N_9596,N_9535);
nand U10220 (N_10220,N_9832,N_9197);
nor U10221 (N_10221,N_9830,N_9199);
or U10222 (N_10222,N_9236,N_9921);
nand U10223 (N_10223,N_9324,N_9126);
and U10224 (N_10224,N_9621,N_9359);
nor U10225 (N_10225,N_9043,N_9463);
and U10226 (N_10226,N_9705,N_9335);
xnor U10227 (N_10227,N_9133,N_9566);
or U10228 (N_10228,N_9631,N_9469);
nand U10229 (N_10229,N_9751,N_9332);
and U10230 (N_10230,N_9390,N_9007);
xnor U10231 (N_10231,N_9493,N_9467);
xor U10232 (N_10232,N_9158,N_9820);
nor U10233 (N_10233,N_9592,N_9402);
and U10234 (N_10234,N_9447,N_9660);
nand U10235 (N_10235,N_9673,N_9434);
xnor U10236 (N_10236,N_9518,N_9553);
or U10237 (N_10237,N_9952,N_9371);
xnor U10238 (N_10238,N_9727,N_9977);
or U10239 (N_10239,N_9481,N_9972);
xnor U10240 (N_10240,N_9552,N_9650);
or U10241 (N_10241,N_9145,N_9607);
nor U10242 (N_10242,N_9869,N_9735);
nor U10243 (N_10243,N_9066,N_9253);
nor U10244 (N_10244,N_9311,N_9020);
nand U10245 (N_10245,N_9767,N_9699);
or U10246 (N_10246,N_9827,N_9979);
or U10247 (N_10247,N_9422,N_9874);
nand U10248 (N_10248,N_9529,N_9966);
or U10249 (N_10249,N_9080,N_9157);
or U10250 (N_10250,N_9525,N_9877);
xnor U10251 (N_10251,N_9794,N_9454);
nor U10252 (N_10252,N_9602,N_9978);
xnor U10253 (N_10253,N_9260,N_9757);
xnor U10254 (N_10254,N_9362,N_9817);
and U10255 (N_10255,N_9572,N_9774);
and U10256 (N_10256,N_9146,N_9652);
xnor U10257 (N_10257,N_9768,N_9099);
or U10258 (N_10258,N_9259,N_9513);
nor U10259 (N_10259,N_9995,N_9116);
or U10260 (N_10260,N_9230,N_9708);
and U10261 (N_10261,N_9742,N_9312);
nor U10262 (N_10262,N_9011,N_9239);
nand U10263 (N_10263,N_9796,N_9219);
and U10264 (N_10264,N_9785,N_9611);
and U10265 (N_10265,N_9797,N_9155);
or U10266 (N_10266,N_9033,N_9273);
nor U10267 (N_10267,N_9549,N_9728);
xor U10268 (N_10268,N_9716,N_9651);
or U10269 (N_10269,N_9003,N_9726);
or U10270 (N_10270,N_9135,N_9936);
xor U10271 (N_10271,N_9627,N_9559);
or U10272 (N_10272,N_9533,N_9267);
nor U10273 (N_10273,N_9094,N_9924);
nor U10274 (N_10274,N_9623,N_9275);
nand U10275 (N_10275,N_9455,N_9682);
xor U10276 (N_10276,N_9442,N_9637);
or U10277 (N_10277,N_9409,N_9154);
xnor U10278 (N_10278,N_9302,N_9903);
and U10279 (N_10279,N_9202,N_9957);
or U10280 (N_10280,N_9010,N_9420);
and U10281 (N_10281,N_9683,N_9863);
nand U10282 (N_10282,N_9075,N_9375);
nor U10283 (N_10283,N_9974,N_9802);
or U10284 (N_10284,N_9514,N_9717);
nand U10285 (N_10285,N_9923,N_9670);
and U10286 (N_10286,N_9119,N_9404);
or U10287 (N_10287,N_9223,N_9249);
or U10288 (N_10288,N_9787,N_9810);
nor U10289 (N_10289,N_9531,N_9776);
or U10290 (N_10290,N_9471,N_9539);
xor U10291 (N_10291,N_9214,N_9521);
nand U10292 (N_10292,N_9247,N_9456);
xor U10293 (N_10293,N_9084,N_9265);
nand U10294 (N_10294,N_9709,N_9613);
xnor U10295 (N_10295,N_9852,N_9564);
or U10296 (N_10296,N_9487,N_9905);
and U10297 (N_10297,N_9429,N_9761);
and U10298 (N_10298,N_9039,N_9948);
or U10299 (N_10299,N_9604,N_9102);
and U10300 (N_10300,N_9241,N_9998);
or U10301 (N_10301,N_9254,N_9217);
and U10302 (N_10302,N_9445,N_9106);
nand U10303 (N_10303,N_9263,N_9189);
nor U10304 (N_10304,N_9926,N_9653);
nor U10305 (N_10305,N_9519,N_9399);
xor U10306 (N_10306,N_9255,N_9320);
xnor U10307 (N_10307,N_9131,N_9860);
or U10308 (N_10308,N_9778,N_9971);
nor U10309 (N_10309,N_9348,N_9415);
or U10310 (N_10310,N_9301,N_9702);
nor U10311 (N_10311,N_9194,N_9413);
xor U10312 (N_10312,N_9095,N_9915);
and U10313 (N_10313,N_9294,N_9628);
nor U10314 (N_10314,N_9468,N_9969);
nand U10315 (N_10315,N_9638,N_9453);
xnor U10316 (N_10316,N_9428,N_9216);
or U10317 (N_10317,N_9569,N_9542);
or U10318 (N_10318,N_9641,N_9112);
xor U10319 (N_10319,N_9803,N_9198);
nor U10320 (N_10320,N_9565,N_9222);
xor U10321 (N_10321,N_9680,N_9457);
nand U10322 (N_10322,N_9715,N_9272);
xor U10323 (N_10323,N_9793,N_9988);
xnor U10324 (N_10324,N_9125,N_9900);
nand U10325 (N_10325,N_9823,N_9274);
nor U10326 (N_10326,N_9114,N_9833);
and U10327 (N_10327,N_9176,N_9436);
nor U10328 (N_10328,N_9098,N_9234);
and U10329 (N_10329,N_9339,N_9662);
xnor U10330 (N_10330,N_9755,N_9861);
nand U10331 (N_10331,N_9373,N_9885);
xnor U10332 (N_10332,N_9654,N_9750);
nor U10333 (N_10333,N_9184,N_9001);
and U10334 (N_10334,N_9989,N_9711);
nand U10335 (N_10335,N_9668,N_9693);
xnor U10336 (N_10336,N_9288,N_9908);
nor U10337 (N_10337,N_9200,N_9875);
nand U10338 (N_10338,N_9169,N_9884);
xnor U10339 (N_10339,N_9997,N_9814);
or U10340 (N_10340,N_9034,N_9919);
xnor U10341 (N_10341,N_9078,N_9117);
and U10342 (N_10342,N_9700,N_9991);
nor U10343 (N_10343,N_9435,N_9502);
xor U10344 (N_10344,N_9686,N_9177);
xnor U10345 (N_10345,N_9647,N_9284);
nor U10346 (N_10346,N_9351,N_9784);
xor U10347 (N_10347,N_9777,N_9244);
or U10348 (N_10348,N_9261,N_9208);
nand U10349 (N_10349,N_9477,N_9985);
and U10350 (N_10350,N_9252,N_9472);
and U10351 (N_10351,N_9626,N_9166);
nand U10352 (N_10352,N_9053,N_9337);
nor U10353 (N_10353,N_9328,N_9367);
nand U10354 (N_10354,N_9465,N_9878);
xor U10355 (N_10355,N_9183,N_9303);
xor U10356 (N_10356,N_9928,N_9961);
xor U10357 (N_10357,N_9380,N_9338);
nand U10358 (N_10358,N_9004,N_9152);
and U10359 (N_10359,N_9738,N_9656);
nand U10360 (N_10360,N_9340,N_9505);
or U10361 (N_10361,N_9486,N_9175);
nor U10362 (N_10362,N_9855,N_9822);
nor U10363 (N_10363,N_9674,N_9887);
nand U10364 (N_10364,N_9594,N_9313);
and U10365 (N_10365,N_9221,N_9904);
nor U10366 (N_10366,N_9798,N_9238);
and U10367 (N_10367,N_9403,N_9824);
nor U10368 (N_10368,N_9132,N_9492);
and U10369 (N_10369,N_9270,N_9285);
nor U10370 (N_10370,N_9432,N_9005);
nand U10371 (N_10371,N_9006,N_9289);
nand U10372 (N_10372,N_9586,N_9695);
xnor U10373 (N_10373,N_9841,N_9305);
nand U10374 (N_10374,N_9879,N_9847);
xnor U10375 (N_10375,N_9792,N_9473);
and U10376 (N_10376,N_9946,N_9681);
or U10377 (N_10377,N_9865,N_9913);
xnor U10378 (N_10378,N_9046,N_9085);
xor U10379 (N_10379,N_9547,N_9510);
xnor U10380 (N_10380,N_9296,N_9568);
xnor U10381 (N_10381,N_9074,N_9139);
and U10382 (N_10382,N_9191,N_9639);
and U10383 (N_10383,N_9495,N_9498);
nand U10384 (N_10384,N_9317,N_9437);
nor U10385 (N_10385,N_9901,N_9308);
nand U10386 (N_10386,N_9891,N_9876);
nor U10387 (N_10387,N_9019,N_9678);
or U10388 (N_10388,N_9405,N_9425);
nand U10389 (N_10389,N_9496,N_9555);
nand U10390 (N_10390,N_9658,N_9406);
nor U10391 (N_10391,N_9426,N_9330);
and U10392 (N_10392,N_9327,N_9366);
nor U10393 (N_10393,N_9756,N_9483);
and U10394 (N_10394,N_9922,N_9890);
nor U10395 (N_10395,N_9563,N_9584);
nand U10396 (N_10396,N_9617,N_9086);
xnor U10397 (N_10397,N_9331,N_9608);
and U10398 (N_10398,N_9635,N_9316);
nand U10399 (N_10399,N_9939,N_9732);
nor U10400 (N_10400,N_9129,N_9504);
and U10401 (N_10401,N_9063,N_9060);
nand U10402 (N_10402,N_9423,N_9730);
nor U10403 (N_10403,N_9113,N_9731);
and U10404 (N_10404,N_9574,N_9411);
and U10405 (N_10405,N_9691,N_9110);
nand U10406 (N_10406,N_9292,N_9306);
and U10407 (N_10407,N_9204,N_9872);
xnor U10408 (N_10408,N_9534,N_9089);
xnor U10409 (N_10409,N_9612,N_9986);
nor U10410 (N_10410,N_9839,N_9182);
xnor U10411 (N_10411,N_9856,N_9233);
nor U10412 (N_10412,N_9657,N_9050);
nor U10413 (N_10413,N_9137,N_9964);
nand U10414 (N_10414,N_9577,N_9314);
nand U10415 (N_10415,N_9056,N_9758);
nor U10416 (N_10416,N_9744,N_9920);
and U10417 (N_10417,N_9013,N_9721);
or U10418 (N_10418,N_9115,N_9955);
and U10419 (N_10419,N_9350,N_9557);
nor U10420 (N_10420,N_9291,N_9076);
nand U10421 (N_10421,N_9368,N_9044);
xnor U10422 (N_10422,N_9008,N_9251);
and U10423 (N_10423,N_9377,N_9142);
or U10424 (N_10424,N_9451,N_9925);
or U10425 (N_10425,N_9174,N_9384);
or U10426 (N_10426,N_9766,N_9501);
xnor U10427 (N_10427,N_9347,N_9181);
and U10428 (N_10428,N_9930,N_9770);
or U10429 (N_10429,N_9918,N_9130);
or U10430 (N_10430,N_9829,N_9775);
nor U10431 (N_10431,N_9588,N_9047);
or U10432 (N_10432,N_9950,N_9128);
nor U10433 (N_10433,N_9993,N_9665);
xnor U10434 (N_10434,N_9070,N_9754);
nand U10435 (N_10435,N_9818,N_9632);
nor U10436 (N_10436,N_9023,N_9578);
and U10437 (N_10437,N_9092,N_9655);
nor U10438 (N_10438,N_9346,N_9688);
xnor U10439 (N_10439,N_9213,N_9279);
xor U10440 (N_10440,N_9211,N_9894);
xnor U10441 (N_10441,N_9560,N_9398);
nor U10442 (N_10442,N_9703,N_9172);
or U10443 (N_10443,N_9945,N_9035);
or U10444 (N_10444,N_9706,N_9836);
and U10445 (N_10445,N_9748,N_9851);
xnor U10446 (N_10446,N_9548,N_9149);
nor U10447 (N_10447,N_9834,N_9120);
nor U10448 (N_10448,N_9724,N_9321);
or U10449 (N_10449,N_9645,N_9037);
or U10450 (N_10450,N_9235,N_9161);
nor U10451 (N_10451,N_9910,N_9740);
nand U10452 (N_10452,N_9134,N_9813);
xor U10453 (N_10453,N_9069,N_9277);
nor U10454 (N_10454,N_9173,N_9508);
nand U10455 (N_10455,N_9271,N_9065);
nand U10456 (N_10456,N_9541,N_9585);
and U10457 (N_10457,N_9002,N_9528);
nor U10458 (N_10458,N_9336,N_9148);
xnor U10459 (N_10459,N_9479,N_9982);
nor U10460 (N_10460,N_9932,N_9156);
nor U10461 (N_10461,N_9960,N_9916);
and U10462 (N_10462,N_9520,N_9980);
nand U10463 (N_10463,N_9369,N_9517);
or U10464 (N_10464,N_9804,N_9698);
nand U10465 (N_10465,N_9687,N_9769);
nand U10466 (N_10466,N_9973,N_9601);
nand U10467 (N_10467,N_9772,N_9391);
nand U10468 (N_10468,N_9150,N_9248);
nor U10469 (N_10469,N_9509,N_9147);
xor U10470 (N_10470,N_9269,N_9636);
xnor U10471 (N_10471,N_9990,N_9124);
and U10472 (N_10472,N_9575,N_9138);
nand U10473 (N_10473,N_9397,N_9806);
nor U10474 (N_10474,N_9512,N_9941);
nand U10475 (N_10475,N_9583,N_9041);
nand U10476 (N_10476,N_9760,N_9917);
xnor U10477 (N_10477,N_9103,N_9418);
and U10478 (N_10478,N_9109,N_9326);
nand U10479 (N_10479,N_9205,N_9051);
or U10480 (N_10480,N_9057,N_9490);
and U10481 (N_10481,N_9021,N_9381);
xor U10482 (N_10482,N_9107,N_9746);
or U10483 (N_10483,N_9077,N_9951);
and U10484 (N_10484,N_9762,N_9868);
or U10485 (N_10485,N_9178,N_9970);
nor U10486 (N_10486,N_9959,N_9571);
nand U10487 (N_10487,N_9225,N_9609);
nand U10488 (N_10488,N_9068,N_9491);
or U10489 (N_10489,N_9661,N_9417);
and U10490 (N_10490,N_9849,N_9689);
nor U10491 (N_10491,N_9853,N_9845);
nor U10492 (N_10492,N_9815,N_9032);
or U10493 (N_10493,N_9914,N_9659);
and U10494 (N_10494,N_9024,N_9895);
xnor U10495 (N_10495,N_9424,N_9215);
nand U10496 (N_10496,N_9268,N_9899);
or U10497 (N_10497,N_9669,N_9304);
nor U10498 (N_10498,N_9016,N_9224);
or U10499 (N_10499,N_9480,N_9118);
nor U10500 (N_10500,N_9579,N_9859);
nor U10501 (N_10501,N_9276,N_9541);
xor U10502 (N_10502,N_9010,N_9449);
nor U10503 (N_10503,N_9102,N_9493);
and U10504 (N_10504,N_9357,N_9337);
nor U10505 (N_10505,N_9516,N_9337);
nand U10506 (N_10506,N_9268,N_9182);
and U10507 (N_10507,N_9298,N_9938);
nand U10508 (N_10508,N_9851,N_9416);
and U10509 (N_10509,N_9246,N_9717);
nor U10510 (N_10510,N_9604,N_9468);
nor U10511 (N_10511,N_9000,N_9604);
xor U10512 (N_10512,N_9835,N_9907);
or U10513 (N_10513,N_9564,N_9995);
and U10514 (N_10514,N_9879,N_9702);
or U10515 (N_10515,N_9162,N_9361);
and U10516 (N_10516,N_9304,N_9924);
nor U10517 (N_10517,N_9482,N_9463);
or U10518 (N_10518,N_9133,N_9123);
nor U10519 (N_10519,N_9734,N_9884);
nor U10520 (N_10520,N_9878,N_9206);
nand U10521 (N_10521,N_9295,N_9438);
nand U10522 (N_10522,N_9105,N_9882);
or U10523 (N_10523,N_9381,N_9149);
and U10524 (N_10524,N_9808,N_9368);
xnor U10525 (N_10525,N_9075,N_9500);
xor U10526 (N_10526,N_9723,N_9322);
nor U10527 (N_10527,N_9754,N_9496);
and U10528 (N_10528,N_9817,N_9878);
or U10529 (N_10529,N_9717,N_9805);
xor U10530 (N_10530,N_9817,N_9630);
and U10531 (N_10531,N_9130,N_9828);
nor U10532 (N_10532,N_9065,N_9996);
or U10533 (N_10533,N_9649,N_9971);
or U10534 (N_10534,N_9709,N_9293);
nand U10535 (N_10535,N_9390,N_9500);
or U10536 (N_10536,N_9469,N_9074);
and U10537 (N_10537,N_9104,N_9774);
and U10538 (N_10538,N_9759,N_9793);
xnor U10539 (N_10539,N_9945,N_9659);
and U10540 (N_10540,N_9646,N_9271);
xor U10541 (N_10541,N_9144,N_9091);
xnor U10542 (N_10542,N_9427,N_9919);
or U10543 (N_10543,N_9654,N_9454);
and U10544 (N_10544,N_9966,N_9836);
nor U10545 (N_10545,N_9867,N_9979);
nor U10546 (N_10546,N_9694,N_9645);
and U10547 (N_10547,N_9914,N_9073);
nor U10548 (N_10548,N_9303,N_9922);
nand U10549 (N_10549,N_9509,N_9340);
or U10550 (N_10550,N_9825,N_9120);
xor U10551 (N_10551,N_9404,N_9406);
nor U10552 (N_10552,N_9465,N_9776);
nor U10553 (N_10553,N_9646,N_9920);
nor U10554 (N_10554,N_9544,N_9756);
xnor U10555 (N_10555,N_9354,N_9062);
and U10556 (N_10556,N_9343,N_9607);
nor U10557 (N_10557,N_9335,N_9552);
xnor U10558 (N_10558,N_9797,N_9668);
nor U10559 (N_10559,N_9078,N_9615);
xor U10560 (N_10560,N_9130,N_9750);
nor U10561 (N_10561,N_9874,N_9413);
xnor U10562 (N_10562,N_9816,N_9519);
nor U10563 (N_10563,N_9334,N_9951);
or U10564 (N_10564,N_9303,N_9636);
nor U10565 (N_10565,N_9866,N_9159);
or U10566 (N_10566,N_9862,N_9387);
nor U10567 (N_10567,N_9465,N_9561);
nand U10568 (N_10568,N_9735,N_9618);
or U10569 (N_10569,N_9553,N_9973);
and U10570 (N_10570,N_9963,N_9242);
nor U10571 (N_10571,N_9199,N_9928);
and U10572 (N_10572,N_9113,N_9354);
or U10573 (N_10573,N_9526,N_9869);
nand U10574 (N_10574,N_9718,N_9493);
nand U10575 (N_10575,N_9170,N_9020);
and U10576 (N_10576,N_9073,N_9165);
and U10577 (N_10577,N_9805,N_9482);
nor U10578 (N_10578,N_9782,N_9498);
or U10579 (N_10579,N_9007,N_9879);
or U10580 (N_10580,N_9805,N_9190);
xor U10581 (N_10581,N_9884,N_9299);
or U10582 (N_10582,N_9638,N_9550);
or U10583 (N_10583,N_9459,N_9218);
nor U10584 (N_10584,N_9175,N_9171);
nand U10585 (N_10585,N_9358,N_9102);
xnor U10586 (N_10586,N_9183,N_9852);
nand U10587 (N_10587,N_9588,N_9041);
or U10588 (N_10588,N_9826,N_9719);
nor U10589 (N_10589,N_9844,N_9473);
xor U10590 (N_10590,N_9870,N_9744);
xnor U10591 (N_10591,N_9080,N_9371);
and U10592 (N_10592,N_9284,N_9296);
and U10593 (N_10593,N_9525,N_9450);
and U10594 (N_10594,N_9311,N_9393);
xor U10595 (N_10595,N_9825,N_9494);
or U10596 (N_10596,N_9399,N_9569);
nand U10597 (N_10597,N_9359,N_9688);
nand U10598 (N_10598,N_9321,N_9189);
nor U10599 (N_10599,N_9388,N_9610);
nand U10600 (N_10600,N_9257,N_9031);
xor U10601 (N_10601,N_9147,N_9696);
or U10602 (N_10602,N_9198,N_9795);
xnor U10603 (N_10603,N_9603,N_9695);
or U10604 (N_10604,N_9442,N_9846);
xor U10605 (N_10605,N_9049,N_9173);
nand U10606 (N_10606,N_9492,N_9973);
nor U10607 (N_10607,N_9470,N_9867);
nand U10608 (N_10608,N_9311,N_9455);
and U10609 (N_10609,N_9767,N_9985);
or U10610 (N_10610,N_9049,N_9638);
or U10611 (N_10611,N_9790,N_9411);
nand U10612 (N_10612,N_9473,N_9125);
nor U10613 (N_10613,N_9539,N_9814);
xnor U10614 (N_10614,N_9254,N_9826);
or U10615 (N_10615,N_9375,N_9939);
xor U10616 (N_10616,N_9127,N_9974);
nand U10617 (N_10617,N_9184,N_9640);
xnor U10618 (N_10618,N_9223,N_9327);
and U10619 (N_10619,N_9799,N_9988);
nand U10620 (N_10620,N_9628,N_9238);
xnor U10621 (N_10621,N_9546,N_9117);
nor U10622 (N_10622,N_9988,N_9769);
and U10623 (N_10623,N_9557,N_9756);
xor U10624 (N_10624,N_9758,N_9232);
or U10625 (N_10625,N_9166,N_9357);
and U10626 (N_10626,N_9467,N_9341);
or U10627 (N_10627,N_9128,N_9125);
nor U10628 (N_10628,N_9293,N_9896);
or U10629 (N_10629,N_9070,N_9293);
and U10630 (N_10630,N_9742,N_9475);
nor U10631 (N_10631,N_9590,N_9124);
or U10632 (N_10632,N_9174,N_9861);
nor U10633 (N_10633,N_9291,N_9398);
nand U10634 (N_10634,N_9911,N_9650);
nand U10635 (N_10635,N_9874,N_9848);
and U10636 (N_10636,N_9084,N_9339);
or U10637 (N_10637,N_9654,N_9096);
nand U10638 (N_10638,N_9124,N_9252);
and U10639 (N_10639,N_9354,N_9551);
xnor U10640 (N_10640,N_9561,N_9890);
nand U10641 (N_10641,N_9682,N_9184);
and U10642 (N_10642,N_9949,N_9406);
and U10643 (N_10643,N_9653,N_9045);
and U10644 (N_10644,N_9070,N_9127);
and U10645 (N_10645,N_9677,N_9239);
or U10646 (N_10646,N_9761,N_9617);
or U10647 (N_10647,N_9084,N_9729);
nand U10648 (N_10648,N_9594,N_9433);
or U10649 (N_10649,N_9907,N_9694);
and U10650 (N_10650,N_9970,N_9792);
or U10651 (N_10651,N_9873,N_9493);
or U10652 (N_10652,N_9812,N_9888);
xor U10653 (N_10653,N_9620,N_9310);
nor U10654 (N_10654,N_9537,N_9131);
nor U10655 (N_10655,N_9415,N_9567);
or U10656 (N_10656,N_9216,N_9735);
nand U10657 (N_10657,N_9386,N_9010);
and U10658 (N_10658,N_9482,N_9170);
and U10659 (N_10659,N_9754,N_9760);
nor U10660 (N_10660,N_9201,N_9449);
nor U10661 (N_10661,N_9538,N_9188);
and U10662 (N_10662,N_9766,N_9162);
xor U10663 (N_10663,N_9839,N_9422);
xor U10664 (N_10664,N_9154,N_9873);
nand U10665 (N_10665,N_9330,N_9918);
and U10666 (N_10666,N_9534,N_9034);
and U10667 (N_10667,N_9844,N_9400);
xnor U10668 (N_10668,N_9399,N_9189);
nand U10669 (N_10669,N_9467,N_9696);
nor U10670 (N_10670,N_9125,N_9674);
and U10671 (N_10671,N_9593,N_9355);
and U10672 (N_10672,N_9392,N_9089);
and U10673 (N_10673,N_9032,N_9021);
or U10674 (N_10674,N_9812,N_9309);
and U10675 (N_10675,N_9468,N_9707);
xor U10676 (N_10676,N_9532,N_9173);
xnor U10677 (N_10677,N_9186,N_9341);
nor U10678 (N_10678,N_9330,N_9388);
nand U10679 (N_10679,N_9015,N_9677);
xor U10680 (N_10680,N_9462,N_9054);
xor U10681 (N_10681,N_9231,N_9333);
nand U10682 (N_10682,N_9617,N_9366);
nand U10683 (N_10683,N_9974,N_9344);
or U10684 (N_10684,N_9672,N_9916);
xnor U10685 (N_10685,N_9606,N_9892);
nor U10686 (N_10686,N_9038,N_9275);
or U10687 (N_10687,N_9486,N_9458);
nor U10688 (N_10688,N_9090,N_9401);
nand U10689 (N_10689,N_9577,N_9033);
or U10690 (N_10690,N_9816,N_9052);
nand U10691 (N_10691,N_9645,N_9629);
nand U10692 (N_10692,N_9878,N_9431);
nor U10693 (N_10693,N_9556,N_9766);
xnor U10694 (N_10694,N_9183,N_9111);
and U10695 (N_10695,N_9358,N_9687);
nor U10696 (N_10696,N_9652,N_9444);
and U10697 (N_10697,N_9797,N_9173);
xor U10698 (N_10698,N_9080,N_9158);
xnor U10699 (N_10699,N_9687,N_9877);
or U10700 (N_10700,N_9995,N_9073);
xor U10701 (N_10701,N_9602,N_9656);
nor U10702 (N_10702,N_9279,N_9432);
and U10703 (N_10703,N_9414,N_9366);
nor U10704 (N_10704,N_9002,N_9992);
and U10705 (N_10705,N_9820,N_9238);
xnor U10706 (N_10706,N_9037,N_9836);
nand U10707 (N_10707,N_9127,N_9824);
xor U10708 (N_10708,N_9732,N_9230);
xnor U10709 (N_10709,N_9546,N_9498);
and U10710 (N_10710,N_9259,N_9290);
xor U10711 (N_10711,N_9067,N_9817);
nand U10712 (N_10712,N_9380,N_9455);
xnor U10713 (N_10713,N_9388,N_9352);
nand U10714 (N_10714,N_9311,N_9397);
nand U10715 (N_10715,N_9395,N_9714);
or U10716 (N_10716,N_9867,N_9333);
xnor U10717 (N_10717,N_9866,N_9309);
nor U10718 (N_10718,N_9573,N_9011);
and U10719 (N_10719,N_9730,N_9775);
xnor U10720 (N_10720,N_9278,N_9344);
and U10721 (N_10721,N_9108,N_9556);
nand U10722 (N_10722,N_9015,N_9212);
xor U10723 (N_10723,N_9497,N_9126);
nand U10724 (N_10724,N_9322,N_9617);
nor U10725 (N_10725,N_9082,N_9449);
nand U10726 (N_10726,N_9775,N_9361);
nor U10727 (N_10727,N_9787,N_9158);
or U10728 (N_10728,N_9195,N_9591);
nand U10729 (N_10729,N_9029,N_9744);
nor U10730 (N_10730,N_9043,N_9159);
xnor U10731 (N_10731,N_9840,N_9950);
or U10732 (N_10732,N_9488,N_9694);
or U10733 (N_10733,N_9871,N_9186);
nor U10734 (N_10734,N_9622,N_9948);
xor U10735 (N_10735,N_9889,N_9550);
xor U10736 (N_10736,N_9395,N_9723);
nor U10737 (N_10737,N_9152,N_9245);
or U10738 (N_10738,N_9568,N_9312);
nand U10739 (N_10739,N_9542,N_9383);
nor U10740 (N_10740,N_9262,N_9497);
and U10741 (N_10741,N_9175,N_9132);
nand U10742 (N_10742,N_9076,N_9566);
nand U10743 (N_10743,N_9373,N_9101);
xnor U10744 (N_10744,N_9576,N_9225);
or U10745 (N_10745,N_9691,N_9479);
nand U10746 (N_10746,N_9514,N_9881);
nor U10747 (N_10747,N_9969,N_9477);
nand U10748 (N_10748,N_9139,N_9646);
and U10749 (N_10749,N_9441,N_9752);
nand U10750 (N_10750,N_9739,N_9017);
and U10751 (N_10751,N_9682,N_9326);
nand U10752 (N_10752,N_9558,N_9320);
nand U10753 (N_10753,N_9197,N_9572);
nor U10754 (N_10754,N_9546,N_9524);
and U10755 (N_10755,N_9546,N_9874);
xor U10756 (N_10756,N_9913,N_9492);
and U10757 (N_10757,N_9488,N_9087);
xor U10758 (N_10758,N_9779,N_9911);
nand U10759 (N_10759,N_9630,N_9458);
nand U10760 (N_10760,N_9421,N_9336);
nand U10761 (N_10761,N_9834,N_9496);
nor U10762 (N_10762,N_9764,N_9393);
nor U10763 (N_10763,N_9452,N_9212);
and U10764 (N_10764,N_9905,N_9717);
and U10765 (N_10765,N_9023,N_9347);
and U10766 (N_10766,N_9211,N_9292);
xnor U10767 (N_10767,N_9128,N_9078);
nand U10768 (N_10768,N_9650,N_9364);
xnor U10769 (N_10769,N_9027,N_9143);
or U10770 (N_10770,N_9402,N_9143);
nor U10771 (N_10771,N_9370,N_9865);
nand U10772 (N_10772,N_9797,N_9258);
and U10773 (N_10773,N_9585,N_9010);
nand U10774 (N_10774,N_9631,N_9385);
and U10775 (N_10775,N_9519,N_9157);
xor U10776 (N_10776,N_9823,N_9418);
nand U10777 (N_10777,N_9217,N_9703);
or U10778 (N_10778,N_9494,N_9253);
nand U10779 (N_10779,N_9255,N_9858);
nor U10780 (N_10780,N_9097,N_9242);
xor U10781 (N_10781,N_9582,N_9656);
xor U10782 (N_10782,N_9147,N_9492);
and U10783 (N_10783,N_9319,N_9017);
xor U10784 (N_10784,N_9936,N_9052);
or U10785 (N_10785,N_9191,N_9680);
xnor U10786 (N_10786,N_9340,N_9779);
nor U10787 (N_10787,N_9429,N_9283);
nor U10788 (N_10788,N_9802,N_9524);
nor U10789 (N_10789,N_9143,N_9433);
or U10790 (N_10790,N_9134,N_9825);
and U10791 (N_10791,N_9380,N_9275);
and U10792 (N_10792,N_9253,N_9407);
and U10793 (N_10793,N_9630,N_9176);
xnor U10794 (N_10794,N_9960,N_9951);
nor U10795 (N_10795,N_9003,N_9671);
or U10796 (N_10796,N_9080,N_9963);
nand U10797 (N_10797,N_9170,N_9957);
or U10798 (N_10798,N_9455,N_9943);
and U10799 (N_10799,N_9769,N_9551);
nand U10800 (N_10800,N_9636,N_9538);
nor U10801 (N_10801,N_9411,N_9083);
and U10802 (N_10802,N_9903,N_9222);
or U10803 (N_10803,N_9664,N_9449);
nor U10804 (N_10804,N_9888,N_9361);
or U10805 (N_10805,N_9819,N_9784);
or U10806 (N_10806,N_9162,N_9772);
or U10807 (N_10807,N_9072,N_9922);
and U10808 (N_10808,N_9885,N_9449);
nor U10809 (N_10809,N_9661,N_9779);
or U10810 (N_10810,N_9796,N_9374);
xnor U10811 (N_10811,N_9044,N_9524);
xor U10812 (N_10812,N_9854,N_9060);
nand U10813 (N_10813,N_9090,N_9076);
nand U10814 (N_10814,N_9911,N_9142);
xnor U10815 (N_10815,N_9080,N_9233);
nand U10816 (N_10816,N_9636,N_9211);
nand U10817 (N_10817,N_9700,N_9314);
xnor U10818 (N_10818,N_9620,N_9639);
or U10819 (N_10819,N_9668,N_9882);
xnor U10820 (N_10820,N_9200,N_9510);
or U10821 (N_10821,N_9241,N_9210);
or U10822 (N_10822,N_9541,N_9907);
or U10823 (N_10823,N_9485,N_9969);
and U10824 (N_10824,N_9433,N_9256);
xnor U10825 (N_10825,N_9523,N_9139);
and U10826 (N_10826,N_9236,N_9071);
nor U10827 (N_10827,N_9455,N_9902);
and U10828 (N_10828,N_9161,N_9060);
xnor U10829 (N_10829,N_9555,N_9710);
xnor U10830 (N_10830,N_9203,N_9372);
xnor U10831 (N_10831,N_9278,N_9229);
and U10832 (N_10832,N_9354,N_9435);
or U10833 (N_10833,N_9461,N_9595);
nor U10834 (N_10834,N_9262,N_9923);
and U10835 (N_10835,N_9061,N_9849);
and U10836 (N_10836,N_9127,N_9500);
nor U10837 (N_10837,N_9717,N_9949);
and U10838 (N_10838,N_9932,N_9903);
nand U10839 (N_10839,N_9204,N_9546);
and U10840 (N_10840,N_9338,N_9468);
or U10841 (N_10841,N_9101,N_9734);
nand U10842 (N_10842,N_9945,N_9516);
xnor U10843 (N_10843,N_9629,N_9775);
nor U10844 (N_10844,N_9774,N_9133);
nand U10845 (N_10845,N_9132,N_9055);
nand U10846 (N_10846,N_9686,N_9840);
nor U10847 (N_10847,N_9557,N_9589);
xnor U10848 (N_10848,N_9554,N_9912);
or U10849 (N_10849,N_9465,N_9717);
and U10850 (N_10850,N_9617,N_9329);
nor U10851 (N_10851,N_9468,N_9479);
and U10852 (N_10852,N_9749,N_9076);
nor U10853 (N_10853,N_9776,N_9976);
or U10854 (N_10854,N_9440,N_9601);
nand U10855 (N_10855,N_9701,N_9346);
and U10856 (N_10856,N_9967,N_9141);
nor U10857 (N_10857,N_9504,N_9503);
or U10858 (N_10858,N_9957,N_9110);
nand U10859 (N_10859,N_9489,N_9900);
nand U10860 (N_10860,N_9619,N_9096);
xnor U10861 (N_10861,N_9437,N_9770);
nor U10862 (N_10862,N_9384,N_9910);
or U10863 (N_10863,N_9275,N_9320);
or U10864 (N_10864,N_9077,N_9974);
and U10865 (N_10865,N_9045,N_9519);
or U10866 (N_10866,N_9782,N_9612);
nand U10867 (N_10867,N_9434,N_9163);
nand U10868 (N_10868,N_9238,N_9878);
or U10869 (N_10869,N_9423,N_9057);
xnor U10870 (N_10870,N_9174,N_9303);
xor U10871 (N_10871,N_9506,N_9774);
and U10872 (N_10872,N_9038,N_9065);
xnor U10873 (N_10873,N_9491,N_9472);
xnor U10874 (N_10874,N_9153,N_9062);
nor U10875 (N_10875,N_9806,N_9144);
nand U10876 (N_10876,N_9331,N_9469);
xor U10877 (N_10877,N_9483,N_9666);
xnor U10878 (N_10878,N_9159,N_9931);
or U10879 (N_10879,N_9073,N_9844);
nand U10880 (N_10880,N_9556,N_9364);
xnor U10881 (N_10881,N_9711,N_9196);
or U10882 (N_10882,N_9352,N_9645);
and U10883 (N_10883,N_9653,N_9922);
nor U10884 (N_10884,N_9578,N_9456);
xnor U10885 (N_10885,N_9366,N_9101);
nand U10886 (N_10886,N_9821,N_9986);
nor U10887 (N_10887,N_9393,N_9478);
xor U10888 (N_10888,N_9783,N_9531);
or U10889 (N_10889,N_9933,N_9335);
nor U10890 (N_10890,N_9081,N_9816);
nor U10891 (N_10891,N_9802,N_9699);
nand U10892 (N_10892,N_9432,N_9107);
and U10893 (N_10893,N_9433,N_9338);
nand U10894 (N_10894,N_9329,N_9661);
and U10895 (N_10895,N_9563,N_9764);
nand U10896 (N_10896,N_9348,N_9812);
xnor U10897 (N_10897,N_9213,N_9677);
or U10898 (N_10898,N_9723,N_9583);
xnor U10899 (N_10899,N_9495,N_9696);
xnor U10900 (N_10900,N_9516,N_9656);
and U10901 (N_10901,N_9308,N_9122);
and U10902 (N_10902,N_9021,N_9632);
xor U10903 (N_10903,N_9821,N_9400);
nand U10904 (N_10904,N_9650,N_9223);
or U10905 (N_10905,N_9094,N_9819);
nor U10906 (N_10906,N_9740,N_9360);
nand U10907 (N_10907,N_9187,N_9224);
nand U10908 (N_10908,N_9359,N_9088);
nor U10909 (N_10909,N_9629,N_9724);
nand U10910 (N_10910,N_9170,N_9401);
or U10911 (N_10911,N_9465,N_9104);
and U10912 (N_10912,N_9119,N_9045);
nand U10913 (N_10913,N_9724,N_9344);
and U10914 (N_10914,N_9561,N_9529);
or U10915 (N_10915,N_9809,N_9054);
nand U10916 (N_10916,N_9733,N_9659);
nor U10917 (N_10917,N_9046,N_9335);
or U10918 (N_10918,N_9279,N_9000);
and U10919 (N_10919,N_9168,N_9621);
and U10920 (N_10920,N_9946,N_9284);
xor U10921 (N_10921,N_9390,N_9282);
and U10922 (N_10922,N_9147,N_9463);
and U10923 (N_10923,N_9066,N_9796);
xnor U10924 (N_10924,N_9913,N_9442);
nand U10925 (N_10925,N_9162,N_9869);
xor U10926 (N_10926,N_9841,N_9227);
xor U10927 (N_10927,N_9814,N_9709);
nor U10928 (N_10928,N_9835,N_9918);
xnor U10929 (N_10929,N_9754,N_9334);
and U10930 (N_10930,N_9695,N_9203);
nand U10931 (N_10931,N_9328,N_9180);
and U10932 (N_10932,N_9142,N_9967);
or U10933 (N_10933,N_9413,N_9290);
xnor U10934 (N_10934,N_9609,N_9361);
nor U10935 (N_10935,N_9691,N_9109);
and U10936 (N_10936,N_9829,N_9104);
or U10937 (N_10937,N_9990,N_9521);
nand U10938 (N_10938,N_9372,N_9449);
and U10939 (N_10939,N_9303,N_9290);
or U10940 (N_10940,N_9807,N_9819);
xnor U10941 (N_10941,N_9407,N_9502);
xor U10942 (N_10942,N_9960,N_9132);
xnor U10943 (N_10943,N_9548,N_9217);
and U10944 (N_10944,N_9477,N_9370);
xor U10945 (N_10945,N_9238,N_9620);
nand U10946 (N_10946,N_9565,N_9882);
nand U10947 (N_10947,N_9028,N_9601);
xor U10948 (N_10948,N_9549,N_9479);
nor U10949 (N_10949,N_9600,N_9392);
xor U10950 (N_10950,N_9731,N_9906);
and U10951 (N_10951,N_9780,N_9331);
and U10952 (N_10952,N_9437,N_9540);
nand U10953 (N_10953,N_9532,N_9614);
xor U10954 (N_10954,N_9936,N_9872);
xor U10955 (N_10955,N_9753,N_9542);
nor U10956 (N_10956,N_9268,N_9490);
nor U10957 (N_10957,N_9511,N_9097);
or U10958 (N_10958,N_9606,N_9826);
nand U10959 (N_10959,N_9295,N_9294);
nand U10960 (N_10960,N_9186,N_9923);
and U10961 (N_10961,N_9200,N_9686);
xor U10962 (N_10962,N_9002,N_9499);
nand U10963 (N_10963,N_9057,N_9628);
nand U10964 (N_10964,N_9552,N_9868);
or U10965 (N_10965,N_9338,N_9432);
nand U10966 (N_10966,N_9208,N_9064);
or U10967 (N_10967,N_9162,N_9877);
nand U10968 (N_10968,N_9131,N_9083);
nand U10969 (N_10969,N_9666,N_9460);
or U10970 (N_10970,N_9893,N_9155);
nand U10971 (N_10971,N_9029,N_9390);
or U10972 (N_10972,N_9513,N_9735);
nand U10973 (N_10973,N_9439,N_9327);
xor U10974 (N_10974,N_9255,N_9696);
nand U10975 (N_10975,N_9256,N_9228);
nand U10976 (N_10976,N_9163,N_9696);
xor U10977 (N_10977,N_9824,N_9308);
nand U10978 (N_10978,N_9391,N_9179);
nand U10979 (N_10979,N_9249,N_9819);
xor U10980 (N_10980,N_9484,N_9429);
xor U10981 (N_10981,N_9042,N_9736);
and U10982 (N_10982,N_9529,N_9889);
or U10983 (N_10983,N_9175,N_9541);
nand U10984 (N_10984,N_9433,N_9400);
or U10985 (N_10985,N_9752,N_9224);
nand U10986 (N_10986,N_9295,N_9235);
xor U10987 (N_10987,N_9978,N_9851);
and U10988 (N_10988,N_9783,N_9187);
or U10989 (N_10989,N_9324,N_9761);
or U10990 (N_10990,N_9042,N_9198);
or U10991 (N_10991,N_9664,N_9707);
and U10992 (N_10992,N_9735,N_9872);
and U10993 (N_10993,N_9328,N_9900);
and U10994 (N_10994,N_9663,N_9462);
nand U10995 (N_10995,N_9390,N_9581);
nand U10996 (N_10996,N_9149,N_9809);
xnor U10997 (N_10997,N_9838,N_9950);
nor U10998 (N_10998,N_9012,N_9447);
or U10999 (N_10999,N_9284,N_9659);
xor U11000 (N_11000,N_10824,N_10594);
nand U11001 (N_11001,N_10672,N_10139);
nor U11002 (N_11002,N_10954,N_10857);
and U11003 (N_11003,N_10840,N_10542);
and U11004 (N_11004,N_10744,N_10298);
or U11005 (N_11005,N_10043,N_10276);
nand U11006 (N_11006,N_10144,N_10736);
nand U11007 (N_11007,N_10914,N_10417);
and U11008 (N_11008,N_10414,N_10749);
or U11009 (N_11009,N_10547,N_10047);
nand U11010 (N_11010,N_10953,N_10738);
xor U11011 (N_11011,N_10131,N_10653);
or U11012 (N_11012,N_10986,N_10784);
or U11013 (N_11013,N_10752,N_10702);
xor U11014 (N_11014,N_10889,N_10141);
or U11015 (N_11015,N_10091,N_10407);
or U11016 (N_11016,N_10393,N_10999);
and U11017 (N_11017,N_10694,N_10516);
and U11018 (N_11018,N_10105,N_10928);
nor U11019 (N_11019,N_10078,N_10778);
or U11020 (N_11020,N_10279,N_10566);
nand U11021 (N_11021,N_10310,N_10274);
xnor U11022 (N_11022,N_10424,N_10696);
nor U11023 (N_11023,N_10419,N_10995);
nor U11024 (N_11024,N_10917,N_10166);
xnor U11025 (N_11025,N_10009,N_10626);
nor U11026 (N_11026,N_10464,N_10774);
and U11027 (N_11027,N_10526,N_10317);
xor U11028 (N_11028,N_10888,N_10447);
xnor U11029 (N_11029,N_10808,N_10941);
nor U11030 (N_11030,N_10190,N_10116);
and U11031 (N_11031,N_10059,N_10266);
and U11032 (N_11032,N_10320,N_10852);
nand U11033 (N_11033,N_10168,N_10234);
and U11034 (N_11034,N_10125,N_10680);
nand U11035 (N_11035,N_10263,N_10201);
nand U11036 (N_11036,N_10783,N_10056);
xor U11037 (N_11037,N_10389,N_10861);
nand U11038 (N_11038,N_10085,N_10289);
nor U11039 (N_11039,N_10466,N_10907);
nand U11040 (N_11040,N_10291,N_10760);
xnor U11041 (N_11041,N_10346,N_10336);
xor U11042 (N_11042,N_10512,N_10037);
nor U11043 (N_11043,N_10379,N_10835);
nor U11044 (N_11044,N_10947,N_10509);
or U11045 (N_11045,N_10032,N_10106);
or U11046 (N_11046,N_10382,N_10571);
nand U11047 (N_11047,N_10202,N_10120);
xnor U11048 (N_11048,N_10016,N_10026);
or U11049 (N_11049,N_10867,N_10442);
and U11050 (N_11050,N_10014,N_10872);
and U11051 (N_11051,N_10136,N_10612);
or U11052 (N_11052,N_10207,N_10874);
or U11053 (N_11053,N_10950,N_10325);
nor U11054 (N_11054,N_10387,N_10648);
nand U11055 (N_11055,N_10756,N_10821);
or U11056 (N_11056,N_10088,N_10747);
nand U11057 (N_11057,N_10918,N_10652);
nand U11058 (N_11058,N_10458,N_10404);
or U11059 (N_11059,N_10212,N_10195);
nor U11060 (N_11060,N_10405,N_10588);
xor U11061 (N_11061,N_10018,N_10904);
nand U11062 (N_11062,N_10965,N_10275);
xnor U11063 (N_11063,N_10455,N_10446);
and U11064 (N_11064,N_10967,N_10997);
nand U11065 (N_11065,N_10795,N_10484);
or U11066 (N_11066,N_10704,N_10870);
and U11067 (N_11067,N_10545,N_10004);
and U11068 (N_11068,N_10988,N_10911);
or U11069 (N_11069,N_10093,N_10340);
and U11070 (N_11070,N_10173,N_10015);
nand U11071 (N_11071,N_10901,N_10748);
nor U11072 (N_11072,N_10506,N_10062);
or U11073 (N_11073,N_10365,N_10300);
nor U11074 (N_11074,N_10277,N_10580);
or U11075 (N_11075,N_10895,N_10332);
or U11076 (N_11076,N_10625,N_10462);
or U11077 (N_11077,N_10705,N_10159);
and U11078 (N_11078,N_10284,N_10853);
or U11079 (N_11079,N_10601,N_10090);
nor U11080 (N_11080,N_10685,N_10330);
nand U11081 (N_11081,N_10724,N_10482);
and U11082 (N_11082,N_10335,N_10347);
xnor U11083 (N_11083,N_10247,N_10589);
xor U11084 (N_11084,N_10735,N_10786);
or U11085 (N_11085,N_10614,N_10563);
or U11086 (N_11086,N_10104,N_10581);
xor U11087 (N_11087,N_10023,N_10540);
xnor U11088 (N_11088,N_10002,N_10497);
or U11089 (N_11089,N_10210,N_10729);
or U11090 (N_11090,N_10025,N_10794);
xor U11091 (N_11091,N_10645,N_10524);
nand U11092 (N_11092,N_10396,N_10945);
or U11093 (N_11093,N_10380,N_10254);
nor U11094 (N_11094,N_10468,N_10802);
nand U11095 (N_11095,N_10372,N_10719);
and U11096 (N_11096,N_10935,N_10480);
and U11097 (N_11097,N_10664,N_10475);
nor U11098 (N_11098,N_10084,N_10005);
nor U11099 (N_11099,N_10113,N_10528);
nand U11100 (N_11100,N_10041,N_10204);
nand U11101 (N_11101,N_10226,N_10651);
and U11102 (N_11102,N_10513,N_10371);
xor U11103 (N_11103,N_10899,N_10145);
and U11104 (N_11104,N_10492,N_10494);
nor U11105 (N_11105,N_10329,N_10514);
and U11106 (N_11106,N_10287,N_10971);
nor U11107 (N_11107,N_10616,N_10679);
and U11108 (N_11108,N_10171,N_10687);
nand U11109 (N_11109,N_10354,N_10903);
nand U11110 (N_11110,N_10011,N_10631);
or U11111 (N_11111,N_10938,N_10040);
and U11112 (N_11112,N_10345,N_10639);
and U11113 (N_11113,N_10314,N_10536);
xnor U11114 (N_11114,N_10553,N_10875);
nor U11115 (N_11115,N_10073,N_10423);
xnor U11116 (N_11116,N_10886,N_10863);
or U11117 (N_11117,N_10017,N_10147);
or U11118 (N_11118,N_10261,N_10946);
or U11119 (N_11119,N_10172,N_10898);
and U11120 (N_11120,N_10211,N_10523);
nor U11121 (N_11121,N_10613,N_10278);
nor U11122 (N_11122,N_10258,N_10080);
or U11123 (N_11123,N_10757,N_10409);
nand U11124 (N_11124,N_10510,N_10481);
xnor U11125 (N_11125,N_10412,N_10418);
nor U11126 (N_11126,N_10871,N_10792);
nand U11127 (N_11127,N_10896,N_10390);
nor U11128 (N_11128,N_10989,N_10909);
and U11129 (N_11129,N_10257,N_10003);
or U11130 (N_11130,N_10913,N_10498);
nor U11131 (N_11131,N_10237,N_10556);
and U11132 (N_11132,N_10877,N_10158);
nor U11133 (N_11133,N_10764,N_10029);
or U11134 (N_11134,N_10829,N_10457);
and U11135 (N_11135,N_10367,N_10101);
and U11136 (N_11136,N_10815,N_10624);
xor U11137 (N_11137,N_10251,N_10855);
nand U11138 (N_11138,N_10187,N_10349);
nand U11139 (N_11139,N_10054,N_10811);
nor U11140 (N_11140,N_10267,N_10772);
xor U11141 (N_11141,N_10008,N_10103);
or U11142 (N_11142,N_10559,N_10420);
nand U11143 (N_11143,N_10638,N_10079);
and U11144 (N_11144,N_10980,N_10595);
nor U11145 (N_11145,N_10565,N_10717);
xnor U11146 (N_11146,N_10681,N_10007);
xnor U11147 (N_11147,N_10642,N_10496);
xnor U11148 (N_11148,N_10842,N_10573);
xor U11149 (N_11149,N_10205,N_10411);
or U11150 (N_11150,N_10578,N_10527);
or U11151 (N_11151,N_10726,N_10939);
or U11152 (N_11152,N_10436,N_10844);
nand U11153 (N_11153,N_10834,N_10908);
and U11154 (N_11154,N_10931,N_10097);
xor U11155 (N_11155,N_10065,N_10926);
and U11156 (N_11156,N_10453,N_10196);
nand U11157 (N_11157,N_10013,N_10323);
xnor U11158 (N_11158,N_10866,N_10699);
xnor U11159 (N_11159,N_10221,N_10940);
nand U11160 (N_11160,N_10100,N_10296);
nand U11161 (N_11161,N_10433,N_10800);
nor U11162 (N_11162,N_10519,N_10000);
xor U11163 (N_11163,N_10948,N_10951);
and U11164 (N_11164,N_10878,N_10958);
nand U11165 (N_11165,N_10845,N_10984);
or U11166 (N_11166,N_10440,N_10334);
nor U11167 (N_11167,N_10596,N_10788);
nor U11168 (N_11168,N_10095,N_10990);
or U11169 (N_11169,N_10444,N_10174);
nor U11170 (N_11170,N_10394,N_10368);
or U11171 (N_11171,N_10071,N_10213);
nor U11172 (N_11172,N_10401,N_10743);
nand U11173 (N_11173,N_10198,N_10768);
nor U11174 (N_11174,N_10331,N_10359);
nand U11175 (N_11175,N_10437,N_10327);
xnor U11176 (N_11176,N_10012,N_10979);
and U11177 (N_11177,N_10698,N_10902);
or U11178 (N_11178,N_10429,N_10203);
nand U11179 (N_11179,N_10552,N_10894);
and U11180 (N_11180,N_10262,N_10021);
and U11181 (N_11181,N_10303,N_10627);
nand U11182 (N_11182,N_10181,N_10683);
nor U11183 (N_11183,N_10236,N_10856);
xnor U11184 (N_11184,N_10813,N_10673);
nand U11185 (N_11185,N_10881,N_10264);
xor U11186 (N_11186,N_10991,N_10434);
nand U11187 (N_11187,N_10508,N_10530);
nand U11188 (N_11188,N_10488,N_10142);
nor U11189 (N_11189,N_10722,N_10255);
or U11190 (N_11190,N_10656,N_10121);
xnor U11191 (N_11191,N_10633,N_10366);
nand U11192 (N_11192,N_10843,N_10750);
xnor U11193 (N_11193,N_10375,N_10583);
xnor U11194 (N_11194,N_10028,N_10241);
and U11195 (N_11195,N_10265,N_10130);
nor U11196 (N_11196,N_10428,N_10677);
xnor U11197 (N_11197,N_10328,N_10848);
nor U11198 (N_11198,N_10030,N_10406);
nor U11199 (N_11199,N_10410,N_10534);
and U11200 (N_11200,N_10819,N_10402);
nor U11201 (N_11201,N_10799,N_10232);
or U11202 (N_11202,N_10322,N_10024);
nand U11203 (N_11203,N_10053,N_10115);
nand U11204 (N_11204,N_10107,N_10427);
nor U11205 (N_11205,N_10117,N_10930);
xnor U11206 (N_11206,N_10200,N_10776);
and U11207 (N_11207,N_10044,N_10543);
nor U11208 (N_11208,N_10932,N_10377);
or U11209 (N_11209,N_10618,N_10055);
and U11210 (N_11210,N_10966,N_10476);
nor U11211 (N_11211,N_10049,N_10165);
nor U11212 (N_11212,N_10532,N_10689);
or U11213 (N_11213,N_10660,N_10269);
or U11214 (N_11214,N_10193,N_10385);
nor U11215 (N_11215,N_10490,N_10910);
xnor U11216 (N_11216,N_10525,N_10827);
nor U11217 (N_11217,N_10803,N_10723);
nand U11218 (N_11218,N_10884,N_10179);
or U11219 (N_11219,N_10228,N_10363);
nand U11220 (N_11220,N_10242,N_10517);
nand U11221 (N_11221,N_10936,N_10176);
nand U11222 (N_11222,N_10491,N_10970);
and U11223 (N_11223,N_10443,N_10880);
nand U11224 (N_11224,N_10841,N_10123);
nor U11225 (N_11225,N_10246,N_10897);
nor U11226 (N_11226,N_10248,N_10692);
xor U11227 (N_11227,N_10146,N_10397);
xor U11228 (N_11228,N_10092,N_10657);
nor U11229 (N_11229,N_10268,N_10189);
nand U11230 (N_11230,N_10956,N_10283);
nor U11231 (N_11231,N_10885,N_10737);
nand U11232 (N_11232,N_10019,N_10152);
nor U11233 (N_11233,N_10533,N_10493);
nand U11234 (N_11234,N_10197,N_10900);
nor U11235 (N_11235,N_10217,N_10658);
or U11236 (N_11236,N_10727,N_10057);
or U11237 (N_11237,N_10782,N_10549);
xor U11238 (N_11238,N_10781,N_10333);
nor U11239 (N_11239,N_10635,N_10229);
nand U11240 (N_11240,N_10319,N_10182);
or U11241 (N_11241,N_10859,N_10157);
and U11242 (N_11242,N_10122,N_10675);
or U11243 (N_11243,N_10511,N_10669);
or U11244 (N_11244,N_10376,N_10826);
nand U11245 (N_11245,N_10169,N_10691);
nor U11246 (N_11246,N_10972,N_10987);
xnor U11247 (N_11247,N_10400,N_10504);
and U11248 (N_11248,N_10592,N_10148);
and U11249 (N_11249,N_10584,N_10887);
and U11250 (N_11250,N_10807,N_10272);
nand U11251 (N_11251,N_10851,N_10127);
nand U11252 (N_11252,N_10598,N_10183);
and U11253 (N_11253,N_10294,N_10609);
or U11254 (N_11254,N_10539,N_10416);
and U11255 (N_11255,N_10108,N_10133);
xor U11256 (N_11256,N_10473,N_10740);
or U11257 (N_11257,N_10288,N_10318);
xnor U11258 (N_11258,N_10864,N_10033);
nand U11259 (N_11259,N_10912,N_10052);
xnor U11260 (N_11260,N_10576,N_10725);
xnor U11261 (N_11261,N_10500,N_10520);
xnor U11262 (N_11262,N_10695,N_10817);
or U11263 (N_11263,N_10273,N_10035);
nor U11264 (N_11264,N_10215,N_10374);
and U11265 (N_11265,N_10304,N_10072);
and U11266 (N_11266,N_10822,N_10070);
or U11267 (N_11267,N_10637,N_10663);
and U11268 (N_11268,N_10688,N_10467);
xor U11269 (N_11269,N_10555,N_10355);
nor U11270 (N_11270,N_10823,N_10378);
or U11271 (N_11271,N_10293,N_10916);
or U11272 (N_11272,N_10569,N_10925);
and U11273 (N_11273,N_10830,N_10759);
nor U11274 (N_11274,N_10531,N_10575);
nor U11275 (N_11275,N_10998,N_10960);
and U11276 (N_11276,N_10191,N_10620);
xor U11277 (N_11277,N_10798,N_10671);
nand U11278 (N_11278,N_10160,N_10083);
nand U11279 (N_11279,N_10067,N_10138);
nor U11280 (N_11280,N_10600,N_10714);
nand U11281 (N_11281,N_10075,N_10306);
and U11282 (N_11282,N_10369,N_10126);
nor U11283 (N_11283,N_10290,N_10828);
nor U11284 (N_11284,N_10321,N_10010);
nand U11285 (N_11285,N_10985,N_10089);
xnor U11286 (N_11286,N_10244,N_10715);
and U11287 (N_11287,N_10413,N_10716);
nand U11288 (N_11288,N_10804,N_10969);
xor U11289 (N_11289,N_10225,N_10312);
and U11290 (N_11290,N_10483,N_10789);
xnor U11291 (N_11291,N_10350,N_10199);
nor U11292 (N_11292,N_10949,N_10461);
or U11293 (N_11293,N_10066,N_10109);
nand U11294 (N_11294,N_10560,N_10621);
nand U11295 (N_11295,N_10707,N_10188);
and U11296 (N_11296,N_10924,N_10118);
nor U11297 (N_11297,N_10114,N_10599);
and U11298 (N_11298,N_10773,N_10362);
or U11299 (N_11299,N_10441,N_10643);
and U11300 (N_11300,N_10432,N_10448);
and U11301 (N_11301,N_10361,N_10479);
nor U11302 (N_11302,N_10352,N_10311);
nor U11303 (N_11303,N_10710,N_10302);
and U11304 (N_11304,N_10602,N_10295);
nand U11305 (N_11305,N_10449,N_10339);
and U11306 (N_11306,N_10622,N_10868);
xor U11307 (N_11307,N_10684,N_10701);
nand U11308 (N_11308,N_10292,N_10944);
or U11309 (N_11309,N_10048,N_10968);
xnor U11310 (N_11310,N_10718,N_10505);
nor U11311 (N_11311,N_10178,N_10006);
nand U11312 (N_11312,N_10537,N_10617);
nand U11313 (N_11313,N_10557,N_10546);
nand U11314 (N_11314,N_10426,N_10765);
xor U11315 (N_11315,N_10838,N_10299);
xor U11316 (N_11316,N_10551,N_10186);
and U11317 (N_11317,N_10810,N_10020);
or U11318 (N_11318,N_10313,N_10156);
nor U11319 (N_11319,N_10422,N_10833);
nand U11320 (N_11320,N_10623,N_10112);
nand U11321 (N_11321,N_10550,N_10143);
nor U11322 (N_11322,N_10129,N_10451);
nand U11323 (N_11323,N_10096,N_10384);
nand U11324 (N_11324,N_10194,N_10544);
nor U11325 (N_11325,N_10670,N_10185);
nand U11326 (N_11326,N_10963,N_10348);
xnor U11327 (N_11327,N_10450,N_10742);
or U11328 (N_11328,N_10356,N_10846);
or U11329 (N_11329,N_10471,N_10570);
and U11330 (N_11330,N_10398,N_10751);
xor U11331 (N_11331,N_10758,N_10713);
nor U11332 (N_11332,N_10102,N_10392);
xor U11333 (N_11333,N_10046,N_10253);
nor U11334 (N_11334,N_10353,N_10240);
xor U11335 (N_11335,N_10515,N_10170);
nand U11336 (N_11336,N_10487,N_10308);
xnor U11337 (N_11337,N_10820,N_10992);
and U11338 (N_11338,N_10892,N_10590);
or U11339 (N_11339,N_10360,N_10252);
and U11340 (N_11340,N_10522,N_10163);
xnor U11341 (N_11341,N_10184,N_10529);
and U11342 (N_11342,N_10796,N_10730);
nor U11343 (N_11343,N_10162,N_10391);
nand U11344 (N_11344,N_10271,N_10386);
nand U11345 (N_11345,N_10587,N_10474);
or U11346 (N_11346,N_10957,N_10809);
nor U11347 (N_11347,N_10250,N_10050);
xnor U11348 (N_11348,N_10847,N_10465);
nor U11349 (N_11349,N_10456,N_10858);
or U11350 (N_11350,N_10001,N_10501);
and U11351 (N_11351,N_10812,N_10469);
nor U11352 (N_11352,N_10978,N_10069);
nor U11353 (N_11353,N_10206,N_10245);
nor U11354 (N_11354,N_10485,N_10955);
xor U11355 (N_11355,N_10216,N_10739);
or U11356 (N_11356,N_10831,N_10927);
nor U11357 (N_11357,N_10068,N_10061);
and U11358 (N_11358,N_10326,N_10720);
nor U11359 (N_11359,N_10630,N_10135);
and U11360 (N_11360,N_10561,N_10733);
xor U11361 (N_11361,N_10430,N_10119);
xor U11362 (N_11362,N_10882,N_10952);
nand U11363 (N_11363,N_10134,N_10825);
nor U11364 (N_11364,N_10666,N_10922);
nand U11365 (N_11365,N_10256,N_10849);
or U11366 (N_11366,N_10585,N_10929);
or U11367 (N_11367,N_10554,N_10341);
xnor U11368 (N_11368,N_10865,N_10604);
nor U11369 (N_11369,N_10439,N_10214);
and U11370 (N_11370,N_10309,N_10793);
and U11371 (N_11371,N_10767,N_10770);
nor U11372 (N_11372,N_10445,N_10883);
xnor U11373 (N_11373,N_10973,N_10507);
xor U11374 (N_11374,N_10316,N_10408);
nand U11375 (N_11375,N_10270,N_10388);
or U11376 (N_11376,N_10593,N_10154);
and U11377 (N_11377,N_10161,N_10734);
and U11378 (N_11378,N_10579,N_10641);
nand U11379 (N_11379,N_10976,N_10399);
or U11380 (N_11380,N_10606,N_10486);
nand U11381 (N_11381,N_10919,N_10654);
nor U11382 (N_11382,N_10087,N_10661);
xnor U11383 (N_11383,N_10285,N_10787);
xnor U11384 (N_11384,N_10674,N_10502);
nor U11385 (N_11385,N_10489,N_10615);
nor U11386 (N_11386,N_10111,N_10086);
nor U11387 (N_11387,N_10063,N_10538);
xnor U11388 (N_11388,N_10132,N_10222);
nor U11389 (N_11389,N_10582,N_10027);
nand U11390 (N_11390,N_10155,N_10470);
xor U11391 (N_11391,N_10876,N_10690);
nand U11392 (N_11392,N_10854,N_10915);
xnor U11393 (N_11393,N_10659,N_10780);
nand U11394 (N_11394,N_10964,N_10706);
nor U11395 (N_11395,N_10634,N_10572);
nand U11396 (N_11396,N_10640,N_10647);
nand U11397 (N_11397,N_10478,N_10777);
nand U11398 (N_11398,N_10682,N_10150);
xnor U11399 (N_11399,N_10220,N_10324);
or U11400 (N_11400,N_10837,N_10337);
or U11401 (N_11401,N_10249,N_10231);
or U11402 (N_11402,N_10064,N_10962);
xnor U11403 (N_11403,N_10728,N_10814);
nor U11404 (N_11404,N_10975,N_10435);
and U11405 (N_11405,N_10632,N_10454);
xnor U11406 (N_11406,N_10574,N_10905);
nor U11407 (N_11407,N_10686,N_10315);
xor U11408 (N_11408,N_10383,N_10438);
nor U11409 (N_11409,N_10094,N_10535);
nor U11410 (N_11410,N_10791,N_10140);
nor U11411 (N_11411,N_10149,N_10610);
and U11412 (N_11412,N_10869,N_10463);
nor U11413 (N_11413,N_10370,N_10564);
nor U11414 (N_11414,N_10961,N_10873);
and U11415 (N_11415,N_10034,N_10472);
nand U11416 (N_11416,N_10790,N_10906);
and U11417 (N_11417,N_10460,N_10137);
nand U11418 (N_11418,N_10208,N_10230);
xor U11419 (N_11419,N_10124,N_10358);
xnor U11420 (N_11420,N_10153,N_10943);
xor U11421 (N_11421,N_10099,N_10151);
nand U11422 (N_11422,N_10636,N_10223);
xnor U11423 (N_11423,N_10974,N_10619);
and U11424 (N_11424,N_10668,N_10459);
nand U11425 (N_11425,N_10771,N_10697);
nor U11426 (N_11426,N_10934,N_10745);
xnor U11427 (N_11427,N_10562,N_10259);
nand U11428 (N_11428,N_10224,N_10766);
nor U11429 (N_11429,N_10243,N_10629);
nor U11430 (N_11430,N_10942,N_10235);
or U11431 (N_11431,N_10541,N_10175);
xor U11432 (N_11432,N_10754,N_10665);
nand U11433 (N_11433,N_10499,N_10923);
and U11434 (N_11434,N_10708,N_10042);
nand U11435 (N_11435,N_10218,N_10721);
and U11436 (N_11436,N_10732,N_10548);
nor U11437 (N_11437,N_10164,N_10395);
xnor U11438 (N_11438,N_10260,N_10503);
or U11439 (N_11439,N_10676,N_10343);
xnor U11440 (N_11440,N_10477,N_10495);
and U11441 (N_11441,N_10238,N_10180);
xor U11442 (N_11442,N_10605,N_10586);
xor U11443 (N_11443,N_10281,N_10058);
or U11444 (N_11444,N_10558,N_10921);
and U11445 (N_11445,N_10879,N_10753);
xnor U11446 (N_11446,N_10342,N_10051);
xnor U11447 (N_11447,N_10649,N_10761);
nand U11448 (N_11448,N_10098,N_10981);
nand U11449 (N_11449,N_10607,N_10805);
nand U11450 (N_11450,N_10818,N_10775);
nor U11451 (N_11451,N_10893,N_10280);
nor U11452 (N_11452,N_10779,N_10650);
or U11453 (N_11453,N_10364,N_10351);
and U11454 (N_11454,N_10801,N_10282);
and U11455 (N_11455,N_10425,N_10806);
and U11456 (N_11456,N_10381,N_10703);
xor U11457 (N_11457,N_10709,N_10628);
nand U11458 (N_11458,N_10693,N_10128);
nor U11459 (N_11459,N_10039,N_10644);
or U11460 (N_11460,N_10239,N_10431);
or U11461 (N_11461,N_10769,N_10577);
or U11462 (N_11462,N_10036,N_10891);
nand U11463 (N_11463,N_10762,N_10357);
xnor U11464 (N_11464,N_10662,N_10755);
and U11465 (N_11465,N_10746,N_10731);
xor U11466 (N_11466,N_10996,N_10301);
or U11467 (N_11467,N_10983,N_10219);
xor U11468 (N_11468,N_10890,N_10038);
or U11469 (N_11469,N_10177,N_10074);
or U11470 (N_11470,N_10031,N_10712);
xor U11471 (N_11471,N_10667,N_10192);
or U11472 (N_11472,N_10700,N_10937);
nor U11473 (N_11473,N_10611,N_10982);
or U11474 (N_11474,N_10045,N_10603);
nor U11475 (N_11475,N_10959,N_10452);
nor U11476 (N_11476,N_10711,N_10518);
or U11477 (N_11477,N_10082,N_10608);
or U11478 (N_11478,N_10836,N_10022);
and U11479 (N_11479,N_10933,N_10167);
nand U11480 (N_11480,N_10832,N_10860);
or U11481 (N_11481,N_10227,N_10977);
nor U11482 (N_11482,N_10305,N_10060);
xnor U11483 (N_11483,N_10597,N_10994);
or U11484 (N_11484,N_10373,N_10678);
xor U11485 (N_11485,N_10307,N_10655);
or U11486 (N_11486,N_10567,N_10763);
xnor U11487 (N_11487,N_10920,N_10403);
nand U11488 (N_11488,N_10286,N_10081);
and U11489 (N_11489,N_10568,N_10741);
or U11490 (N_11490,N_10797,N_10338);
nand U11491 (N_11491,N_10110,N_10297);
and U11492 (N_11492,N_10421,N_10839);
nor U11493 (N_11493,N_10344,N_10646);
nor U11494 (N_11494,N_10415,N_10785);
nand U11495 (N_11495,N_10076,N_10521);
nand U11496 (N_11496,N_10862,N_10850);
nor U11497 (N_11497,N_10816,N_10233);
and U11498 (N_11498,N_10077,N_10209);
and U11499 (N_11499,N_10993,N_10591);
nor U11500 (N_11500,N_10136,N_10200);
nor U11501 (N_11501,N_10567,N_10644);
xor U11502 (N_11502,N_10295,N_10502);
and U11503 (N_11503,N_10742,N_10655);
nand U11504 (N_11504,N_10465,N_10095);
nor U11505 (N_11505,N_10251,N_10420);
nand U11506 (N_11506,N_10868,N_10073);
nand U11507 (N_11507,N_10006,N_10019);
xor U11508 (N_11508,N_10108,N_10304);
or U11509 (N_11509,N_10512,N_10140);
xnor U11510 (N_11510,N_10063,N_10958);
xnor U11511 (N_11511,N_10238,N_10013);
and U11512 (N_11512,N_10702,N_10972);
nor U11513 (N_11513,N_10919,N_10727);
and U11514 (N_11514,N_10530,N_10539);
nor U11515 (N_11515,N_10725,N_10498);
nor U11516 (N_11516,N_10614,N_10877);
nor U11517 (N_11517,N_10044,N_10031);
and U11518 (N_11518,N_10682,N_10505);
nand U11519 (N_11519,N_10600,N_10890);
and U11520 (N_11520,N_10816,N_10655);
nor U11521 (N_11521,N_10141,N_10384);
or U11522 (N_11522,N_10542,N_10959);
and U11523 (N_11523,N_10064,N_10711);
or U11524 (N_11524,N_10049,N_10270);
and U11525 (N_11525,N_10442,N_10852);
and U11526 (N_11526,N_10527,N_10182);
and U11527 (N_11527,N_10923,N_10281);
and U11528 (N_11528,N_10575,N_10953);
and U11529 (N_11529,N_10739,N_10887);
nor U11530 (N_11530,N_10886,N_10098);
xnor U11531 (N_11531,N_10752,N_10353);
nand U11532 (N_11532,N_10003,N_10907);
xnor U11533 (N_11533,N_10950,N_10013);
and U11534 (N_11534,N_10329,N_10331);
nand U11535 (N_11535,N_10355,N_10864);
or U11536 (N_11536,N_10273,N_10854);
or U11537 (N_11537,N_10470,N_10612);
nor U11538 (N_11538,N_10638,N_10952);
or U11539 (N_11539,N_10427,N_10705);
nand U11540 (N_11540,N_10722,N_10039);
and U11541 (N_11541,N_10291,N_10166);
nand U11542 (N_11542,N_10336,N_10361);
or U11543 (N_11543,N_10135,N_10751);
and U11544 (N_11544,N_10538,N_10721);
nor U11545 (N_11545,N_10949,N_10332);
or U11546 (N_11546,N_10519,N_10378);
nand U11547 (N_11547,N_10609,N_10387);
nand U11548 (N_11548,N_10942,N_10622);
nand U11549 (N_11549,N_10657,N_10604);
and U11550 (N_11550,N_10689,N_10238);
xnor U11551 (N_11551,N_10663,N_10561);
nor U11552 (N_11552,N_10349,N_10862);
xnor U11553 (N_11553,N_10416,N_10422);
and U11554 (N_11554,N_10044,N_10672);
xnor U11555 (N_11555,N_10314,N_10243);
xor U11556 (N_11556,N_10679,N_10048);
nor U11557 (N_11557,N_10674,N_10883);
nand U11558 (N_11558,N_10929,N_10997);
nand U11559 (N_11559,N_10780,N_10707);
nor U11560 (N_11560,N_10913,N_10180);
nor U11561 (N_11561,N_10388,N_10718);
or U11562 (N_11562,N_10205,N_10849);
nor U11563 (N_11563,N_10353,N_10899);
nand U11564 (N_11564,N_10076,N_10392);
nand U11565 (N_11565,N_10286,N_10941);
nand U11566 (N_11566,N_10717,N_10905);
nand U11567 (N_11567,N_10568,N_10333);
or U11568 (N_11568,N_10695,N_10503);
xnor U11569 (N_11569,N_10759,N_10809);
or U11570 (N_11570,N_10951,N_10601);
or U11571 (N_11571,N_10124,N_10118);
nor U11572 (N_11572,N_10043,N_10743);
or U11573 (N_11573,N_10940,N_10672);
and U11574 (N_11574,N_10940,N_10237);
nand U11575 (N_11575,N_10954,N_10399);
nor U11576 (N_11576,N_10488,N_10397);
xor U11577 (N_11577,N_10738,N_10436);
nor U11578 (N_11578,N_10934,N_10827);
xnor U11579 (N_11579,N_10110,N_10983);
and U11580 (N_11580,N_10519,N_10911);
xor U11581 (N_11581,N_10032,N_10234);
xor U11582 (N_11582,N_10448,N_10132);
nand U11583 (N_11583,N_10870,N_10365);
or U11584 (N_11584,N_10661,N_10337);
nand U11585 (N_11585,N_10614,N_10018);
or U11586 (N_11586,N_10360,N_10267);
or U11587 (N_11587,N_10157,N_10854);
xnor U11588 (N_11588,N_10642,N_10847);
or U11589 (N_11589,N_10224,N_10330);
or U11590 (N_11590,N_10288,N_10116);
xor U11591 (N_11591,N_10047,N_10052);
nor U11592 (N_11592,N_10519,N_10196);
xor U11593 (N_11593,N_10602,N_10802);
xor U11594 (N_11594,N_10713,N_10266);
xnor U11595 (N_11595,N_10587,N_10343);
or U11596 (N_11596,N_10420,N_10317);
xnor U11597 (N_11597,N_10408,N_10677);
or U11598 (N_11598,N_10022,N_10713);
xor U11599 (N_11599,N_10189,N_10234);
xor U11600 (N_11600,N_10826,N_10298);
nor U11601 (N_11601,N_10943,N_10497);
xor U11602 (N_11602,N_10354,N_10679);
xor U11603 (N_11603,N_10797,N_10971);
xnor U11604 (N_11604,N_10124,N_10744);
nand U11605 (N_11605,N_10951,N_10073);
and U11606 (N_11606,N_10223,N_10955);
nor U11607 (N_11607,N_10453,N_10910);
nand U11608 (N_11608,N_10136,N_10243);
and U11609 (N_11609,N_10758,N_10862);
and U11610 (N_11610,N_10489,N_10108);
nor U11611 (N_11611,N_10847,N_10809);
xor U11612 (N_11612,N_10047,N_10351);
nand U11613 (N_11613,N_10716,N_10480);
xnor U11614 (N_11614,N_10097,N_10509);
or U11615 (N_11615,N_10310,N_10100);
and U11616 (N_11616,N_10857,N_10982);
xnor U11617 (N_11617,N_10797,N_10287);
nand U11618 (N_11618,N_10192,N_10492);
and U11619 (N_11619,N_10334,N_10834);
or U11620 (N_11620,N_10393,N_10611);
or U11621 (N_11621,N_10586,N_10652);
nand U11622 (N_11622,N_10901,N_10613);
or U11623 (N_11623,N_10853,N_10981);
and U11624 (N_11624,N_10105,N_10386);
xor U11625 (N_11625,N_10709,N_10278);
or U11626 (N_11626,N_10491,N_10198);
xor U11627 (N_11627,N_10302,N_10243);
or U11628 (N_11628,N_10198,N_10823);
nor U11629 (N_11629,N_10490,N_10897);
nor U11630 (N_11630,N_10625,N_10321);
nor U11631 (N_11631,N_10328,N_10906);
nand U11632 (N_11632,N_10208,N_10593);
nand U11633 (N_11633,N_10827,N_10642);
and U11634 (N_11634,N_10015,N_10285);
nor U11635 (N_11635,N_10199,N_10223);
or U11636 (N_11636,N_10041,N_10452);
nand U11637 (N_11637,N_10269,N_10553);
and U11638 (N_11638,N_10315,N_10522);
or U11639 (N_11639,N_10101,N_10444);
nand U11640 (N_11640,N_10812,N_10654);
nand U11641 (N_11641,N_10228,N_10335);
nor U11642 (N_11642,N_10442,N_10418);
xor U11643 (N_11643,N_10592,N_10361);
nand U11644 (N_11644,N_10318,N_10364);
nand U11645 (N_11645,N_10668,N_10386);
nor U11646 (N_11646,N_10316,N_10307);
xnor U11647 (N_11647,N_10259,N_10676);
nor U11648 (N_11648,N_10904,N_10153);
nor U11649 (N_11649,N_10955,N_10054);
xor U11650 (N_11650,N_10991,N_10994);
nor U11651 (N_11651,N_10160,N_10937);
nor U11652 (N_11652,N_10324,N_10409);
and U11653 (N_11653,N_10800,N_10676);
and U11654 (N_11654,N_10373,N_10910);
xor U11655 (N_11655,N_10284,N_10238);
nand U11656 (N_11656,N_10136,N_10379);
xnor U11657 (N_11657,N_10827,N_10027);
xnor U11658 (N_11658,N_10974,N_10862);
or U11659 (N_11659,N_10276,N_10515);
or U11660 (N_11660,N_10140,N_10152);
xor U11661 (N_11661,N_10605,N_10784);
or U11662 (N_11662,N_10494,N_10526);
xor U11663 (N_11663,N_10728,N_10426);
nand U11664 (N_11664,N_10756,N_10015);
xnor U11665 (N_11665,N_10245,N_10762);
nor U11666 (N_11666,N_10614,N_10729);
nand U11667 (N_11667,N_10182,N_10158);
and U11668 (N_11668,N_10120,N_10053);
nor U11669 (N_11669,N_10396,N_10432);
nand U11670 (N_11670,N_10476,N_10065);
nand U11671 (N_11671,N_10490,N_10355);
or U11672 (N_11672,N_10603,N_10665);
xnor U11673 (N_11673,N_10997,N_10946);
nor U11674 (N_11674,N_10043,N_10098);
and U11675 (N_11675,N_10240,N_10430);
or U11676 (N_11676,N_10195,N_10078);
or U11677 (N_11677,N_10034,N_10558);
xor U11678 (N_11678,N_10740,N_10613);
nand U11679 (N_11679,N_10277,N_10912);
nor U11680 (N_11680,N_10902,N_10773);
nor U11681 (N_11681,N_10549,N_10412);
xor U11682 (N_11682,N_10425,N_10632);
and U11683 (N_11683,N_10011,N_10915);
and U11684 (N_11684,N_10153,N_10407);
or U11685 (N_11685,N_10890,N_10339);
nor U11686 (N_11686,N_10104,N_10705);
nand U11687 (N_11687,N_10593,N_10283);
nor U11688 (N_11688,N_10241,N_10629);
or U11689 (N_11689,N_10496,N_10542);
nor U11690 (N_11690,N_10726,N_10724);
nor U11691 (N_11691,N_10062,N_10164);
nor U11692 (N_11692,N_10304,N_10875);
and U11693 (N_11693,N_10781,N_10949);
or U11694 (N_11694,N_10194,N_10745);
nand U11695 (N_11695,N_10246,N_10463);
or U11696 (N_11696,N_10269,N_10179);
or U11697 (N_11697,N_10066,N_10063);
nand U11698 (N_11698,N_10955,N_10721);
xor U11699 (N_11699,N_10237,N_10353);
and U11700 (N_11700,N_10597,N_10852);
or U11701 (N_11701,N_10707,N_10587);
and U11702 (N_11702,N_10710,N_10512);
nor U11703 (N_11703,N_10217,N_10768);
nand U11704 (N_11704,N_10324,N_10720);
and U11705 (N_11705,N_10004,N_10813);
and U11706 (N_11706,N_10173,N_10529);
nand U11707 (N_11707,N_10175,N_10971);
nor U11708 (N_11708,N_10776,N_10903);
and U11709 (N_11709,N_10828,N_10829);
and U11710 (N_11710,N_10058,N_10028);
nand U11711 (N_11711,N_10789,N_10999);
or U11712 (N_11712,N_10362,N_10506);
xnor U11713 (N_11713,N_10163,N_10264);
nor U11714 (N_11714,N_10857,N_10161);
nand U11715 (N_11715,N_10431,N_10221);
and U11716 (N_11716,N_10474,N_10630);
nor U11717 (N_11717,N_10087,N_10559);
and U11718 (N_11718,N_10472,N_10947);
xor U11719 (N_11719,N_10079,N_10688);
nand U11720 (N_11720,N_10833,N_10214);
or U11721 (N_11721,N_10801,N_10413);
xor U11722 (N_11722,N_10115,N_10268);
and U11723 (N_11723,N_10414,N_10102);
nor U11724 (N_11724,N_10375,N_10580);
nor U11725 (N_11725,N_10542,N_10112);
xor U11726 (N_11726,N_10057,N_10759);
nand U11727 (N_11727,N_10812,N_10273);
xnor U11728 (N_11728,N_10547,N_10085);
nor U11729 (N_11729,N_10148,N_10759);
nor U11730 (N_11730,N_10396,N_10428);
nor U11731 (N_11731,N_10072,N_10353);
and U11732 (N_11732,N_10606,N_10858);
and U11733 (N_11733,N_10915,N_10342);
nor U11734 (N_11734,N_10734,N_10184);
nor U11735 (N_11735,N_10559,N_10873);
nand U11736 (N_11736,N_10529,N_10921);
and U11737 (N_11737,N_10701,N_10555);
and U11738 (N_11738,N_10871,N_10216);
nand U11739 (N_11739,N_10436,N_10965);
nand U11740 (N_11740,N_10573,N_10582);
nor U11741 (N_11741,N_10242,N_10795);
and U11742 (N_11742,N_10843,N_10297);
or U11743 (N_11743,N_10187,N_10324);
xor U11744 (N_11744,N_10521,N_10845);
nand U11745 (N_11745,N_10514,N_10542);
and U11746 (N_11746,N_10215,N_10945);
xnor U11747 (N_11747,N_10463,N_10475);
or U11748 (N_11748,N_10704,N_10755);
nor U11749 (N_11749,N_10057,N_10878);
nand U11750 (N_11750,N_10259,N_10213);
or U11751 (N_11751,N_10821,N_10365);
nand U11752 (N_11752,N_10745,N_10959);
xor U11753 (N_11753,N_10824,N_10479);
or U11754 (N_11754,N_10231,N_10516);
xor U11755 (N_11755,N_10708,N_10279);
or U11756 (N_11756,N_10490,N_10575);
xor U11757 (N_11757,N_10948,N_10511);
or U11758 (N_11758,N_10901,N_10196);
or U11759 (N_11759,N_10536,N_10281);
xor U11760 (N_11760,N_10992,N_10698);
nor U11761 (N_11761,N_10987,N_10302);
xor U11762 (N_11762,N_10563,N_10670);
nand U11763 (N_11763,N_10753,N_10976);
or U11764 (N_11764,N_10971,N_10669);
nand U11765 (N_11765,N_10431,N_10947);
and U11766 (N_11766,N_10011,N_10556);
xnor U11767 (N_11767,N_10703,N_10415);
nor U11768 (N_11768,N_10432,N_10447);
and U11769 (N_11769,N_10096,N_10103);
nor U11770 (N_11770,N_10357,N_10289);
nand U11771 (N_11771,N_10228,N_10264);
nand U11772 (N_11772,N_10059,N_10717);
nand U11773 (N_11773,N_10560,N_10765);
or U11774 (N_11774,N_10692,N_10469);
nor U11775 (N_11775,N_10882,N_10164);
and U11776 (N_11776,N_10458,N_10640);
nand U11777 (N_11777,N_10983,N_10264);
xnor U11778 (N_11778,N_10674,N_10647);
nor U11779 (N_11779,N_10610,N_10437);
nor U11780 (N_11780,N_10672,N_10763);
nor U11781 (N_11781,N_10049,N_10597);
nor U11782 (N_11782,N_10214,N_10186);
nor U11783 (N_11783,N_10971,N_10016);
or U11784 (N_11784,N_10489,N_10026);
nor U11785 (N_11785,N_10546,N_10063);
or U11786 (N_11786,N_10777,N_10064);
nor U11787 (N_11787,N_10547,N_10406);
or U11788 (N_11788,N_10245,N_10056);
xnor U11789 (N_11789,N_10830,N_10698);
nor U11790 (N_11790,N_10731,N_10933);
xnor U11791 (N_11791,N_10419,N_10846);
nor U11792 (N_11792,N_10277,N_10972);
nor U11793 (N_11793,N_10681,N_10905);
nor U11794 (N_11794,N_10681,N_10803);
nor U11795 (N_11795,N_10552,N_10259);
and U11796 (N_11796,N_10115,N_10830);
nand U11797 (N_11797,N_10320,N_10225);
nand U11798 (N_11798,N_10956,N_10490);
nand U11799 (N_11799,N_10363,N_10726);
and U11800 (N_11800,N_10668,N_10420);
xor U11801 (N_11801,N_10035,N_10405);
nor U11802 (N_11802,N_10699,N_10401);
and U11803 (N_11803,N_10745,N_10403);
nor U11804 (N_11804,N_10260,N_10138);
nor U11805 (N_11805,N_10992,N_10306);
and U11806 (N_11806,N_10110,N_10713);
nand U11807 (N_11807,N_10026,N_10959);
xnor U11808 (N_11808,N_10991,N_10487);
or U11809 (N_11809,N_10746,N_10471);
or U11810 (N_11810,N_10930,N_10995);
and U11811 (N_11811,N_10705,N_10346);
and U11812 (N_11812,N_10039,N_10385);
xnor U11813 (N_11813,N_10211,N_10186);
and U11814 (N_11814,N_10990,N_10691);
xor U11815 (N_11815,N_10458,N_10365);
or U11816 (N_11816,N_10627,N_10951);
and U11817 (N_11817,N_10392,N_10962);
nand U11818 (N_11818,N_10576,N_10222);
nand U11819 (N_11819,N_10612,N_10522);
nand U11820 (N_11820,N_10695,N_10230);
xnor U11821 (N_11821,N_10142,N_10442);
nor U11822 (N_11822,N_10668,N_10762);
or U11823 (N_11823,N_10575,N_10134);
and U11824 (N_11824,N_10595,N_10602);
and U11825 (N_11825,N_10702,N_10626);
xor U11826 (N_11826,N_10074,N_10772);
or U11827 (N_11827,N_10996,N_10098);
and U11828 (N_11828,N_10427,N_10106);
nand U11829 (N_11829,N_10133,N_10962);
or U11830 (N_11830,N_10909,N_10287);
nor U11831 (N_11831,N_10890,N_10639);
nand U11832 (N_11832,N_10353,N_10964);
and U11833 (N_11833,N_10815,N_10250);
or U11834 (N_11834,N_10753,N_10030);
xnor U11835 (N_11835,N_10842,N_10991);
and U11836 (N_11836,N_10871,N_10421);
xnor U11837 (N_11837,N_10254,N_10873);
or U11838 (N_11838,N_10929,N_10227);
or U11839 (N_11839,N_10445,N_10742);
nand U11840 (N_11840,N_10391,N_10198);
xnor U11841 (N_11841,N_10666,N_10777);
nand U11842 (N_11842,N_10858,N_10537);
or U11843 (N_11843,N_10351,N_10903);
and U11844 (N_11844,N_10060,N_10643);
and U11845 (N_11845,N_10246,N_10736);
nand U11846 (N_11846,N_10130,N_10439);
nor U11847 (N_11847,N_10994,N_10748);
nor U11848 (N_11848,N_10353,N_10961);
and U11849 (N_11849,N_10236,N_10583);
xnor U11850 (N_11850,N_10148,N_10551);
nor U11851 (N_11851,N_10372,N_10563);
or U11852 (N_11852,N_10617,N_10877);
nand U11853 (N_11853,N_10729,N_10912);
or U11854 (N_11854,N_10360,N_10855);
or U11855 (N_11855,N_10049,N_10860);
nor U11856 (N_11856,N_10322,N_10668);
nand U11857 (N_11857,N_10455,N_10166);
xor U11858 (N_11858,N_10259,N_10873);
nor U11859 (N_11859,N_10916,N_10693);
or U11860 (N_11860,N_10547,N_10545);
or U11861 (N_11861,N_10293,N_10671);
nor U11862 (N_11862,N_10174,N_10726);
nor U11863 (N_11863,N_10999,N_10756);
or U11864 (N_11864,N_10626,N_10144);
or U11865 (N_11865,N_10010,N_10769);
nor U11866 (N_11866,N_10912,N_10433);
nor U11867 (N_11867,N_10686,N_10554);
and U11868 (N_11868,N_10149,N_10854);
xnor U11869 (N_11869,N_10534,N_10592);
and U11870 (N_11870,N_10782,N_10693);
nor U11871 (N_11871,N_10270,N_10215);
xnor U11872 (N_11872,N_10214,N_10167);
nand U11873 (N_11873,N_10587,N_10325);
or U11874 (N_11874,N_10350,N_10637);
nand U11875 (N_11875,N_10658,N_10554);
and U11876 (N_11876,N_10034,N_10466);
nor U11877 (N_11877,N_10353,N_10180);
and U11878 (N_11878,N_10443,N_10040);
nor U11879 (N_11879,N_10905,N_10041);
or U11880 (N_11880,N_10068,N_10752);
xnor U11881 (N_11881,N_10079,N_10534);
nand U11882 (N_11882,N_10794,N_10501);
xnor U11883 (N_11883,N_10747,N_10482);
nor U11884 (N_11884,N_10017,N_10936);
nand U11885 (N_11885,N_10973,N_10582);
xnor U11886 (N_11886,N_10311,N_10996);
or U11887 (N_11887,N_10107,N_10722);
nor U11888 (N_11888,N_10707,N_10518);
xor U11889 (N_11889,N_10327,N_10288);
nor U11890 (N_11890,N_10127,N_10133);
and U11891 (N_11891,N_10778,N_10052);
nand U11892 (N_11892,N_10829,N_10568);
or U11893 (N_11893,N_10724,N_10099);
xnor U11894 (N_11894,N_10447,N_10381);
xnor U11895 (N_11895,N_10837,N_10075);
nor U11896 (N_11896,N_10487,N_10591);
xnor U11897 (N_11897,N_10508,N_10738);
nor U11898 (N_11898,N_10604,N_10483);
and U11899 (N_11899,N_10921,N_10116);
xor U11900 (N_11900,N_10097,N_10866);
and U11901 (N_11901,N_10404,N_10200);
nor U11902 (N_11902,N_10365,N_10922);
and U11903 (N_11903,N_10612,N_10891);
and U11904 (N_11904,N_10292,N_10203);
xor U11905 (N_11905,N_10003,N_10198);
xor U11906 (N_11906,N_10799,N_10360);
nor U11907 (N_11907,N_10714,N_10481);
and U11908 (N_11908,N_10851,N_10203);
nor U11909 (N_11909,N_10653,N_10129);
and U11910 (N_11910,N_10696,N_10956);
xor U11911 (N_11911,N_10538,N_10778);
nor U11912 (N_11912,N_10678,N_10256);
xor U11913 (N_11913,N_10783,N_10607);
xor U11914 (N_11914,N_10506,N_10179);
nand U11915 (N_11915,N_10506,N_10170);
nor U11916 (N_11916,N_10478,N_10843);
or U11917 (N_11917,N_10059,N_10440);
and U11918 (N_11918,N_10888,N_10353);
and U11919 (N_11919,N_10682,N_10015);
nand U11920 (N_11920,N_10821,N_10268);
or U11921 (N_11921,N_10386,N_10152);
and U11922 (N_11922,N_10032,N_10007);
or U11923 (N_11923,N_10949,N_10901);
or U11924 (N_11924,N_10763,N_10907);
nand U11925 (N_11925,N_10318,N_10443);
and U11926 (N_11926,N_10389,N_10981);
xor U11927 (N_11927,N_10971,N_10092);
xor U11928 (N_11928,N_10065,N_10118);
and U11929 (N_11929,N_10866,N_10775);
nor U11930 (N_11930,N_10951,N_10408);
or U11931 (N_11931,N_10349,N_10182);
or U11932 (N_11932,N_10142,N_10761);
xor U11933 (N_11933,N_10917,N_10920);
or U11934 (N_11934,N_10614,N_10483);
xnor U11935 (N_11935,N_10141,N_10915);
nor U11936 (N_11936,N_10717,N_10952);
nor U11937 (N_11937,N_10470,N_10237);
and U11938 (N_11938,N_10460,N_10496);
or U11939 (N_11939,N_10561,N_10444);
or U11940 (N_11940,N_10871,N_10930);
and U11941 (N_11941,N_10361,N_10666);
xnor U11942 (N_11942,N_10284,N_10941);
xor U11943 (N_11943,N_10909,N_10538);
xnor U11944 (N_11944,N_10732,N_10187);
or U11945 (N_11945,N_10805,N_10052);
or U11946 (N_11946,N_10745,N_10254);
and U11947 (N_11947,N_10987,N_10438);
or U11948 (N_11948,N_10581,N_10071);
and U11949 (N_11949,N_10031,N_10977);
xnor U11950 (N_11950,N_10284,N_10321);
or U11951 (N_11951,N_10679,N_10599);
or U11952 (N_11952,N_10656,N_10231);
and U11953 (N_11953,N_10520,N_10502);
nor U11954 (N_11954,N_10445,N_10613);
nand U11955 (N_11955,N_10236,N_10598);
nand U11956 (N_11956,N_10681,N_10864);
nor U11957 (N_11957,N_10343,N_10780);
xor U11958 (N_11958,N_10403,N_10953);
nor U11959 (N_11959,N_10406,N_10293);
and U11960 (N_11960,N_10137,N_10044);
or U11961 (N_11961,N_10215,N_10494);
or U11962 (N_11962,N_10941,N_10822);
xnor U11963 (N_11963,N_10884,N_10087);
nand U11964 (N_11964,N_10258,N_10013);
or U11965 (N_11965,N_10691,N_10768);
nand U11966 (N_11966,N_10271,N_10887);
nand U11967 (N_11967,N_10002,N_10146);
nor U11968 (N_11968,N_10090,N_10176);
xor U11969 (N_11969,N_10885,N_10399);
nor U11970 (N_11970,N_10326,N_10129);
nor U11971 (N_11971,N_10396,N_10239);
nand U11972 (N_11972,N_10036,N_10521);
and U11973 (N_11973,N_10638,N_10205);
nor U11974 (N_11974,N_10519,N_10095);
nand U11975 (N_11975,N_10721,N_10382);
nand U11976 (N_11976,N_10627,N_10856);
nor U11977 (N_11977,N_10746,N_10836);
nand U11978 (N_11978,N_10265,N_10596);
or U11979 (N_11979,N_10178,N_10571);
nand U11980 (N_11980,N_10355,N_10040);
or U11981 (N_11981,N_10702,N_10882);
nand U11982 (N_11982,N_10622,N_10819);
nand U11983 (N_11983,N_10876,N_10112);
nor U11984 (N_11984,N_10368,N_10737);
and U11985 (N_11985,N_10332,N_10395);
nor U11986 (N_11986,N_10910,N_10355);
or U11987 (N_11987,N_10751,N_10869);
nor U11988 (N_11988,N_10937,N_10526);
or U11989 (N_11989,N_10043,N_10051);
or U11990 (N_11990,N_10447,N_10069);
nor U11991 (N_11991,N_10031,N_10964);
xor U11992 (N_11992,N_10818,N_10351);
nand U11993 (N_11993,N_10349,N_10538);
or U11994 (N_11994,N_10407,N_10461);
nor U11995 (N_11995,N_10226,N_10562);
and U11996 (N_11996,N_10957,N_10695);
or U11997 (N_11997,N_10055,N_10322);
or U11998 (N_11998,N_10388,N_10381);
xor U11999 (N_11999,N_10509,N_10184);
nand U12000 (N_12000,N_11581,N_11559);
xor U12001 (N_12001,N_11982,N_11359);
nor U12002 (N_12002,N_11826,N_11278);
xor U12003 (N_12003,N_11180,N_11532);
nor U12004 (N_12004,N_11763,N_11160);
and U12005 (N_12005,N_11034,N_11661);
xnor U12006 (N_12006,N_11777,N_11530);
and U12007 (N_12007,N_11063,N_11209);
xnor U12008 (N_12008,N_11322,N_11634);
xnor U12009 (N_12009,N_11702,N_11939);
nand U12010 (N_12010,N_11593,N_11156);
nor U12011 (N_12011,N_11103,N_11269);
or U12012 (N_12012,N_11750,N_11219);
and U12013 (N_12013,N_11338,N_11473);
xor U12014 (N_12014,N_11493,N_11766);
nand U12015 (N_12015,N_11543,N_11005);
nand U12016 (N_12016,N_11980,N_11778);
nor U12017 (N_12017,N_11587,N_11635);
nand U12018 (N_12018,N_11310,N_11296);
and U12019 (N_12019,N_11628,N_11946);
nand U12020 (N_12020,N_11110,N_11508);
xnor U12021 (N_12021,N_11050,N_11298);
nand U12022 (N_12022,N_11347,N_11011);
xor U12023 (N_12023,N_11645,N_11061);
nand U12024 (N_12024,N_11455,N_11267);
and U12025 (N_12025,N_11868,N_11080);
xor U12026 (N_12026,N_11496,N_11447);
nand U12027 (N_12027,N_11453,N_11921);
nor U12028 (N_12028,N_11669,N_11290);
xor U12029 (N_12029,N_11124,N_11520);
or U12030 (N_12030,N_11206,N_11190);
or U12031 (N_12031,N_11188,N_11606);
nor U12032 (N_12032,N_11069,N_11875);
nor U12033 (N_12033,N_11402,N_11734);
nand U12034 (N_12034,N_11392,N_11500);
and U12035 (N_12035,N_11933,N_11154);
and U12036 (N_12036,N_11991,N_11886);
or U12037 (N_12037,N_11884,N_11627);
and U12038 (N_12038,N_11118,N_11531);
xnor U12039 (N_12039,N_11812,N_11772);
nor U12040 (N_12040,N_11566,N_11243);
and U12041 (N_12041,N_11689,N_11273);
xor U12042 (N_12042,N_11687,N_11230);
xor U12043 (N_12043,N_11987,N_11995);
xnor U12044 (N_12044,N_11705,N_11315);
and U12045 (N_12045,N_11744,N_11348);
nand U12046 (N_12046,N_11856,N_11096);
or U12047 (N_12047,N_11014,N_11994);
nor U12048 (N_12048,N_11091,N_11458);
or U12049 (N_12049,N_11607,N_11226);
or U12050 (N_12050,N_11914,N_11984);
xnor U12051 (N_12051,N_11907,N_11625);
or U12052 (N_12052,N_11108,N_11346);
or U12053 (N_12053,N_11730,N_11603);
xnor U12054 (N_12054,N_11125,N_11311);
or U12055 (N_12055,N_11442,N_11563);
and U12056 (N_12056,N_11053,N_11105);
or U12057 (N_12057,N_11275,N_11268);
or U12058 (N_12058,N_11706,N_11174);
and U12059 (N_12059,N_11748,N_11102);
or U12060 (N_12060,N_11800,N_11715);
or U12061 (N_12061,N_11840,N_11522);
or U12062 (N_12062,N_11421,N_11942);
or U12063 (N_12063,N_11406,N_11420);
nand U12064 (N_12064,N_11758,N_11138);
xor U12065 (N_12065,N_11584,N_11039);
or U12066 (N_12066,N_11414,N_11131);
nand U12067 (N_12067,N_11617,N_11207);
and U12068 (N_12068,N_11895,N_11221);
and U12069 (N_12069,N_11242,N_11943);
nand U12070 (N_12070,N_11880,N_11787);
nor U12071 (N_12071,N_11743,N_11650);
xor U12072 (N_12072,N_11478,N_11900);
xnor U12073 (N_12073,N_11764,N_11197);
nand U12074 (N_12074,N_11577,N_11250);
xor U12075 (N_12075,N_11858,N_11874);
or U12076 (N_12076,N_11057,N_11934);
and U12077 (N_12077,N_11133,N_11860);
or U12078 (N_12078,N_11229,N_11854);
xor U12079 (N_12079,N_11780,N_11461);
and U12080 (N_12080,N_11595,N_11353);
nand U12081 (N_12081,N_11232,N_11010);
xnor U12082 (N_12082,N_11888,N_11396);
or U12083 (N_12083,N_11788,N_11967);
and U12084 (N_12084,N_11572,N_11477);
and U12085 (N_12085,N_11379,N_11345);
nand U12086 (N_12086,N_11537,N_11383);
and U12087 (N_12087,N_11799,N_11123);
and U12088 (N_12088,N_11996,N_11470);
nor U12089 (N_12089,N_11968,N_11594);
and U12090 (N_12090,N_11699,N_11899);
and U12091 (N_12091,N_11240,N_11279);
nand U12092 (N_12092,N_11046,N_11893);
and U12093 (N_12093,N_11802,N_11241);
and U12094 (N_12094,N_11926,N_11360);
nor U12095 (N_12095,N_11312,N_11507);
or U12096 (N_12096,N_11717,N_11641);
xor U12097 (N_12097,N_11244,N_11239);
and U12098 (N_12098,N_11382,N_11032);
nand U12099 (N_12099,N_11388,N_11159);
and U12100 (N_12100,N_11525,N_11284);
xor U12101 (N_12101,N_11342,N_11412);
or U12102 (N_12102,N_11803,N_11300);
and U12103 (N_12103,N_11936,N_11785);
and U12104 (N_12104,N_11601,N_11055);
or U12105 (N_12105,N_11375,N_11998);
nor U12106 (N_12106,N_11134,N_11839);
xnor U12107 (N_12107,N_11847,N_11505);
or U12108 (N_12108,N_11077,N_11618);
nor U12109 (N_12109,N_11686,N_11115);
nand U12110 (N_12110,N_11947,N_11695);
or U12111 (N_12111,N_11527,N_11341);
and U12112 (N_12112,N_11700,N_11970);
and U12113 (N_12113,N_11747,N_11426);
nor U12114 (N_12114,N_11724,N_11539);
nor U12115 (N_12115,N_11517,N_11042);
nor U12116 (N_12116,N_11691,N_11490);
and U12117 (N_12117,N_11815,N_11562);
nand U12118 (N_12118,N_11088,N_11983);
xnor U12119 (N_12119,N_11664,N_11407);
or U12120 (N_12120,N_11541,N_11609);
nor U12121 (N_12121,N_11830,N_11574);
xnor U12122 (N_12122,N_11150,N_11701);
nand U12123 (N_12123,N_11148,N_11481);
nand U12124 (N_12124,N_11621,N_11885);
or U12125 (N_12125,N_11806,N_11979);
or U12126 (N_12126,N_11155,N_11684);
nand U12127 (N_12127,N_11390,N_11344);
or U12128 (N_12128,N_11896,N_11521);
nand U12129 (N_12129,N_11114,N_11018);
nand U12130 (N_12130,N_11578,N_11674);
nor U12131 (N_12131,N_11660,N_11203);
and U12132 (N_12132,N_11638,N_11678);
and U12133 (N_12133,N_11633,N_11923);
and U12134 (N_12134,N_11350,N_11090);
nor U12135 (N_12135,N_11357,N_11876);
or U12136 (N_12136,N_11327,N_11252);
or U12137 (N_12137,N_11164,N_11266);
nand U12138 (N_12138,N_11172,N_11765);
xor U12139 (N_12139,N_11690,N_11857);
and U12140 (N_12140,N_11280,N_11928);
xor U12141 (N_12141,N_11040,N_11189);
and U12142 (N_12142,N_11126,N_11746);
or U12143 (N_12143,N_11408,N_11973);
or U12144 (N_12144,N_11043,N_11718);
and U12145 (N_12145,N_11460,N_11963);
nor U12146 (N_12146,N_11065,N_11445);
nor U12147 (N_12147,N_11277,N_11903);
and U12148 (N_12148,N_11852,N_11865);
and U12149 (N_12149,N_11703,N_11072);
or U12150 (N_12150,N_11540,N_11450);
and U12151 (N_12151,N_11654,N_11051);
nor U12152 (N_12152,N_11986,N_11683);
nand U12153 (N_12153,N_11146,N_11086);
or U12154 (N_12154,N_11413,N_11073);
nand U12155 (N_12155,N_11644,N_11104);
or U12156 (N_12156,N_11319,N_11902);
nor U12157 (N_12157,N_11049,N_11978);
nand U12158 (N_12158,N_11200,N_11380);
xnor U12159 (N_12159,N_11120,N_11567);
and U12160 (N_12160,N_11851,N_11931);
nand U12161 (N_12161,N_11579,N_11231);
or U12162 (N_12162,N_11526,N_11637);
xor U12163 (N_12163,N_11246,N_11948);
or U12164 (N_12164,N_11165,N_11871);
and U12165 (N_12165,N_11391,N_11711);
and U12166 (N_12166,N_11951,N_11590);
nand U12167 (N_12167,N_11261,N_11598);
and U12168 (N_12168,N_11916,N_11837);
nand U12169 (N_12169,N_11211,N_11938);
xor U12170 (N_12170,N_11247,N_11504);
xor U12171 (N_12171,N_11013,N_11666);
xnor U12172 (N_12172,N_11332,N_11845);
or U12173 (N_12173,N_11652,N_11836);
nor U12174 (N_12174,N_11047,N_11728);
nand U12175 (N_12175,N_11889,N_11707);
or U12176 (N_12176,N_11622,N_11992);
and U12177 (N_12177,N_11575,N_11769);
xnor U12178 (N_12178,N_11472,N_11565);
nand U12179 (N_12179,N_11591,N_11135);
or U12180 (N_12180,N_11642,N_11542);
nand U12181 (N_12181,N_11514,N_11873);
or U12182 (N_12182,N_11217,N_11173);
nand U12183 (N_12183,N_11283,N_11007);
nor U12184 (N_12184,N_11499,N_11999);
nand U12185 (N_12185,N_11761,N_11615);
or U12186 (N_12186,N_11552,N_11810);
nor U12187 (N_12187,N_11553,N_11685);
nand U12188 (N_12188,N_11651,N_11941);
nand U12189 (N_12189,N_11774,N_11805);
nand U12190 (N_12190,N_11592,N_11869);
nor U12191 (N_12191,N_11523,N_11440);
and U12192 (N_12192,N_11356,N_11670);
nor U12193 (N_12193,N_11658,N_11820);
or U12194 (N_12194,N_11849,N_11457);
or U12195 (N_12195,N_11509,N_11632);
xnor U12196 (N_12196,N_11227,N_11887);
or U12197 (N_12197,N_11629,N_11516);
and U12198 (N_12198,N_11254,N_11988);
nor U12199 (N_12199,N_11913,N_11479);
nor U12200 (N_12200,N_11966,N_11038);
nor U12201 (N_12201,N_11100,N_11835);
and U12202 (N_12202,N_11194,N_11956);
or U12203 (N_12203,N_11130,N_11149);
and U12204 (N_12204,N_11688,N_11178);
or U12205 (N_12205,N_11435,N_11117);
nor U12206 (N_12206,N_11404,N_11367);
or U12207 (N_12207,N_11289,N_11804);
nand U12208 (N_12208,N_11872,N_11850);
nor U12209 (N_12209,N_11693,N_11544);
and U12210 (N_12210,N_11604,N_11258);
and U12211 (N_12211,N_11399,N_11897);
xor U12212 (N_12212,N_11841,N_11220);
nor U12213 (N_12213,N_11909,N_11430);
xnor U12214 (N_12214,N_11397,N_11078);
nand U12215 (N_12215,N_11955,N_11535);
nor U12216 (N_12216,N_11433,N_11709);
nor U12217 (N_12217,N_11816,N_11656);
or U12218 (N_12218,N_11827,N_11486);
nor U12219 (N_12219,N_11422,N_11557);
xor U12220 (N_12220,N_11681,N_11832);
xnor U12221 (N_12221,N_11225,N_11952);
or U12222 (N_12222,N_11253,N_11972);
and U12223 (N_12223,N_11713,N_11671);
nor U12224 (N_12224,N_11151,N_11639);
nor U12225 (N_12225,N_11503,N_11613);
and U12226 (N_12226,N_11299,N_11119);
xnor U12227 (N_12227,N_11331,N_11580);
or U12228 (N_12228,N_11771,N_11270);
nor U12229 (N_12229,N_11121,N_11364);
xor U12230 (N_12230,N_11704,N_11494);
nor U12231 (N_12231,N_11001,N_11663);
and U12232 (N_12232,N_11838,N_11546);
or U12233 (N_12233,N_11533,N_11791);
nor U12234 (N_12234,N_11265,N_11294);
and U12235 (N_12235,N_11009,N_11198);
nand U12236 (N_12236,N_11245,N_11263);
nand U12237 (N_12237,N_11989,N_11030);
and U12238 (N_12238,N_11843,N_11890);
xnor U12239 (N_12239,N_11662,N_11175);
nand U12240 (N_12240,N_11462,N_11679);
or U12241 (N_12241,N_11302,N_11395);
and U12242 (N_12242,N_11997,N_11292);
or U12243 (N_12243,N_11186,N_11630);
or U12244 (N_12244,N_11818,N_11547);
nand U12245 (N_12245,N_11511,N_11793);
nor U12246 (N_12246,N_11716,N_11111);
and U12247 (N_12247,N_11976,N_11466);
nand U12248 (N_12248,N_11081,N_11855);
xnor U12249 (N_12249,N_11449,N_11436);
nor U12250 (N_12250,N_11068,N_11285);
and U12251 (N_12251,N_11035,N_11834);
or U12252 (N_12252,N_11811,N_11441);
and U12253 (N_12253,N_11616,N_11667);
and U12254 (N_12254,N_11853,N_11288);
xnor U12255 (N_12255,N_11021,N_11176);
and U12256 (N_12256,N_11372,N_11352);
or U12257 (N_12257,N_11714,N_11048);
and U12258 (N_12258,N_11095,N_11583);
or U12259 (N_12259,N_11904,N_11410);
nand U12260 (N_12260,N_11318,N_11153);
nand U12261 (N_12261,N_11293,N_11554);
or U12262 (N_12262,N_11415,N_11191);
or U12263 (N_12263,N_11325,N_11306);
nand U12264 (N_12264,N_11323,N_11949);
nor U12265 (N_12265,N_11624,N_11798);
or U12266 (N_12266,N_11783,N_11958);
nand U12267 (N_12267,N_11981,N_11476);
or U12268 (N_12268,N_11251,N_11668);
xor U12269 (N_12269,N_11141,N_11614);
xor U12270 (N_12270,N_11281,N_11427);
nor U12271 (N_12271,N_11147,N_11321);
xnor U12272 (N_12272,N_11745,N_11673);
nor U12273 (N_12273,N_11394,N_11093);
and U12274 (N_12274,N_11193,N_11037);
xnor U12275 (N_12275,N_11927,N_11376);
nand U12276 (N_12276,N_11894,N_11074);
nor U12277 (N_12277,N_11158,N_11431);
xnor U12278 (N_12278,N_11287,N_11937);
nand U12279 (N_12279,N_11045,N_11424);
nand U12280 (N_12280,N_11400,N_11256);
and U12281 (N_12281,N_11255,N_11085);
nand U12282 (N_12282,N_11107,N_11401);
and U12283 (N_12283,N_11861,N_11501);
nand U12284 (N_12284,N_11612,N_11682);
nor U12285 (N_12285,N_11218,N_11932);
nor U12286 (N_12286,N_11731,N_11792);
nand U12287 (N_12287,N_11089,N_11732);
and U12288 (N_12288,N_11863,N_11215);
xor U12289 (N_12289,N_11564,N_11127);
or U12290 (N_12290,N_11064,N_11677);
or U12291 (N_12291,N_11463,N_11112);
xor U12292 (N_12292,N_11161,N_11944);
or U12293 (N_12293,N_11586,N_11099);
or U12294 (N_12294,N_11597,N_11528);
nand U12295 (N_12295,N_11512,N_11170);
nor U12296 (N_12296,N_11060,N_11719);
and U12297 (N_12297,N_11444,N_11735);
xor U12298 (N_12298,N_11398,N_11729);
and U12299 (N_12299,N_11454,N_11483);
nor U12300 (N_12300,N_11482,N_11672);
nand U12301 (N_12301,N_11762,N_11432);
nor U12302 (N_12302,N_11727,N_11092);
nand U12303 (N_12303,N_11751,N_11741);
nor U12304 (N_12304,N_11495,N_11881);
xnor U12305 (N_12305,N_11301,N_11545);
nor U12306 (N_12306,N_11201,N_11740);
or U12307 (N_12307,N_11066,N_11680);
or U12308 (N_12308,N_11710,N_11692);
or U12309 (N_12309,N_11469,N_11877);
nor U12310 (N_12310,N_11824,N_11752);
nand U12311 (N_12311,N_11862,N_11825);
and U12312 (N_12312,N_11600,N_11882);
nand U12313 (N_12313,N_11665,N_11317);
or U12314 (N_12314,N_11184,N_11846);
nor U12315 (N_12315,N_11801,N_11142);
nor U12316 (N_12316,N_11384,N_11451);
or U12317 (N_12317,N_11343,N_11106);
xnor U12318 (N_12318,N_11696,N_11821);
xor U12319 (N_12319,N_11419,N_11468);
xnor U12320 (N_12320,N_11721,N_11599);
and U12321 (N_12321,N_11646,N_11456);
and U12322 (N_12322,N_11171,N_11029);
and U12323 (N_12323,N_11233,N_11202);
and U12324 (N_12324,N_11286,N_11183);
xor U12325 (N_12325,N_11738,N_11498);
and U12326 (N_12326,N_11262,N_11291);
nor U12327 (N_12327,N_11974,N_11097);
and U12328 (N_12328,N_11326,N_11339);
xnor U12329 (N_12329,N_11789,N_11140);
nor U12330 (N_12330,N_11879,N_11524);
or U12331 (N_12331,N_11238,N_11878);
or U12332 (N_12332,N_11082,N_11259);
nand U12333 (N_12333,N_11708,N_11538);
nand U12334 (N_12334,N_11519,N_11272);
and U12335 (N_12335,N_11844,N_11019);
nor U12336 (N_12336,N_11712,N_11316);
nor U12337 (N_12337,N_11675,N_11823);
and U12338 (N_12338,N_11136,N_11403);
nor U12339 (N_12339,N_11075,N_11487);
nor U12340 (N_12340,N_11276,N_11726);
nor U12341 (N_12341,N_11378,N_11320);
nor U12342 (N_12342,N_11919,N_11859);
or U12343 (N_12343,N_11373,N_11328);
and U12344 (N_12344,N_11767,N_11964);
xor U12345 (N_12345,N_11725,N_11362);
xnor U12346 (N_12346,N_11083,N_11475);
xnor U12347 (N_12347,N_11797,N_11977);
and U12348 (N_12348,N_11129,N_11168);
xnor U12349 (N_12349,N_11502,N_11182);
and U12350 (N_12350,N_11417,N_11814);
or U12351 (N_12351,N_11636,N_11015);
xnor U12352 (N_12352,N_11739,N_11790);
or U12353 (N_12353,N_11784,N_11969);
nor U12354 (N_12354,N_11733,N_11585);
or U12355 (N_12355,N_11393,N_11961);
nand U12356 (N_12356,N_11016,N_11355);
xnor U12357 (N_12357,N_11782,N_11779);
nor U12358 (N_12358,N_11409,N_11358);
nor U12359 (N_12359,N_11349,N_11303);
nor U12360 (N_12360,N_11084,N_11169);
xnor U12361 (N_12361,N_11550,N_11602);
and U12362 (N_12362,N_11781,N_11167);
nand U12363 (N_12363,N_11137,N_11489);
nand U12364 (N_12364,N_11930,N_11822);
and U12365 (N_12365,N_11901,N_11199);
nand U12366 (N_12366,N_11467,N_11759);
nand U12367 (N_12367,N_11381,N_11305);
and U12368 (N_12368,N_11560,N_11145);
nor U12369 (N_12369,N_11027,N_11054);
or U12370 (N_12370,N_11883,N_11000);
and U12371 (N_12371,N_11236,N_11918);
nor U12372 (N_12372,N_11813,N_11143);
or U12373 (N_12373,N_11480,N_11534);
or U12374 (N_12374,N_11891,N_11611);
nor U12375 (N_12375,N_11518,N_11549);
nand U12376 (N_12376,N_11443,N_11492);
nand U12377 (N_12377,N_11570,N_11370);
and U12378 (N_12378,N_11058,N_11589);
or U12379 (N_12379,N_11561,N_11079);
or U12380 (N_12380,N_11012,N_11573);
and U12381 (N_12381,N_11271,N_11337);
nand U12382 (N_12382,N_11794,N_11529);
nor U12383 (N_12383,N_11697,N_11274);
and U12384 (N_12384,N_11329,N_11488);
nand U12385 (N_12385,N_11006,N_11760);
or U12386 (N_12386,N_11959,N_11649);
nand U12387 (N_12387,N_11309,N_11389);
and U12388 (N_12388,N_11101,N_11336);
xor U12389 (N_12389,N_11333,N_11647);
xnor U12390 (N_12390,N_11556,N_11925);
nor U12391 (N_12391,N_11179,N_11062);
nor U12392 (N_12392,N_11551,N_11228);
nor U12393 (N_12393,N_11620,N_11437);
or U12394 (N_12394,N_11770,N_11922);
and U12395 (N_12395,N_11950,N_11605);
or U12396 (N_12396,N_11210,N_11304);
nand U12397 (N_12397,N_11898,N_11915);
and U12398 (N_12398,N_11631,N_11911);
nor U12399 (N_12399,N_11354,N_11571);
nand U12400 (N_12400,N_11087,N_11536);
xor U12401 (N_12401,N_11828,N_11335);
nor U12402 (N_12402,N_11643,N_11222);
and U12403 (N_12403,N_11387,N_11216);
nand U12404 (N_12404,N_11212,N_11736);
xor U12405 (N_12405,N_11474,N_11204);
or U12406 (N_12406,N_11829,N_11870);
and U12407 (N_12407,N_11558,N_11753);
nor U12408 (N_12408,N_11205,N_11807);
or U12409 (N_12409,N_11513,N_11003);
and U12410 (N_12410,N_11548,N_11340);
nand U12411 (N_12411,N_11448,N_11369);
and U12412 (N_12412,N_11723,N_11425);
or U12413 (N_12413,N_11640,N_11192);
nand U12414 (N_12414,N_11768,N_11749);
nor U12415 (N_12415,N_11195,N_11036);
or U12416 (N_12416,N_11386,N_11659);
nand U12417 (N_12417,N_11313,N_11737);
nand U12418 (N_12418,N_11076,N_11908);
xor U12419 (N_12419,N_11910,N_11608);
or U12420 (N_12420,N_11248,N_11059);
xnor U12421 (N_12421,N_11177,N_11510);
and U12422 (N_12422,N_11439,N_11428);
nor U12423 (N_12423,N_11960,N_11459);
nand U12424 (N_12424,N_11945,N_11754);
xnor U12425 (N_12425,N_11831,N_11795);
nor U12426 (N_12426,N_11993,N_11985);
or U12427 (N_12427,N_11257,N_11166);
and U12428 (N_12428,N_11022,N_11623);
and U12429 (N_12429,N_11905,N_11940);
nand U12430 (N_12430,N_11906,N_11004);
xor U12431 (N_12431,N_11416,N_11314);
and U12432 (N_12432,N_11775,N_11497);
nand U12433 (N_12433,N_11582,N_11892);
nand U12434 (N_12434,N_11866,N_11363);
xnor U12435 (N_12435,N_11223,N_11917);
or U12436 (N_12436,N_11366,N_11626);
and U12437 (N_12437,N_11653,N_11965);
nand U12438 (N_12438,N_11957,N_11438);
or U12439 (N_12439,N_11864,N_11308);
nand U12440 (N_12440,N_11098,N_11377);
and U12441 (N_12441,N_11755,N_11423);
nor U12442 (N_12442,N_11776,N_11307);
and U12443 (N_12443,N_11260,N_11935);
xnor U12444 (N_12444,N_11044,N_11786);
and U12445 (N_12445,N_11405,N_11070);
nand U12446 (N_12446,N_11020,N_11187);
nand U12447 (N_12447,N_11374,N_11596);
and U12448 (N_12448,N_11295,N_11282);
nor U12449 (N_12449,N_11452,N_11722);
nand U12450 (N_12450,N_11773,N_11757);
nor U12451 (N_12451,N_11742,N_11411);
and U12452 (N_12452,N_11555,N_11576);
nor U12453 (N_12453,N_11485,N_11234);
and U12454 (N_12454,N_11471,N_11181);
nor U12455 (N_12455,N_11196,N_11023);
nor U12456 (N_12456,N_11610,N_11334);
nor U12457 (N_12457,N_11031,N_11157);
nand U12458 (N_12458,N_11676,N_11214);
nor U12459 (N_12459,N_11954,N_11867);
or U12460 (N_12460,N_11657,N_11208);
xnor U12461 (N_12461,N_11144,N_11185);
nand U12462 (N_12462,N_11975,N_11213);
nor U12463 (N_12463,N_11953,N_11506);
or U12464 (N_12464,N_11152,N_11264);
nand U12465 (N_12465,N_11052,N_11162);
xor U12466 (N_12466,N_11515,N_11026);
xnor U12467 (N_12467,N_11163,N_11324);
xor U12468 (N_12468,N_11809,N_11971);
or U12469 (N_12469,N_11429,N_11446);
and U12470 (N_12470,N_11028,N_11132);
xnor U12471 (N_12471,N_11464,N_11017);
nand U12472 (N_12472,N_11122,N_11235);
xor U12473 (N_12473,N_11833,N_11385);
and U12474 (N_12474,N_11371,N_11920);
nor U12475 (N_12475,N_11588,N_11249);
nand U12476 (N_12476,N_11924,N_11067);
nor U12477 (N_12477,N_11698,N_11116);
xor U12478 (N_12478,N_11024,N_11361);
nand U12479 (N_12479,N_11655,N_11796);
nor U12480 (N_12480,N_11962,N_11368);
nor U12481 (N_12481,N_11297,N_11694);
xnor U12482 (N_12482,N_11929,N_11139);
and U12483 (N_12483,N_11756,N_11434);
or U12484 (N_12484,N_11109,N_11365);
xor U12485 (N_12485,N_11819,N_11990);
and U12486 (N_12486,N_11720,N_11071);
or U12487 (N_12487,N_11568,N_11237);
xor U12488 (N_12488,N_11330,N_11484);
xnor U12489 (N_12489,N_11808,N_11817);
nand U12490 (N_12490,N_11842,N_11224);
xnor U12491 (N_12491,N_11056,N_11491);
xor U12492 (N_12492,N_11418,N_11113);
and U12493 (N_12493,N_11025,N_11569);
nor U12494 (N_12494,N_11094,N_11033);
and U12495 (N_12495,N_11002,N_11848);
nor U12496 (N_12496,N_11619,N_11648);
or U12497 (N_12497,N_11128,N_11041);
xor U12498 (N_12498,N_11465,N_11008);
xnor U12499 (N_12499,N_11912,N_11351);
nand U12500 (N_12500,N_11986,N_11406);
and U12501 (N_12501,N_11350,N_11492);
or U12502 (N_12502,N_11620,N_11557);
and U12503 (N_12503,N_11817,N_11725);
xor U12504 (N_12504,N_11601,N_11392);
xor U12505 (N_12505,N_11418,N_11245);
nand U12506 (N_12506,N_11722,N_11718);
or U12507 (N_12507,N_11454,N_11804);
nor U12508 (N_12508,N_11600,N_11677);
or U12509 (N_12509,N_11839,N_11189);
and U12510 (N_12510,N_11245,N_11810);
or U12511 (N_12511,N_11835,N_11237);
nand U12512 (N_12512,N_11054,N_11116);
xor U12513 (N_12513,N_11719,N_11203);
or U12514 (N_12514,N_11975,N_11073);
nand U12515 (N_12515,N_11236,N_11180);
nand U12516 (N_12516,N_11850,N_11917);
or U12517 (N_12517,N_11059,N_11386);
and U12518 (N_12518,N_11040,N_11279);
and U12519 (N_12519,N_11318,N_11347);
nand U12520 (N_12520,N_11521,N_11090);
nand U12521 (N_12521,N_11156,N_11915);
nand U12522 (N_12522,N_11606,N_11122);
nor U12523 (N_12523,N_11395,N_11806);
nand U12524 (N_12524,N_11951,N_11418);
nor U12525 (N_12525,N_11258,N_11887);
nor U12526 (N_12526,N_11451,N_11469);
or U12527 (N_12527,N_11543,N_11994);
or U12528 (N_12528,N_11357,N_11410);
nor U12529 (N_12529,N_11642,N_11323);
or U12530 (N_12530,N_11817,N_11222);
nor U12531 (N_12531,N_11991,N_11636);
nand U12532 (N_12532,N_11961,N_11891);
or U12533 (N_12533,N_11541,N_11851);
xnor U12534 (N_12534,N_11847,N_11264);
nand U12535 (N_12535,N_11761,N_11728);
and U12536 (N_12536,N_11466,N_11983);
nand U12537 (N_12537,N_11717,N_11813);
xor U12538 (N_12538,N_11995,N_11649);
xor U12539 (N_12539,N_11757,N_11000);
nor U12540 (N_12540,N_11215,N_11053);
and U12541 (N_12541,N_11096,N_11267);
and U12542 (N_12542,N_11677,N_11982);
nand U12543 (N_12543,N_11985,N_11839);
xnor U12544 (N_12544,N_11245,N_11223);
nor U12545 (N_12545,N_11720,N_11164);
nor U12546 (N_12546,N_11753,N_11910);
xnor U12547 (N_12547,N_11651,N_11557);
and U12548 (N_12548,N_11545,N_11599);
or U12549 (N_12549,N_11142,N_11582);
or U12550 (N_12550,N_11003,N_11751);
nand U12551 (N_12551,N_11859,N_11242);
and U12552 (N_12552,N_11070,N_11482);
nand U12553 (N_12553,N_11469,N_11830);
nand U12554 (N_12554,N_11076,N_11674);
nor U12555 (N_12555,N_11411,N_11060);
xor U12556 (N_12556,N_11289,N_11749);
nand U12557 (N_12557,N_11249,N_11438);
or U12558 (N_12558,N_11655,N_11814);
and U12559 (N_12559,N_11796,N_11374);
nor U12560 (N_12560,N_11820,N_11969);
or U12561 (N_12561,N_11528,N_11744);
xor U12562 (N_12562,N_11874,N_11294);
or U12563 (N_12563,N_11120,N_11048);
nand U12564 (N_12564,N_11389,N_11624);
xor U12565 (N_12565,N_11026,N_11205);
nand U12566 (N_12566,N_11194,N_11991);
nor U12567 (N_12567,N_11070,N_11081);
xor U12568 (N_12568,N_11620,N_11308);
nand U12569 (N_12569,N_11447,N_11716);
nand U12570 (N_12570,N_11089,N_11344);
xor U12571 (N_12571,N_11109,N_11413);
nor U12572 (N_12572,N_11437,N_11068);
nand U12573 (N_12573,N_11979,N_11503);
or U12574 (N_12574,N_11897,N_11259);
nor U12575 (N_12575,N_11386,N_11699);
or U12576 (N_12576,N_11463,N_11108);
nand U12577 (N_12577,N_11422,N_11008);
and U12578 (N_12578,N_11199,N_11631);
and U12579 (N_12579,N_11958,N_11982);
xnor U12580 (N_12580,N_11439,N_11729);
xnor U12581 (N_12581,N_11053,N_11913);
or U12582 (N_12582,N_11606,N_11864);
nor U12583 (N_12583,N_11429,N_11461);
nor U12584 (N_12584,N_11995,N_11871);
and U12585 (N_12585,N_11972,N_11413);
xor U12586 (N_12586,N_11963,N_11468);
xor U12587 (N_12587,N_11477,N_11359);
nor U12588 (N_12588,N_11419,N_11151);
nand U12589 (N_12589,N_11100,N_11979);
and U12590 (N_12590,N_11269,N_11000);
nor U12591 (N_12591,N_11029,N_11434);
nor U12592 (N_12592,N_11915,N_11150);
nor U12593 (N_12593,N_11322,N_11746);
nand U12594 (N_12594,N_11274,N_11003);
nor U12595 (N_12595,N_11656,N_11665);
xor U12596 (N_12596,N_11430,N_11470);
xor U12597 (N_12597,N_11366,N_11065);
or U12598 (N_12598,N_11517,N_11616);
nor U12599 (N_12599,N_11487,N_11828);
nor U12600 (N_12600,N_11893,N_11527);
and U12601 (N_12601,N_11718,N_11974);
nor U12602 (N_12602,N_11004,N_11577);
nand U12603 (N_12603,N_11247,N_11506);
and U12604 (N_12604,N_11379,N_11603);
and U12605 (N_12605,N_11685,N_11511);
and U12606 (N_12606,N_11407,N_11258);
nand U12607 (N_12607,N_11245,N_11442);
and U12608 (N_12608,N_11216,N_11019);
nor U12609 (N_12609,N_11386,N_11538);
nand U12610 (N_12610,N_11658,N_11654);
or U12611 (N_12611,N_11987,N_11203);
nor U12612 (N_12612,N_11092,N_11806);
or U12613 (N_12613,N_11947,N_11068);
nand U12614 (N_12614,N_11282,N_11842);
nor U12615 (N_12615,N_11631,N_11514);
xnor U12616 (N_12616,N_11207,N_11901);
and U12617 (N_12617,N_11507,N_11462);
and U12618 (N_12618,N_11554,N_11451);
nand U12619 (N_12619,N_11392,N_11268);
nand U12620 (N_12620,N_11736,N_11002);
nand U12621 (N_12621,N_11699,N_11712);
or U12622 (N_12622,N_11104,N_11276);
nor U12623 (N_12623,N_11901,N_11982);
nor U12624 (N_12624,N_11632,N_11338);
xnor U12625 (N_12625,N_11659,N_11752);
nand U12626 (N_12626,N_11014,N_11083);
or U12627 (N_12627,N_11063,N_11992);
and U12628 (N_12628,N_11330,N_11246);
xnor U12629 (N_12629,N_11821,N_11004);
and U12630 (N_12630,N_11258,N_11418);
xnor U12631 (N_12631,N_11316,N_11212);
nand U12632 (N_12632,N_11216,N_11105);
or U12633 (N_12633,N_11246,N_11488);
and U12634 (N_12634,N_11740,N_11369);
and U12635 (N_12635,N_11778,N_11047);
or U12636 (N_12636,N_11127,N_11951);
or U12637 (N_12637,N_11072,N_11655);
xnor U12638 (N_12638,N_11626,N_11961);
xor U12639 (N_12639,N_11607,N_11471);
or U12640 (N_12640,N_11681,N_11393);
xnor U12641 (N_12641,N_11362,N_11402);
and U12642 (N_12642,N_11332,N_11363);
and U12643 (N_12643,N_11750,N_11811);
nand U12644 (N_12644,N_11795,N_11779);
nor U12645 (N_12645,N_11313,N_11046);
and U12646 (N_12646,N_11345,N_11654);
nor U12647 (N_12647,N_11916,N_11501);
and U12648 (N_12648,N_11273,N_11603);
or U12649 (N_12649,N_11179,N_11504);
or U12650 (N_12650,N_11376,N_11892);
and U12651 (N_12651,N_11764,N_11995);
nor U12652 (N_12652,N_11001,N_11017);
nand U12653 (N_12653,N_11938,N_11344);
or U12654 (N_12654,N_11026,N_11343);
nor U12655 (N_12655,N_11306,N_11977);
and U12656 (N_12656,N_11769,N_11062);
nand U12657 (N_12657,N_11164,N_11187);
nand U12658 (N_12658,N_11434,N_11457);
and U12659 (N_12659,N_11604,N_11404);
nand U12660 (N_12660,N_11505,N_11280);
and U12661 (N_12661,N_11018,N_11981);
or U12662 (N_12662,N_11186,N_11916);
xnor U12663 (N_12663,N_11261,N_11900);
nand U12664 (N_12664,N_11588,N_11308);
nor U12665 (N_12665,N_11116,N_11274);
and U12666 (N_12666,N_11834,N_11566);
xnor U12667 (N_12667,N_11980,N_11287);
and U12668 (N_12668,N_11571,N_11696);
or U12669 (N_12669,N_11401,N_11861);
xor U12670 (N_12670,N_11826,N_11627);
nor U12671 (N_12671,N_11092,N_11118);
and U12672 (N_12672,N_11707,N_11272);
nand U12673 (N_12673,N_11311,N_11728);
xor U12674 (N_12674,N_11754,N_11281);
xor U12675 (N_12675,N_11618,N_11403);
nand U12676 (N_12676,N_11358,N_11698);
xnor U12677 (N_12677,N_11919,N_11340);
xor U12678 (N_12678,N_11145,N_11946);
or U12679 (N_12679,N_11732,N_11233);
nor U12680 (N_12680,N_11869,N_11999);
nor U12681 (N_12681,N_11865,N_11947);
xor U12682 (N_12682,N_11845,N_11932);
nand U12683 (N_12683,N_11035,N_11168);
nand U12684 (N_12684,N_11385,N_11443);
nor U12685 (N_12685,N_11635,N_11631);
or U12686 (N_12686,N_11713,N_11517);
and U12687 (N_12687,N_11350,N_11234);
nand U12688 (N_12688,N_11530,N_11560);
nor U12689 (N_12689,N_11003,N_11488);
xnor U12690 (N_12690,N_11461,N_11068);
or U12691 (N_12691,N_11632,N_11475);
and U12692 (N_12692,N_11621,N_11886);
nor U12693 (N_12693,N_11844,N_11296);
nand U12694 (N_12694,N_11177,N_11986);
or U12695 (N_12695,N_11434,N_11665);
or U12696 (N_12696,N_11222,N_11766);
or U12697 (N_12697,N_11723,N_11872);
or U12698 (N_12698,N_11801,N_11080);
nand U12699 (N_12699,N_11897,N_11286);
nor U12700 (N_12700,N_11019,N_11976);
nor U12701 (N_12701,N_11026,N_11482);
xor U12702 (N_12702,N_11544,N_11926);
and U12703 (N_12703,N_11508,N_11949);
and U12704 (N_12704,N_11171,N_11032);
xor U12705 (N_12705,N_11491,N_11236);
and U12706 (N_12706,N_11299,N_11943);
or U12707 (N_12707,N_11065,N_11670);
nor U12708 (N_12708,N_11900,N_11776);
or U12709 (N_12709,N_11173,N_11228);
nor U12710 (N_12710,N_11980,N_11446);
nand U12711 (N_12711,N_11564,N_11348);
xnor U12712 (N_12712,N_11185,N_11637);
and U12713 (N_12713,N_11706,N_11754);
nand U12714 (N_12714,N_11560,N_11748);
and U12715 (N_12715,N_11515,N_11937);
xor U12716 (N_12716,N_11485,N_11681);
or U12717 (N_12717,N_11620,N_11348);
nand U12718 (N_12718,N_11598,N_11572);
xnor U12719 (N_12719,N_11205,N_11413);
nor U12720 (N_12720,N_11353,N_11615);
xnor U12721 (N_12721,N_11835,N_11297);
and U12722 (N_12722,N_11999,N_11737);
nor U12723 (N_12723,N_11069,N_11634);
nand U12724 (N_12724,N_11809,N_11436);
and U12725 (N_12725,N_11567,N_11434);
and U12726 (N_12726,N_11356,N_11621);
or U12727 (N_12727,N_11653,N_11838);
nand U12728 (N_12728,N_11891,N_11919);
or U12729 (N_12729,N_11901,N_11008);
xor U12730 (N_12730,N_11684,N_11295);
or U12731 (N_12731,N_11828,N_11825);
and U12732 (N_12732,N_11690,N_11373);
or U12733 (N_12733,N_11880,N_11081);
xnor U12734 (N_12734,N_11922,N_11820);
or U12735 (N_12735,N_11163,N_11861);
nor U12736 (N_12736,N_11849,N_11518);
and U12737 (N_12737,N_11760,N_11579);
nand U12738 (N_12738,N_11954,N_11518);
xnor U12739 (N_12739,N_11346,N_11185);
or U12740 (N_12740,N_11485,N_11897);
nor U12741 (N_12741,N_11333,N_11400);
and U12742 (N_12742,N_11774,N_11261);
or U12743 (N_12743,N_11191,N_11419);
nor U12744 (N_12744,N_11840,N_11568);
and U12745 (N_12745,N_11130,N_11259);
or U12746 (N_12746,N_11454,N_11526);
nor U12747 (N_12747,N_11034,N_11674);
and U12748 (N_12748,N_11030,N_11511);
nor U12749 (N_12749,N_11821,N_11150);
xor U12750 (N_12750,N_11700,N_11341);
or U12751 (N_12751,N_11529,N_11423);
nor U12752 (N_12752,N_11649,N_11647);
and U12753 (N_12753,N_11017,N_11978);
and U12754 (N_12754,N_11405,N_11674);
nand U12755 (N_12755,N_11456,N_11252);
nand U12756 (N_12756,N_11133,N_11077);
xor U12757 (N_12757,N_11859,N_11309);
xnor U12758 (N_12758,N_11282,N_11173);
and U12759 (N_12759,N_11891,N_11739);
or U12760 (N_12760,N_11679,N_11233);
nor U12761 (N_12761,N_11724,N_11790);
and U12762 (N_12762,N_11876,N_11309);
nand U12763 (N_12763,N_11805,N_11229);
xnor U12764 (N_12764,N_11313,N_11088);
nand U12765 (N_12765,N_11202,N_11353);
or U12766 (N_12766,N_11657,N_11386);
nand U12767 (N_12767,N_11647,N_11734);
nor U12768 (N_12768,N_11425,N_11075);
xnor U12769 (N_12769,N_11215,N_11658);
and U12770 (N_12770,N_11374,N_11127);
or U12771 (N_12771,N_11622,N_11011);
xor U12772 (N_12772,N_11415,N_11809);
xnor U12773 (N_12773,N_11437,N_11720);
nand U12774 (N_12774,N_11611,N_11922);
or U12775 (N_12775,N_11243,N_11057);
xnor U12776 (N_12776,N_11662,N_11358);
xor U12777 (N_12777,N_11751,N_11336);
xor U12778 (N_12778,N_11276,N_11362);
and U12779 (N_12779,N_11138,N_11892);
nand U12780 (N_12780,N_11154,N_11316);
nand U12781 (N_12781,N_11979,N_11641);
or U12782 (N_12782,N_11127,N_11556);
or U12783 (N_12783,N_11164,N_11907);
and U12784 (N_12784,N_11930,N_11827);
nor U12785 (N_12785,N_11467,N_11548);
or U12786 (N_12786,N_11842,N_11836);
and U12787 (N_12787,N_11654,N_11006);
nor U12788 (N_12788,N_11467,N_11653);
nor U12789 (N_12789,N_11825,N_11351);
nand U12790 (N_12790,N_11887,N_11870);
xor U12791 (N_12791,N_11155,N_11715);
and U12792 (N_12792,N_11014,N_11349);
or U12793 (N_12793,N_11610,N_11908);
or U12794 (N_12794,N_11555,N_11227);
or U12795 (N_12795,N_11719,N_11394);
or U12796 (N_12796,N_11199,N_11275);
and U12797 (N_12797,N_11370,N_11017);
xor U12798 (N_12798,N_11219,N_11849);
or U12799 (N_12799,N_11380,N_11214);
nor U12800 (N_12800,N_11641,N_11420);
xnor U12801 (N_12801,N_11777,N_11423);
nand U12802 (N_12802,N_11141,N_11919);
nand U12803 (N_12803,N_11593,N_11170);
nand U12804 (N_12804,N_11458,N_11258);
or U12805 (N_12805,N_11714,N_11836);
xnor U12806 (N_12806,N_11020,N_11459);
xor U12807 (N_12807,N_11749,N_11852);
and U12808 (N_12808,N_11271,N_11634);
nand U12809 (N_12809,N_11663,N_11734);
nor U12810 (N_12810,N_11863,N_11610);
and U12811 (N_12811,N_11193,N_11262);
or U12812 (N_12812,N_11321,N_11511);
and U12813 (N_12813,N_11277,N_11911);
nand U12814 (N_12814,N_11658,N_11127);
or U12815 (N_12815,N_11438,N_11476);
nor U12816 (N_12816,N_11607,N_11543);
and U12817 (N_12817,N_11965,N_11945);
nor U12818 (N_12818,N_11285,N_11377);
nor U12819 (N_12819,N_11512,N_11480);
xor U12820 (N_12820,N_11765,N_11001);
xnor U12821 (N_12821,N_11924,N_11336);
or U12822 (N_12822,N_11966,N_11945);
xor U12823 (N_12823,N_11481,N_11373);
nor U12824 (N_12824,N_11311,N_11165);
xor U12825 (N_12825,N_11999,N_11722);
nand U12826 (N_12826,N_11080,N_11686);
and U12827 (N_12827,N_11618,N_11444);
nor U12828 (N_12828,N_11393,N_11616);
and U12829 (N_12829,N_11209,N_11720);
or U12830 (N_12830,N_11976,N_11534);
or U12831 (N_12831,N_11061,N_11639);
nand U12832 (N_12832,N_11036,N_11700);
xnor U12833 (N_12833,N_11124,N_11470);
xor U12834 (N_12834,N_11035,N_11151);
and U12835 (N_12835,N_11440,N_11928);
or U12836 (N_12836,N_11699,N_11392);
nor U12837 (N_12837,N_11614,N_11070);
nand U12838 (N_12838,N_11978,N_11538);
and U12839 (N_12839,N_11514,N_11781);
xor U12840 (N_12840,N_11728,N_11697);
nor U12841 (N_12841,N_11099,N_11836);
nand U12842 (N_12842,N_11863,N_11786);
and U12843 (N_12843,N_11748,N_11817);
xnor U12844 (N_12844,N_11606,N_11426);
or U12845 (N_12845,N_11485,N_11299);
or U12846 (N_12846,N_11812,N_11185);
or U12847 (N_12847,N_11881,N_11814);
and U12848 (N_12848,N_11181,N_11635);
nand U12849 (N_12849,N_11093,N_11554);
or U12850 (N_12850,N_11348,N_11356);
xor U12851 (N_12851,N_11332,N_11162);
xor U12852 (N_12852,N_11488,N_11769);
nor U12853 (N_12853,N_11998,N_11141);
nand U12854 (N_12854,N_11816,N_11313);
nand U12855 (N_12855,N_11230,N_11465);
xor U12856 (N_12856,N_11182,N_11290);
nand U12857 (N_12857,N_11432,N_11451);
nand U12858 (N_12858,N_11375,N_11108);
nand U12859 (N_12859,N_11295,N_11492);
or U12860 (N_12860,N_11491,N_11956);
or U12861 (N_12861,N_11768,N_11556);
nor U12862 (N_12862,N_11441,N_11255);
nand U12863 (N_12863,N_11949,N_11731);
and U12864 (N_12864,N_11497,N_11072);
nor U12865 (N_12865,N_11149,N_11194);
xnor U12866 (N_12866,N_11124,N_11707);
xor U12867 (N_12867,N_11123,N_11020);
nor U12868 (N_12868,N_11994,N_11056);
xor U12869 (N_12869,N_11310,N_11319);
and U12870 (N_12870,N_11313,N_11864);
xor U12871 (N_12871,N_11259,N_11461);
or U12872 (N_12872,N_11624,N_11622);
or U12873 (N_12873,N_11202,N_11420);
and U12874 (N_12874,N_11155,N_11733);
nor U12875 (N_12875,N_11106,N_11088);
nand U12876 (N_12876,N_11189,N_11095);
nor U12877 (N_12877,N_11460,N_11079);
nand U12878 (N_12878,N_11343,N_11571);
or U12879 (N_12879,N_11852,N_11252);
nor U12880 (N_12880,N_11853,N_11995);
nand U12881 (N_12881,N_11596,N_11538);
xnor U12882 (N_12882,N_11314,N_11939);
nor U12883 (N_12883,N_11862,N_11994);
or U12884 (N_12884,N_11098,N_11147);
nor U12885 (N_12885,N_11113,N_11724);
nand U12886 (N_12886,N_11079,N_11507);
nand U12887 (N_12887,N_11764,N_11842);
nand U12888 (N_12888,N_11435,N_11478);
nand U12889 (N_12889,N_11671,N_11609);
nand U12890 (N_12890,N_11195,N_11566);
and U12891 (N_12891,N_11363,N_11455);
or U12892 (N_12892,N_11230,N_11626);
xnor U12893 (N_12893,N_11882,N_11739);
xor U12894 (N_12894,N_11283,N_11646);
xnor U12895 (N_12895,N_11497,N_11266);
and U12896 (N_12896,N_11764,N_11996);
or U12897 (N_12897,N_11399,N_11703);
or U12898 (N_12898,N_11814,N_11017);
nand U12899 (N_12899,N_11498,N_11936);
nand U12900 (N_12900,N_11747,N_11975);
xnor U12901 (N_12901,N_11182,N_11012);
nor U12902 (N_12902,N_11960,N_11654);
xor U12903 (N_12903,N_11765,N_11277);
xnor U12904 (N_12904,N_11963,N_11485);
xor U12905 (N_12905,N_11031,N_11459);
xnor U12906 (N_12906,N_11442,N_11242);
and U12907 (N_12907,N_11579,N_11063);
and U12908 (N_12908,N_11714,N_11126);
and U12909 (N_12909,N_11350,N_11669);
or U12910 (N_12910,N_11866,N_11060);
nand U12911 (N_12911,N_11841,N_11722);
and U12912 (N_12912,N_11780,N_11230);
and U12913 (N_12913,N_11143,N_11131);
xnor U12914 (N_12914,N_11889,N_11318);
nor U12915 (N_12915,N_11338,N_11453);
xnor U12916 (N_12916,N_11553,N_11284);
nor U12917 (N_12917,N_11710,N_11758);
nand U12918 (N_12918,N_11195,N_11416);
nand U12919 (N_12919,N_11141,N_11043);
or U12920 (N_12920,N_11996,N_11551);
and U12921 (N_12921,N_11447,N_11790);
and U12922 (N_12922,N_11766,N_11312);
nor U12923 (N_12923,N_11169,N_11719);
or U12924 (N_12924,N_11287,N_11911);
nand U12925 (N_12925,N_11461,N_11231);
nor U12926 (N_12926,N_11015,N_11863);
and U12927 (N_12927,N_11551,N_11390);
xnor U12928 (N_12928,N_11082,N_11438);
nand U12929 (N_12929,N_11758,N_11081);
and U12930 (N_12930,N_11996,N_11033);
and U12931 (N_12931,N_11479,N_11921);
nor U12932 (N_12932,N_11321,N_11160);
nand U12933 (N_12933,N_11209,N_11786);
xor U12934 (N_12934,N_11433,N_11847);
or U12935 (N_12935,N_11451,N_11401);
and U12936 (N_12936,N_11343,N_11157);
nand U12937 (N_12937,N_11088,N_11694);
or U12938 (N_12938,N_11056,N_11683);
and U12939 (N_12939,N_11026,N_11851);
and U12940 (N_12940,N_11600,N_11773);
nor U12941 (N_12941,N_11120,N_11879);
nand U12942 (N_12942,N_11163,N_11175);
and U12943 (N_12943,N_11575,N_11046);
or U12944 (N_12944,N_11659,N_11739);
nor U12945 (N_12945,N_11458,N_11197);
nand U12946 (N_12946,N_11716,N_11819);
or U12947 (N_12947,N_11888,N_11519);
xor U12948 (N_12948,N_11465,N_11484);
nor U12949 (N_12949,N_11288,N_11458);
nand U12950 (N_12950,N_11882,N_11090);
and U12951 (N_12951,N_11757,N_11296);
nor U12952 (N_12952,N_11151,N_11374);
nor U12953 (N_12953,N_11699,N_11911);
nor U12954 (N_12954,N_11339,N_11931);
xnor U12955 (N_12955,N_11997,N_11117);
or U12956 (N_12956,N_11083,N_11094);
nor U12957 (N_12957,N_11179,N_11015);
xor U12958 (N_12958,N_11512,N_11904);
xor U12959 (N_12959,N_11282,N_11172);
nor U12960 (N_12960,N_11354,N_11435);
xor U12961 (N_12961,N_11855,N_11983);
nand U12962 (N_12962,N_11754,N_11015);
nand U12963 (N_12963,N_11460,N_11546);
nand U12964 (N_12964,N_11077,N_11322);
nand U12965 (N_12965,N_11658,N_11122);
and U12966 (N_12966,N_11011,N_11513);
nor U12967 (N_12967,N_11714,N_11908);
or U12968 (N_12968,N_11006,N_11484);
nand U12969 (N_12969,N_11034,N_11381);
or U12970 (N_12970,N_11583,N_11336);
nor U12971 (N_12971,N_11385,N_11317);
and U12972 (N_12972,N_11950,N_11152);
xor U12973 (N_12973,N_11142,N_11398);
or U12974 (N_12974,N_11478,N_11716);
nor U12975 (N_12975,N_11577,N_11816);
and U12976 (N_12976,N_11199,N_11681);
or U12977 (N_12977,N_11223,N_11581);
and U12978 (N_12978,N_11997,N_11586);
nand U12979 (N_12979,N_11491,N_11082);
nor U12980 (N_12980,N_11328,N_11474);
and U12981 (N_12981,N_11325,N_11132);
or U12982 (N_12982,N_11048,N_11092);
and U12983 (N_12983,N_11976,N_11329);
nand U12984 (N_12984,N_11725,N_11020);
or U12985 (N_12985,N_11196,N_11195);
nand U12986 (N_12986,N_11382,N_11437);
nand U12987 (N_12987,N_11294,N_11896);
or U12988 (N_12988,N_11455,N_11935);
nand U12989 (N_12989,N_11880,N_11470);
xor U12990 (N_12990,N_11680,N_11307);
and U12991 (N_12991,N_11933,N_11666);
nand U12992 (N_12992,N_11533,N_11121);
xnor U12993 (N_12993,N_11883,N_11977);
nor U12994 (N_12994,N_11974,N_11413);
and U12995 (N_12995,N_11488,N_11298);
or U12996 (N_12996,N_11058,N_11996);
nor U12997 (N_12997,N_11537,N_11248);
nand U12998 (N_12998,N_11462,N_11329);
or U12999 (N_12999,N_11423,N_11904);
nor U13000 (N_13000,N_12979,N_12113);
nand U13001 (N_13001,N_12073,N_12642);
and U13002 (N_13002,N_12904,N_12859);
xnor U13003 (N_13003,N_12052,N_12489);
nor U13004 (N_13004,N_12107,N_12567);
and U13005 (N_13005,N_12829,N_12883);
nand U13006 (N_13006,N_12893,N_12830);
and U13007 (N_13007,N_12026,N_12190);
nor U13008 (N_13008,N_12901,N_12668);
and U13009 (N_13009,N_12866,N_12771);
nor U13010 (N_13010,N_12416,N_12229);
xor U13011 (N_13011,N_12576,N_12903);
xnor U13012 (N_13012,N_12290,N_12695);
and U13013 (N_13013,N_12943,N_12592);
or U13014 (N_13014,N_12178,N_12206);
or U13015 (N_13015,N_12264,N_12101);
nand U13016 (N_13016,N_12594,N_12498);
nor U13017 (N_13017,N_12602,N_12837);
xor U13018 (N_13018,N_12855,N_12126);
xnor U13019 (N_13019,N_12089,N_12329);
and U13020 (N_13020,N_12817,N_12388);
xnor U13021 (N_13021,N_12554,N_12856);
and U13022 (N_13022,N_12300,N_12608);
nand U13023 (N_13023,N_12906,N_12352);
xnor U13024 (N_13024,N_12278,N_12078);
or U13025 (N_13025,N_12560,N_12044);
nand U13026 (N_13026,N_12442,N_12670);
nand U13027 (N_13027,N_12994,N_12680);
and U13028 (N_13028,N_12372,N_12435);
or U13029 (N_13029,N_12623,N_12114);
nor U13030 (N_13030,N_12854,N_12577);
and U13031 (N_13031,N_12848,N_12985);
nand U13032 (N_13032,N_12010,N_12143);
nand U13033 (N_13033,N_12796,N_12378);
nor U13034 (N_13034,N_12481,N_12952);
and U13035 (N_13035,N_12539,N_12007);
and U13036 (N_13036,N_12675,N_12415);
nand U13037 (N_13037,N_12452,N_12136);
and U13038 (N_13038,N_12925,N_12125);
xnor U13039 (N_13039,N_12768,N_12050);
nor U13040 (N_13040,N_12786,N_12934);
xnor U13041 (N_13041,N_12860,N_12946);
nor U13042 (N_13042,N_12355,N_12558);
nand U13043 (N_13043,N_12729,N_12016);
xnor U13044 (N_13044,N_12940,N_12566);
nor U13045 (N_13045,N_12248,N_12028);
nand U13046 (N_13046,N_12779,N_12978);
xnor U13047 (N_13047,N_12165,N_12487);
or U13048 (N_13048,N_12317,N_12595);
xnor U13049 (N_13049,N_12490,N_12845);
nor U13050 (N_13050,N_12041,N_12606);
or U13051 (N_13051,N_12531,N_12534);
nand U13052 (N_13052,N_12631,N_12621);
xnor U13053 (N_13053,N_12221,N_12493);
nor U13054 (N_13054,N_12256,N_12699);
xor U13055 (N_13055,N_12155,N_12214);
nor U13056 (N_13056,N_12792,N_12599);
or U13057 (N_13057,N_12981,N_12331);
xnor U13058 (N_13058,N_12755,N_12931);
or U13059 (N_13059,N_12239,N_12316);
nand U13060 (N_13060,N_12156,N_12822);
nor U13061 (N_13061,N_12243,N_12718);
or U13062 (N_13062,N_12582,N_12789);
and U13063 (N_13063,N_12158,N_12207);
and U13064 (N_13064,N_12162,N_12289);
nand U13065 (N_13065,N_12501,N_12080);
xnor U13066 (N_13066,N_12068,N_12432);
or U13067 (N_13067,N_12613,N_12227);
xnor U13068 (N_13068,N_12223,N_12879);
nor U13069 (N_13069,N_12488,N_12077);
nand U13070 (N_13070,N_12431,N_12094);
or U13071 (N_13071,N_12141,N_12169);
xor U13072 (N_13072,N_12787,N_12987);
nand U13073 (N_13073,N_12698,N_12793);
nor U13074 (N_13074,N_12122,N_12970);
and U13075 (N_13075,N_12980,N_12087);
nor U13076 (N_13076,N_12543,N_12656);
nand U13077 (N_13077,N_12701,N_12466);
nor U13078 (N_13078,N_12727,N_12739);
nor U13079 (N_13079,N_12253,N_12968);
or U13080 (N_13080,N_12051,N_12622);
nand U13081 (N_13081,N_12537,N_12453);
and U13082 (N_13082,N_12425,N_12526);
nand U13083 (N_13083,N_12395,N_12332);
xnor U13084 (N_13084,N_12111,N_12942);
and U13085 (N_13085,N_12760,N_12836);
nand U13086 (N_13086,N_12882,N_12439);
xnor U13087 (N_13087,N_12540,N_12579);
nor U13088 (N_13088,N_12008,N_12957);
xor U13089 (N_13089,N_12049,N_12059);
or U13090 (N_13090,N_12939,N_12034);
nor U13091 (N_13091,N_12651,N_12853);
nor U13092 (N_13092,N_12387,N_12693);
nor U13093 (N_13093,N_12447,N_12632);
nand U13094 (N_13094,N_12174,N_12495);
and U13095 (N_13095,N_12884,N_12319);
xnor U13096 (N_13096,N_12983,N_12163);
and U13097 (N_13097,N_12139,N_12724);
or U13098 (N_13098,N_12605,N_12688);
nor U13099 (N_13099,N_12508,N_12524);
xnor U13100 (N_13100,N_12468,N_12285);
nor U13101 (N_13101,N_12090,N_12711);
xor U13102 (N_13102,N_12475,N_12330);
xor U13103 (N_13103,N_12694,N_12177);
nor U13104 (N_13104,N_12669,N_12210);
and U13105 (N_13105,N_12652,N_12963);
or U13106 (N_13106,N_12861,N_12244);
nand U13107 (N_13107,N_12639,N_12536);
xnor U13108 (N_13108,N_12772,N_12857);
nor U13109 (N_13109,N_12231,N_12245);
xor U13110 (N_13110,N_12828,N_12144);
nor U13111 (N_13111,N_12572,N_12671);
nor U13112 (N_13112,N_12851,N_12785);
and U13113 (N_13113,N_12635,N_12216);
nand U13114 (N_13114,N_12507,N_12203);
nand U13115 (N_13115,N_12871,N_12017);
nor U13116 (N_13116,N_12265,N_12810);
or U13117 (N_13117,N_12133,N_12304);
nor U13118 (N_13118,N_12287,N_12607);
nand U13119 (N_13119,N_12192,N_12862);
or U13120 (N_13120,N_12804,N_12657);
nand U13121 (N_13121,N_12018,N_12011);
xor U13122 (N_13122,N_12436,N_12181);
nand U13123 (N_13123,N_12972,N_12091);
xnor U13124 (N_13124,N_12166,N_12198);
nand U13125 (N_13125,N_12234,N_12847);
or U13126 (N_13126,N_12058,N_12267);
and U13127 (N_13127,N_12948,N_12926);
xor U13128 (N_13128,N_12662,N_12914);
nor U13129 (N_13129,N_12782,N_12868);
or U13130 (N_13130,N_12708,N_12081);
xor U13131 (N_13131,N_12037,N_12917);
and U13132 (N_13132,N_12767,N_12341);
xor U13133 (N_13133,N_12348,N_12315);
xor U13134 (N_13134,N_12411,N_12528);
or U13135 (N_13135,N_12544,N_12676);
or U13136 (N_13136,N_12298,N_12975);
and U13137 (N_13137,N_12308,N_12412);
nor U13138 (N_13138,N_12263,N_12811);
and U13139 (N_13139,N_12032,N_12532);
nand U13140 (N_13140,N_12824,N_12658);
nand U13141 (N_13141,N_12219,N_12197);
nand U13142 (N_13142,N_12097,N_12413);
or U13143 (N_13143,N_12428,N_12993);
and U13144 (N_13144,N_12681,N_12715);
nand U13145 (N_13145,N_12106,N_12805);
or U13146 (N_13146,N_12434,N_12825);
xor U13147 (N_13147,N_12795,N_12641);
or U13148 (N_13148,N_12838,N_12719);
xor U13149 (N_13149,N_12600,N_12677);
or U13150 (N_13150,N_12800,N_12405);
or U13151 (N_13151,N_12842,N_12124);
xnor U13152 (N_13152,N_12320,N_12874);
nor U13153 (N_13153,N_12679,N_12741);
nor U13154 (N_13154,N_12687,N_12057);
nand U13155 (N_13155,N_12328,N_12846);
and U13156 (N_13156,N_12568,N_12246);
xor U13157 (N_13157,N_12515,N_12104);
and U13158 (N_13158,N_12464,N_12312);
or U13159 (N_13159,N_12003,N_12826);
nor U13160 (N_13160,N_12305,N_12184);
and U13161 (N_13161,N_12773,N_12259);
nor U13162 (N_13162,N_12459,N_12752);
and U13163 (N_13163,N_12306,N_12645);
or U13164 (N_13164,N_12344,N_12474);
nor U13165 (N_13165,N_12666,N_12438);
and U13166 (N_13166,N_12483,N_12953);
nor U13167 (N_13167,N_12182,N_12019);
nand U13168 (N_13168,N_12685,N_12504);
or U13169 (N_13169,N_12189,N_12761);
nand U13170 (N_13170,N_12086,N_12697);
nor U13171 (N_13171,N_12923,N_12974);
xnor U13172 (N_13172,N_12938,N_12102);
or U13173 (N_13173,N_12581,N_12870);
nor U13174 (N_13174,N_12247,N_12816);
nand U13175 (N_13175,N_12397,N_12311);
or U13176 (N_13176,N_12295,N_12281);
xor U13177 (N_13177,N_12716,N_12261);
xor U13178 (N_13178,N_12389,N_12471);
and U13179 (N_13179,N_12364,N_12462);
nand U13180 (N_13180,N_12910,N_12712);
xnor U13181 (N_13181,N_12170,N_12218);
nor U13182 (N_13182,N_12888,N_12840);
and U13183 (N_13183,N_12650,N_12835);
nor U13184 (N_13184,N_12033,N_12947);
nand U13185 (N_13185,N_12250,N_12626);
nand U13186 (N_13186,N_12457,N_12375);
xor U13187 (N_13187,N_12895,N_12160);
or U13188 (N_13188,N_12777,N_12873);
nor U13189 (N_13189,N_12790,N_12065);
or U13190 (N_13190,N_12900,N_12056);
nor U13191 (N_13191,N_12713,N_12643);
nor U13192 (N_13192,N_12343,N_12665);
nand U13193 (N_13193,N_12120,N_12340);
and U13194 (N_13194,N_12396,N_12575);
nand U13195 (N_13195,N_12588,N_12990);
nor U13196 (N_13196,N_12337,N_12750);
xor U13197 (N_13197,N_12597,N_12615);
nand U13198 (N_13198,N_12744,N_12776);
nor U13199 (N_13199,N_12187,N_12527);
nor U13200 (N_13200,N_12446,N_12730);
xor U13201 (N_13201,N_12691,N_12808);
nor U13202 (N_13202,N_12885,N_12201);
nand U13203 (N_13203,N_12318,N_12284);
nor U13204 (N_13204,N_12110,N_12492);
or U13205 (N_13205,N_12754,N_12271);
and U13206 (N_13206,N_12633,N_12092);
nand U13207 (N_13207,N_12458,N_12421);
and U13208 (N_13208,N_12027,N_12580);
xnor U13209 (N_13209,N_12302,N_12031);
nand U13210 (N_13210,N_12944,N_12757);
nor U13211 (N_13211,N_12054,N_12272);
and U13212 (N_13212,N_12927,N_12038);
and U13213 (N_13213,N_12732,N_12047);
xnor U13214 (N_13214,N_12976,N_12408);
nor U13215 (N_13215,N_12103,N_12132);
xor U13216 (N_13216,N_12722,N_12589);
nor U13217 (N_13217,N_12908,N_12237);
nand U13218 (N_13218,N_12911,N_12630);
nor U13219 (N_13219,N_12749,N_12445);
xor U13220 (N_13220,N_12076,N_12273);
nand U13221 (N_13221,N_12366,N_12313);
xnor U13222 (N_13222,N_12074,N_12276);
xor U13223 (N_13223,N_12570,N_12516);
and U13224 (N_13224,N_12533,N_12919);
or U13225 (N_13225,N_12401,N_12105);
and U13226 (N_13226,N_12819,N_12646);
nand U13227 (N_13227,N_12996,N_12678);
and U13228 (N_13228,N_12707,N_12959);
nor U13229 (N_13229,N_12001,N_12061);
and U13230 (N_13230,N_12145,N_12999);
and U13231 (N_13231,N_12867,N_12154);
xnor U13232 (N_13232,N_12989,N_12128);
nand U13233 (N_13233,N_12562,N_12299);
or U13234 (N_13234,N_12735,N_12083);
nor U13235 (N_13235,N_12479,N_12283);
or U13236 (N_13236,N_12035,N_12067);
or U13237 (N_13237,N_12053,N_12213);
xnor U13238 (N_13238,N_12202,N_12486);
nand U13239 (N_13239,N_12894,N_12444);
and U13240 (N_13240,N_12303,N_12071);
nand U13241 (N_13241,N_12880,N_12667);
xor U13242 (N_13242,N_12945,N_12941);
and U13243 (N_13243,N_12381,N_12541);
or U13244 (N_13244,N_12359,N_12004);
and U13245 (N_13245,N_12150,N_12199);
nand U13246 (N_13246,N_12881,N_12907);
nor U13247 (N_13247,N_12045,N_12046);
xor U13248 (N_13248,N_12557,N_12598);
nor U13249 (N_13249,N_12021,N_12610);
nand U13250 (N_13250,N_12358,N_12733);
nand U13251 (N_13251,N_12494,N_12356);
nand U13252 (N_13252,N_12322,N_12241);
or U13253 (N_13253,N_12200,N_12036);
and U13254 (N_13254,N_12503,N_12039);
or U13255 (N_13255,N_12876,N_12763);
and U13256 (N_13256,N_12255,N_12960);
and U13257 (N_13257,N_12801,N_12638);
nor U13258 (N_13258,N_12357,N_12254);
and U13259 (N_13259,N_12628,N_12758);
xnor U13260 (N_13260,N_12618,N_12393);
nor U13261 (N_13261,N_12406,N_12585);
xor U13262 (N_13262,N_12386,N_12781);
xor U13263 (N_13263,N_12673,N_12916);
nand U13264 (N_13264,N_12173,N_12085);
nand U13265 (N_13265,N_12921,N_12653);
and U13266 (N_13266,N_12286,N_12522);
xor U13267 (N_13267,N_12686,N_12188);
xor U13268 (N_13268,N_12042,N_12417);
nand U13269 (N_13269,N_12784,N_12151);
nand U13270 (N_13270,N_12998,N_12672);
nand U13271 (N_13271,N_12731,N_12877);
nor U13272 (N_13272,N_12814,N_12043);
and U13273 (N_13273,N_12561,N_12753);
and U13274 (N_13274,N_12832,N_12186);
or U13275 (N_13275,N_12865,N_12211);
nand U13276 (N_13276,N_12482,N_12291);
or U13277 (N_13277,N_12084,N_12335);
and U13278 (N_13278,N_12721,N_12740);
xnor U13279 (N_13279,N_12280,N_12529);
or U13280 (N_13280,N_12629,N_12909);
xnor U13281 (N_13281,N_12193,N_12756);
nand U13282 (N_13282,N_12232,N_12725);
nor U13283 (N_13283,N_12022,N_12692);
nand U13284 (N_13284,N_12456,N_12469);
nor U13285 (N_13285,N_12933,N_12121);
nand U13286 (N_13286,N_12889,N_12726);
and U13287 (N_13287,N_12346,N_12172);
nand U13288 (N_13288,N_12611,N_12765);
nor U13289 (N_13289,N_12831,N_12684);
nor U13290 (N_13290,N_12858,N_12799);
xor U13291 (N_13291,N_12325,N_12728);
nand U13292 (N_13292,N_12924,N_12478);
xnor U13293 (N_13293,N_12863,N_12511);
xnor U13294 (N_13294,N_12555,N_12269);
nor U13295 (N_13295,N_12368,N_12260);
and U13296 (N_13296,N_12194,N_12183);
nand U13297 (N_13297,N_12205,N_12342);
or U13298 (N_13298,N_12209,N_12890);
and U13299 (N_13299,N_12336,N_12377);
nor U13300 (N_13300,N_12918,N_12204);
or U13301 (N_13301,N_12950,N_12887);
or U13302 (N_13302,N_12109,N_12292);
nor U13303 (N_13303,N_12545,N_12005);
and U13304 (N_13304,N_12228,N_12440);
or U13305 (N_13305,N_12400,N_12324);
nand U13306 (N_13306,N_12794,N_12360);
xnor U13307 (N_13307,N_12461,N_12149);
xnor U13308 (N_13308,N_12282,N_12778);
nand U13309 (N_13309,N_12674,N_12556);
xor U13310 (N_13310,N_12079,N_12617);
xnor U13311 (N_13311,N_12689,N_12803);
nand U13312 (N_13312,N_12820,N_12683);
nor U13313 (N_13313,N_12118,N_12573);
or U13314 (N_13314,N_12547,N_12326);
nor U13315 (N_13315,N_12896,N_12029);
and U13316 (N_13316,N_12171,N_12775);
and U13317 (N_13317,N_12798,N_12463);
or U13318 (N_13318,N_12659,N_12624);
nor U13319 (N_13319,N_12376,N_12815);
nor U13320 (N_13320,N_12929,N_12593);
xor U13321 (N_13321,N_12473,N_12590);
xor U13322 (N_13322,N_12899,N_12637);
xnor U13323 (N_13323,N_12964,N_12423);
xor U13324 (N_13324,N_12578,N_12382);
xor U13325 (N_13325,N_12099,N_12958);
xor U13326 (N_13326,N_12802,N_12864);
and U13327 (N_13327,N_12644,N_12982);
and U13328 (N_13328,N_12485,N_12745);
xnor U13329 (N_13329,N_12069,N_12497);
and U13330 (N_13330,N_12649,N_12362);
nor U13331 (N_13331,N_12410,N_12850);
xnor U13332 (N_13332,N_12000,N_12394);
nor U13333 (N_13333,N_12361,N_12409);
nand U13334 (N_13334,N_12971,N_12384);
nor U13335 (N_13335,N_12168,N_12986);
nand U13336 (N_13336,N_12640,N_12966);
and U13337 (N_13337,N_12129,N_12220);
xnor U13338 (N_13338,N_12791,N_12098);
or U13339 (N_13339,N_12454,N_12743);
nor U13340 (N_13340,N_12912,N_12130);
and U13341 (N_13341,N_12604,N_12212);
and U13342 (N_13342,N_12552,N_12620);
xor U13343 (N_13343,N_12852,N_12821);
and U13344 (N_13344,N_12152,N_12723);
xnor U13345 (N_13345,N_12339,N_12932);
and U13346 (N_13346,N_12517,N_12235);
nand U13347 (N_13347,N_12878,N_12140);
nand U13348 (N_13348,N_12157,N_12574);
nand U13349 (N_13349,N_12013,N_12569);
nor U13350 (N_13350,N_12634,N_12233);
nor U13351 (N_13351,N_12751,N_12663);
xnor U13352 (N_13352,N_12738,N_12208);
and U13353 (N_13353,N_12759,N_12661);
nand U13354 (N_13354,N_12512,N_12430);
or U13355 (N_13355,N_12530,N_12818);
nand U13356 (N_13356,N_12175,N_12748);
nand U13357 (N_13357,N_12612,N_12040);
or U13358 (N_13358,N_12403,N_12108);
xnor U13359 (N_13359,N_12238,N_12437);
nor U13360 (N_13360,N_12258,N_12134);
and U13361 (N_13361,N_12353,N_12636);
nand U13362 (N_13362,N_12424,N_12519);
and U13363 (N_13363,N_12060,N_12823);
xor U13364 (N_13364,N_12843,N_12350);
nor U13365 (N_13365,N_12892,N_12737);
nand U13366 (N_13366,N_12294,N_12465);
or U13367 (N_13367,N_12402,N_12138);
or U13368 (N_13368,N_12048,N_12700);
or U13369 (N_13369,N_12812,N_12967);
nor U13370 (N_13370,N_12277,N_12928);
nand U13371 (N_13371,N_12135,N_12391);
nor U13372 (N_13372,N_12023,N_12296);
and U13373 (N_13373,N_12100,N_12525);
or U13374 (N_13374,N_12167,N_12915);
nor U13375 (N_13375,N_12770,N_12849);
nand U13376 (N_13376,N_12546,N_12654);
or U13377 (N_13377,N_12995,N_12538);
or U13378 (N_13378,N_12734,N_12806);
and U13379 (N_13379,N_12476,N_12147);
nor U13380 (N_13380,N_12648,N_12148);
or U13381 (N_13381,N_12905,N_12327);
nand U13382 (N_13382,N_12509,N_12137);
xnor U13383 (N_13383,N_12603,N_12809);
xor U13384 (N_13384,N_12288,N_12704);
or U13385 (N_13385,N_12392,N_12553);
and U13386 (N_13386,N_12309,N_12176);
xnor U13387 (N_13387,N_12742,N_12467);
and U13388 (N_13388,N_12965,N_12872);
or U13389 (N_13389,N_12380,N_12523);
and U13390 (N_13390,N_12764,N_12333);
xor U13391 (N_13391,N_12370,N_12780);
nand U13392 (N_13392,N_12429,N_12420);
or U13393 (N_13393,N_12601,N_12185);
xor U13394 (N_13394,N_12559,N_12591);
xor U13395 (N_13395,N_12922,N_12690);
or U13396 (N_13396,N_12030,N_12345);
and U13397 (N_13397,N_12844,N_12146);
nand U13398 (N_13398,N_12788,N_12472);
xnor U13399 (N_13399,N_12379,N_12609);
xnor U13400 (N_13400,N_12902,N_12564);
or U13401 (N_13401,N_12619,N_12450);
and U13402 (N_13402,N_12002,N_12935);
nor U13403 (N_13403,N_12955,N_12123);
nor U13404 (N_13404,N_12647,N_12706);
nand U13405 (N_13405,N_12596,N_12367);
or U13406 (N_13406,N_12180,N_12949);
nor U13407 (N_13407,N_12012,N_12349);
xnor U13408 (N_13408,N_12913,N_12127);
and U13409 (N_13409,N_12548,N_12009);
nand U13410 (N_13410,N_12937,N_12072);
xnor U13411 (N_13411,N_12191,N_12584);
nand U13412 (N_13412,N_12164,N_12398);
nand U13413 (N_13413,N_12310,N_12696);
nand U13414 (N_13414,N_12627,N_12520);
xor U13415 (N_13415,N_12660,N_12470);
and U13416 (N_13416,N_12371,N_12954);
nor U13417 (N_13417,N_12427,N_12682);
or U13418 (N_13418,N_12338,N_12390);
and U13419 (N_13419,N_12433,N_12020);
or U13420 (N_13420,N_12441,N_12354);
and U13421 (N_13421,N_12351,N_12015);
nand U13422 (N_13422,N_12702,N_12897);
nor U13423 (N_13423,N_12369,N_12586);
or U13424 (N_13424,N_12119,N_12230);
nor U13425 (N_13425,N_12484,N_12518);
nor U13426 (N_13426,N_12251,N_12196);
xor U13427 (N_13427,N_12321,N_12962);
or U13428 (N_13428,N_12797,N_12833);
and U13429 (N_13429,N_12703,N_12563);
and U13430 (N_13430,N_12542,N_12502);
nor U13431 (N_13431,N_12116,N_12066);
or U13432 (N_13432,N_12279,N_12014);
xnor U13433 (N_13433,N_12616,N_12153);
nand U13434 (N_13434,N_12274,N_12500);
or U13435 (N_13435,N_12514,N_12070);
xnor U13436 (N_13436,N_12082,N_12813);
nor U13437 (N_13437,N_12774,N_12951);
or U13438 (N_13438,N_12736,N_12024);
nor U13439 (N_13439,N_12807,N_12549);
nand U13440 (N_13440,N_12055,N_12249);
xor U13441 (N_13441,N_12025,N_12268);
nor U13442 (N_13442,N_12385,N_12977);
xnor U13443 (N_13443,N_12571,N_12095);
and U13444 (N_13444,N_12834,N_12093);
and U13445 (N_13445,N_12480,N_12323);
and U13446 (N_13446,N_12006,N_12717);
nor U13447 (N_13447,N_12404,N_12293);
nor U13448 (N_13448,N_12969,N_12841);
or U13449 (N_13449,N_12891,N_12997);
nand U13450 (N_13450,N_12224,N_12550);
nor U13451 (N_13451,N_12875,N_12215);
or U13452 (N_13452,N_12365,N_12088);
or U13453 (N_13453,N_12827,N_12297);
and U13454 (N_13454,N_12383,N_12710);
and U13455 (N_13455,N_12499,N_12448);
or U13456 (N_13456,N_12614,N_12920);
xor U13457 (N_13457,N_12449,N_12535);
xor U13458 (N_13458,N_12422,N_12886);
xor U13459 (N_13459,N_12222,N_12992);
and U13460 (N_13460,N_12363,N_12374);
xor U13461 (N_13461,N_12240,N_12956);
xnor U13462 (N_13462,N_12505,N_12347);
xnor U13463 (N_13463,N_12451,N_12115);
xnor U13464 (N_13464,N_12266,N_12491);
or U13465 (N_13465,N_12869,N_12112);
and U13466 (N_13466,N_12314,N_12510);
nand U13467 (N_13467,N_12625,N_12307);
and U13468 (N_13468,N_12839,N_12655);
xnor U13469 (N_13469,N_12513,N_12988);
nand U13470 (N_13470,N_12746,N_12195);
nand U13471 (N_13471,N_12063,N_12783);
and U13472 (N_13472,N_12496,N_12226);
nand U13473 (N_13473,N_12418,N_12275);
nor U13474 (N_13474,N_12709,N_12301);
or U13475 (N_13475,N_12984,N_12407);
xor U13476 (N_13476,N_12521,N_12714);
or U13477 (N_13477,N_12443,N_12460);
and U13478 (N_13478,N_12414,N_12506);
nor U13479 (N_13479,N_12762,N_12257);
or U13480 (N_13480,N_12991,N_12426);
or U13481 (N_13481,N_12064,N_12075);
nand U13482 (N_13482,N_12930,N_12705);
nor U13483 (N_13483,N_12455,N_12096);
and U13484 (N_13484,N_12747,N_12252);
nand U13485 (N_13485,N_12769,N_12477);
nand U13486 (N_13486,N_12587,N_12262);
xnor U13487 (N_13487,N_12664,N_12142);
nand U13488 (N_13488,N_12062,N_12131);
xnor U13489 (N_13489,N_12720,N_12936);
and U13490 (N_13490,N_12551,N_12117);
nand U13491 (N_13491,N_12973,N_12225);
nor U13492 (N_13492,N_12270,N_12898);
or U13493 (N_13493,N_12161,N_12159);
nor U13494 (N_13494,N_12334,N_12373);
and U13495 (N_13495,N_12217,N_12419);
xor U13496 (N_13496,N_12242,N_12565);
nor U13497 (N_13497,N_12766,N_12179);
nor U13498 (N_13498,N_12399,N_12961);
and U13499 (N_13499,N_12236,N_12583);
nor U13500 (N_13500,N_12549,N_12531);
xor U13501 (N_13501,N_12852,N_12381);
xor U13502 (N_13502,N_12251,N_12343);
and U13503 (N_13503,N_12357,N_12436);
nor U13504 (N_13504,N_12621,N_12660);
and U13505 (N_13505,N_12377,N_12299);
xnor U13506 (N_13506,N_12177,N_12865);
and U13507 (N_13507,N_12660,N_12391);
and U13508 (N_13508,N_12089,N_12343);
nor U13509 (N_13509,N_12098,N_12457);
nor U13510 (N_13510,N_12693,N_12934);
and U13511 (N_13511,N_12849,N_12473);
xor U13512 (N_13512,N_12040,N_12435);
xnor U13513 (N_13513,N_12342,N_12449);
nor U13514 (N_13514,N_12063,N_12650);
xnor U13515 (N_13515,N_12599,N_12077);
nor U13516 (N_13516,N_12091,N_12716);
and U13517 (N_13517,N_12503,N_12530);
xnor U13518 (N_13518,N_12840,N_12367);
and U13519 (N_13519,N_12187,N_12218);
nor U13520 (N_13520,N_12108,N_12579);
nor U13521 (N_13521,N_12102,N_12694);
and U13522 (N_13522,N_12306,N_12506);
nand U13523 (N_13523,N_12380,N_12780);
nor U13524 (N_13524,N_12234,N_12233);
xnor U13525 (N_13525,N_12129,N_12630);
and U13526 (N_13526,N_12893,N_12581);
or U13527 (N_13527,N_12134,N_12518);
or U13528 (N_13528,N_12108,N_12700);
and U13529 (N_13529,N_12286,N_12425);
and U13530 (N_13530,N_12588,N_12289);
nor U13531 (N_13531,N_12153,N_12648);
nand U13532 (N_13532,N_12393,N_12172);
xor U13533 (N_13533,N_12582,N_12466);
and U13534 (N_13534,N_12368,N_12940);
nand U13535 (N_13535,N_12244,N_12704);
or U13536 (N_13536,N_12512,N_12305);
and U13537 (N_13537,N_12472,N_12902);
or U13538 (N_13538,N_12577,N_12882);
nor U13539 (N_13539,N_12222,N_12009);
nor U13540 (N_13540,N_12098,N_12711);
or U13541 (N_13541,N_12358,N_12739);
nor U13542 (N_13542,N_12642,N_12111);
and U13543 (N_13543,N_12898,N_12935);
or U13544 (N_13544,N_12065,N_12483);
nand U13545 (N_13545,N_12732,N_12291);
nand U13546 (N_13546,N_12392,N_12500);
or U13547 (N_13547,N_12281,N_12211);
nor U13548 (N_13548,N_12638,N_12847);
nor U13549 (N_13549,N_12656,N_12947);
or U13550 (N_13550,N_12369,N_12672);
xor U13551 (N_13551,N_12911,N_12893);
and U13552 (N_13552,N_12537,N_12870);
or U13553 (N_13553,N_12473,N_12043);
nor U13554 (N_13554,N_12513,N_12850);
and U13555 (N_13555,N_12253,N_12714);
xor U13556 (N_13556,N_12237,N_12268);
xnor U13557 (N_13557,N_12498,N_12771);
and U13558 (N_13558,N_12460,N_12319);
or U13559 (N_13559,N_12673,N_12131);
nor U13560 (N_13560,N_12566,N_12367);
and U13561 (N_13561,N_12410,N_12840);
and U13562 (N_13562,N_12224,N_12453);
and U13563 (N_13563,N_12801,N_12472);
xnor U13564 (N_13564,N_12102,N_12309);
or U13565 (N_13565,N_12116,N_12491);
nand U13566 (N_13566,N_12663,N_12065);
xor U13567 (N_13567,N_12940,N_12398);
nand U13568 (N_13568,N_12371,N_12302);
nand U13569 (N_13569,N_12354,N_12004);
nor U13570 (N_13570,N_12626,N_12918);
xnor U13571 (N_13571,N_12876,N_12766);
xnor U13572 (N_13572,N_12583,N_12941);
xor U13573 (N_13573,N_12372,N_12359);
nand U13574 (N_13574,N_12854,N_12805);
or U13575 (N_13575,N_12626,N_12111);
nor U13576 (N_13576,N_12652,N_12348);
xor U13577 (N_13577,N_12809,N_12645);
nor U13578 (N_13578,N_12216,N_12221);
nand U13579 (N_13579,N_12869,N_12426);
and U13580 (N_13580,N_12013,N_12231);
nor U13581 (N_13581,N_12999,N_12290);
nand U13582 (N_13582,N_12343,N_12954);
xnor U13583 (N_13583,N_12678,N_12771);
nor U13584 (N_13584,N_12807,N_12904);
xor U13585 (N_13585,N_12669,N_12667);
or U13586 (N_13586,N_12045,N_12668);
nor U13587 (N_13587,N_12981,N_12602);
or U13588 (N_13588,N_12727,N_12807);
and U13589 (N_13589,N_12546,N_12498);
and U13590 (N_13590,N_12077,N_12388);
nor U13591 (N_13591,N_12871,N_12079);
xnor U13592 (N_13592,N_12044,N_12555);
nor U13593 (N_13593,N_12367,N_12880);
nand U13594 (N_13594,N_12509,N_12879);
nor U13595 (N_13595,N_12212,N_12924);
nand U13596 (N_13596,N_12158,N_12611);
or U13597 (N_13597,N_12185,N_12255);
nand U13598 (N_13598,N_12670,N_12588);
and U13599 (N_13599,N_12931,N_12552);
nand U13600 (N_13600,N_12055,N_12005);
nand U13601 (N_13601,N_12035,N_12021);
nand U13602 (N_13602,N_12674,N_12727);
nand U13603 (N_13603,N_12555,N_12196);
nor U13604 (N_13604,N_12818,N_12723);
nand U13605 (N_13605,N_12265,N_12699);
nand U13606 (N_13606,N_12335,N_12657);
and U13607 (N_13607,N_12701,N_12300);
and U13608 (N_13608,N_12513,N_12152);
or U13609 (N_13609,N_12259,N_12550);
and U13610 (N_13610,N_12660,N_12247);
xor U13611 (N_13611,N_12888,N_12770);
or U13612 (N_13612,N_12130,N_12995);
and U13613 (N_13613,N_12025,N_12393);
xnor U13614 (N_13614,N_12759,N_12571);
xnor U13615 (N_13615,N_12395,N_12768);
and U13616 (N_13616,N_12697,N_12539);
or U13617 (N_13617,N_12522,N_12263);
xnor U13618 (N_13618,N_12054,N_12947);
or U13619 (N_13619,N_12523,N_12368);
nand U13620 (N_13620,N_12099,N_12137);
nand U13621 (N_13621,N_12554,N_12808);
xnor U13622 (N_13622,N_12284,N_12247);
or U13623 (N_13623,N_12368,N_12821);
xor U13624 (N_13624,N_12931,N_12004);
nand U13625 (N_13625,N_12977,N_12822);
nor U13626 (N_13626,N_12357,N_12726);
and U13627 (N_13627,N_12923,N_12539);
nor U13628 (N_13628,N_12221,N_12065);
and U13629 (N_13629,N_12376,N_12407);
xor U13630 (N_13630,N_12111,N_12780);
or U13631 (N_13631,N_12733,N_12629);
nor U13632 (N_13632,N_12227,N_12356);
xnor U13633 (N_13633,N_12002,N_12996);
and U13634 (N_13634,N_12277,N_12591);
nor U13635 (N_13635,N_12314,N_12219);
xnor U13636 (N_13636,N_12498,N_12000);
nor U13637 (N_13637,N_12973,N_12598);
xor U13638 (N_13638,N_12606,N_12686);
nor U13639 (N_13639,N_12691,N_12455);
nand U13640 (N_13640,N_12955,N_12815);
and U13641 (N_13641,N_12646,N_12822);
and U13642 (N_13642,N_12215,N_12925);
xor U13643 (N_13643,N_12076,N_12679);
nor U13644 (N_13644,N_12912,N_12323);
nand U13645 (N_13645,N_12381,N_12201);
xor U13646 (N_13646,N_12267,N_12113);
nand U13647 (N_13647,N_12403,N_12951);
xnor U13648 (N_13648,N_12188,N_12919);
and U13649 (N_13649,N_12552,N_12200);
nor U13650 (N_13650,N_12826,N_12564);
or U13651 (N_13651,N_12395,N_12721);
xnor U13652 (N_13652,N_12383,N_12957);
nor U13653 (N_13653,N_12029,N_12932);
nand U13654 (N_13654,N_12815,N_12855);
nand U13655 (N_13655,N_12747,N_12642);
nand U13656 (N_13656,N_12694,N_12422);
and U13657 (N_13657,N_12421,N_12873);
xnor U13658 (N_13658,N_12560,N_12883);
or U13659 (N_13659,N_12561,N_12998);
xnor U13660 (N_13660,N_12744,N_12577);
nor U13661 (N_13661,N_12347,N_12787);
nor U13662 (N_13662,N_12379,N_12364);
and U13663 (N_13663,N_12262,N_12618);
xor U13664 (N_13664,N_12664,N_12329);
and U13665 (N_13665,N_12666,N_12447);
nand U13666 (N_13666,N_12988,N_12494);
xor U13667 (N_13667,N_12499,N_12701);
or U13668 (N_13668,N_12060,N_12056);
nor U13669 (N_13669,N_12053,N_12498);
nor U13670 (N_13670,N_12657,N_12361);
nand U13671 (N_13671,N_12231,N_12981);
nand U13672 (N_13672,N_12236,N_12289);
xnor U13673 (N_13673,N_12172,N_12031);
nand U13674 (N_13674,N_12762,N_12605);
nor U13675 (N_13675,N_12781,N_12207);
and U13676 (N_13676,N_12251,N_12187);
nor U13677 (N_13677,N_12231,N_12001);
nor U13678 (N_13678,N_12972,N_12179);
and U13679 (N_13679,N_12822,N_12401);
or U13680 (N_13680,N_12578,N_12505);
or U13681 (N_13681,N_12515,N_12259);
nor U13682 (N_13682,N_12643,N_12137);
and U13683 (N_13683,N_12114,N_12045);
nand U13684 (N_13684,N_12009,N_12094);
and U13685 (N_13685,N_12007,N_12990);
nor U13686 (N_13686,N_12504,N_12733);
and U13687 (N_13687,N_12114,N_12634);
nor U13688 (N_13688,N_12377,N_12087);
nor U13689 (N_13689,N_12790,N_12970);
or U13690 (N_13690,N_12196,N_12161);
nand U13691 (N_13691,N_12614,N_12033);
nor U13692 (N_13692,N_12099,N_12577);
xor U13693 (N_13693,N_12830,N_12491);
nor U13694 (N_13694,N_12784,N_12174);
nor U13695 (N_13695,N_12505,N_12360);
nand U13696 (N_13696,N_12508,N_12552);
nand U13697 (N_13697,N_12798,N_12531);
xnor U13698 (N_13698,N_12451,N_12519);
xnor U13699 (N_13699,N_12589,N_12182);
or U13700 (N_13700,N_12930,N_12245);
nor U13701 (N_13701,N_12963,N_12366);
xnor U13702 (N_13702,N_12635,N_12704);
or U13703 (N_13703,N_12322,N_12833);
and U13704 (N_13704,N_12764,N_12157);
nand U13705 (N_13705,N_12241,N_12090);
nor U13706 (N_13706,N_12983,N_12174);
nor U13707 (N_13707,N_12926,N_12479);
or U13708 (N_13708,N_12622,N_12355);
xor U13709 (N_13709,N_12567,N_12575);
nor U13710 (N_13710,N_12210,N_12524);
or U13711 (N_13711,N_12568,N_12060);
or U13712 (N_13712,N_12918,N_12862);
and U13713 (N_13713,N_12922,N_12827);
and U13714 (N_13714,N_12249,N_12589);
and U13715 (N_13715,N_12952,N_12846);
and U13716 (N_13716,N_12874,N_12239);
nor U13717 (N_13717,N_12719,N_12722);
and U13718 (N_13718,N_12731,N_12603);
nor U13719 (N_13719,N_12684,N_12208);
and U13720 (N_13720,N_12381,N_12650);
xnor U13721 (N_13721,N_12426,N_12904);
xor U13722 (N_13722,N_12405,N_12555);
nand U13723 (N_13723,N_12601,N_12341);
nor U13724 (N_13724,N_12422,N_12835);
xnor U13725 (N_13725,N_12217,N_12761);
or U13726 (N_13726,N_12217,N_12915);
xnor U13727 (N_13727,N_12094,N_12840);
and U13728 (N_13728,N_12524,N_12882);
or U13729 (N_13729,N_12515,N_12527);
nand U13730 (N_13730,N_12177,N_12875);
nand U13731 (N_13731,N_12557,N_12325);
xnor U13732 (N_13732,N_12037,N_12551);
xor U13733 (N_13733,N_12505,N_12559);
xor U13734 (N_13734,N_12082,N_12882);
nor U13735 (N_13735,N_12752,N_12943);
nand U13736 (N_13736,N_12679,N_12494);
or U13737 (N_13737,N_12917,N_12891);
and U13738 (N_13738,N_12049,N_12629);
and U13739 (N_13739,N_12759,N_12094);
nor U13740 (N_13740,N_12488,N_12850);
or U13741 (N_13741,N_12649,N_12327);
nand U13742 (N_13742,N_12871,N_12579);
and U13743 (N_13743,N_12293,N_12673);
xor U13744 (N_13744,N_12318,N_12898);
nand U13745 (N_13745,N_12326,N_12997);
or U13746 (N_13746,N_12655,N_12667);
or U13747 (N_13747,N_12282,N_12160);
and U13748 (N_13748,N_12979,N_12628);
xnor U13749 (N_13749,N_12718,N_12948);
nand U13750 (N_13750,N_12988,N_12526);
nor U13751 (N_13751,N_12145,N_12228);
and U13752 (N_13752,N_12409,N_12510);
nor U13753 (N_13753,N_12266,N_12089);
nor U13754 (N_13754,N_12850,N_12430);
nand U13755 (N_13755,N_12478,N_12200);
or U13756 (N_13756,N_12758,N_12545);
nand U13757 (N_13757,N_12343,N_12337);
or U13758 (N_13758,N_12420,N_12313);
and U13759 (N_13759,N_12815,N_12162);
and U13760 (N_13760,N_12974,N_12566);
nor U13761 (N_13761,N_12532,N_12318);
xor U13762 (N_13762,N_12510,N_12887);
and U13763 (N_13763,N_12407,N_12406);
and U13764 (N_13764,N_12261,N_12313);
nand U13765 (N_13765,N_12081,N_12664);
or U13766 (N_13766,N_12918,N_12467);
xnor U13767 (N_13767,N_12315,N_12723);
or U13768 (N_13768,N_12169,N_12923);
or U13769 (N_13769,N_12548,N_12938);
and U13770 (N_13770,N_12001,N_12349);
nor U13771 (N_13771,N_12002,N_12215);
xor U13772 (N_13772,N_12713,N_12317);
and U13773 (N_13773,N_12203,N_12350);
or U13774 (N_13774,N_12919,N_12626);
nand U13775 (N_13775,N_12840,N_12697);
nand U13776 (N_13776,N_12988,N_12396);
and U13777 (N_13777,N_12556,N_12399);
and U13778 (N_13778,N_12316,N_12147);
nand U13779 (N_13779,N_12966,N_12092);
and U13780 (N_13780,N_12995,N_12476);
xnor U13781 (N_13781,N_12023,N_12243);
and U13782 (N_13782,N_12184,N_12272);
nand U13783 (N_13783,N_12458,N_12418);
nor U13784 (N_13784,N_12800,N_12473);
or U13785 (N_13785,N_12933,N_12500);
nand U13786 (N_13786,N_12156,N_12845);
and U13787 (N_13787,N_12912,N_12947);
xnor U13788 (N_13788,N_12085,N_12087);
or U13789 (N_13789,N_12197,N_12040);
xor U13790 (N_13790,N_12419,N_12126);
xor U13791 (N_13791,N_12235,N_12625);
xor U13792 (N_13792,N_12878,N_12900);
or U13793 (N_13793,N_12698,N_12854);
nand U13794 (N_13794,N_12586,N_12067);
or U13795 (N_13795,N_12185,N_12293);
or U13796 (N_13796,N_12009,N_12765);
nand U13797 (N_13797,N_12845,N_12417);
or U13798 (N_13798,N_12914,N_12450);
nor U13799 (N_13799,N_12898,N_12656);
or U13800 (N_13800,N_12517,N_12642);
xnor U13801 (N_13801,N_12662,N_12026);
or U13802 (N_13802,N_12447,N_12437);
xor U13803 (N_13803,N_12722,N_12631);
or U13804 (N_13804,N_12994,N_12578);
nand U13805 (N_13805,N_12430,N_12729);
and U13806 (N_13806,N_12851,N_12709);
nor U13807 (N_13807,N_12206,N_12873);
nor U13808 (N_13808,N_12810,N_12361);
or U13809 (N_13809,N_12627,N_12079);
nand U13810 (N_13810,N_12263,N_12370);
or U13811 (N_13811,N_12972,N_12756);
nand U13812 (N_13812,N_12974,N_12621);
nand U13813 (N_13813,N_12602,N_12100);
nand U13814 (N_13814,N_12533,N_12316);
or U13815 (N_13815,N_12957,N_12832);
nand U13816 (N_13816,N_12304,N_12590);
xor U13817 (N_13817,N_12661,N_12543);
or U13818 (N_13818,N_12034,N_12201);
nand U13819 (N_13819,N_12937,N_12251);
or U13820 (N_13820,N_12667,N_12185);
xnor U13821 (N_13821,N_12233,N_12055);
xor U13822 (N_13822,N_12104,N_12455);
nand U13823 (N_13823,N_12301,N_12675);
nor U13824 (N_13824,N_12575,N_12815);
and U13825 (N_13825,N_12087,N_12907);
nor U13826 (N_13826,N_12263,N_12866);
nand U13827 (N_13827,N_12519,N_12138);
nand U13828 (N_13828,N_12835,N_12481);
nor U13829 (N_13829,N_12717,N_12911);
xor U13830 (N_13830,N_12283,N_12176);
and U13831 (N_13831,N_12927,N_12988);
or U13832 (N_13832,N_12350,N_12999);
and U13833 (N_13833,N_12958,N_12915);
nor U13834 (N_13834,N_12596,N_12674);
or U13835 (N_13835,N_12348,N_12649);
nor U13836 (N_13836,N_12131,N_12761);
nand U13837 (N_13837,N_12030,N_12684);
and U13838 (N_13838,N_12583,N_12676);
or U13839 (N_13839,N_12934,N_12023);
and U13840 (N_13840,N_12296,N_12490);
nor U13841 (N_13841,N_12766,N_12193);
nand U13842 (N_13842,N_12294,N_12534);
or U13843 (N_13843,N_12057,N_12963);
nor U13844 (N_13844,N_12483,N_12159);
nor U13845 (N_13845,N_12150,N_12484);
or U13846 (N_13846,N_12333,N_12069);
nand U13847 (N_13847,N_12756,N_12133);
and U13848 (N_13848,N_12368,N_12580);
and U13849 (N_13849,N_12401,N_12504);
nor U13850 (N_13850,N_12586,N_12205);
or U13851 (N_13851,N_12238,N_12891);
xor U13852 (N_13852,N_12965,N_12011);
and U13853 (N_13853,N_12336,N_12479);
xor U13854 (N_13854,N_12840,N_12456);
and U13855 (N_13855,N_12184,N_12416);
or U13856 (N_13856,N_12742,N_12031);
nand U13857 (N_13857,N_12009,N_12697);
or U13858 (N_13858,N_12903,N_12863);
and U13859 (N_13859,N_12825,N_12902);
or U13860 (N_13860,N_12994,N_12668);
and U13861 (N_13861,N_12416,N_12603);
or U13862 (N_13862,N_12094,N_12884);
and U13863 (N_13863,N_12090,N_12850);
nor U13864 (N_13864,N_12330,N_12024);
nor U13865 (N_13865,N_12971,N_12265);
or U13866 (N_13866,N_12033,N_12451);
nor U13867 (N_13867,N_12457,N_12501);
xnor U13868 (N_13868,N_12924,N_12897);
and U13869 (N_13869,N_12143,N_12580);
and U13870 (N_13870,N_12487,N_12832);
nor U13871 (N_13871,N_12778,N_12592);
nor U13872 (N_13872,N_12040,N_12919);
xnor U13873 (N_13873,N_12603,N_12996);
or U13874 (N_13874,N_12866,N_12181);
xor U13875 (N_13875,N_12957,N_12917);
nand U13876 (N_13876,N_12530,N_12247);
or U13877 (N_13877,N_12311,N_12126);
nand U13878 (N_13878,N_12164,N_12033);
and U13879 (N_13879,N_12903,N_12583);
nor U13880 (N_13880,N_12393,N_12915);
xnor U13881 (N_13881,N_12474,N_12982);
or U13882 (N_13882,N_12606,N_12262);
nand U13883 (N_13883,N_12187,N_12078);
nand U13884 (N_13884,N_12595,N_12983);
xnor U13885 (N_13885,N_12079,N_12982);
and U13886 (N_13886,N_12831,N_12277);
xor U13887 (N_13887,N_12100,N_12998);
nor U13888 (N_13888,N_12934,N_12366);
and U13889 (N_13889,N_12995,N_12330);
nand U13890 (N_13890,N_12857,N_12558);
nand U13891 (N_13891,N_12932,N_12595);
xor U13892 (N_13892,N_12511,N_12372);
nand U13893 (N_13893,N_12694,N_12956);
nor U13894 (N_13894,N_12631,N_12932);
or U13895 (N_13895,N_12129,N_12532);
xor U13896 (N_13896,N_12345,N_12437);
nor U13897 (N_13897,N_12260,N_12002);
nor U13898 (N_13898,N_12590,N_12142);
xor U13899 (N_13899,N_12523,N_12906);
or U13900 (N_13900,N_12938,N_12875);
or U13901 (N_13901,N_12357,N_12094);
nand U13902 (N_13902,N_12773,N_12086);
and U13903 (N_13903,N_12031,N_12801);
and U13904 (N_13904,N_12689,N_12343);
or U13905 (N_13905,N_12473,N_12191);
nor U13906 (N_13906,N_12448,N_12236);
or U13907 (N_13907,N_12988,N_12193);
xor U13908 (N_13908,N_12719,N_12904);
nor U13909 (N_13909,N_12804,N_12701);
xnor U13910 (N_13910,N_12582,N_12463);
nand U13911 (N_13911,N_12903,N_12737);
nor U13912 (N_13912,N_12038,N_12141);
nand U13913 (N_13913,N_12672,N_12691);
xnor U13914 (N_13914,N_12399,N_12375);
nand U13915 (N_13915,N_12606,N_12702);
and U13916 (N_13916,N_12732,N_12066);
and U13917 (N_13917,N_12995,N_12474);
nand U13918 (N_13918,N_12692,N_12031);
and U13919 (N_13919,N_12343,N_12699);
and U13920 (N_13920,N_12285,N_12673);
and U13921 (N_13921,N_12948,N_12180);
nand U13922 (N_13922,N_12918,N_12248);
or U13923 (N_13923,N_12561,N_12097);
xnor U13924 (N_13924,N_12992,N_12469);
xor U13925 (N_13925,N_12097,N_12745);
and U13926 (N_13926,N_12945,N_12067);
nand U13927 (N_13927,N_12079,N_12305);
and U13928 (N_13928,N_12483,N_12150);
and U13929 (N_13929,N_12017,N_12174);
nor U13930 (N_13930,N_12664,N_12207);
and U13931 (N_13931,N_12255,N_12416);
xor U13932 (N_13932,N_12923,N_12633);
nor U13933 (N_13933,N_12916,N_12081);
or U13934 (N_13934,N_12793,N_12814);
and U13935 (N_13935,N_12935,N_12176);
and U13936 (N_13936,N_12567,N_12273);
nor U13937 (N_13937,N_12917,N_12033);
nor U13938 (N_13938,N_12494,N_12663);
or U13939 (N_13939,N_12101,N_12435);
xnor U13940 (N_13940,N_12240,N_12861);
xnor U13941 (N_13941,N_12863,N_12181);
nor U13942 (N_13942,N_12349,N_12287);
xnor U13943 (N_13943,N_12632,N_12343);
nand U13944 (N_13944,N_12300,N_12652);
nand U13945 (N_13945,N_12389,N_12526);
nand U13946 (N_13946,N_12506,N_12681);
xnor U13947 (N_13947,N_12031,N_12202);
xor U13948 (N_13948,N_12455,N_12892);
xnor U13949 (N_13949,N_12859,N_12093);
or U13950 (N_13950,N_12758,N_12492);
or U13951 (N_13951,N_12559,N_12310);
xnor U13952 (N_13952,N_12277,N_12795);
nor U13953 (N_13953,N_12070,N_12682);
xor U13954 (N_13954,N_12923,N_12722);
or U13955 (N_13955,N_12714,N_12602);
nand U13956 (N_13956,N_12823,N_12176);
nand U13957 (N_13957,N_12785,N_12750);
xor U13958 (N_13958,N_12763,N_12099);
xor U13959 (N_13959,N_12844,N_12760);
nor U13960 (N_13960,N_12203,N_12868);
xnor U13961 (N_13961,N_12310,N_12195);
nand U13962 (N_13962,N_12150,N_12117);
nor U13963 (N_13963,N_12788,N_12246);
nor U13964 (N_13964,N_12526,N_12055);
nor U13965 (N_13965,N_12755,N_12751);
and U13966 (N_13966,N_12954,N_12568);
and U13967 (N_13967,N_12606,N_12751);
or U13968 (N_13968,N_12480,N_12254);
and U13969 (N_13969,N_12925,N_12435);
nand U13970 (N_13970,N_12418,N_12915);
nand U13971 (N_13971,N_12680,N_12037);
nor U13972 (N_13972,N_12911,N_12502);
xnor U13973 (N_13973,N_12916,N_12562);
nand U13974 (N_13974,N_12966,N_12237);
nand U13975 (N_13975,N_12793,N_12416);
xor U13976 (N_13976,N_12430,N_12187);
or U13977 (N_13977,N_12926,N_12903);
nor U13978 (N_13978,N_12590,N_12189);
and U13979 (N_13979,N_12411,N_12786);
or U13980 (N_13980,N_12281,N_12434);
nand U13981 (N_13981,N_12367,N_12945);
nor U13982 (N_13982,N_12418,N_12048);
xnor U13983 (N_13983,N_12411,N_12184);
nor U13984 (N_13984,N_12241,N_12927);
or U13985 (N_13985,N_12652,N_12301);
nor U13986 (N_13986,N_12777,N_12728);
and U13987 (N_13987,N_12287,N_12686);
xnor U13988 (N_13988,N_12563,N_12006);
nor U13989 (N_13989,N_12364,N_12801);
xor U13990 (N_13990,N_12051,N_12595);
and U13991 (N_13991,N_12433,N_12369);
nand U13992 (N_13992,N_12224,N_12861);
nor U13993 (N_13993,N_12857,N_12423);
nor U13994 (N_13994,N_12270,N_12021);
xnor U13995 (N_13995,N_12115,N_12226);
nor U13996 (N_13996,N_12410,N_12908);
xor U13997 (N_13997,N_12728,N_12219);
and U13998 (N_13998,N_12940,N_12336);
nand U13999 (N_13999,N_12133,N_12358);
and U14000 (N_14000,N_13147,N_13158);
and U14001 (N_14001,N_13439,N_13737);
nand U14002 (N_14002,N_13132,N_13687);
or U14003 (N_14003,N_13528,N_13004);
and U14004 (N_14004,N_13465,N_13875);
nor U14005 (N_14005,N_13005,N_13759);
nand U14006 (N_14006,N_13643,N_13275);
nor U14007 (N_14007,N_13827,N_13518);
or U14008 (N_14008,N_13848,N_13935);
or U14009 (N_14009,N_13671,N_13870);
nor U14010 (N_14010,N_13694,N_13812);
nor U14011 (N_14011,N_13548,N_13809);
nor U14012 (N_14012,N_13762,N_13562);
xor U14013 (N_14013,N_13222,N_13735);
nor U14014 (N_14014,N_13788,N_13586);
xor U14015 (N_14015,N_13311,N_13955);
or U14016 (N_14016,N_13183,N_13137);
xor U14017 (N_14017,N_13422,N_13871);
xnor U14018 (N_14018,N_13866,N_13313);
or U14019 (N_14019,N_13908,N_13393);
nand U14020 (N_14020,N_13302,N_13757);
nor U14021 (N_14021,N_13987,N_13516);
and U14022 (N_14022,N_13801,N_13943);
nor U14023 (N_14023,N_13052,N_13717);
nor U14024 (N_14024,N_13670,N_13392);
or U14025 (N_14025,N_13751,N_13403);
and U14026 (N_14026,N_13780,N_13909);
nor U14027 (N_14027,N_13248,N_13127);
or U14028 (N_14028,N_13122,N_13542);
xor U14029 (N_14029,N_13881,N_13773);
or U14030 (N_14030,N_13649,N_13854);
xnor U14031 (N_14031,N_13497,N_13188);
nand U14032 (N_14032,N_13981,N_13842);
xor U14033 (N_14033,N_13769,N_13993);
and U14034 (N_14034,N_13511,N_13262);
or U14035 (N_14035,N_13416,N_13829);
or U14036 (N_14036,N_13556,N_13772);
xor U14037 (N_14037,N_13195,N_13309);
or U14038 (N_14038,N_13090,N_13216);
xor U14039 (N_14039,N_13035,N_13808);
nor U14040 (N_14040,N_13153,N_13464);
or U14041 (N_14041,N_13844,N_13891);
nor U14042 (N_14042,N_13106,N_13790);
or U14043 (N_14043,N_13830,N_13385);
nand U14044 (N_14044,N_13240,N_13488);
or U14045 (N_14045,N_13595,N_13269);
or U14046 (N_14046,N_13194,N_13331);
nor U14047 (N_14047,N_13657,N_13133);
nand U14048 (N_14048,N_13710,N_13683);
xnor U14049 (N_14049,N_13894,N_13878);
nand U14050 (N_14050,N_13159,N_13040);
and U14051 (N_14051,N_13430,N_13903);
or U14052 (N_14052,N_13089,N_13980);
nor U14053 (N_14053,N_13550,N_13921);
nor U14054 (N_14054,N_13959,N_13524);
nand U14055 (N_14055,N_13641,N_13371);
and U14056 (N_14056,N_13951,N_13152);
nor U14057 (N_14057,N_13006,N_13287);
xnor U14058 (N_14058,N_13324,N_13249);
or U14059 (N_14059,N_13644,N_13811);
nor U14060 (N_14060,N_13274,N_13702);
or U14061 (N_14061,N_13372,N_13294);
or U14062 (N_14062,N_13437,N_13614);
and U14063 (N_14063,N_13964,N_13858);
xor U14064 (N_14064,N_13869,N_13938);
or U14065 (N_14065,N_13983,N_13362);
xnor U14066 (N_14066,N_13631,N_13902);
and U14067 (N_14067,N_13696,N_13950);
xnor U14068 (N_14068,N_13017,N_13030);
nor U14069 (N_14069,N_13927,N_13303);
and U14070 (N_14070,N_13241,N_13230);
xor U14071 (N_14071,N_13297,N_13920);
and U14072 (N_14072,N_13092,N_13620);
xor U14073 (N_14073,N_13148,N_13621);
nand U14074 (N_14074,N_13117,N_13859);
xnor U14075 (N_14075,N_13380,N_13304);
xnor U14076 (N_14076,N_13863,N_13387);
xor U14077 (N_14077,N_13658,N_13554);
and U14078 (N_14078,N_13049,N_13892);
nor U14079 (N_14079,N_13744,N_13190);
or U14080 (N_14080,N_13697,N_13023);
or U14081 (N_14081,N_13642,N_13491);
or U14082 (N_14082,N_13507,N_13342);
nand U14083 (N_14083,N_13896,N_13399);
nand U14084 (N_14084,N_13748,N_13666);
and U14085 (N_14085,N_13397,N_13532);
nor U14086 (N_14086,N_13982,N_13637);
nor U14087 (N_14087,N_13754,N_13058);
and U14088 (N_14088,N_13967,N_13296);
xor U14089 (N_14089,N_13746,N_13700);
xnor U14090 (N_14090,N_13953,N_13170);
and U14091 (N_14091,N_13600,N_13119);
xor U14092 (N_14092,N_13025,N_13822);
and U14093 (N_14093,N_13501,N_13413);
and U14094 (N_14094,N_13623,N_13229);
nor U14095 (N_14095,N_13057,N_13165);
or U14096 (N_14096,N_13479,N_13618);
or U14097 (N_14097,N_13599,N_13468);
and U14098 (N_14098,N_13319,N_13584);
and U14099 (N_14099,N_13143,N_13734);
nor U14100 (N_14100,N_13651,N_13013);
or U14101 (N_14101,N_13062,N_13374);
and U14102 (N_14102,N_13745,N_13779);
xor U14103 (N_14103,N_13610,N_13617);
and U14104 (N_14104,N_13952,N_13008);
nand U14105 (N_14105,N_13555,N_13227);
nand U14106 (N_14106,N_13984,N_13087);
nor U14107 (N_14107,N_13794,N_13765);
nand U14108 (N_14108,N_13708,N_13003);
or U14109 (N_14109,N_13312,N_13034);
xor U14110 (N_14110,N_13290,N_13237);
nand U14111 (N_14111,N_13091,N_13922);
and U14112 (N_14112,N_13277,N_13455);
or U14113 (N_14113,N_13791,N_13458);
and U14114 (N_14114,N_13865,N_13690);
xnor U14115 (N_14115,N_13031,N_13574);
xor U14116 (N_14116,N_13815,N_13919);
nor U14117 (N_14117,N_13077,N_13925);
or U14118 (N_14118,N_13376,N_13820);
nand U14119 (N_14119,N_13454,N_13583);
nor U14120 (N_14120,N_13345,N_13002);
or U14121 (N_14121,N_13300,N_13207);
xor U14122 (N_14122,N_13024,N_13598);
or U14123 (N_14123,N_13720,N_13853);
xnor U14124 (N_14124,N_13019,N_13536);
nand U14125 (N_14125,N_13270,N_13814);
xor U14126 (N_14126,N_13064,N_13322);
and U14127 (N_14127,N_13381,N_13601);
xnor U14128 (N_14128,N_13793,N_13564);
xnor U14129 (N_14129,N_13818,N_13774);
nor U14130 (N_14130,N_13699,N_13966);
xor U14131 (N_14131,N_13906,N_13945);
and U14132 (N_14132,N_13428,N_13405);
or U14133 (N_14133,N_13572,N_13415);
or U14134 (N_14134,N_13560,N_13423);
and U14135 (N_14135,N_13351,N_13293);
xnor U14136 (N_14136,N_13101,N_13440);
nand U14137 (N_14137,N_13292,N_13149);
or U14138 (N_14138,N_13756,N_13168);
xor U14139 (N_14139,N_13299,N_13884);
or U14140 (N_14140,N_13893,N_13817);
xnor U14141 (N_14141,N_13496,N_13676);
nand U14142 (N_14142,N_13068,N_13418);
nor U14143 (N_14143,N_13862,N_13931);
nor U14144 (N_14144,N_13608,N_13934);
or U14145 (N_14145,N_13315,N_13050);
and U14146 (N_14146,N_13459,N_13732);
nand U14147 (N_14147,N_13653,N_13961);
nor U14148 (N_14148,N_13037,N_13924);
or U14149 (N_14149,N_13721,N_13219);
or U14150 (N_14150,N_13272,N_13460);
or U14151 (N_14151,N_13590,N_13047);
and U14152 (N_14152,N_13969,N_13016);
nor U14153 (N_14153,N_13786,N_13897);
and U14154 (N_14154,N_13729,N_13174);
and U14155 (N_14155,N_13861,N_13531);
xnor U14156 (N_14156,N_13962,N_13674);
or U14157 (N_14157,N_13226,N_13355);
and U14158 (N_14158,N_13263,N_13755);
or U14159 (N_14159,N_13273,N_13557);
and U14160 (N_14160,N_13807,N_13014);
nor U14161 (N_14161,N_13154,N_13974);
xnor U14162 (N_14162,N_13916,N_13346);
nand U14163 (N_14163,N_13402,N_13802);
and U14164 (N_14164,N_13481,N_13466);
nand U14165 (N_14165,N_13112,N_13752);
nor U14166 (N_14166,N_13494,N_13484);
xnor U14167 (N_14167,N_13205,N_13736);
nor U14168 (N_14168,N_13514,N_13010);
xnor U14169 (N_14169,N_13487,N_13787);
and U14170 (N_14170,N_13225,N_13761);
and U14171 (N_14171,N_13510,N_13912);
and U14172 (N_14172,N_13760,N_13360);
or U14173 (N_14173,N_13677,N_13076);
or U14174 (N_14174,N_13072,N_13026);
xor U14175 (N_14175,N_13622,N_13043);
xor U14176 (N_14176,N_13999,N_13289);
and U14177 (N_14177,N_13123,N_13840);
or U14178 (N_14178,N_13180,N_13832);
or U14179 (N_14179,N_13138,N_13410);
or U14180 (N_14180,N_13395,N_13389);
or U14181 (N_14181,N_13509,N_13976);
or U14182 (N_14182,N_13452,N_13094);
or U14183 (N_14183,N_13992,N_13711);
and U14184 (N_14184,N_13558,N_13940);
nor U14185 (N_14185,N_13989,N_13145);
xnor U14186 (N_14186,N_13692,N_13575);
nand U14187 (N_14187,N_13379,N_13831);
xor U14188 (N_14188,N_13053,N_13502);
xor U14189 (N_14189,N_13224,N_13255);
or U14190 (N_14190,N_13204,N_13877);
or U14191 (N_14191,N_13704,N_13171);
or U14192 (N_14192,N_13730,N_13682);
nand U14193 (N_14193,N_13963,N_13334);
and U14194 (N_14194,N_13933,N_13135);
nor U14195 (N_14195,N_13941,N_13740);
or U14196 (N_14196,N_13580,N_13100);
nand U14197 (N_14197,N_13107,N_13472);
or U14198 (N_14198,N_13321,N_13475);
nand U14199 (N_14199,N_13178,N_13517);
nand U14200 (N_14200,N_13626,N_13446);
nand U14201 (N_14201,N_13177,N_13088);
xnor U14202 (N_14202,N_13445,N_13160);
nand U14203 (N_14203,N_13500,N_13505);
or U14204 (N_14204,N_13672,N_13099);
and U14205 (N_14205,N_13797,N_13256);
nand U14206 (N_14206,N_13725,N_13607);
nor U14207 (N_14207,N_13689,N_13232);
or U14208 (N_14208,N_13427,N_13343);
nand U14209 (N_14209,N_13753,N_13563);
nand U14210 (N_14210,N_13664,N_13104);
or U14211 (N_14211,N_13714,N_13946);
xor U14212 (N_14212,N_13566,N_13639);
nor U14213 (N_14213,N_13038,N_13476);
or U14214 (N_14214,N_13553,N_13675);
xnor U14215 (N_14215,N_13471,N_13184);
nand U14216 (N_14216,N_13930,N_13115);
nand U14217 (N_14217,N_13882,N_13377);
or U14218 (N_14218,N_13162,N_13582);
and U14219 (N_14219,N_13680,N_13245);
nor U14220 (N_14220,N_13084,N_13490);
nor U14221 (N_14221,N_13552,N_13911);
nand U14222 (N_14222,N_13108,N_13235);
nor U14223 (N_14223,N_13246,N_13824);
nor U14224 (N_14224,N_13394,N_13495);
or U14225 (N_14225,N_13286,N_13383);
nor U14226 (N_14226,N_13977,N_13698);
nor U14227 (N_14227,N_13356,N_13095);
nand U14228 (N_14228,N_13202,N_13937);
xnor U14229 (N_14229,N_13126,N_13073);
xor U14230 (N_14230,N_13526,N_13450);
nand U14231 (N_14231,N_13492,N_13872);
nor U14232 (N_14232,N_13200,N_13763);
nor U14233 (N_14233,N_13265,N_13571);
nor U14234 (N_14234,N_13485,N_13910);
nand U14235 (N_14235,N_13731,N_13267);
xor U14236 (N_14236,N_13388,N_13662);
nand U14237 (N_14237,N_13705,N_13268);
xor U14238 (N_14238,N_13358,N_13109);
nor U14239 (N_14239,N_13520,N_13400);
and U14240 (N_14240,N_13193,N_13357);
or U14241 (N_14241,N_13596,N_13546);
and U14242 (N_14242,N_13396,N_13474);
or U14243 (N_14243,N_13142,N_13783);
xor U14244 (N_14244,N_13244,N_13463);
nand U14245 (N_14245,N_13619,N_13486);
or U14246 (N_14246,N_13764,N_13201);
or U14247 (N_14247,N_13291,N_13523);
or U14248 (N_14248,N_13578,N_13917);
nor U14249 (N_14249,N_13074,N_13602);
nand U14250 (N_14250,N_13960,N_13914);
or U14251 (N_14251,N_13443,N_13498);
nand U14252 (N_14252,N_13684,N_13991);
and U14253 (N_14253,N_13071,N_13363);
and U14254 (N_14254,N_13723,N_13703);
or U14255 (N_14255,N_13873,N_13747);
nor U14256 (N_14256,N_13134,N_13979);
or U14257 (N_14257,N_13067,N_13738);
or U14258 (N_14258,N_13968,N_13741);
xor U14259 (N_14259,N_13477,N_13885);
or U14260 (N_14260,N_13625,N_13654);
nand U14261 (N_14261,N_13965,N_13581);
nand U14262 (N_14262,N_13776,N_13172);
nand U14263 (N_14263,N_13281,N_13176);
nor U14264 (N_14264,N_13923,N_13904);
nand U14265 (N_14265,N_13789,N_13668);
nand U14266 (N_14266,N_13469,N_13295);
or U14267 (N_14267,N_13796,N_13775);
nor U14268 (N_14268,N_13570,N_13407);
and U14269 (N_14269,N_13627,N_13918);
xnor U14270 (N_14270,N_13988,N_13606);
or U14271 (N_14271,N_13929,N_13533);
or U14272 (N_14272,N_13144,N_13887);
or U14273 (N_14273,N_13522,N_13352);
xor U14274 (N_14274,N_13534,N_13915);
or U14275 (N_14275,N_13196,N_13181);
nor U14276 (N_14276,N_13425,N_13185);
or U14277 (N_14277,N_13280,N_13199);
nand U14278 (N_14278,N_13856,N_13766);
or U14279 (N_14279,N_13549,N_13260);
or U14280 (N_14280,N_13417,N_13628);
or U14281 (N_14281,N_13409,N_13022);
nor U14282 (N_14282,N_13886,N_13335);
and U14283 (N_14283,N_13480,N_13573);
or U14284 (N_14284,N_13715,N_13333);
or U14285 (N_14285,N_13800,N_13206);
or U14286 (N_14286,N_13613,N_13868);
and U14287 (N_14287,N_13792,N_13855);
or U14288 (N_14288,N_13799,N_13308);
nor U14289 (N_14289,N_13364,N_13384);
or U14290 (N_14290,N_13434,N_13949);
nor U14291 (N_14291,N_13585,N_13332);
nor U14292 (N_14292,N_13771,N_13130);
or U14293 (N_14293,N_13667,N_13883);
xor U14294 (N_14294,N_13743,N_13841);
or U14295 (N_14295,N_13932,N_13161);
or U14296 (N_14296,N_13768,N_13718);
nor U14297 (N_14297,N_13326,N_13650);
xnor U14298 (N_14298,N_13412,N_13124);
or U14299 (N_14299,N_13630,N_13944);
xnor U14300 (N_14300,N_13447,N_13102);
and U14301 (N_14301,N_13042,N_13239);
or U14302 (N_14302,N_13592,N_13876);
xnor U14303 (N_14303,N_13603,N_13347);
or U14304 (N_14304,N_13231,N_13661);
nor U14305 (N_14305,N_13182,N_13954);
nor U14306 (N_14306,N_13985,N_13990);
nand U14307 (N_14307,N_13691,N_13836);
or U14308 (N_14308,N_13640,N_13709);
nor U14309 (N_14309,N_13852,N_13189);
nand U14310 (N_14310,N_13591,N_13320);
xnor U14311 (N_14311,N_13995,N_13850);
and U14312 (N_14312,N_13438,N_13568);
and U14313 (N_14313,N_13323,N_13093);
and U14314 (N_14314,N_13139,N_13164);
or U14315 (N_14315,N_13879,N_13544);
nand U14316 (N_14316,N_13656,N_13449);
nand U14317 (N_14317,N_13328,N_13398);
nand U14318 (N_14318,N_13411,N_13939);
nor U14319 (N_14319,N_13825,N_13338);
and U14320 (N_14320,N_13513,N_13847);
and U14321 (N_14321,N_13118,N_13215);
xor U14322 (N_14322,N_13901,N_13359);
or U14323 (N_14323,N_13436,N_13724);
xnor U14324 (N_14324,N_13758,N_13027);
xor U14325 (N_14325,N_13616,N_13344);
xor U14326 (N_14326,N_13673,N_13096);
nor U14327 (N_14327,N_13365,N_13493);
and U14328 (N_14328,N_13947,N_13713);
xor U14329 (N_14329,N_13261,N_13426);
or U14330 (N_14330,N_13905,N_13781);
xnor U14331 (N_14331,N_13098,N_13431);
nor U14332 (N_14332,N_13997,N_13210);
or U14333 (N_14333,N_13382,N_13803);
nand U14334 (N_14334,N_13305,N_13624);
nand U14335 (N_14335,N_13712,N_13361);
nor U14336 (N_14336,N_13530,N_13066);
or U14337 (N_14337,N_13048,N_13685);
nor U14338 (N_14338,N_13634,N_13131);
nor U14339 (N_14339,N_13462,N_13233);
nor U14340 (N_14340,N_13259,N_13001);
and U14341 (N_14341,N_13442,N_13795);
nand U14342 (N_14342,N_13543,N_13061);
nand U14343 (N_14343,N_13111,N_13678);
or U14344 (N_14344,N_13083,N_13688);
xor U14345 (N_14345,N_13128,N_13565);
or U14346 (N_14346,N_13041,N_13898);
xor U14347 (N_14347,N_13167,N_13369);
and U14348 (N_14348,N_13593,N_13310);
or U14349 (N_14349,N_13508,N_13318);
xor U14350 (N_14350,N_13065,N_13354);
and U14351 (N_14351,N_13819,N_13701);
xnor U14352 (N_14352,N_13629,N_13806);
xnor U14353 (N_14353,N_13838,N_13253);
or U14354 (N_14354,N_13470,N_13551);
xnor U14355 (N_14355,N_13032,N_13867);
nand U14356 (N_14356,N_13081,N_13849);
xnor U14357 (N_14357,N_13538,N_13972);
xnor U14358 (N_14358,N_13742,N_13424);
nand U14359 (N_14359,N_13519,N_13012);
xnor U14360 (N_14360,N_13021,N_13928);
or U14361 (N_14361,N_13009,N_13136);
or U14362 (N_14362,N_13151,N_13186);
and U14363 (N_14363,N_13414,N_13957);
xnor U14364 (N_14364,N_13316,N_13638);
xor U14365 (N_14365,N_13218,N_13155);
nand U14366 (N_14366,N_13956,N_13429);
nor U14367 (N_14367,N_13288,N_13217);
xnor U14368 (N_14368,N_13611,N_13597);
xor U14369 (N_14369,N_13489,N_13282);
xnor U14370 (N_14370,N_13660,N_13039);
and U14371 (N_14371,N_13913,N_13577);
or U14372 (N_14372,N_13615,N_13998);
nand U14373 (N_14373,N_13579,N_13541);
or U14374 (N_14374,N_13604,N_13266);
nor U14375 (N_14375,N_13512,N_13843);
xor U14376 (N_14376,N_13521,N_13069);
or U14377 (N_14377,N_13453,N_13329);
nor U14378 (N_14378,N_13834,N_13432);
nand U14379 (N_14379,N_13045,N_13234);
xnor U14380 (N_14380,N_13527,N_13051);
and U14381 (N_14381,N_13238,N_13539);
or U14382 (N_14382,N_13173,N_13301);
nor U14383 (N_14383,N_13353,N_13279);
nand U14384 (N_14384,N_13845,N_13340);
nand U14385 (N_14385,N_13733,N_13191);
nand U14386 (N_14386,N_13408,N_13113);
and U14387 (N_14387,N_13813,N_13105);
nand U14388 (N_14388,N_13895,N_13576);
nand U14389 (N_14389,N_13907,N_13327);
nand U14390 (N_14390,N_13341,N_13116);
xor U14391 (N_14391,N_13350,N_13278);
nand U14392 (N_14392,N_13816,N_13970);
xnor U14393 (N_14393,N_13444,N_13007);
xnor U14394 (N_14394,N_13686,N_13015);
xnor U14395 (N_14395,N_13257,N_13749);
and U14396 (N_14396,N_13545,N_13647);
nor U14397 (N_14397,N_13864,N_13276);
and U14398 (N_14398,N_13140,N_13652);
or U14399 (N_14399,N_13996,N_13314);
nor U14400 (N_14400,N_13635,N_13254);
xor U14401 (N_14401,N_13285,N_13055);
nor U14402 (N_14402,N_13589,N_13837);
nor U14403 (N_14403,N_13243,N_13846);
xor U14404 (N_14404,N_13889,N_13125);
xnor U14405 (N_14405,N_13448,N_13080);
nor U14406 (N_14406,N_13419,N_13663);
nor U14407 (N_14407,N_13778,N_13659);
or U14408 (N_14408,N_13726,N_13420);
nand U14409 (N_14409,N_13063,N_13823);
nand U14410 (N_14410,N_13942,N_13456);
nand U14411 (N_14411,N_13537,N_13587);
nand U14412 (N_14412,N_13665,N_13679);
or U14413 (N_14413,N_13994,N_13441);
nor U14414 (N_14414,N_13208,N_13750);
or U14415 (N_14415,N_13782,N_13636);
nand U14416 (N_14416,N_13525,N_13075);
xor U14417 (N_14417,N_13567,N_13503);
nand U14418 (N_14418,N_13366,N_13605);
and U14419 (N_14419,N_13421,N_13146);
nor U14420 (N_14420,N_13298,N_13060);
nand U14421 (N_14421,N_13478,N_13569);
or U14422 (N_14422,N_13633,N_13223);
nor U14423 (N_14423,N_13857,N_13888);
nor U14424 (N_14424,N_13336,N_13317);
nand U14425 (N_14425,N_13461,N_13169);
nand U14426 (N_14426,N_13784,N_13540);
nor U14427 (N_14427,N_13805,N_13515);
xnor U14428 (N_14428,N_13406,N_13722);
and U14429 (N_14429,N_13390,N_13833);
xor U14430 (N_14430,N_13258,N_13044);
nor U14431 (N_14431,N_13046,N_13059);
and U14432 (N_14432,N_13214,N_13264);
or U14433 (N_14433,N_13375,N_13900);
or U14434 (N_14434,N_13349,N_13307);
and U14435 (N_14435,N_13054,N_13499);
or U14436 (N_14436,N_13588,N_13810);
and U14437 (N_14437,N_13777,N_13086);
and U14438 (N_14438,N_13719,N_13826);
xnor U14439 (N_14439,N_13284,N_13804);
xor U14440 (N_14440,N_13727,N_13975);
nor U14441 (N_14441,N_13890,N_13860);
or U14442 (N_14442,N_13029,N_13020);
and U14443 (N_14443,N_13211,N_13283);
or U14444 (N_14444,N_13669,N_13120);
or U14445 (N_14445,N_13958,N_13110);
nor U14446 (N_14446,N_13785,N_13767);
nor U14447 (N_14447,N_13348,N_13150);
nor U14448 (N_14448,N_13166,N_13391);
xor U14449 (N_14449,N_13197,N_13175);
nor U14450 (N_14450,N_13213,N_13609);
nor U14451 (N_14451,N_13504,N_13078);
nand U14452 (N_14452,N_13011,N_13561);
xor U14453 (N_14453,N_13482,N_13645);
nor U14454 (N_14454,N_13252,N_13018);
and U14455 (N_14455,N_13798,N_13559);
and U14456 (N_14456,N_13457,N_13473);
xnor U14457 (N_14457,N_13835,N_13250);
nand U14458 (N_14458,N_13114,N_13220);
and U14459 (N_14459,N_13986,N_13706);
nand U14460 (N_14460,N_13451,N_13236);
nand U14461 (N_14461,N_13228,N_13695);
nand U14462 (N_14462,N_13693,N_13156);
nor U14463 (N_14463,N_13655,N_13547);
or U14464 (N_14464,N_13936,N_13079);
nor U14465 (N_14465,N_13378,N_13404);
nor U14466 (N_14466,N_13247,N_13121);
and U14467 (N_14467,N_13971,N_13163);
nand U14468 (N_14468,N_13028,N_13271);
or U14469 (N_14469,N_13056,N_13612);
nor U14470 (N_14470,N_13212,N_13097);
nand U14471 (N_14471,N_13203,N_13337);
or U14472 (N_14472,N_13251,N_13839);
and U14473 (N_14473,N_13036,N_13594);
or U14474 (N_14474,N_13141,N_13103);
and U14475 (N_14475,N_13535,N_13851);
or U14476 (N_14476,N_13728,N_13033);
nand U14477 (N_14477,N_13401,N_13467);
nand U14478 (N_14478,N_13435,N_13198);
xnor U14479 (N_14479,N_13325,N_13828);
nor U14480 (N_14480,N_13529,N_13221);
and U14481 (N_14481,N_13821,N_13948);
nor U14482 (N_14482,N_13926,N_13506);
nor U14483 (N_14483,N_13070,N_13433);
xor U14484 (N_14484,N_13899,N_13880);
xnor U14485 (N_14485,N_13483,N_13874);
nand U14486 (N_14486,N_13000,N_13973);
nor U14487 (N_14487,N_13368,N_13157);
nor U14488 (N_14488,N_13739,N_13632);
nand U14489 (N_14489,N_13648,N_13306);
nor U14490 (N_14490,N_13187,N_13716);
and U14491 (N_14491,N_13707,N_13085);
nor U14492 (N_14492,N_13082,N_13681);
xnor U14493 (N_14493,N_13646,N_13367);
and U14494 (N_14494,N_13242,N_13179);
nor U14495 (N_14495,N_13192,N_13209);
xnor U14496 (N_14496,N_13370,N_13373);
or U14497 (N_14497,N_13978,N_13129);
and U14498 (N_14498,N_13386,N_13339);
xnor U14499 (N_14499,N_13330,N_13770);
nor U14500 (N_14500,N_13966,N_13681);
xnor U14501 (N_14501,N_13939,N_13916);
and U14502 (N_14502,N_13811,N_13657);
or U14503 (N_14503,N_13756,N_13266);
xor U14504 (N_14504,N_13433,N_13254);
xor U14505 (N_14505,N_13012,N_13861);
nor U14506 (N_14506,N_13723,N_13821);
xor U14507 (N_14507,N_13283,N_13545);
nand U14508 (N_14508,N_13789,N_13759);
or U14509 (N_14509,N_13059,N_13396);
or U14510 (N_14510,N_13704,N_13163);
or U14511 (N_14511,N_13191,N_13087);
xnor U14512 (N_14512,N_13604,N_13479);
nor U14513 (N_14513,N_13135,N_13067);
xor U14514 (N_14514,N_13069,N_13601);
nor U14515 (N_14515,N_13415,N_13120);
or U14516 (N_14516,N_13246,N_13196);
nand U14517 (N_14517,N_13871,N_13339);
or U14518 (N_14518,N_13824,N_13425);
xor U14519 (N_14519,N_13480,N_13738);
or U14520 (N_14520,N_13829,N_13551);
and U14521 (N_14521,N_13839,N_13198);
nor U14522 (N_14522,N_13594,N_13096);
and U14523 (N_14523,N_13523,N_13220);
xor U14524 (N_14524,N_13738,N_13823);
nand U14525 (N_14525,N_13212,N_13239);
nor U14526 (N_14526,N_13408,N_13960);
nand U14527 (N_14527,N_13696,N_13413);
nor U14528 (N_14528,N_13172,N_13110);
nor U14529 (N_14529,N_13317,N_13379);
xnor U14530 (N_14530,N_13495,N_13967);
or U14531 (N_14531,N_13063,N_13054);
or U14532 (N_14532,N_13505,N_13906);
and U14533 (N_14533,N_13774,N_13043);
and U14534 (N_14534,N_13597,N_13717);
and U14535 (N_14535,N_13569,N_13846);
nor U14536 (N_14536,N_13885,N_13582);
nor U14537 (N_14537,N_13368,N_13064);
nand U14538 (N_14538,N_13040,N_13963);
nor U14539 (N_14539,N_13174,N_13431);
nor U14540 (N_14540,N_13540,N_13624);
xnor U14541 (N_14541,N_13585,N_13101);
or U14542 (N_14542,N_13834,N_13934);
nor U14543 (N_14543,N_13583,N_13283);
and U14544 (N_14544,N_13168,N_13785);
or U14545 (N_14545,N_13652,N_13046);
nand U14546 (N_14546,N_13685,N_13010);
or U14547 (N_14547,N_13800,N_13531);
or U14548 (N_14548,N_13667,N_13531);
or U14549 (N_14549,N_13698,N_13107);
or U14550 (N_14550,N_13566,N_13627);
nor U14551 (N_14551,N_13746,N_13255);
nor U14552 (N_14552,N_13881,N_13036);
and U14553 (N_14553,N_13565,N_13829);
or U14554 (N_14554,N_13205,N_13772);
nand U14555 (N_14555,N_13387,N_13834);
or U14556 (N_14556,N_13065,N_13735);
or U14557 (N_14557,N_13893,N_13985);
nor U14558 (N_14558,N_13357,N_13767);
xor U14559 (N_14559,N_13456,N_13538);
xnor U14560 (N_14560,N_13743,N_13279);
or U14561 (N_14561,N_13421,N_13038);
xor U14562 (N_14562,N_13153,N_13335);
nand U14563 (N_14563,N_13981,N_13853);
nor U14564 (N_14564,N_13795,N_13028);
nand U14565 (N_14565,N_13595,N_13961);
nor U14566 (N_14566,N_13539,N_13232);
nand U14567 (N_14567,N_13224,N_13623);
nand U14568 (N_14568,N_13914,N_13881);
nor U14569 (N_14569,N_13482,N_13527);
nand U14570 (N_14570,N_13789,N_13827);
or U14571 (N_14571,N_13865,N_13849);
and U14572 (N_14572,N_13307,N_13080);
and U14573 (N_14573,N_13256,N_13600);
xor U14574 (N_14574,N_13910,N_13259);
and U14575 (N_14575,N_13206,N_13236);
nand U14576 (N_14576,N_13635,N_13306);
nand U14577 (N_14577,N_13667,N_13012);
xnor U14578 (N_14578,N_13973,N_13345);
and U14579 (N_14579,N_13553,N_13485);
xnor U14580 (N_14580,N_13430,N_13266);
nor U14581 (N_14581,N_13883,N_13193);
and U14582 (N_14582,N_13621,N_13054);
nor U14583 (N_14583,N_13448,N_13669);
nand U14584 (N_14584,N_13637,N_13814);
nor U14585 (N_14585,N_13928,N_13439);
nand U14586 (N_14586,N_13800,N_13710);
nor U14587 (N_14587,N_13564,N_13149);
and U14588 (N_14588,N_13578,N_13767);
and U14589 (N_14589,N_13071,N_13141);
xor U14590 (N_14590,N_13214,N_13891);
nand U14591 (N_14591,N_13580,N_13247);
xor U14592 (N_14592,N_13114,N_13573);
or U14593 (N_14593,N_13131,N_13276);
and U14594 (N_14594,N_13351,N_13020);
and U14595 (N_14595,N_13073,N_13889);
or U14596 (N_14596,N_13508,N_13335);
xor U14597 (N_14597,N_13760,N_13152);
nand U14598 (N_14598,N_13075,N_13244);
nand U14599 (N_14599,N_13607,N_13596);
and U14600 (N_14600,N_13112,N_13155);
nor U14601 (N_14601,N_13994,N_13737);
or U14602 (N_14602,N_13578,N_13664);
xnor U14603 (N_14603,N_13703,N_13705);
nor U14604 (N_14604,N_13457,N_13090);
nor U14605 (N_14605,N_13845,N_13036);
or U14606 (N_14606,N_13093,N_13555);
nor U14607 (N_14607,N_13863,N_13105);
nor U14608 (N_14608,N_13905,N_13153);
or U14609 (N_14609,N_13172,N_13614);
and U14610 (N_14610,N_13251,N_13106);
nor U14611 (N_14611,N_13914,N_13980);
nor U14612 (N_14612,N_13215,N_13328);
nor U14613 (N_14613,N_13056,N_13699);
nor U14614 (N_14614,N_13307,N_13381);
and U14615 (N_14615,N_13487,N_13197);
and U14616 (N_14616,N_13534,N_13746);
nand U14617 (N_14617,N_13818,N_13740);
nand U14618 (N_14618,N_13043,N_13453);
nand U14619 (N_14619,N_13192,N_13865);
nand U14620 (N_14620,N_13924,N_13207);
and U14621 (N_14621,N_13668,N_13125);
or U14622 (N_14622,N_13376,N_13830);
or U14623 (N_14623,N_13607,N_13874);
nor U14624 (N_14624,N_13694,N_13983);
xnor U14625 (N_14625,N_13477,N_13163);
nand U14626 (N_14626,N_13530,N_13945);
nand U14627 (N_14627,N_13858,N_13540);
xnor U14628 (N_14628,N_13441,N_13178);
or U14629 (N_14629,N_13054,N_13473);
nand U14630 (N_14630,N_13692,N_13347);
or U14631 (N_14631,N_13483,N_13529);
and U14632 (N_14632,N_13774,N_13209);
nand U14633 (N_14633,N_13908,N_13596);
nor U14634 (N_14634,N_13199,N_13131);
nor U14635 (N_14635,N_13716,N_13878);
and U14636 (N_14636,N_13156,N_13147);
nand U14637 (N_14637,N_13683,N_13718);
nor U14638 (N_14638,N_13823,N_13275);
xnor U14639 (N_14639,N_13420,N_13113);
xor U14640 (N_14640,N_13312,N_13968);
xnor U14641 (N_14641,N_13329,N_13240);
or U14642 (N_14642,N_13969,N_13059);
or U14643 (N_14643,N_13854,N_13155);
nand U14644 (N_14644,N_13044,N_13049);
nor U14645 (N_14645,N_13774,N_13977);
xor U14646 (N_14646,N_13831,N_13198);
xnor U14647 (N_14647,N_13751,N_13908);
and U14648 (N_14648,N_13786,N_13031);
nand U14649 (N_14649,N_13132,N_13666);
and U14650 (N_14650,N_13939,N_13749);
and U14651 (N_14651,N_13497,N_13321);
xnor U14652 (N_14652,N_13572,N_13200);
and U14653 (N_14653,N_13677,N_13916);
or U14654 (N_14654,N_13318,N_13189);
and U14655 (N_14655,N_13943,N_13847);
nor U14656 (N_14656,N_13782,N_13615);
nand U14657 (N_14657,N_13674,N_13539);
or U14658 (N_14658,N_13471,N_13884);
nor U14659 (N_14659,N_13487,N_13067);
xor U14660 (N_14660,N_13182,N_13588);
nor U14661 (N_14661,N_13623,N_13707);
nand U14662 (N_14662,N_13942,N_13415);
xor U14663 (N_14663,N_13041,N_13182);
nand U14664 (N_14664,N_13887,N_13480);
or U14665 (N_14665,N_13719,N_13276);
nor U14666 (N_14666,N_13172,N_13239);
xnor U14667 (N_14667,N_13674,N_13706);
or U14668 (N_14668,N_13444,N_13547);
nand U14669 (N_14669,N_13019,N_13569);
xnor U14670 (N_14670,N_13653,N_13465);
nand U14671 (N_14671,N_13042,N_13067);
nand U14672 (N_14672,N_13980,N_13881);
xnor U14673 (N_14673,N_13835,N_13076);
and U14674 (N_14674,N_13874,N_13156);
or U14675 (N_14675,N_13943,N_13890);
and U14676 (N_14676,N_13211,N_13009);
nor U14677 (N_14677,N_13955,N_13799);
nor U14678 (N_14678,N_13440,N_13774);
or U14679 (N_14679,N_13138,N_13238);
nor U14680 (N_14680,N_13878,N_13640);
nand U14681 (N_14681,N_13408,N_13103);
nand U14682 (N_14682,N_13346,N_13448);
and U14683 (N_14683,N_13199,N_13641);
xor U14684 (N_14684,N_13049,N_13293);
xnor U14685 (N_14685,N_13147,N_13484);
and U14686 (N_14686,N_13651,N_13112);
nand U14687 (N_14687,N_13264,N_13789);
and U14688 (N_14688,N_13929,N_13337);
xnor U14689 (N_14689,N_13665,N_13526);
or U14690 (N_14690,N_13841,N_13233);
nor U14691 (N_14691,N_13820,N_13795);
xnor U14692 (N_14692,N_13860,N_13904);
and U14693 (N_14693,N_13052,N_13987);
nand U14694 (N_14694,N_13704,N_13658);
nor U14695 (N_14695,N_13906,N_13220);
and U14696 (N_14696,N_13050,N_13758);
or U14697 (N_14697,N_13637,N_13769);
and U14698 (N_14698,N_13307,N_13486);
nor U14699 (N_14699,N_13968,N_13635);
nor U14700 (N_14700,N_13547,N_13633);
and U14701 (N_14701,N_13588,N_13529);
nand U14702 (N_14702,N_13683,N_13298);
or U14703 (N_14703,N_13300,N_13512);
nor U14704 (N_14704,N_13418,N_13531);
nand U14705 (N_14705,N_13532,N_13643);
or U14706 (N_14706,N_13608,N_13629);
or U14707 (N_14707,N_13410,N_13519);
or U14708 (N_14708,N_13525,N_13193);
or U14709 (N_14709,N_13436,N_13639);
or U14710 (N_14710,N_13468,N_13215);
nand U14711 (N_14711,N_13616,N_13517);
or U14712 (N_14712,N_13187,N_13519);
xnor U14713 (N_14713,N_13137,N_13964);
xor U14714 (N_14714,N_13370,N_13279);
and U14715 (N_14715,N_13338,N_13856);
nand U14716 (N_14716,N_13527,N_13702);
or U14717 (N_14717,N_13637,N_13587);
or U14718 (N_14718,N_13690,N_13048);
nand U14719 (N_14719,N_13203,N_13980);
nand U14720 (N_14720,N_13082,N_13583);
nand U14721 (N_14721,N_13844,N_13538);
or U14722 (N_14722,N_13158,N_13545);
xor U14723 (N_14723,N_13677,N_13451);
or U14724 (N_14724,N_13740,N_13072);
xnor U14725 (N_14725,N_13184,N_13066);
nand U14726 (N_14726,N_13330,N_13203);
and U14727 (N_14727,N_13494,N_13645);
nor U14728 (N_14728,N_13641,N_13756);
nand U14729 (N_14729,N_13581,N_13032);
nand U14730 (N_14730,N_13959,N_13951);
or U14731 (N_14731,N_13667,N_13654);
and U14732 (N_14732,N_13064,N_13173);
xor U14733 (N_14733,N_13843,N_13600);
xor U14734 (N_14734,N_13562,N_13925);
nand U14735 (N_14735,N_13149,N_13513);
xnor U14736 (N_14736,N_13886,N_13319);
nand U14737 (N_14737,N_13351,N_13828);
and U14738 (N_14738,N_13699,N_13849);
nand U14739 (N_14739,N_13865,N_13966);
nor U14740 (N_14740,N_13870,N_13295);
or U14741 (N_14741,N_13151,N_13695);
nand U14742 (N_14742,N_13747,N_13020);
and U14743 (N_14743,N_13656,N_13429);
nand U14744 (N_14744,N_13289,N_13224);
xnor U14745 (N_14745,N_13676,N_13812);
nand U14746 (N_14746,N_13964,N_13506);
nand U14747 (N_14747,N_13252,N_13837);
nand U14748 (N_14748,N_13806,N_13340);
or U14749 (N_14749,N_13205,N_13512);
xor U14750 (N_14750,N_13333,N_13927);
nor U14751 (N_14751,N_13158,N_13965);
xnor U14752 (N_14752,N_13646,N_13907);
or U14753 (N_14753,N_13385,N_13382);
nand U14754 (N_14754,N_13748,N_13725);
xor U14755 (N_14755,N_13395,N_13313);
nor U14756 (N_14756,N_13767,N_13897);
or U14757 (N_14757,N_13187,N_13002);
nor U14758 (N_14758,N_13698,N_13844);
nor U14759 (N_14759,N_13407,N_13393);
and U14760 (N_14760,N_13055,N_13234);
nor U14761 (N_14761,N_13684,N_13089);
nand U14762 (N_14762,N_13720,N_13030);
and U14763 (N_14763,N_13016,N_13581);
nor U14764 (N_14764,N_13976,N_13595);
xor U14765 (N_14765,N_13103,N_13049);
nand U14766 (N_14766,N_13825,N_13859);
nand U14767 (N_14767,N_13155,N_13608);
xnor U14768 (N_14768,N_13654,N_13608);
nand U14769 (N_14769,N_13979,N_13678);
xor U14770 (N_14770,N_13110,N_13003);
and U14771 (N_14771,N_13013,N_13525);
nand U14772 (N_14772,N_13365,N_13069);
or U14773 (N_14773,N_13644,N_13692);
xor U14774 (N_14774,N_13527,N_13025);
nor U14775 (N_14775,N_13745,N_13118);
xnor U14776 (N_14776,N_13494,N_13214);
or U14777 (N_14777,N_13847,N_13077);
xnor U14778 (N_14778,N_13922,N_13862);
or U14779 (N_14779,N_13311,N_13224);
xnor U14780 (N_14780,N_13078,N_13251);
and U14781 (N_14781,N_13505,N_13741);
xor U14782 (N_14782,N_13283,N_13601);
xnor U14783 (N_14783,N_13133,N_13480);
or U14784 (N_14784,N_13634,N_13087);
and U14785 (N_14785,N_13767,N_13518);
and U14786 (N_14786,N_13522,N_13173);
or U14787 (N_14787,N_13755,N_13402);
nor U14788 (N_14788,N_13964,N_13205);
nor U14789 (N_14789,N_13877,N_13628);
nor U14790 (N_14790,N_13152,N_13586);
and U14791 (N_14791,N_13639,N_13717);
nand U14792 (N_14792,N_13939,N_13155);
or U14793 (N_14793,N_13119,N_13188);
and U14794 (N_14794,N_13180,N_13645);
xnor U14795 (N_14795,N_13974,N_13259);
or U14796 (N_14796,N_13678,N_13512);
nor U14797 (N_14797,N_13541,N_13137);
xnor U14798 (N_14798,N_13944,N_13701);
nand U14799 (N_14799,N_13582,N_13692);
nand U14800 (N_14800,N_13433,N_13672);
or U14801 (N_14801,N_13962,N_13811);
or U14802 (N_14802,N_13273,N_13640);
nand U14803 (N_14803,N_13135,N_13379);
xor U14804 (N_14804,N_13045,N_13694);
or U14805 (N_14805,N_13802,N_13573);
nand U14806 (N_14806,N_13515,N_13787);
and U14807 (N_14807,N_13265,N_13509);
and U14808 (N_14808,N_13432,N_13448);
or U14809 (N_14809,N_13380,N_13050);
nand U14810 (N_14810,N_13470,N_13766);
or U14811 (N_14811,N_13374,N_13741);
nor U14812 (N_14812,N_13901,N_13720);
nand U14813 (N_14813,N_13234,N_13591);
xnor U14814 (N_14814,N_13936,N_13594);
and U14815 (N_14815,N_13150,N_13623);
nor U14816 (N_14816,N_13855,N_13637);
nor U14817 (N_14817,N_13887,N_13140);
or U14818 (N_14818,N_13889,N_13959);
and U14819 (N_14819,N_13820,N_13743);
nor U14820 (N_14820,N_13539,N_13462);
nand U14821 (N_14821,N_13500,N_13099);
xor U14822 (N_14822,N_13683,N_13119);
nor U14823 (N_14823,N_13897,N_13694);
or U14824 (N_14824,N_13598,N_13409);
nand U14825 (N_14825,N_13422,N_13452);
and U14826 (N_14826,N_13782,N_13778);
nor U14827 (N_14827,N_13902,N_13006);
or U14828 (N_14828,N_13865,N_13084);
nor U14829 (N_14829,N_13298,N_13393);
xnor U14830 (N_14830,N_13362,N_13985);
and U14831 (N_14831,N_13036,N_13538);
xnor U14832 (N_14832,N_13401,N_13637);
nor U14833 (N_14833,N_13431,N_13609);
or U14834 (N_14834,N_13265,N_13291);
nand U14835 (N_14835,N_13418,N_13895);
nand U14836 (N_14836,N_13073,N_13282);
xor U14837 (N_14837,N_13700,N_13673);
and U14838 (N_14838,N_13304,N_13783);
and U14839 (N_14839,N_13143,N_13365);
and U14840 (N_14840,N_13064,N_13938);
and U14841 (N_14841,N_13409,N_13680);
nand U14842 (N_14842,N_13579,N_13405);
nand U14843 (N_14843,N_13885,N_13299);
xor U14844 (N_14844,N_13077,N_13034);
and U14845 (N_14845,N_13535,N_13239);
or U14846 (N_14846,N_13787,N_13594);
nand U14847 (N_14847,N_13630,N_13005);
nand U14848 (N_14848,N_13988,N_13948);
or U14849 (N_14849,N_13027,N_13286);
nand U14850 (N_14850,N_13300,N_13025);
or U14851 (N_14851,N_13190,N_13538);
nand U14852 (N_14852,N_13462,N_13574);
xnor U14853 (N_14853,N_13404,N_13086);
nand U14854 (N_14854,N_13306,N_13426);
nor U14855 (N_14855,N_13691,N_13794);
nand U14856 (N_14856,N_13251,N_13630);
nor U14857 (N_14857,N_13858,N_13029);
or U14858 (N_14858,N_13942,N_13536);
xor U14859 (N_14859,N_13256,N_13883);
nand U14860 (N_14860,N_13089,N_13358);
nand U14861 (N_14861,N_13612,N_13911);
or U14862 (N_14862,N_13214,N_13723);
and U14863 (N_14863,N_13802,N_13763);
xor U14864 (N_14864,N_13920,N_13498);
or U14865 (N_14865,N_13893,N_13234);
and U14866 (N_14866,N_13332,N_13231);
xor U14867 (N_14867,N_13647,N_13576);
xor U14868 (N_14868,N_13518,N_13657);
or U14869 (N_14869,N_13817,N_13206);
xnor U14870 (N_14870,N_13414,N_13917);
nand U14871 (N_14871,N_13141,N_13133);
and U14872 (N_14872,N_13573,N_13476);
nor U14873 (N_14873,N_13893,N_13242);
or U14874 (N_14874,N_13397,N_13529);
nor U14875 (N_14875,N_13128,N_13667);
xnor U14876 (N_14876,N_13015,N_13169);
nand U14877 (N_14877,N_13341,N_13085);
xnor U14878 (N_14878,N_13285,N_13417);
xor U14879 (N_14879,N_13360,N_13571);
and U14880 (N_14880,N_13373,N_13139);
nor U14881 (N_14881,N_13357,N_13342);
and U14882 (N_14882,N_13960,N_13760);
nor U14883 (N_14883,N_13972,N_13029);
nand U14884 (N_14884,N_13904,N_13423);
nor U14885 (N_14885,N_13708,N_13131);
xnor U14886 (N_14886,N_13972,N_13614);
and U14887 (N_14887,N_13198,N_13635);
xnor U14888 (N_14888,N_13443,N_13652);
nand U14889 (N_14889,N_13755,N_13712);
nand U14890 (N_14890,N_13013,N_13972);
nor U14891 (N_14891,N_13911,N_13455);
nor U14892 (N_14892,N_13722,N_13818);
nor U14893 (N_14893,N_13773,N_13872);
xnor U14894 (N_14894,N_13865,N_13809);
and U14895 (N_14895,N_13782,N_13113);
nand U14896 (N_14896,N_13367,N_13704);
xnor U14897 (N_14897,N_13697,N_13534);
and U14898 (N_14898,N_13835,N_13588);
and U14899 (N_14899,N_13245,N_13069);
nand U14900 (N_14900,N_13093,N_13251);
or U14901 (N_14901,N_13020,N_13813);
and U14902 (N_14902,N_13959,N_13794);
or U14903 (N_14903,N_13703,N_13345);
and U14904 (N_14904,N_13281,N_13275);
and U14905 (N_14905,N_13445,N_13199);
or U14906 (N_14906,N_13999,N_13528);
nor U14907 (N_14907,N_13798,N_13627);
xnor U14908 (N_14908,N_13960,N_13025);
and U14909 (N_14909,N_13299,N_13673);
or U14910 (N_14910,N_13300,N_13483);
or U14911 (N_14911,N_13889,N_13884);
xor U14912 (N_14912,N_13521,N_13989);
and U14913 (N_14913,N_13160,N_13575);
and U14914 (N_14914,N_13165,N_13210);
and U14915 (N_14915,N_13293,N_13383);
nor U14916 (N_14916,N_13281,N_13879);
nand U14917 (N_14917,N_13761,N_13781);
nand U14918 (N_14918,N_13552,N_13693);
or U14919 (N_14919,N_13108,N_13950);
or U14920 (N_14920,N_13602,N_13004);
or U14921 (N_14921,N_13419,N_13960);
xnor U14922 (N_14922,N_13744,N_13440);
nor U14923 (N_14923,N_13849,N_13157);
or U14924 (N_14924,N_13904,N_13700);
and U14925 (N_14925,N_13404,N_13991);
nor U14926 (N_14926,N_13993,N_13131);
nor U14927 (N_14927,N_13563,N_13328);
nor U14928 (N_14928,N_13759,N_13779);
nor U14929 (N_14929,N_13382,N_13742);
or U14930 (N_14930,N_13689,N_13640);
xnor U14931 (N_14931,N_13282,N_13633);
or U14932 (N_14932,N_13703,N_13916);
nor U14933 (N_14933,N_13815,N_13945);
or U14934 (N_14934,N_13195,N_13836);
nand U14935 (N_14935,N_13265,N_13746);
or U14936 (N_14936,N_13062,N_13828);
nand U14937 (N_14937,N_13793,N_13279);
and U14938 (N_14938,N_13095,N_13469);
or U14939 (N_14939,N_13642,N_13054);
nor U14940 (N_14940,N_13401,N_13732);
or U14941 (N_14941,N_13195,N_13498);
nand U14942 (N_14942,N_13686,N_13649);
or U14943 (N_14943,N_13261,N_13927);
nor U14944 (N_14944,N_13631,N_13549);
and U14945 (N_14945,N_13904,N_13032);
xnor U14946 (N_14946,N_13242,N_13436);
and U14947 (N_14947,N_13822,N_13856);
nand U14948 (N_14948,N_13035,N_13952);
nand U14949 (N_14949,N_13339,N_13054);
and U14950 (N_14950,N_13842,N_13747);
nand U14951 (N_14951,N_13097,N_13720);
or U14952 (N_14952,N_13070,N_13414);
xor U14953 (N_14953,N_13450,N_13030);
or U14954 (N_14954,N_13503,N_13241);
or U14955 (N_14955,N_13855,N_13626);
xnor U14956 (N_14956,N_13553,N_13060);
xor U14957 (N_14957,N_13002,N_13026);
nor U14958 (N_14958,N_13395,N_13250);
nor U14959 (N_14959,N_13707,N_13605);
and U14960 (N_14960,N_13475,N_13699);
and U14961 (N_14961,N_13602,N_13807);
nand U14962 (N_14962,N_13001,N_13796);
or U14963 (N_14963,N_13197,N_13975);
nand U14964 (N_14964,N_13753,N_13390);
nor U14965 (N_14965,N_13385,N_13296);
xor U14966 (N_14966,N_13591,N_13729);
and U14967 (N_14967,N_13814,N_13411);
nor U14968 (N_14968,N_13790,N_13093);
and U14969 (N_14969,N_13415,N_13612);
nand U14970 (N_14970,N_13181,N_13901);
nand U14971 (N_14971,N_13936,N_13890);
and U14972 (N_14972,N_13465,N_13783);
nand U14973 (N_14973,N_13536,N_13072);
nor U14974 (N_14974,N_13667,N_13377);
or U14975 (N_14975,N_13378,N_13289);
or U14976 (N_14976,N_13095,N_13577);
xnor U14977 (N_14977,N_13086,N_13598);
nand U14978 (N_14978,N_13114,N_13401);
xor U14979 (N_14979,N_13487,N_13438);
xnor U14980 (N_14980,N_13874,N_13637);
xnor U14981 (N_14981,N_13364,N_13085);
nand U14982 (N_14982,N_13800,N_13844);
xnor U14983 (N_14983,N_13157,N_13832);
nand U14984 (N_14984,N_13404,N_13370);
and U14985 (N_14985,N_13178,N_13194);
nor U14986 (N_14986,N_13257,N_13060);
or U14987 (N_14987,N_13288,N_13769);
xor U14988 (N_14988,N_13068,N_13060);
nor U14989 (N_14989,N_13700,N_13816);
or U14990 (N_14990,N_13383,N_13216);
and U14991 (N_14991,N_13966,N_13038);
or U14992 (N_14992,N_13926,N_13998);
xor U14993 (N_14993,N_13823,N_13210);
xnor U14994 (N_14994,N_13270,N_13611);
nand U14995 (N_14995,N_13377,N_13947);
xor U14996 (N_14996,N_13205,N_13266);
xor U14997 (N_14997,N_13356,N_13975);
nor U14998 (N_14998,N_13591,N_13661);
nand U14999 (N_14999,N_13200,N_13749);
and U15000 (N_15000,N_14840,N_14139);
nor U15001 (N_15001,N_14624,N_14220);
nand U15002 (N_15002,N_14989,N_14902);
or U15003 (N_15003,N_14424,N_14962);
nand U15004 (N_15004,N_14213,N_14505);
xnor U15005 (N_15005,N_14644,N_14049);
xor U15006 (N_15006,N_14948,N_14843);
and U15007 (N_15007,N_14630,N_14861);
nor U15008 (N_15008,N_14282,N_14390);
nand U15009 (N_15009,N_14541,N_14971);
nor U15010 (N_15010,N_14702,N_14090);
nor U15011 (N_15011,N_14946,N_14279);
and U15012 (N_15012,N_14781,N_14397);
xor U15013 (N_15013,N_14046,N_14918);
and U15014 (N_15014,N_14242,N_14799);
xor U15015 (N_15015,N_14006,N_14952);
nand U15016 (N_15016,N_14357,N_14637);
xor U15017 (N_15017,N_14504,N_14115);
xor U15018 (N_15018,N_14113,N_14267);
and U15019 (N_15019,N_14784,N_14371);
and U15020 (N_15020,N_14647,N_14565);
xor U15021 (N_15021,N_14980,N_14634);
or U15022 (N_15022,N_14848,N_14506);
xnor U15023 (N_15023,N_14523,N_14244);
xnor U15024 (N_15024,N_14804,N_14581);
and U15025 (N_15025,N_14414,N_14496);
nand U15026 (N_15026,N_14274,N_14193);
nor U15027 (N_15027,N_14407,N_14863);
or U15028 (N_15028,N_14502,N_14923);
nor U15029 (N_15029,N_14064,N_14803);
nand U15030 (N_15030,N_14806,N_14256);
nor U15031 (N_15031,N_14159,N_14105);
nand U15032 (N_15032,N_14755,N_14930);
xnor U15033 (N_15033,N_14034,N_14566);
xnor U15034 (N_15034,N_14199,N_14321);
nand U15035 (N_15035,N_14628,N_14188);
and U15036 (N_15036,N_14040,N_14073);
nand U15037 (N_15037,N_14104,N_14540);
or U15038 (N_15038,N_14751,N_14617);
and U15039 (N_15039,N_14068,N_14154);
nand U15040 (N_15040,N_14999,N_14698);
nor U15041 (N_15041,N_14223,N_14697);
nand U15042 (N_15042,N_14163,N_14347);
nor U15043 (N_15043,N_14680,N_14783);
nor U15044 (N_15044,N_14873,N_14607);
nand U15045 (N_15045,N_14036,N_14805);
or U15046 (N_15046,N_14706,N_14704);
and U15047 (N_15047,N_14892,N_14079);
nor U15048 (N_15048,N_14091,N_14016);
nor U15049 (N_15049,N_14968,N_14981);
xnor U15050 (N_15050,N_14658,N_14310);
nand U15051 (N_15051,N_14136,N_14820);
nor U15052 (N_15052,N_14531,N_14621);
nor U15053 (N_15053,N_14524,N_14395);
nand U15054 (N_15054,N_14828,N_14731);
nand U15055 (N_15055,N_14898,N_14983);
nand U15056 (N_15056,N_14536,N_14479);
nor U15057 (N_15057,N_14233,N_14998);
nand U15058 (N_15058,N_14945,N_14168);
nor U15059 (N_15059,N_14343,N_14782);
xnor U15060 (N_15060,N_14076,N_14430);
nor U15061 (N_15061,N_14421,N_14281);
xor U15062 (N_15062,N_14827,N_14956);
xnor U15063 (N_15063,N_14556,N_14004);
nor U15064 (N_15064,N_14285,N_14023);
nand U15065 (N_15065,N_14398,N_14676);
or U15066 (N_15066,N_14186,N_14675);
and U15067 (N_15067,N_14598,N_14082);
and U15068 (N_15068,N_14965,N_14450);
and U15069 (N_15069,N_14942,N_14544);
xor U15070 (N_15070,N_14775,N_14022);
and U15071 (N_15071,N_14974,N_14319);
xor U15072 (N_15072,N_14548,N_14694);
or U15073 (N_15073,N_14099,N_14575);
xnor U15074 (N_15074,N_14405,N_14530);
nor U15075 (N_15075,N_14570,N_14741);
xor U15076 (N_15076,N_14733,N_14916);
xnor U15077 (N_15077,N_14273,N_14060);
or U15078 (N_15078,N_14786,N_14175);
and U15079 (N_15079,N_14525,N_14486);
xor U15080 (N_15080,N_14609,N_14065);
xor U15081 (N_15081,N_14802,N_14287);
nand U15082 (N_15082,N_14846,N_14276);
nor U15083 (N_15083,N_14203,N_14976);
nor U15084 (N_15084,N_14101,N_14222);
or U15085 (N_15085,N_14423,N_14355);
nor U15086 (N_15086,N_14686,N_14173);
or U15087 (N_15087,N_14742,N_14312);
nor U15088 (N_15088,N_14263,N_14960);
nor U15089 (N_15089,N_14318,N_14042);
nor U15090 (N_15090,N_14917,N_14161);
or U15091 (N_15091,N_14257,N_14937);
or U15092 (N_15092,N_14869,N_14009);
nor U15093 (N_15093,N_14206,N_14472);
xor U15094 (N_15094,N_14176,N_14533);
and U15095 (N_15095,N_14526,N_14158);
or U15096 (N_15096,N_14798,N_14789);
and U15097 (N_15097,N_14765,N_14227);
nand U15098 (N_15098,N_14709,N_14850);
or U15099 (N_15099,N_14895,N_14514);
xnor U15100 (N_15100,N_14370,N_14773);
nor U15101 (N_15101,N_14132,N_14026);
nand U15102 (N_15102,N_14054,N_14857);
and U15103 (N_15103,N_14238,N_14084);
xnor U15104 (N_15104,N_14551,N_14237);
xor U15105 (N_15105,N_14756,N_14467);
or U15106 (N_15106,N_14547,N_14564);
nand U15107 (N_15107,N_14392,N_14074);
nand U15108 (N_15108,N_14679,N_14109);
xnor U15109 (N_15109,N_14305,N_14500);
nand U15110 (N_15110,N_14979,N_14627);
nor U15111 (N_15111,N_14126,N_14520);
nand U15112 (N_15112,N_14640,N_14604);
xor U15113 (N_15113,N_14954,N_14482);
or U15114 (N_15114,N_14182,N_14382);
or U15115 (N_15115,N_14134,N_14133);
or U15116 (N_15116,N_14164,N_14428);
nor U15117 (N_15117,N_14881,N_14476);
and U15118 (N_15118,N_14631,N_14934);
or U15119 (N_15119,N_14330,N_14075);
xnor U15120 (N_15120,N_14352,N_14183);
or U15121 (N_15121,N_14872,N_14118);
and U15122 (N_15122,N_14757,N_14668);
and U15123 (N_15123,N_14744,N_14247);
nand U15124 (N_15124,N_14125,N_14893);
nand U15125 (N_15125,N_14448,N_14130);
or U15126 (N_15126,N_14991,N_14859);
and U15127 (N_15127,N_14933,N_14599);
or U15128 (N_15128,N_14573,N_14653);
or U15129 (N_15129,N_14057,N_14453);
nor U15130 (N_15130,N_14290,N_14418);
nand U15131 (N_15131,N_14532,N_14995);
or U15132 (N_15132,N_14320,N_14822);
nor U15133 (N_15133,N_14089,N_14928);
or U15134 (N_15134,N_14224,N_14807);
xnor U15135 (N_15135,N_14762,N_14093);
nor U15136 (N_15136,N_14294,N_14334);
or U15137 (N_15137,N_14379,N_14791);
nor U15138 (N_15138,N_14816,N_14384);
or U15139 (N_15139,N_14162,N_14953);
nand U15140 (N_15140,N_14323,N_14100);
or U15141 (N_15141,N_14077,N_14205);
nand U15142 (N_15142,N_14568,N_14303);
nor U15143 (N_15143,N_14339,N_14521);
nor U15144 (N_15144,N_14584,N_14292);
and U15145 (N_15145,N_14550,N_14826);
xnor U15146 (N_15146,N_14411,N_14255);
or U15147 (N_15147,N_14179,N_14510);
xor U15148 (N_15148,N_14723,N_14272);
nor U15149 (N_15149,N_14880,N_14487);
nor U15150 (N_15150,N_14817,N_14906);
nor U15151 (N_15151,N_14024,N_14462);
nor U15152 (N_15152,N_14071,N_14335);
nand U15153 (N_15153,N_14813,N_14854);
and U15154 (N_15154,N_14660,N_14608);
xor U15155 (N_15155,N_14322,N_14864);
and U15156 (N_15156,N_14684,N_14777);
and U15157 (N_15157,N_14908,N_14473);
and U15158 (N_15158,N_14663,N_14459);
and U15159 (N_15159,N_14687,N_14830);
nor U15160 (N_15160,N_14410,N_14198);
xor U15161 (N_15161,N_14844,N_14885);
nand U15162 (N_15162,N_14468,N_14715);
nand U15163 (N_15163,N_14589,N_14248);
or U15164 (N_15164,N_14776,N_14127);
nand U15165 (N_15165,N_14221,N_14963);
or U15166 (N_15166,N_14094,N_14443);
nor U15167 (N_15167,N_14062,N_14020);
nor U15168 (N_15168,N_14085,N_14559);
and U15169 (N_15169,N_14216,N_14574);
or U15170 (N_15170,N_14420,N_14612);
nor U15171 (N_15171,N_14236,N_14416);
or U15172 (N_15172,N_14152,N_14920);
xnor U15173 (N_15173,N_14780,N_14011);
or U15174 (N_15174,N_14461,N_14157);
or U15175 (N_15175,N_14261,N_14674);
xnor U15176 (N_15176,N_14340,N_14047);
or U15177 (N_15177,N_14904,N_14717);
and U15178 (N_15178,N_14138,N_14571);
nor U15179 (N_15179,N_14485,N_14797);
xnor U15180 (N_15180,N_14265,N_14700);
xor U15181 (N_15181,N_14737,N_14795);
or U15182 (N_15182,N_14761,N_14309);
and U15183 (N_15183,N_14695,N_14240);
and U15184 (N_15184,N_14545,N_14311);
xnor U15185 (N_15185,N_14386,N_14650);
xnor U15186 (N_15186,N_14122,N_14929);
and U15187 (N_15187,N_14048,N_14790);
xor U15188 (N_15188,N_14033,N_14217);
nor U15189 (N_15189,N_14639,N_14897);
nor U15190 (N_15190,N_14317,N_14728);
nand U15191 (N_15191,N_14116,N_14483);
and U15192 (N_15192,N_14110,N_14388);
nand U15193 (N_15193,N_14160,N_14484);
nor U15194 (N_15194,N_14678,N_14189);
xor U15195 (N_15195,N_14764,N_14181);
nor U15196 (N_15196,N_14517,N_14909);
nand U15197 (N_15197,N_14345,N_14856);
nand U15198 (N_15198,N_14325,N_14901);
and U15199 (N_15199,N_14560,N_14452);
nand U15200 (N_15200,N_14529,N_14539);
nor U15201 (N_15201,N_14131,N_14470);
and U15202 (N_15202,N_14375,N_14996);
nand U15203 (N_15203,N_14595,N_14124);
or U15204 (N_15204,N_14800,N_14977);
nand U15205 (N_15205,N_14824,N_14554);
nor U15206 (N_15206,N_14839,N_14825);
xnor U15207 (N_15207,N_14625,N_14734);
xor U15208 (N_15208,N_14596,N_14249);
and U15209 (N_15209,N_14088,N_14787);
nand U15210 (N_15210,N_14368,N_14754);
xor U15211 (N_15211,N_14832,N_14030);
or U15212 (N_15212,N_14315,N_14886);
nor U15213 (N_15213,N_14950,N_14117);
and U15214 (N_15214,N_14391,N_14726);
and U15215 (N_15215,N_14597,N_14014);
xor U15216 (N_15216,N_14427,N_14264);
or U15217 (N_15217,N_14149,N_14618);
and U15218 (N_15218,N_14689,N_14810);
nand U15219 (N_15219,N_14936,N_14070);
nor U15220 (N_15220,N_14254,N_14210);
or U15221 (N_15221,N_14501,N_14739);
nor U15222 (N_15222,N_14356,N_14972);
nand U15223 (N_15223,N_14364,N_14150);
nand U15224 (N_15224,N_14600,N_14577);
nand U15225 (N_15225,N_14050,N_14767);
or U15226 (N_15226,N_14809,N_14446);
xnor U15227 (N_15227,N_14900,N_14636);
xor U15228 (N_15228,N_14727,N_14646);
nand U15229 (N_15229,N_14997,N_14835);
nand U15230 (N_15230,N_14590,N_14141);
or U15231 (N_15231,N_14447,N_14667);
nand U15232 (N_15232,N_14670,N_14387);
xnor U15233 (N_15233,N_14629,N_14449);
and U15234 (N_15234,N_14578,N_14092);
nor U15235 (N_15235,N_14927,N_14992);
nor U15236 (N_15236,N_14135,N_14415);
and U15237 (N_15237,N_14669,N_14400);
and U15238 (N_15238,N_14656,N_14383);
and U15239 (N_15239,N_14185,N_14019);
xor U15240 (N_15240,N_14569,N_14114);
and U15241 (N_15241,N_14284,N_14988);
nor U15242 (N_15242,N_14013,N_14747);
or U15243 (N_15243,N_14299,N_14711);
xnor U15244 (N_15244,N_14592,N_14978);
nor U15245 (N_15245,N_14729,N_14426);
nor U15246 (N_15246,N_14393,N_14402);
xnor U15247 (N_15247,N_14632,N_14984);
nand U15248 (N_15248,N_14177,N_14701);
xnor U15249 (N_15249,N_14353,N_14492);
and U15250 (N_15250,N_14337,N_14466);
nor U15251 (N_15251,N_14278,N_14774);
nor U15252 (N_15252,N_14812,N_14376);
nand U15253 (N_15253,N_14833,N_14507);
or U15254 (N_15254,N_14932,N_14855);
xnor U15255 (N_15255,N_14685,N_14987);
nor U15256 (N_15256,N_14601,N_14534);
or U15257 (N_15257,N_14202,N_14245);
xnor U15258 (N_15258,N_14419,N_14852);
xnor U15259 (N_15259,N_14041,N_14713);
or U15260 (N_15260,N_14377,N_14488);
nor U15261 (N_15261,N_14029,N_14921);
nand U15262 (N_15262,N_14753,N_14829);
nand U15263 (N_15263,N_14940,N_14061);
xnor U15264 (N_15264,N_14924,N_14563);
or U15265 (N_15265,N_14403,N_14912);
and U15266 (N_15266,N_14437,N_14329);
nand U15267 (N_15267,N_14170,N_14925);
and U15268 (N_15268,N_14032,N_14591);
or U15269 (N_15269,N_14435,N_14148);
nor U15270 (N_15270,N_14616,N_14553);
nor U15271 (N_15271,N_14858,N_14831);
and U15272 (N_15272,N_14288,N_14128);
and U15273 (N_15273,N_14230,N_14439);
and U15274 (N_15274,N_14301,N_14518);
and U15275 (N_15275,N_14688,N_14045);
xor U15276 (N_15276,N_14745,N_14259);
or U15277 (N_15277,N_14796,N_14588);
nor U15278 (N_15278,N_14635,N_14280);
nand U15279 (N_15279,N_14474,N_14973);
nor U15280 (N_15280,N_14404,N_14326);
xnor U15281 (N_15281,N_14365,N_14044);
nand U15282 (N_15282,N_14174,N_14772);
nor U15283 (N_15283,N_14622,N_14381);
or U15284 (N_15284,N_14253,N_14888);
and U15285 (N_15285,N_14313,N_14643);
nand U15286 (N_15286,N_14759,N_14958);
or U15287 (N_15287,N_14231,N_14884);
nor U15288 (N_15288,N_14102,N_14481);
nor U15289 (N_15289,N_14055,N_14673);
nand U15290 (N_15290,N_14095,N_14915);
xor U15291 (N_15291,N_14511,N_14655);
and U15292 (N_15292,N_14811,N_14519);
nor U15293 (N_15293,N_14362,N_14516);
or U15294 (N_15294,N_14870,N_14750);
nand U15295 (N_15295,N_14043,N_14196);
xnor U15296 (N_15296,N_14209,N_14666);
and U15297 (N_15297,N_14191,N_14620);
nand U15298 (N_15298,N_14769,N_14037);
and U15299 (N_15299,N_14982,N_14342);
xnor U15300 (N_15300,N_14192,N_14328);
or U15301 (N_15301,N_14211,N_14096);
and U15302 (N_15302,N_14718,N_14241);
nor U15303 (N_15303,N_14293,N_14059);
nor U15304 (N_15304,N_14296,N_14542);
xnor U15305 (N_15305,N_14779,N_14576);
xnor U15306 (N_15306,N_14178,N_14478);
and U15307 (N_15307,N_14583,N_14025);
or U15308 (N_15308,N_14513,N_14067);
nor U15309 (N_15309,N_14369,N_14106);
nand U15310 (N_15310,N_14166,N_14939);
and U15311 (N_15311,N_14010,N_14801);
nand U15312 (N_15312,N_14842,N_14367);
or U15313 (N_15313,N_14465,N_14103);
and U15314 (N_15314,N_14003,N_14585);
or U15315 (N_15315,N_14018,N_14012);
nand U15316 (N_15316,N_14072,N_14648);
and U15317 (N_15317,N_14732,N_14582);
and U15318 (N_15318,N_14808,N_14232);
or U15319 (N_15319,N_14911,N_14615);
and U15320 (N_15320,N_14868,N_14875);
and U15321 (N_15321,N_14794,N_14155);
xor U15322 (N_15322,N_14056,N_14137);
nor U15323 (N_15323,N_14926,N_14195);
xnor U15324 (N_15324,N_14306,N_14495);
nand U15325 (N_15325,N_14603,N_14957);
nor U15326 (N_15326,N_14611,N_14735);
or U15327 (N_15327,N_14683,N_14552);
or U15328 (N_15328,N_14749,N_14295);
nor U15329 (N_15329,N_14691,N_14063);
and U15330 (N_15330,N_14580,N_14112);
nor U15331 (N_15331,N_14538,N_14455);
and U15332 (N_15332,N_14699,N_14457);
nor U15333 (N_15333,N_14922,N_14144);
nand U15334 (N_15334,N_14165,N_14720);
and U15335 (N_15335,N_14746,N_14944);
and U15336 (N_15336,N_14184,N_14866);
and U15337 (N_15337,N_14119,N_14008);
xor U15338 (N_15338,N_14454,N_14360);
xnor U15339 (N_15339,N_14374,N_14587);
or U15340 (N_15340,N_14194,N_14899);
nor U15341 (N_15341,N_14234,N_14031);
nand U15342 (N_15342,N_14436,N_14664);
and U15343 (N_15343,N_14494,N_14823);
nand U15344 (N_15344,N_14270,N_14406);
and U15345 (N_15345,N_14187,N_14662);
nor U15346 (N_15346,N_14725,N_14000);
and U15347 (N_15347,N_14266,N_14693);
xnor U15348 (N_15348,N_14425,N_14949);
nor U15349 (N_15349,N_14432,N_14017);
xnor U15350 (N_15350,N_14336,N_14304);
xor U15351 (N_15351,N_14308,N_14298);
and U15352 (N_15352,N_14681,N_14878);
or U15353 (N_15353,N_14503,N_14409);
and U15354 (N_15354,N_14887,N_14417);
nor U15355 (N_15355,N_14834,N_14277);
nor U15356 (N_15356,N_14359,N_14378);
nor U15357 (N_15357,N_14002,N_14035);
and U15358 (N_15358,N_14366,N_14324);
nor U15359 (N_15359,N_14412,N_14275);
nor U15360 (N_15360,N_14258,N_14225);
or U15361 (N_15361,N_14204,N_14349);
nand U15362 (N_15362,N_14350,N_14837);
xnor U15363 (N_15363,N_14964,N_14431);
or U15364 (N_15364,N_14867,N_14229);
or U15365 (N_15365,N_14348,N_14219);
and U15366 (N_15366,N_14993,N_14120);
or U15367 (N_15367,N_14738,N_14760);
and U15368 (N_15368,N_14297,N_14730);
and U15369 (N_15369,N_14876,N_14172);
nand U15370 (N_15370,N_14586,N_14201);
and U15371 (N_15371,N_14849,N_14508);
xor U15372 (N_15372,N_14527,N_14385);
or U15373 (N_15373,N_14338,N_14879);
or U15374 (N_15374,N_14140,N_14951);
nor U15375 (N_15375,N_14327,N_14373);
and U15376 (N_15376,N_14705,N_14243);
or U15377 (N_15377,N_14907,N_14719);
xor U15378 (N_15378,N_14471,N_14086);
and U15379 (N_15379,N_14151,N_14792);
xor U15380 (N_15380,N_14399,N_14561);
and U15381 (N_15381,N_14708,N_14235);
xnor U15382 (N_15382,N_14053,N_14143);
or U15383 (N_15383,N_14358,N_14434);
or U15384 (N_15384,N_14847,N_14260);
nor U15385 (N_15385,N_14111,N_14558);
xor U15386 (N_15386,N_14543,N_14522);
or U15387 (N_15387,N_14252,N_14372);
xor U15388 (N_15388,N_14218,N_14671);
and U15389 (N_15389,N_14363,N_14793);
or U15390 (N_15390,N_14758,N_14905);
nand U15391 (N_15391,N_14696,N_14672);
xnor U15392 (N_15392,N_14712,N_14351);
nor U15393 (N_15393,N_14147,N_14959);
xor U15394 (N_15394,N_14475,N_14028);
or U15395 (N_15395,N_14642,N_14142);
or U15396 (N_15396,N_14943,N_14610);
nand U15397 (N_15397,N_14641,N_14722);
nand U15398 (N_15398,N_14682,N_14052);
xor U15399 (N_15399,N_14919,N_14557);
nand U15400 (N_15400,N_14931,N_14380);
xor U15401 (N_15401,N_14080,N_14903);
and U15402 (N_15402,N_14314,N_14066);
nand U15403 (N_15403,N_14562,N_14785);
or U15404 (N_15404,N_14354,N_14480);
nand U15405 (N_15405,N_14724,N_14572);
or U15406 (N_15406,N_14955,N_14489);
nor U15407 (N_15407,N_14845,N_14200);
xnor U15408 (N_15408,N_14967,N_14707);
or U15409 (N_15409,N_14768,N_14307);
or U15410 (N_15410,N_14442,N_14458);
and U15411 (N_15411,N_14528,N_14862);
and U15412 (N_15412,N_14877,N_14394);
and U15413 (N_15413,N_14771,N_14069);
nand U15414 (N_15414,N_14821,N_14251);
or U15415 (N_15415,N_14208,N_14078);
nand U15416 (N_15416,N_14081,N_14891);
nor U15417 (N_15417,N_14039,N_14770);
or U15418 (N_15418,N_14499,N_14645);
xnor U15419 (N_15419,N_14167,N_14910);
nor U15420 (N_15420,N_14605,N_14456);
or U15421 (N_15421,N_14422,N_14890);
xnor U15422 (N_15422,N_14537,N_14703);
and U15423 (N_15423,N_14512,N_14190);
nand U15424 (N_15424,N_14269,N_14108);
and U15425 (N_15425,N_14652,N_14654);
or U15426 (N_15426,N_14021,N_14291);
xor U15427 (N_15427,N_14638,N_14815);
or U15428 (N_15428,N_14752,N_14649);
nor U15429 (N_15429,N_14659,N_14567);
xor U15430 (N_15430,N_14626,N_14316);
or U15431 (N_15431,N_14129,N_14464);
nor U15432 (N_15432,N_14961,N_14440);
nand U15433 (N_15433,N_14994,N_14226);
or U15434 (N_15434,N_14361,N_14289);
nand U15435 (N_15435,N_14493,N_14246);
xnor U15436 (N_15436,N_14346,N_14438);
nor U15437 (N_15437,N_14123,N_14509);
or U15438 (N_15438,N_14740,N_14087);
xor U15439 (N_15439,N_14677,N_14491);
xor U15440 (N_15440,N_14874,N_14083);
and U15441 (N_15441,N_14549,N_14180);
nand U15442 (N_15442,N_14433,N_14990);
or U15443 (N_15443,N_14515,N_14214);
and U15444 (N_15444,N_14853,N_14896);
nor U15445 (N_15445,N_14710,N_14743);
or U15446 (N_15446,N_14286,N_14778);
or U15447 (N_15447,N_14935,N_14171);
nor U15448 (N_15448,N_14239,N_14207);
nor U15449 (N_15449,N_14250,N_14889);
xor U15450 (N_15450,N_14766,N_14146);
or U15451 (N_15451,N_14215,N_14300);
nand U15452 (N_15452,N_14692,N_14788);
and U15453 (N_15453,N_14107,N_14121);
or U15454 (N_15454,N_14763,N_14015);
nor U15455 (N_15455,N_14614,N_14005);
xnor U15456 (N_15456,N_14490,N_14001);
nand U15457 (N_15457,N_14593,N_14341);
nand U15458 (N_15458,N_14156,N_14714);
and U15459 (N_15459,N_14441,N_14651);
nor U15460 (N_15460,N_14058,N_14332);
and U15461 (N_15461,N_14871,N_14451);
xnor U15462 (N_15462,N_14413,N_14097);
xor U15463 (N_15463,N_14445,N_14098);
and U15464 (N_15464,N_14613,N_14819);
or U15465 (N_15465,N_14331,N_14665);
nor U15466 (N_15466,N_14283,N_14401);
xnor U15467 (N_15467,N_14623,N_14941);
nand U15468 (N_15468,N_14619,N_14721);
and U15469 (N_15469,N_14497,N_14302);
and U15470 (N_15470,N_14814,N_14027);
or U15471 (N_15471,N_14271,N_14579);
nor U15472 (N_15472,N_14546,N_14606);
nand U15473 (N_15473,N_14818,N_14836);
or U15474 (N_15474,N_14396,N_14555);
nor U15475 (N_15475,N_14633,N_14882);
xnor U15476 (N_15476,N_14038,N_14838);
and U15477 (N_15477,N_14716,N_14748);
nor U15478 (N_15478,N_14966,N_14736);
and U15479 (N_15479,N_14602,N_14947);
nand U15480 (N_15480,N_14268,N_14051);
or U15481 (N_15481,N_14262,N_14938);
nor U15482 (N_15482,N_14851,N_14970);
or U15483 (N_15483,N_14333,N_14894);
nand U15484 (N_15484,N_14477,N_14986);
nand U15485 (N_15485,N_14429,N_14408);
xor U15486 (N_15486,N_14153,N_14883);
nand U15487 (N_15487,N_14145,N_14169);
or U15488 (N_15488,N_14969,N_14228);
xor U15489 (N_15489,N_14535,N_14212);
or U15490 (N_15490,N_14460,N_14498);
nor U15491 (N_15491,N_14975,N_14661);
or U15492 (N_15492,N_14344,N_14197);
and U15493 (N_15493,N_14469,N_14657);
or U15494 (N_15494,N_14865,N_14913);
and U15495 (N_15495,N_14690,N_14594);
nor U15496 (N_15496,N_14914,N_14389);
nand U15497 (N_15497,N_14985,N_14860);
and U15498 (N_15498,N_14841,N_14463);
nor U15499 (N_15499,N_14007,N_14444);
nand U15500 (N_15500,N_14090,N_14328);
nand U15501 (N_15501,N_14900,N_14721);
or U15502 (N_15502,N_14293,N_14807);
or U15503 (N_15503,N_14851,N_14130);
nand U15504 (N_15504,N_14999,N_14279);
nand U15505 (N_15505,N_14826,N_14998);
xnor U15506 (N_15506,N_14730,N_14790);
and U15507 (N_15507,N_14679,N_14098);
or U15508 (N_15508,N_14556,N_14150);
nor U15509 (N_15509,N_14514,N_14054);
nand U15510 (N_15510,N_14272,N_14514);
and U15511 (N_15511,N_14063,N_14134);
and U15512 (N_15512,N_14284,N_14966);
nand U15513 (N_15513,N_14523,N_14162);
and U15514 (N_15514,N_14989,N_14396);
or U15515 (N_15515,N_14830,N_14816);
and U15516 (N_15516,N_14504,N_14035);
or U15517 (N_15517,N_14219,N_14639);
xor U15518 (N_15518,N_14433,N_14647);
nor U15519 (N_15519,N_14084,N_14758);
or U15520 (N_15520,N_14821,N_14142);
or U15521 (N_15521,N_14055,N_14144);
xnor U15522 (N_15522,N_14583,N_14831);
or U15523 (N_15523,N_14705,N_14416);
nor U15524 (N_15524,N_14111,N_14821);
or U15525 (N_15525,N_14087,N_14502);
nor U15526 (N_15526,N_14092,N_14845);
nand U15527 (N_15527,N_14724,N_14776);
nand U15528 (N_15528,N_14623,N_14654);
xnor U15529 (N_15529,N_14754,N_14855);
xnor U15530 (N_15530,N_14578,N_14907);
nand U15531 (N_15531,N_14703,N_14678);
xor U15532 (N_15532,N_14926,N_14839);
or U15533 (N_15533,N_14963,N_14456);
nor U15534 (N_15534,N_14380,N_14379);
nand U15535 (N_15535,N_14012,N_14111);
or U15536 (N_15536,N_14045,N_14059);
xor U15537 (N_15537,N_14240,N_14942);
xor U15538 (N_15538,N_14894,N_14062);
or U15539 (N_15539,N_14761,N_14495);
or U15540 (N_15540,N_14276,N_14982);
or U15541 (N_15541,N_14028,N_14459);
and U15542 (N_15542,N_14126,N_14568);
or U15543 (N_15543,N_14176,N_14211);
and U15544 (N_15544,N_14776,N_14425);
or U15545 (N_15545,N_14617,N_14170);
and U15546 (N_15546,N_14438,N_14347);
and U15547 (N_15547,N_14820,N_14006);
nand U15548 (N_15548,N_14972,N_14631);
and U15549 (N_15549,N_14491,N_14601);
or U15550 (N_15550,N_14381,N_14879);
and U15551 (N_15551,N_14148,N_14190);
nor U15552 (N_15552,N_14652,N_14706);
nand U15553 (N_15553,N_14850,N_14827);
and U15554 (N_15554,N_14565,N_14331);
and U15555 (N_15555,N_14083,N_14153);
and U15556 (N_15556,N_14571,N_14076);
nor U15557 (N_15557,N_14996,N_14754);
nand U15558 (N_15558,N_14734,N_14597);
nand U15559 (N_15559,N_14564,N_14458);
nor U15560 (N_15560,N_14775,N_14475);
nor U15561 (N_15561,N_14935,N_14963);
nor U15562 (N_15562,N_14803,N_14350);
nor U15563 (N_15563,N_14499,N_14137);
and U15564 (N_15564,N_14781,N_14873);
nand U15565 (N_15565,N_14025,N_14885);
xnor U15566 (N_15566,N_14418,N_14515);
nand U15567 (N_15567,N_14652,N_14623);
or U15568 (N_15568,N_14970,N_14425);
nor U15569 (N_15569,N_14728,N_14347);
or U15570 (N_15570,N_14837,N_14255);
xor U15571 (N_15571,N_14111,N_14549);
nand U15572 (N_15572,N_14689,N_14055);
and U15573 (N_15573,N_14985,N_14354);
nor U15574 (N_15574,N_14853,N_14823);
nand U15575 (N_15575,N_14743,N_14236);
nand U15576 (N_15576,N_14078,N_14513);
nand U15577 (N_15577,N_14915,N_14593);
nand U15578 (N_15578,N_14948,N_14904);
or U15579 (N_15579,N_14589,N_14836);
nor U15580 (N_15580,N_14542,N_14252);
nor U15581 (N_15581,N_14101,N_14907);
nor U15582 (N_15582,N_14783,N_14910);
or U15583 (N_15583,N_14371,N_14347);
xor U15584 (N_15584,N_14821,N_14648);
nor U15585 (N_15585,N_14787,N_14364);
or U15586 (N_15586,N_14297,N_14570);
nand U15587 (N_15587,N_14293,N_14528);
nand U15588 (N_15588,N_14361,N_14804);
or U15589 (N_15589,N_14568,N_14676);
and U15590 (N_15590,N_14747,N_14182);
nand U15591 (N_15591,N_14550,N_14447);
nand U15592 (N_15592,N_14174,N_14474);
and U15593 (N_15593,N_14827,N_14215);
nand U15594 (N_15594,N_14517,N_14499);
or U15595 (N_15595,N_14090,N_14847);
and U15596 (N_15596,N_14209,N_14682);
nor U15597 (N_15597,N_14605,N_14225);
and U15598 (N_15598,N_14984,N_14806);
nand U15599 (N_15599,N_14852,N_14892);
and U15600 (N_15600,N_14868,N_14225);
and U15601 (N_15601,N_14835,N_14548);
nand U15602 (N_15602,N_14472,N_14637);
nand U15603 (N_15603,N_14438,N_14513);
nor U15604 (N_15604,N_14212,N_14013);
xnor U15605 (N_15605,N_14742,N_14337);
and U15606 (N_15606,N_14562,N_14093);
and U15607 (N_15607,N_14771,N_14151);
xnor U15608 (N_15608,N_14526,N_14175);
and U15609 (N_15609,N_14383,N_14447);
nand U15610 (N_15610,N_14513,N_14899);
nor U15611 (N_15611,N_14680,N_14110);
and U15612 (N_15612,N_14125,N_14739);
xor U15613 (N_15613,N_14229,N_14052);
nand U15614 (N_15614,N_14651,N_14382);
and U15615 (N_15615,N_14284,N_14575);
and U15616 (N_15616,N_14493,N_14599);
or U15617 (N_15617,N_14243,N_14170);
and U15618 (N_15618,N_14588,N_14768);
xnor U15619 (N_15619,N_14364,N_14303);
xnor U15620 (N_15620,N_14093,N_14272);
xor U15621 (N_15621,N_14242,N_14818);
nor U15622 (N_15622,N_14673,N_14355);
and U15623 (N_15623,N_14121,N_14740);
or U15624 (N_15624,N_14844,N_14227);
xnor U15625 (N_15625,N_14833,N_14198);
or U15626 (N_15626,N_14272,N_14838);
xnor U15627 (N_15627,N_14322,N_14631);
and U15628 (N_15628,N_14311,N_14171);
and U15629 (N_15629,N_14678,N_14677);
nand U15630 (N_15630,N_14745,N_14224);
and U15631 (N_15631,N_14923,N_14455);
or U15632 (N_15632,N_14640,N_14122);
or U15633 (N_15633,N_14067,N_14975);
and U15634 (N_15634,N_14206,N_14763);
or U15635 (N_15635,N_14782,N_14792);
and U15636 (N_15636,N_14800,N_14092);
xnor U15637 (N_15637,N_14944,N_14601);
or U15638 (N_15638,N_14280,N_14682);
nand U15639 (N_15639,N_14948,N_14807);
nor U15640 (N_15640,N_14436,N_14867);
nor U15641 (N_15641,N_14923,N_14388);
nand U15642 (N_15642,N_14909,N_14902);
or U15643 (N_15643,N_14492,N_14773);
nand U15644 (N_15644,N_14984,N_14456);
and U15645 (N_15645,N_14710,N_14087);
nor U15646 (N_15646,N_14498,N_14664);
or U15647 (N_15647,N_14397,N_14700);
or U15648 (N_15648,N_14971,N_14049);
and U15649 (N_15649,N_14748,N_14303);
xnor U15650 (N_15650,N_14682,N_14758);
and U15651 (N_15651,N_14057,N_14178);
or U15652 (N_15652,N_14294,N_14802);
and U15653 (N_15653,N_14339,N_14032);
xor U15654 (N_15654,N_14350,N_14878);
xnor U15655 (N_15655,N_14022,N_14522);
xor U15656 (N_15656,N_14291,N_14952);
xnor U15657 (N_15657,N_14863,N_14768);
or U15658 (N_15658,N_14452,N_14879);
nand U15659 (N_15659,N_14823,N_14159);
xor U15660 (N_15660,N_14549,N_14803);
and U15661 (N_15661,N_14229,N_14615);
xor U15662 (N_15662,N_14145,N_14023);
nor U15663 (N_15663,N_14768,N_14861);
or U15664 (N_15664,N_14695,N_14117);
or U15665 (N_15665,N_14724,N_14564);
nor U15666 (N_15666,N_14210,N_14974);
nor U15667 (N_15667,N_14637,N_14036);
xnor U15668 (N_15668,N_14430,N_14585);
xnor U15669 (N_15669,N_14984,N_14630);
and U15670 (N_15670,N_14481,N_14478);
nand U15671 (N_15671,N_14279,N_14430);
nor U15672 (N_15672,N_14498,N_14780);
and U15673 (N_15673,N_14673,N_14670);
nand U15674 (N_15674,N_14743,N_14105);
and U15675 (N_15675,N_14869,N_14555);
or U15676 (N_15676,N_14553,N_14639);
xor U15677 (N_15677,N_14063,N_14927);
nor U15678 (N_15678,N_14416,N_14272);
xor U15679 (N_15679,N_14476,N_14299);
and U15680 (N_15680,N_14163,N_14349);
or U15681 (N_15681,N_14793,N_14364);
nor U15682 (N_15682,N_14422,N_14232);
xor U15683 (N_15683,N_14355,N_14327);
or U15684 (N_15684,N_14177,N_14725);
nand U15685 (N_15685,N_14154,N_14534);
or U15686 (N_15686,N_14727,N_14444);
and U15687 (N_15687,N_14792,N_14968);
or U15688 (N_15688,N_14295,N_14361);
nor U15689 (N_15689,N_14438,N_14758);
xnor U15690 (N_15690,N_14913,N_14171);
xnor U15691 (N_15691,N_14322,N_14693);
nand U15692 (N_15692,N_14623,N_14846);
xor U15693 (N_15693,N_14417,N_14943);
nand U15694 (N_15694,N_14020,N_14358);
xor U15695 (N_15695,N_14077,N_14995);
or U15696 (N_15696,N_14462,N_14165);
and U15697 (N_15697,N_14193,N_14708);
xor U15698 (N_15698,N_14479,N_14253);
xor U15699 (N_15699,N_14601,N_14375);
nor U15700 (N_15700,N_14906,N_14054);
or U15701 (N_15701,N_14784,N_14877);
nor U15702 (N_15702,N_14535,N_14825);
and U15703 (N_15703,N_14872,N_14885);
nand U15704 (N_15704,N_14369,N_14930);
nand U15705 (N_15705,N_14827,N_14046);
or U15706 (N_15706,N_14313,N_14842);
and U15707 (N_15707,N_14630,N_14635);
xnor U15708 (N_15708,N_14538,N_14084);
and U15709 (N_15709,N_14310,N_14617);
nand U15710 (N_15710,N_14913,N_14943);
nor U15711 (N_15711,N_14091,N_14089);
nor U15712 (N_15712,N_14003,N_14202);
or U15713 (N_15713,N_14651,N_14321);
and U15714 (N_15714,N_14128,N_14637);
nand U15715 (N_15715,N_14724,N_14645);
or U15716 (N_15716,N_14979,N_14352);
xnor U15717 (N_15717,N_14985,N_14438);
xor U15718 (N_15718,N_14044,N_14360);
nor U15719 (N_15719,N_14457,N_14547);
nor U15720 (N_15720,N_14615,N_14889);
xor U15721 (N_15721,N_14207,N_14793);
xnor U15722 (N_15722,N_14558,N_14232);
nand U15723 (N_15723,N_14582,N_14208);
nor U15724 (N_15724,N_14995,N_14187);
or U15725 (N_15725,N_14243,N_14873);
and U15726 (N_15726,N_14556,N_14840);
nand U15727 (N_15727,N_14945,N_14848);
nand U15728 (N_15728,N_14943,N_14892);
xor U15729 (N_15729,N_14006,N_14858);
nand U15730 (N_15730,N_14290,N_14931);
xor U15731 (N_15731,N_14564,N_14365);
nand U15732 (N_15732,N_14026,N_14720);
nand U15733 (N_15733,N_14545,N_14704);
nor U15734 (N_15734,N_14324,N_14358);
nor U15735 (N_15735,N_14136,N_14069);
and U15736 (N_15736,N_14998,N_14529);
xor U15737 (N_15737,N_14787,N_14075);
nand U15738 (N_15738,N_14503,N_14103);
nor U15739 (N_15739,N_14982,N_14375);
xnor U15740 (N_15740,N_14715,N_14518);
and U15741 (N_15741,N_14175,N_14402);
and U15742 (N_15742,N_14313,N_14041);
nand U15743 (N_15743,N_14143,N_14633);
and U15744 (N_15744,N_14791,N_14851);
nor U15745 (N_15745,N_14644,N_14903);
and U15746 (N_15746,N_14298,N_14134);
xnor U15747 (N_15747,N_14863,N_14595);
and U15748 (N_15748,N_14854,N_14738);
nand U15749 (N_15749,N_14976,N_14171);
or U15750 (N_15750,N_14998,N_14302);
or U15751 (N_15751,N_14078,N_14527);
and U15752 (N_15752,N_14897,N_14561);
or U15753 (N_15753,N_14274,N_14614);
nand U15754 (N_15754,N_14465,N_14985);
nor U15755 (N_15755,N_14202,N_14904);
or U15756 (N_15756,N_14929,N_14120);
nor U15757 (N_15757,N_14678,N_14629);
nand U15758 (N_15758,N_14889,N_14959);
nand U15759 (N_15759,N_14725,N_14250);
nor U15760 (N_15760,N_14913,N_14059);
or U15761 (N_15761,N_14119,N_14767);
and U15762 (N_15762,N_14836,N_14084);
or U15763 (N_15763,N_14460,N_14589);
and U15764 (N_15764,N_14841,N_14266);
nor U15765 (N_15765,N_14216,N_14043);
nand U15766 (N_15766,N_14605,N_14736);
or U15767 (N_15767,N_14979,N_14428);
nand U15768 (N_15768,N_14217,N_14976);
or U15769 (N_15769,N_14919,N_14825);
or U15770 (N_15770,N_14178,N_14395);
nand U15771 (N_15771,N_14317,N_14568);
and U15772 (N_15772,N_14807,N_14240);
or U15773 (N_15773,N_14688,N_14601);
and U15774 (N_15774,N_14292,N_14130);
xor U15775 (N_15775,N_14935,N_14172);
or U15776 (N_15776,N_14430,N_14710);
xor U15777 (N_15777,N_14192,N_14879);
and U15778 (N_15778,N_14894,N_14291);
xnor U15779 (N_15779,N_14490,N_14572);
nor U15780 (N_15780,N_14776,N_14958);
nand U15781 (N_15781,N_14768,N_14247);
xnor U15782 (N_15782,N_14278,N_14257);
xnor U15783 (N_15783,N_14519,N_14906);
nor U15784 (N_15784,N_14870,N_14009);
and U15785 (N_15785,N_14131,N_14654);
xnor U15786 (N_15786,N_14082,N_14492);
and U15787 (N_15787,N_14543,N_14011);
and U15788 (N_15788,N_14555,N_14611);
nand U15789 (N_15789,N_14299,N_14399);
xnor U15790 (N_15790,N_14536,N_14015);
and U15791 (N_15791,N_14680,N_14946);
xnor U15792 (N_15792,N_14540,N_14775);
nand U15793 (N_15793,N_14339,N_14592);
xor U15794 (N_15794,N_14530,N_14187);
or U15795 (N_15795,N_14392,N_14425);
nor U15796 (N_15796,N_14906,N_14121);
nand U15797 (N_15797,N_14219,N_14539);
and U15798 (N_15798,N_14305,N_14968);
and U15799 (N_15799,N_14759,N_14638);
nand U15800 (N_15800,N_14098,N_14109);
and U15801 (N_15801,N_14650,N_14981);
and U15802 (N_15802,N_14875,N_14357);
or U15803 (N_15803,N_14634,N_14012);
nand U15804 (N_15804,N_14890,N_14108);
nor U15805 (N_15805,N_14846,N_14119);
or U15806 (N_15806,N_14035,N_14898);
nor U15807 (N_15807,N_14130,N_14689);
nand U15808 (N_15808,N_14148,N_14438);
nand U15809 (N_15809,N_14569,N_14436);
and U15810 (N_15810,N_14497,N_14226);
xor U15811 (N_15811,N_14067,N_14663);
nand U15812 (N_15812,N_14551,N_14710);
nand U15813 (N_15813,N_14690,N_14670);
nand U15814 (N_15814,N_14115,N_14059);
nand U15815 (N_15815,N_14343,N_14929);
or U15816 (N_15816,N_14886,N_14013);
xnor U15817 (N_15817,N_14618,N_14866);
nand U15818 (N_15818,N_14683,N_14660);
nand U15819 (N_15819,N_14137,N_14547);
nor U15820 (N_15820,N_14417,N_14540);
and U15821 (N_15821,N_14285,N_14103);
or U15822 (N_15822,N_14913,N_14661);
nor U15823 (N_15823,N_14029,N_14120);
nor U15824 (N_15824,N_14977,N_14448);
or U15825 (N_15825,N_14777,N_14216);
or U15826 (N_15826,N_14798,N_14548);
and U15827 (N_15827,N_14874,N_14492);
or U15828 (N_15828,N_14656,N_14379);
xnor U15829 (N_15829,N_14926,N_14260);
nor U15830 (N_15830,N_14854,N_14573);
xor U15831 (N_15831,N_14307,N_14128);
nor U15832 (N_15832,N_14630,N_14001);
nor U15833 (N_15833,N_14372,N_14407);
or U15834 (N_15834,N_14061,N_14462);
or U15835 (N_15835,N_14061,N_14707);
nand U15836 (N_15836,N_14861,N_14908);
nor U15837 (N_15837,N_14802,N_14656);
or U15838 (N_15838,N_14953,N_14130);
xor U15839 (N_15839,N_14058,N_14974);
xnor U15840 (N_15840,N_14489,N_14253);
nand U15841 (N_15841,N_14932,N_14287);
nand U15842 (N_15842,N_14931,N_14838);
and U15843 (N_15843,N_14294,N_14078);
nand U15844 (N_15844,N_14589,N_14939);
and U15845 (N_15845,N_14820,N_14527);
xor U15846 (N_15846,N_14765,N_14450);
xor U15847 (N_15847,N_14930,N_14621);
nor U15848 (N_15848,N_14870,N_14738);
nand U15849 (N_15849,N_14924,N_14060);
nand U15850 (N_15850,N_14688,N_14414);
xnor U15851 (N_15851,N_14485,N_14417);
and U15852 (N_15852,N_14839,N_14373);
and U15853 (N_15853,N_14066,N_14840);
or U15854 (N_15854,N_14657,N_14865);
or U15855 (N_15855,N_14976,N_14400);
and U15856 (N_15856,N_14449,N_14251);
or U15857 (N_15857,N_14603,N_14136);
xor U15858 (N_15858,N_14282,N_14720);
or U15859 (N_15859,N_14635,N_14473);
xor U15860 (N_15860,N_14763,N_14157);
nor U15861 (N_15861,N_14048,N_14389);
nand U15862 (N_15862,N_14052,N_14719);
and U15863 (N_15863,N_14452,N_14213);
nor U15864 (N_15864,N_14340,N_14731);
and U15865 (N_15865,N_14769,N_14573);
or U15866 (N_15866,N_14398,N_14439);
nand U15867 (N_15867,N_14387,N_14694);
nand U15868 (N_15868,N_14458,N_14003);
and U15869 (N_15869,N_14048,N_14958);
and U15870 (N_15870,N_14359,N_14894);
xnor U15871 (N_15871,N_14774,N_14265);
and U15872 (N_15872,N_14129,N_14619);
nor U15873 (N_15873,N_14671,N_14024);
nor U15874 (N_15874,N_14636,N_14546);
or U15875 (N_15875,N_14975,N_14139);
and U15876 (N_15876,N_14598,N_14896);
xor U15877 (N_15877,N_14776,N_14722);
xnor U15878 (N_15878,N_14128,N_14517);
nor U15879 (N_15879,N_14192,N_14124);
nor U15880 (N_15880,N_14941,N_14123);
nand U15881 (N_15881,N_14483,N_14505);
and U15882 (N_15882,N_14632,N_14019);
nor U15883 (N_15883,N_14320,N_14803);
nand U15884 (N_15884,N_14407,N_14381);
nand U15885 (N_15885,N_14049,N_14464);
and U15886 (N_15886,N_14351,N_14826);
or U15887 (N_15887,N_14835,N_14790);
nand U15888 (N_15888,N_14176,N_14894);
nand U15889 (N_15889,N_14119,N_14512);
nand U15890 (N_15890,N_14337,N_14777);
or U15891 (N_15891,N_14093,N_14284);
or U15892 (N_15892,N_14795,N_14091);
or U15893 (N_15893,N_14321,N_14527);
or U15894 (N_15894,N_14402,N_14980);
nand U15895 (N_15895,N_14757,N_14784);
or U15896 (N_15896,N_14357,N_14081);
nand U15897 (N_15897,N_14288,N_14580);
nor U15898 (N_15898,N_14557,N_14055);
nand U15899 (N_15899,N_14316,N_14286);
and U15900 (N_15900,N_14360,N_14155);
or U15901 (N_15901,N_14938,N_14966);
or U15902 (N_15902,N_14469,N_14003);
and U15903 (N_15903,N_14864,N_14075);
and U15904 (N_15904,N_14700,N_14230);
nand U15905 (N_15905,N_14599,N_14420);
xnor U15906 (N_15906,N_14212,N_14441);
xnor U15907 (N_15907,N_14972,N_14876);
nand U15908 (N_15908,N_14138,N_14075);
or U15909 (N_15909,N_14353,N_14212);
nand U15910 (N_15910,N_14063,N_14301);
or U15911 (N_15911,N_14983,N_14907);
or U15912 (N_15912,N_14198,N_14922);
and U15913 (N_15913,N_14842,N_14266);
xnor U15914 (N_15914,N_14925,N_14131);
nor U15915 (N_15915,N_14848,N_14593);
nor U15916 (N_15916,N_14042,N_14253);
or U15917 (N_15917,N_14655,N_14792);
xor U15918 (N_15918,N_14331,N_14594);
nand U15919 (N_15919,N_14518,N_14382);
xnor U15920 (N_15920,N_14413,N_14383);
and U15921 (N_15921,N_14858,N_14889);
and U15922 (N_15922,N_14493,N_14102);
nand U15923 (N_15923,N_14328,N_14901);
xnor U15924 (N_15924,N_14827,N_14948);
nand U15925 (N_15925,N_14506,N_14370);
nand U15926 (N_15926,N_14103,N_14272);
and U15927 (N_15927,N_14088,N_14092);
or U15928 (N_15928,N_14482,N_14860);
xnor U15929 (N_15929,N_14719,N_14638);
xnor U15930 (N_15930,N_14324,N_14111);
nor U15931 (N_15931,N_14828,N_14378);
nor U15932 (N_15932,N_14632,N_14555);
xnor U15933 (N_15933,N_14640,N_14057);
nand U15934 (N_15934,N_14281,N_14406);
nand U15935 (N_15935,N_14136,N_14736);
or U15936 (N_15936,N_14477,N_14005);
and U15937 (N_15937,N_14310,N_14696);
nor U15938 (N_15938,N_14451,N_14456);
and U15939 (N_15939,N_14227,N_14075);
xnor U15940 (N_15940,N_14439,N_14787);
nand U15941 (N_15941,N_14593,N_14321);
xnor U15942 (N_15942,N_14552,N_14738);
and U15943 (N_15943,N_14440,N_14572);
or U15944 (N_15944,N_14782,N_14098);
and U15945 (N_15945,N_14119,N_14892);
or U15946 (N_15946,N_14516,N_14921);
nand U15947 (N_15947,N_14397,N_14337);
nand U15948 (N_15948,N_14637,N_14418);
xnor U15949 (N_15949,N_14377,N_14497);
and U15950 (N_15950,N_14448,N_14464);
nand U15951 (N_15951,N_14274,N_14925);
or U15952 (N_15952,N_14401,N_14782);
or U15953 (N_15953,N_14010,N_14632);
or U15954 (N_15954,N_14808,N_14914);
nor U15955 (N_15955,N_14603,N_14031);
or U15956 (N_15956,N_14671,N_14420);
and U15957 (N_15957,N_14090,N_14673);
and U15958 (N_15958,N_14153,N_14220);
nand U15959 (N_15959,N_14004,N_14200);
nor U15960 (N_15960,N_14827,N_14981);
nand U15961 (N_15961,N_14507,N_14116);
or U15962 (N_15962,N_14596,N_14880);
nor U15963 (N_15963,N_14263,N_14419);
nand U15964 (N_15964,N_14169,N_14265);
nand U15965 (N_15965,N_14504,N_14975);
xor U15966 (N_15966,N_14861,N_14806);
or U15967 (N_15967,N_14755,N_14036);
xnor U15968 (N_15968,N_14579,N_14569);
nor U15969 (N_15969,N_14202,N_14093);
xnor U15970 (N_15970,N_14517,N_14368);
or U15971 (N_15971,N_14235,N_14145);
and U15972 (N_15972,N_14084,N_14068);
nor U15973 (N_15973,N_14385,N_14375);
or U15974 (N_15974,N_14120,N_14581);
xnor U15975 (N_15975,N_14222,N_14910);
and U15976 (N_15976,N_14746,N_14522);
and U15977 (N_15977,N_14425,N_14282);
xor U15978 (N_15978,N_14114,N_14080);
and U15979 (N_15979,N_14715,N_14187);
and U15980 (N_15980,N_14868,N_14753);
and U15981 (N_15981,N_14841,N_14526);
nand U15982 (N_15982,N_14347,N_14318);
nand U15983 (N_15983,N_14452,N_14872);
xnor U15984 (N_15984,N_14701,N_14601);
nor U15985 (N_15985,N_14658,N_14346);
nor U15986 (N_15986,N_14705,N_14658);
nand U15987 (N_15987,N_14722,N_14383);
nor U15988 (N_15988,N_14459,N_14495);
nor U15989 (N_15989,N_14629,N_14811);
and U15990 (N_15990,N_14662,N_14104);
xnor U15991 (N_15991,N_14203,N_14302);
xor U15992 (N_15992,N_14402,N_14756);
and U15993 (N_15993,N_14367,N_14630);
xor U15994 (N_15994,N_14863,N_14908);
xor U15995 (N_15995,N_14404,N_14076);
xnor U15996 (N_15996,N_14033,N_14486);
nor U15997 (N_15997,N_14147,N_14422);
xnor U15998 (N_15998,N_14322,N_14750);
nor U15999 (N_15999,N_14163,N_14342);
nor U16000 (N_16000,N_15456,N_15294);
xnor U16001 (N_16001,N_15139,N_15233);
xor U16002 (N_16002,N_15940,N_15025);
or U16003 (N_16003,N_15527,N_15167);
nand U16004 (N_16004,N_15767,N_15994);
nor U16005 (N_16005,N_15726,N_15566);
or U16006 (N_16006,N_15946,N_15452);
nand U16007 (N_16007,N_15161,N_15772);
and U16008 (N_16008,N_15895,N_15819);
and U16009 (N_16009,N_15902,N_15311);
and U16010 (N_16010,N_15461,N_15255);
nor U16011 (N_16011,N_15427,N_15990);
and U16012 (N_16012,N_15251,N_15371);
nand U16013 (N_16013,N_15069,N_15288);
xnor U16014 (N_16014,N_15389,N_15567);
nand U16015 (N_16015,N_15221,N_15017);
nor U16016 (N_16016,N_15958,N_15220);
and U16017 (N_16017,N_15812,N_15876);
or U16018 (N_16018,N_15290,N_15103);
and U16019 (N_16019,N_15591,N_15287);
and U16020 (N_16020,N_15827,N_15367);
nand U16021 (N_16021,N_15935,N_15753);
nor U16022 (N_16022,N_15119,N_15628);
nor U16023 (N_16023,N_15655,N_15621);
and U16024 (N_16024,N_15576,N_15612);
nand U16025 (N_16025,N_15916,N_15387);
and U16026 (N_16026,N_15084,N_15455);
or U16027 (N_16027,N_15690,N_15085);
nand U16028 (N_16028,N_15260,N_15900);
or U16029 (N_16029,N_15128,N_15903);
nand U16030 (N_16030,N_15569,N_15337);
xnor U16031 (N_16031,N_15425,N_15875);
xnor U16032 (N_16032,N_15829,N_15604);
or U16033 (N_16033,N_15988,N_15140);
xor U16034 (N_16034,N_15402,N_15750);
nand U16035 (N_16035,N_15888,N_15626);
and U16036 (N_16036,N_15963,N_15265);
or U16037 (N_16037,N_15634,N_15667);
nor U16038 (N_16038,N_15151,N_15385);
nand U16039 (N_16039,N_15465,N_15633);
nor U16040 (N_16040,N_15196,N_15226);
nand U16041 (N_16041,N_15511,N_15577);
or U16042 (N_16042,N_15172,N_15152);
or U16043 (N_16043,N_15663,N_15163);
nor U16044 (N_16044,N_15516,N_15598);
xor U16045 (N_16045,N_15399,N_15378);
xnor U16046 (N_16046,N_15679,N_15477);
or U16047 (N_16047,N_15955,N_15973);
nor U16048 (N_16048,N_15227,N_15266);
and U16049 (N_16049,N_15885,N_15334);
nand U16050 (N_16050,N_15118,N_15354);
and U16051 (N_16051,N_15659,N_15929);
and U16052 (N_16052,N_15324,N_15507);
nor U16053 (N_16053,N_15045,N_15433);
nor U16054 (N_16054,N_15510,N_15018);
nand U16055 (N_16055,N_15966,N_15215);
nand U16056 (N_16056,N_15114,N_15107);
nand U16057 (N_16057,N_15780,N_15478);
nor U16058 (N_16058,N_15579,N_15432);
and U16059 (N_16059,N_15373,N_15609);
nor U16060 (N_16060,N_15559,N_15654);
nor U16061 (N_16061,N_15896,N_15155);
or U16062 (N_16062,N_15773,N_15382);
nand U16063 (N_16063,N_15438,N_15785);
and U16064 (N_16064,N_15380,N_15209);
nor U16065 (N_16065,N_15968,N_15436);
and U16066 (N_16066,N_15732,N_15312);
xor U16067 (N_16067,N_15999,N_15374);
or U16068 (N_16068,N_15586,N_15201);
and U16069 (N_16069,N_15719,N_15755);
xor U16070 (N_16070,N_15638,N_15415);
xor U16071 (N_16071,N_15470,N_15774);
xnor U16072 (N_16072,N_15141,N_15684);
nor U16073 (N_16073,N_15596,N_15820);
and U16074 (N_16074,N_15234,N_15906);
nor U16075 (N_16075,N_15713,N_15463);
nor U16076 (N_16076,N_15872,N_15942);
or U16077 (N_16077,N_15602,N_15693);
or U16078 (N_16078,N_15762,N_15049);
nor U16079 (N_16079,N_15351,N_15519);
nor U16080 (N_16080,N_15967,N_15701);
nor U16081 (N_16081,N_15618,N_15611);
nand U16082 (N_16082,N_15176,N_15008);
nand U16083 (N_16083,N_15318,N_15131);
xnor U16084 (N_16084,N_15802,N_15299);
nand U16085 (N_16085,N_15801,N_15570);
or U16086 (N_16086,N_15120,N_15460);
xnor U16087 (N_16087,N_15093,N_15745);
or U16088 (N_16088,N_15068,N_15995);
xor U16089 (N_16089,N_15959,N_15817);
xor U16090 (N_16090,N_15216,N_15147);
nor U16091 (N_16091,N_15664,N_15206);
xnor U16092 (N_16092,N_15178,N_15945);
and U16093 (N_16093,N_15855,N_15349);
xnor U16094 (N_16094,N_15353,N_15582);
and U16095 (N_16095,N_15081,N_15024);
nor U16096 (N_16096,N_15080,N_15866);
and U16097 (N_16097,N_15082,N_15286);
xor U16098 (N_16098,N_15962,N_15584);
nand U16099 (N_16099,N_15742,N_15744);
xnor U16100 (N_16100,N_15957,N_15792);
nand U16101 (N_16101,N_15270,N_15708);
or U16102 (N_16102,N_15170,N_15165);
xor U16103 (N_16103,N_15077,N_15471);
nand U16104 (N_16104,N_15256,N_15169);
nand U16105 (N_16105,N_15106,N_15149);
nor U16106 (N_16106,N_15394,N_15188);
xor U16107 (N_16107,N_15769,N_15211);
xor U16108 (N_16108,N_15052,N_15834);
nor U16109 (N_16109,N_15901,N_15859);
nand U16110 (N_16110,N_15558,N_15410);
or U16111 (N_16111,N_15295,N_15891);
nor U16112 (N_16112,N_15530,N_15273);
xnor U16113 (N_16113,N_15203,N_15243);
or U16114 (N_16114,N_15102,N_15258);
nor U16115 (N_16115,N_15696,N_15327);
nand U16116 (N_16116,N_15800,N_15662);
xnor U16117 (N_16117,N_15212,N_15113);
nor U16118 (N_16118,N_15056,N_15392);
or U16119 (N_16119,N_15884,N_15244);
nand U16120 (N_16120,N_15092,N_15445);
xnor U16121 (N_16121,N_15498,N_15706);
xor U16122 (N_16122,N_15756,N_15793);
or U16123 (N_16123,N_15549,N_15200);
nand U16124 (N_16124,N_15187,N_15036);
nor U16125 (N_16125,N_15557,N_15937);
or U16126 (N_16126,N_15849,N_15766);
nand U16127 (N_16127,N_15043,N_15926);
nor U16128 (N_16128,N_15006,N_15013);
and U16129 (N_16129,N_15741,N_15504);
nand U16130 (N_16130,N_15646,N_15649);
nand U16131 (N_16131,N_15457,N_15669);
xor U16132 (N_16132,N_15593,N_15112);
nand U16133 (N_16133,N_15019,N_15788);
nor U16134 (N_16134,N_15276,N_15225);
and U16135 (N_16135,N_15562,N_15279);
and U16136 (N_16136,N_15489,N_15466);
and U16137 (N_16137,N_15459,N_15403);
and U16138 (N_16138,N_15386,N_15365);
nand U16139 (N_16139,N_15987,N_15127);
or U16140 (N_16140,N_15871,N_15309);
xnor U16141 (N_16141,N_15998,N_15674);
nand U16142 (N_16142,N_15631,N_15641);
xor U16143 (N_16143,N_15997,N_15924);
xor U16144 (N_16144,N_15525,N_15429);
nand U16145 (N_16145,N_15217,N_15449);
or U16146 (N_16146,N_15850,N_15921);
and U16147 (N_16147,N_15556,N_15363);
or U16148 (N_16148,N_15978,N_15330);
and U16149 (N_16149,N_15236,N_15761);
and U16150 (N_16150,N_15032,N_15063);
nor U16151 (N_16151,N_15359,N_15135);
and U16152 (N_16152,N_15707,N_15199);
nand U16153 (N_16153,N_15893,N_15301);
nand U16154 (N_16154,N_15676,N_15880);
nor U16155 (N_16155,N_15914,N_15689);
or U16156 (N_16156,N_15985,N_15542);
nand U16157 (N_16157,N_15828,N_15458);
nand U16158 (N_16158,N_15191,N_15336);
or U16159 (N_16159,N_15691,N_15718);
or U16160 (N_16160,N_15600,N_15253);
nand U16161 (N_16161,N_15033,N_15765);
and U16162 (N_16162,N_15627,N_15796);
or U16163 (N_16163,N_15815,N_15160);
xnor U16164 (N_16164,N_15502,N_15908);
or U16165 (N_16165,N_15381,N_15551);
xnor U16166 (N_16166,N_15848,N_15541);
xor U16167 (N_16167,N_15061,N_15770);
and U16168 (N_16168,N_15954,N_15736);
nand U16169 (N_16169,N_15971,N_15364);
xnor U16170 (N_16170,N_15450,N_15682);
nor U16171 (N_16171,N_15144,N_15843);
nand U16172 (N_16172,N_15710,N_15038);
and U16173 (N_16173,N_15090,N_15768);
xor U16174 (N_16174,N_15347,N_15307);
nand U16175 (N_16175,N_15435,N_15687);
nor U16176 (N_16176,N_15305,N_15254);
or U16177 (N_16177,N_15317,N_15430);
or U16178 (N_16178,N_15976,N_15007);
nor U16179 (N_16179,N_15269,N_15874);
nor U16180 (N_16180,N_15821,N_15731);
or U16181 (N_16181,N_15192,N_15688);
nor U16182 (N_16182,N_15132,N_15300);
nor U16183 (N_16183,N_15372,N_15657);
or U16184 (N_16184,N_15016,N_15915);
nor U16185 (N_16185,N_15503,N_15931);
and U16186 (N_16186,N_15314,N_15514);
and U16187 (N_16187,N_15228,N_15845);
or U16188 (N_16188,N_15179,N_15614);
nor U16189 (N_16189,N_15520,N_15791);
xnor U16190 (N_16190,N_15292,N_15099);
nor U16191 (N_16191,N_15580,N_15224);
nand U16192 (N_16192,N_15238,N_15934);
or U16193 (N_16193,N_15360,N_15042);
or U16194 (N_16194,N_15062,N_15037);
xor U16195 (N_16195,N_15029,N_15974);
or U16196 (N_16196,N_15342,N_15775);
nor U16197 (N_16197,N_15705,N_15020);
and U16198 (N_16198,N_15677,N_15341);
nand U16199 (N_16199,N_15724,N_15095);
nor U16200 (N_16200,N_15248,N_15572);
nor U16201 (N_16201,N_15700,N_15804);
nand U16202 (N_16202,N_15441,N_15362);
nand U16203 (N_16203,N_15923,N_15345);
nand U16204 (N_16204,N_15001,N_15574);
nand U16205 (N_16205,N_15004,N_15488);
and U16206 (N_16206,N_15658,N_15535);
and U16207 (N_16207,N_15331,N_15428);
nor U16208 (N_16208,N_15421,N_15146);
xor U16209 (N_16209,N_15840,N_15259);
xnor U16210 (N_16210,N_15715,N_15492);
xnor U16211 (N_16211,N_15328,N_15501);
nand U16212 (N_16212,N_15297,N_15853);
nand U16213 (N_16213,N_15547,N_15332);
xor U16214 (N_16214,N_15599,N_15608);
or U16215 (N_16215,N_15247,N_15668);
xnor U16216 (N_16216,N_15518,N_15264);
or U16217 (N_16217,N_15133,N_15193);
nand U16218 (N_16218,N_15806,N_15473);
nor U16219 (N_16219,N_15182,N_15832);
or U16220 (N_16220,N_15422,N_15961);
nand U16221 (N_16221,N_15404,N_15833);
or U16222 (N_16222,N_15537,N_15747);
and U16223 (N_16223,N_15936,N_15407);
xor U16224 (N_16224,N_15740,N_15304);
xor U16225 (N_16225,N_15075,N_15350);
nand U16226 (N_16226,N_15920,N_15396);
nor U16227 (N_16227,N_15565,N_15078);
or U16228 (N_16228,N_15015,N_15048);
or U16229 (N_16229,N_15656,N_15469);
nor U16230 (N_16230,N_15245,N_15841);
nand U16231 (N_16231,N_15343,N_15219);
or U16232 (N_16232,N_15948,N_15794);
xnor U16233 (N_16233,N_15010,N_15623);
xnor U16234 (N_16234,N_15285,N_15100);
xnor U16235 (N_16235,N_15035,N_15733);
xnor U16236 (N_16236,N_15440,N_15088);
nand U16237 (N_16237,N_15922,N_15607);
nand U16238 (N_16238,N_15027,N_15298);
and U16239 (N_16239,N_15861,N_15698);
and U16240 (N_16240,N_15091,N_15130);
and U16241 (N_16241,N_15418,N_15323);
or U16242 (N_16242,N_15970,N_15413);
xor U16243 (N_16243,N_15969,N_15057);
and U16244 (N_16244,N_15252,N_15390);
or U16245 (N_16245,N_15695,N_15003);
nor U16246 (N_16246,N_15808,N_15417);
nand U16247 (N_16247,N_15158,N_15499);
nor U16248 (N_16248,N_15526,N_15122);
or U16249 (N_16249,N_15790,N_15678);
xnor U16250 (N_16250,N_15778,N_15814);
or U16251 (N_16251,N_15882,N_15272);
or U16252 (N_16252,N_15506,N_15560);
nand U16253 (N_16253,N_15239,N_15727);
nand U16254 (N_16254,N_15605,N_15751);
and U16255 (N_16255,N_15714,N_15065);
nor U16256 (N_16256,N_15748,N_15344);
or U16257 (N_16257,N_15860,N_15781);
xor U16258 (N_16258,N_15313,N_15447);
nor U16259 (N_16259,N_15493,N_15616);
and U16260 (N_16260,N_15391,N_15624);
nor U16261 (N_16261,N_15729,N_15643);
xnor U16262 (N_16262,N_15758,N_15864);
xor U16263 (N_16263,N_15284,N_15666);
and U16264 (N_16264,N_15865,N_15613);
or U16265 (N_16265,N_15097,N_15597);
nor U16266 (N_16266,N_15189,N_15280);
or U16267 (N_16267,N_15811,N_15379);
xnor U16268 (N_16268,N_15907,N_15975);
and U16269 (N_16269,N_15933,N_15564);
nand U16270 (N_16270,N_15759,N_15321);
xor U16271 (N_16271,N_15249,N_15303);
xor U16272 (N_16272,N_15156,N_15699);
or U16273 (N_16273,N_15494,N_15326);
xnor U16274 (N_16274,N_15476,N_15738);
nor U16275 (N_16275,N_15086,N_15947);
and U16276 (N_16276,N_15568,N_15070);
xnor U16277 (N_16277,N_15645,N_15355);
xor U16278 (N_16278,N_15480,N_15198);
nand U16279 (N_16279,N_15782,N_15316);
xor U16280 (N_16280,N_15870,N_15743);
and U16281 (N_16281,N_15980,N_15771);
nor U16282 (N_16282,N_15508,N_15873);
and U16283 (N_16283,N_15358,N_15983);
and U16284 (N_16284,N_15513,N_15944);
or U16285 (N_16285,N_15898,N_15322);
nor U16286 (N_16286,N_15938,N_15484);
xor U16287 (N_16287,N_15240,N_15237);
nand U16288 (N_16288,N_15137,N_15384);
and U16289 (N_16289,N_15683,N_15651);
or U16290 (N_16290,N_15777,N_15680);
nand U16291 (N_16291,N_15889,N_15482);
nor U16292 (N_16292,N_15992,N_15573);
nor U16293 (N_16293,N_15401,N_15487);
or U16294 (N_16294,N_15592,N_15515);
nand U16295 (N_16295,N_15746,N_15431);
xnor U16296 (N_16296,N_15474,N_15416);
and U16297 (N_16297,N_15340,N_15545);
nor U16298 (N_16298,N_15411,N_15606);
xor U16299 (N_16299,N_15125,N_15185);
or U16300 (N_16300,N_15022,N_15528);
nor U16301 (N_16301,N_15563,N_15356);
and U16302 (N_16302,N_15617,N_15282);
and U16303 (N_16303,N_15448,N_15670);
or U16304 (N_16304,N_15105,N_15712);
nor U16305 (N_16305,N_15619,N_15797);
xor U16306 (N_16306,N_15087,N_15293);
and U16307 (N_16307,N_15846,N_15171);
nor U16308 (N_16308,N_15660,N_15723);
or U16309 (N_16309,N_15405,N_15419);
xnor U16310 (N_16310,N_15055,N_15590);
nand U16311 (N_16311,N_15148,N_15752);
and U16312 (N_16312,N_15928,N_15485);
and U16313 (N_16313,N_15462,N_15021);
and U16314 (N_16314,N_15857,N_15074);
and U16315 (N_16315,N_15737,N_15177);
nor U16316 (N_16316,N_15338,N_15277);
nor U16317 (N_16317,N_15764,N_15325);
nand U16318 (N_16318,N_15468,N_15012);
and U16319 (N_16319,N_15868,N_15138);
xor U16320 (N_16320,N_15588,N_15539);
nor U16321 (N_16321,N_15129,N_15000);
nand U16322 (N_16322,N_15826,N_15686);
or U16323 (N_16323,N_15863,N_15296);
nand U16324 (N_16324,N_15939,N_15979);
xnor U16325 (N_16325,N_15960,N_15496);
nand U16326 (N_16326,N_15538,N_15058);
xnor U16327 (N_16327,N_15472,N_15420);
nand U16328 (N_16328,N_15630,N_15034);
xnor U16329 (N_16329,N_15175,N_15434);
nor U16330 (N_16330,N_15986,N_15205);
nor U16331 (N_16331,N_15809,N_15534);
or U16332 (N_16332,N_15366,N_15134);
or U16333 (N_16333,N_15877,N_15283);
nand U16334 (N_16334,N_15635,N_15375);
nor U16335 (N_16335,N_15453,N_15076);
nand U16336 (N_16336,N_15991,N_15716);
or U16337 (N_16337,N_15072,N_15544);
or U16338 (N_16338,N_15842,N_15704);
and U16339 (N_16339,N_15524,N_15319);
xor U16340 (N_16340,N_15483,N_15423);
nor U16341 (N_16341,N_15589,N_15500);
and U16342 (N_16342,N_15368,N_15208);
nand U16343 (N_16343,N_15642,N_15509);
xor U16344 (N_16344,N_15553,N_15536);
or U16345 (N_16345,N_15333,N_15951);
nor U16346 (N_16346,N_15028,N_15023);
or U16347 (N_16347,N_15867,N_15787);
nor U16348 (N_16348,N_15823,N_15972);
or U16349 (N_16349,N_15835,N_15444);
nand U16350 (N_16350,N_15879,N_15104);
xnor U16351 (N_16351,N_15847,N_15388);
nand U16352 (N_16352,N_15913,N_15490);
and U16353 (N_16353,N_15648,N_15681);
nor U16354 (N_16354,N_15281,N_15153);
nand U16355 (N_16355,N_15763,N_15862);
and U16356 (N_16356,N_15210,N_15836);
nor U16357 (N_16357,N_15442,N_15395);
nor U16358 (N_16358,N_15230,N_15703);
xor U16359 (N_16359,N_15625,N_15202);
and U16360 (N_16360,N_15308,N_15552);
or U16361 (N_16361,N_15143,N_15533);
xor U16362 (N_16362,N_15250,N_15734);
xor U16363 (N_16363,N_15692,N_15181);
and U16364 (N_16364,N_15858,N_15014);
and U16365 (N_16365,N_15094,N_15117);
xor U16366 (N_16366,N_15917,N_15523);
nand U16367 (N_16367,N_15408,N_15571);
or U16368 (N_16368,N_15339,N_15813);
and U16369 (N_16369,N_15517,N_15886);
nand U16370 (N_16370,N_15702,N_15798);
nor U16371 (N_16371,N_15952,N_15096);
nand U16372 (N_16372,N_15838,N_15451);
nand U16373 (N_16373,N_15044,N_15894);
and U16374 (N_16374,N_15241,N_15041);
nor U16375 (N_16375,N_15910,N_15110);
and U16376 (N_16376,N_15807,N_15174);
xnor U16377 (N_16377,N_15982,N_15760);
or U16378 (N_16378,N_15142,N_15437);
and U16379 (N_16379,N_15443,N_15267);
nor U16380 (N_16380,N_15213,N_15109);
nor U16381 (N_16381,N_15186,N_15831);
nor U16382 (N_16382,N_15837,N_15890);
nand U16383 (N_16383,N_15825,N_15464);
xor U16384 (N_16384,N_15720,N_15652);
nor U16385 (N_16385,N_15673,N_15050);
or U16386 (N_16386,N_15830,N_15932);
nor U16387 (N_16387,N_15810,N_15479);
nor U16388 (N_16388,N_15291,N_15124);
and U16389 (N_16389,N_15370,N_15818);
or U16390 (N_16390,N_15357,N_15783);
and U16391 (N_16391,N_15603,N_15166);
nand U16392 (N_16392,N_15799,N_15984);
nor U16393 (N_16393,N_15905,N_15650);
xor U16394 (N_16394,N_15030,N_15439);
and U16395 (N_16395,N_15786,N_15735);
nor U16396 (N_16396,N_15529,N_15709);
nor U16397 (N_16397,N_15505,N_15989);
xor U16398 (N_16398,N_15795,N_15730);
xor U16399 (N_16399,N_15521,N_15497);
or U16400 (N_16400,N_15400,N_15981);
and U16401 (N_16401,N_15190,N_15066);
xor U16402 (N_16402,N_15587,N_15383);
xnor U16403 (N_16403,N_15661,N_15851);
xor U16404 (N_16404,N_15377,N_15263);
xnor U16405 (N_16405,N_15197,N_15111);
xor U16406 (N_16406,N_15491,N_15930);
nor U16407 (N_16407,N_15610,N_15150);
or U16408 (N_16408,N_15671,N_15306);
or U16409 (N_16409,N_15168,N_15047);
and U16410 (N_16410,N_15647,N_15904);
and U16411 (N_16411,N_15543,N_15145);
nand U16412 (N_16412,N_15594,N_15002);
or U16413 (N_16413,N_15329,N_15222);
and U16414 (N_16414,N_15546,N_15912);
xnor U16415 (N_16415,N_15622,N_15031);
nand U16416 (N_16416,N_15925,N_15776);
nand U16417 (N_16417,N_15426,N_15214);
nand U16418 (N_16418,N_15629,N_15136);
xnor U16419 (N_16419,N_15060,N_15721);
and U16420 (N_16420,N_15512,N_15852);
or U16421 (N_16421,N_15369,N_15672);
or U16422 (N_16422,N_15026,N_15412);
nor U16423 (N_16423,N_15725,N_15722);
nor U16424 (N_16424,N_15274,N_15949);
or U16425 (N_16425,N_15278,N_15685);
or U16426 (N_16426,N_15640,N_15011);
nand U16427 (N_16427,N_15899,N_15675);
and U16428 (N_16428,N_15918,N_15157);
xor U16429 (N_16429,N_15839,N_15071);
nor U16430 (N_16430,N_15059,N_15261);
or U16431 (N_16431,N_15079,N_15183);
or U16432 (N_16432,N_15257,N_15009);
nor U16433 (N_16433,N_15115,N_15854);
or U16434 (N_16434,N_15089,N_15194);
or U16435 (N_16435,N_15054,N_15414);
or U16436 (N_16436,N_15583,N_15154);
xor U16437 (N_16437,N_15927,N_15601);
nand U16438 (N_16438,N_15126,N_15361);
and U16439 (N_16439,N_15346,N_15262);
and U16440 (N_16440,N_15824,N_15943);
xnor U16441 (N_16441,N_15531,N_15856);
nor U16442 (N_16442,N_15653,N_15953);
nand U16443 (N_16443,N_15711,N_15098);
nor U16444 (N_16444,N_15548,N_15749);
xnor U16445 (N_16445,N_15554,N_15941);
xor U16446 (N_16446,N_15615,N_15207);
xor U16447 (N_16447,N_15878,N_15310);
xnor U16448 (N_16448,N_15467,N_15869);
nand U16449 (N_16449,N_15881,N_15204);
or U16450 (N_16450,N_15632,N_15406);
and U16451 (N_16451,N_15789,N_15805);
nor U16452 (N_16452,N_15897,N_15522);
and U16453 (N_16453,N_15578,N_15779);
nand U16454 (N_16454,N_15246,N_15784);
nand U16455 (N_16455,N_15540,N_15116);
nand U16456 (N_16456,N_15739,N_15302);
or U16457 (N_16457,N_15620,N_15040);
and U16458 (N_16458,N_15039,N_15993);
nand U16459 (N_16459,N_15486,N_15816);
or U16460 (N_16460,N_15231,N_15376);
nor U16461 (N_16461,N_15398,N_15561);
xnor U16462 (N_16462,N_15575,N_15352);
nand U16463 (N_16463,N_15639,N_15956);
nand U16464 (N_16464,N_15424,N_15108);
or U16465 (N_16465,N_15051,N_15046);
or U16466 (N_16466,N_15757,N_15996);
nand U16467 (N_16467,N_15595,N_15911);
xnor U16468 (N_16468,N_15173,N_15064);
or U16469 (N_16469,N_15315,N_15235);
and U16470 (N_16470,N_15446,N_15101);
xnor U16471 (N_16471,N_15164,N_15242);
or U16472 (N_16472,N_15348,N_15005);
xor U16473 (N_16473,N_15909,N_15803);
and U16474 (N_16474,N_15697,N_15887);
xor U16475 (N_16475,N_15180,N_15159);
xnor U16476 (N_16476,N_15083,N_15665);
nand U16477 (N_16477,N_15532,N_15644);
nor U16478 (N_16478,N_15844,N_15229);
xnor U16479 (N_16479,N_15585,N_15550);
and U16480 (N_16480,N_15073,N_15409);
nand U16481 (N_16481,N_15475,N_15232);
nand U16482 (N_16482,N_15950,N_15754);
and U16483 (N_16483,N_15964,N_15555);
nor U16484 (N_16484,N_15694,N_15919);
and U16485 (N_16485,N_15162,N_15397);
or U16486 (N_16486,N_15320,N_15275);
and U16487 (N_16487,N_15067,N_15123);
or U16488 (N_16488,N_15053,N_15636);
nand U16489 (N_16489,N_15223,N_15481);
nand U16490 (N_16490,N_15977,N_15728);
nor U16491 (N_16491,N_15637,N_15892);
and U16492 (N_16492,N_15289,N_15495);
nor U16493 (N_16493,N_15218,N_15271);
and U16494 (N_16494,N_15454,N_15822);
or U16495 (N_16495,N_15268,N_15195);
xor U16496 (N_16496,N_15965,N_15335);
xor U16497 (N_16497,N_15883,N_15121);
or U16498 (N_16498,N_15581,N_15393);
and U16499 (N_16499,N_15184,N_15717);
nand U16500 (N_16500,N_15852,N_15333);
or U16501 (N_16501,N_15062,N_15327);
nand U16502 (N_16502,N_15461,N_15503);
and U16503 (N_16503,N_15119,N_15092);
xor U16504 (N_16504,N_15234,N_15593);
and U16505 (N_16505,N_15353,N_15689);
or U16506 (N_16506,N_15407,N_15119);
nor U16507 (N_16507,N_15353,N_15735);
or U16508 (N_16508,N_15861,N_15001);
nor U16509 (N_16509,N_15207,N_15536);
and U16510 (N_16510,N_15629,N_15190);
or U16511 (N_16511,N_15146,N_15205);
and U16512 (N_16512,N_15499,N_15702);
and U16513 (N_16513,N_15207,N_15251);
nand U16514 (N_16514,N_15789,N_15515);
or U16515 (N_16515,N_15466,N_15524);
nand U16516 (N_16516,N_15344,N_15232);
and U16517 (N_16517,N_15079,N_15294);
or U16518 (N_16518,N_15695,N_15036);
and U16519 (N_16519,N_15184,N_15064);
nand U16520 (N_16520,N_15692,N_15542);
nand U16521 (N_16521,N_15350,N_15852);
nand U16522 (N_16522,N_15042,N_15934);
nor U16523 (N_16523,N_15154,N_15274);
nor U16524 (N_16524,N_15074,N_15001);
and U16525 (N_16525,N_15595,N_15822);
and U16526 (N_16526,N_15351,N_15109);
and U16527 (N_16527,N_15956,N_15708);
and U16528 (N_16528,N_15867,N_15561);
and U16529 (N_16529,N_15443,N_15487);
xor U16530 (N_16530,N_15390,N_15197);
xnor U16531 (N_16531,N_15595,N_15976);
or U16532 (N_16532,N_15985,N_15284);
nor U16533 (N_16533,N_15597,N_15987);
or U16534 (N_16534,N_15101,N_15877);
or U16535 (N_16535,N_15132,N_15338);
nor U16536 (N_16536,N_15119,N_15499);
and U16537 (N_16537,N_15034,N_15639);
nand U16538 (N_16538,N_15302,N_15053);
nor U16539 (N_16539,N_15030,N_15468);
nor U16540 (N_16540,N_15978,N_15215);
and U16541 (N_16541,N_15668,N_15440);
and U16542 (N_16542,N_15421,N_15901);
nor U16543 (N_16543,N_15164,N_15414);
nor U16544 (N_16544,N_15205,N_15248);
nand U16545 (N_16545,N_15405,N_15210);
and U16546 (N_16546,N_15261,N_15857);
and U16547 (N_16547,N_15030,N_15118);
nand U16548 (N_16548,N_15747,N_15602);
nand U16549 (N_16549,N_15068,N_15522);
nor U16550 (N_16550,N_15198,N_15641);
xor U16551 (N_16551,N_15017,N_15493);
and U16552 (N_16552,N_15678,N_15642);
or U16553 (N_16553,N_15132,N_15161);
nand U16554 (N_16554,N_15527,N_15307);
nand U16555 (N_16555,N_15298,N_15958);
and U16556 (N_16556,N_15131,N_15110);
nor U16557 (N_16557,N_15982,N_15147);
and U16558 (N_16558,N_15094,N_15751);
nor U16559 (N_16559,N_15623,N_15528);
nand U16560 (N_16560,N_15628,N_15237);
nor U16561 (N_16561,N_15376,N_15499);
and U16562 (N_16562,N_15149,N_15494);
nor U16563 (N_16563,N_15062,N_15002);
or U16564 (N_16564,N_15671,N_15088);
nor U16565 (N_16565,N_15400,N_15231);
and U16566 (N_16566,N_15601,N_15117);
nor U16567 (N_16567,N_15879,N_15744);
and U16568 (N_16568,N_15994,N_15828);
xnor U16569 (N_16569,N_15679,N_15652);
and U16570 (N_16570,N_15227,N_15040);
nor U16571 (N_16571,N_15259,N_15704);
nor U16572 (N_16572,N_15526,N_15248);
and U16573 (N_16573,N_15991,N_15456);
nand U16574 (N_16574,N_15746,N_15387);
and U16575 (N_16575,N_15990,N_15968);
nor U16576 (N_16576,N_15658,N_15889);
xnor U16577 (N_16577,N_15126,N_15210);
nor U16578 (N_16578,N_15212,N_15915);
nand U16579 (N_16579,N_15339,N_15623);
and U16580 (N_16580,N_15078,N_15840);
nor U16581 (N_16581,N_15238,N_15729);
or U16582 (N_16582,N_15373,N_15800);
nand U16583 (N_16583,N_15120,N_15167);
nand U16584 (N_16584,N_15684,N_15250);
or U16585 (N_16585,N_15166,N_15393);
or U16586 (N_16586,N_15099,N_15596);
nor U16587 (N_16587,N_15824,N_15991);
nand U16588 (N_16588,N_15732,N_15061);
and U16589 (N_16589,N_15367,N_15028);
and U16590 (N_16590,N_15159,N_15606);
nor U16591 (N_16591,N_15407,N_15805);
or U16592 (N_16592,N_15723,N_15142);
nand U16593 (N_16593,N_15918,N_15353);
nand U16594 (N_16594,N_15237,N_15193);
or U16595 (N_16595,N_15834,N_15874);
and U16596 (N_16596,N_15215,N_15014);
or U16597 (N_16597,N_15629,N_15792);
or U16598 (N_16598,N_15221,N_15743);
nor U16599 (N_16599,N_15717,N_15210);
xnor U16600 (N_16600,N_15231,N_15872);
and U16601 (N_16601,N_15541,N_15588);
and U16602 (N_16602,N_15103,N_15639);
or U16603 (N_16603,N_15651,N_15921);
xor U16604 (N_16604,N_15896,N_15662);
or U16605 (N_16605,N_15916,N_15626);
xnor U16606 (N_16606,N_15285,N_15653);
and U16607 (N_16607,N_15545,N_15006);
xnor U16608 (N_16608,N_15387,N_15430);
and U16609 (N_16609,N_15650,N_15993);
nand U16610 (N_16610,N_15688,N_15709);
or U16611 (N_16611,N_15116,N_15703);
and U16612 (N_16612,N_15498,N_15028);
nand U16613 (N_16613,N_15368,N_15161);
nand U16614 (N_16614,N_15997,N_15670);
nand U16615 (N_16615,N_15595,N_15023);
nor U16616 (N_16616,N_15744,N_15413);
or U16617 (N_16617,N_15812,N_15295);
xnor U16618 (N_16618,N_15970,N_15075);
nand U16619 (N_16619,N_15516,N_15986);
or U16620 (N_16620,N_15981,N_15470);
xnor U16621 (N_16621,N_15885,N_15279);
xor U16622 (N_16622,N_15839,N_15683);
nand U16623 (N_16623,N_15666,N_15751);
nand U16624 (N_16624,N_15960,N_15784);
xor U16625 (N_16625,N_15731,N_15524);
or U16626 (N_16626,N_15588,N_15345);
and U16627 (N_16627,N_15120,N_15954);
and U16628 (N_16628,N_15770,N_15297);
and U16629 (N_16629,N_15707,N_15032);
nor U16630 (N_16630,N_15677,N_15750);
nand U16631 (N_16631,N_15897,N_15074);
and U16632 (N_16632,N_15429,N_15387);
nand U16633 (N_16633,N_15786,N_15077);
and U16634 (N_16634,N_15456,N_15487);
nor U16635 (N_16635,N_15184,N_15333);
and U16636 (N_16636,N_15744,N_15647);
xnor U16637 (N_16637,N_15312,N_15805);
xor U16638 (N_16638,N_15785,N_15679);
nor U16639 (N_16639,N_15764,N_15259);
or U16640 (N_16640,N_15111,N_15138);
or U16641 (N_16641,N_15626,N_15277);
or U16642 (N_16642,N_15148,N_15664);
xor U16643 (N_16643,N_15902,N_15699);
nor U16644 (N_16644,N_15584,N_15443);
xor U16645 (N_16645,N_15933,N_15770);
nand U16646 (N_16646,N_15988,N_15463);
or U16647 (N_16647,N_15671,N_15327);
or U16648 (N_16648,N_15011,N_15556);
or U16649 (N_16649,N_15848,N_15354);
nand U16650 (N_16650,N_15494,N_15413);
and U16651 (N_16651,N_15497,N_15677);
and U16652 (N_16652,N_15304,N_15580);
and U16653 (N_16653,N_15660,N_15943);
and U16654 (N_16654,N_15684,N_15748);
nand U16655 (N_16655,N_15482,N_15749);
xor U16656 (N_16656,N_15376,N_15167);
or U16657 (N_16657,N_15611,N_15255);
xor U16658 (N_16658,N_15971,N_15858);
nor U16659 (N_16659,N_15884,N_15541);
nor U16660 (N_16660,N_15933,N_15421);
nand U16661 (N_16661,N_15690,N_15535);
or U16662 (N_16662,N_15946,N_15814);
or U16663 (N_16663,N_15558,N_15754);
nand U16664 (N_16664,N_15239,N_15555);
nand U16665 (N_16665,N_15979,N_15543);
xnor U16666 (N_16666,N_15650,N_15131);
xor U16667 (N_16667,N_15396,N_15611);
or U16668 (N_16668,N_15480,N_15185);
and U16669 (N_16669,N_15606,N_15374);
xor U16670 (N_16670,N_15391,N_15033);
or U16671 (N_16671,N_15932,N_15892);
or U16672 (N_16672,N_15319,N_15159);
nor U16673 (N_16673,N_15841,N_15683);
or U16674 (N_16674,N_15612,N_15646);
nor U16675 (N_16675,N_15064,N_15818);
xnor U16676 (N_16676,N_15400,N_15625);
nand U16677 (N_16677,N_15790,N_15321);
nand U16678 (N_16678,N_15598,N_15676);
or U16679 (N_16679,N_15464,N_15165);
and U16680 (N_16680,N_15793,N_15851);
and U16681 (N_16681,N_15145,N_15763);
nand U16682 (N_16682,N_15626,N_15923);
nor U16683 (N_16683,N_15677,N_15061);
nor U16684 (N_16684,N_15401,N_15915);
nor U16685 (N_16685,N_15443,N_15702);
nor U16686 (N_16686,N_15080,N_15154);
xor U16687 (N_16687,N_15787,N_15927);
xnor U16688 (N_16688,N_15429,N_15900);
xor U16689 (N_16689,N_15175,N_15633);
nor U16690 (N_16690,N_15039,N_15727);
or U16691 (N_16691,N_15829,N_15008);
nor U16692 (N_16692,N_15005,N_15718);
xnor U16693 (N_16693,N_15848,N_15619);
xnor U16694 (N_16694,N_15665,N_15681);
xnor U16695 (N_16695,N_15354,N_15921);
and U16696 (N_16696,N_15279,N_15049);
nor U16697 (N_16697,N_15653,N_15497);
or U16698 (N_16698,N_15468,N_15221);
and U16699 (N_16699,N_15579,N_15143);
and U16700 (N_16700,N_15047,N_15052);
and U16701 (N_16701,N_15651,N_15417);
or U16702 (N_16702,N_15655,N_15431);
nand U16703 (N_16703,N_15161,N_15839);
or U16704 (N_16704,N_15408,N_15162);
or U16705 (N_16705,N_15720,N_15587);
nor U16706 (N_16706,N_15351,N_15246);
nor U16707 (N_16707,N_15740,N_15080);
nand U16708 (N_16708,N_15593,N_15429);
nand U16709 (N_16709,N_15116,N_15920);
and U16710 (N_16710,N_15754,N_15362);
or U16711 (N_16711,N_15594,N_15360);
and U16712 (N_16712,N_15902,N_15161);
nand U16713 (N_16713,N_15760,N_15320);
or U16714 (N_16714,N_15015,N_15643);
nand U16715 (N_16715,N_15518,N_15002);
or U16716 (N_16716,N_15557,N_15464);
nor U16717 (N_16717,N_15984,N_15201);
nor U16718 (N_16718,N_15869,N_15651);
nand U16719 (N_16719,N_15165,N_15224);
and U16720 (N_16720,N_15734,N_15304);
nand U16721 (N_16721,N_15169,N_15628);
or U16722 (N_16722,N_15151,N_15807);
nor U16723 (N_16723,N_15955,N_15585);
nand U16724 (N_16724,N_15553,N_15346);
nor U16725 (N_16725,N_15288,N_15845);
xor U16726 (N_16726,N_15231,N_15177);
and U16727 (N_16727,N_15376,N_15697);
or U16728 (N_16728,N_15775,N_15130);
or U16729 (N_16729,N_15241,N_15093);
and U16730 (N_16730,N_15349,N_15552);
xnor U16731 (N_16731,N_15978,N_15241);
nor U16732 (N_16732,N_15164,N_15844);
nand U16733 (N_16733,N_15800,N_15943);
nor U16734 (N_16734,N_15778,N_15178);
nor U16735 (N_16735,N_15312,N_15423);
nand U16736 (N_16736,N_15366,N_15822);
xor U16737 (N_16737,N_15749,N_15066);
nand U16738 (N_16738,N_15628,N_15418);
nand U16739 (N_16739,N_15712,N_15623);
and U16740 (N_16740,N_15686,N_15424);
xor U16741 (N_16741,N_15643,N_15461);
or U16742 (N_16742,N_15481,N_15285);
or U16743 (N_16743,N_15925,N_15552);
xnor U16744 (N_16744,N_15821,N_15645);
or U16745 (N_16745,N_15350,N_15993);
xor U16746 (N_16746,N_15665,N_15400);
and U16747 (N_16747,N_15435,N_15417);
or U16748 (N_16748,N_15704,N_15937);
nor U16749 (N_16749,N_15465,N_15044);
nor U16750 (N_16750,N_15104,N_15181);
and U16751 (N_16751,N_15112,N_15143);
xnor U16752 (N_16752,N_15327,N_15905);
or U16753 (N_16753,N_15268,N_15626);
xnor U16754 (N_16754,N_15729,N_15663);
nor U16755 (N_16755,N_15021,N_15437);
nor U16756 (N_16756,N_15156,N_15186);
xnor U16757 (N_16757,N_15639,N_15542);
nand U16758 (N_16758,N_15023,N_15268);
nand U16759 (N_16759,N_15977,N_15120);
and U16760 (N_16760,N_15692,N_15125);
nor U16761 (N_16761,N_15066,N_15473);
or U16762 (N_16762,N_15131,N_15468);
and U16763 (N_16763,N_15966,N_15783);
or U16764 (N_16764,N_15568,N_15311);
nor U16765 (N_16765,N_15770,N_15202);
nor U16766 (N_16766,N_15046,N_15785);
nand U16767 (N_16767,N_15795,N_15499);
xnor U16768 (N_16768,N_15597,N_15167);
xnor U16769 (N_16769,N_15072,N_15328);
nand U16770 (N_16770,N_15433,N_15159);
and U16771 (N_16771,N_15693,N_15294);
and U16772 (N_16772,N_15856,N_15602);
xnor U16773 (N_16773,N_15205,N_15551);
and U16774 (N_16774,N_15107,N_15778);
and U16775 (N_16775,N_15704,N_15479);
xnor U16776 (N_16776,N_15101,N_15769);
or U16777 (N_16777,N_15582,N_15502);
xnor U16778 (N_16778,N_15874,N_15400);
nor U16779 (N_16779,N_15154,N_15684);
xnor U16780 (N_16780,N_15274,N_15501);
or U16781 (N_16781,N_15340,N_15428);
nor U16782 (N_16782,N_15239,N_15535);
or U16783 (N_16783,N_15003,N_15454);
nor U16784 (N_16784,N_15299,N_15319);
or U16785 (N_16785,N_15355,N_15651);
nor U16786 (N_16786,N_15757,N_15260);
nor U16787 (N_16787,N_15740,N_15038);
xor U16788 (N_16788,N_15558,N_15643);
xor U16789 (N_16789,N_15441,N_15690);
and U16790 (N_16790,N_15173,N_15676);
xnor U16791 (N_16791,N_15315,N_15928);
nand U16792 (N_16792,N_15035,N_15657);
xor U16793 (N_16793,N_15828,N_15388);
or U16794 (N_16794,N_15901,N_15082);
nor U16795 (N_16795,N_15022,N_15703);
nand U16796 (N_16796,N_15366,N_15123);
nor U16797 (N_16797,N_15206,N_15790);
and U16798 (N_16798,N_15862,N_15665);
nand U16799 (N_16799,N_15380,N_15394);
xor U16800 (N_16800,N_15868,N_15996);
xor U16801 (N_16801,N_15519,N_15676);
nand U16802 (N_16802,N_15413,N_15969);
nand U16803 (N_16803,N_15603,N_15772);
and U16804 (N_16804,N_15063,N_15292);
nand U16805 (N_16805,N_15325,N_15272);
xnor U16806 (N_16806,N_15017,N_15752);
nand U16807 (N_16807,N_15130,N_15170);
and U16808 (N_16808,N_15313,N_15713);
or U16809 (N_16809,N_15459,N_15149);
or U16810 (N_16810,N_15006,N_15086);
xor U16811 (N_16811,N_15770,N_15049);
or U16812 (N_16812,N_15106,N_15417);
nand U16813 (N_16813,N_15937,N_15628);
and U16814 (N_16814,N_15945,N_15699);
nand U16815 (N_16815,N_15312,N_15875);
nor U16816 (N_16816,N_15180,N_15911);
nand U16817 (N_16817,N_15053,N_15547);
or U16818 (N_16818,N_15448,N_15703);
or U16819 (N_16819,N_15596,N_15682);
nor U16820 (N_16820,N_15276,N_15650);
nand U16821 (N_16821,N_15905,N_15902);
nand U16822 (N_16822,N_15762,N_15334);
nor U16823 (N_16823,N_15500,N_15368);
or U16824 (N_16824,N_15829,N_15137);
or U16825 (N_16825,N_15525,N_15310);
xor U16826 (N_16826,N_15666,N_15497);
nor U16827 (N_16827,N_15027,N_15714);
nor U16828 (N_16828,N_15698,N_15206);
nor U16829 (N_16829,N_15821,N_15531);
and U16830 (N_16830,N_15049,N_15865);
xor U16831 (N_16831,N_15877,N_15349);
xnor U16832 (N_16832,N_15961,N_15183);
nor U16833 (N_16833,N_15687,N_15366);
xnor U16834 (N_16834,N_15745,N_15542);
nor U16835 (N_16835,N_15267,N_15241);
or U16836 (N_16836,N_15428,N_15199);
nor U16837 (N_16837,N_15113,N_15785);
xnor U16838 (N_16838,N_15867,N_15614);
nor U16839 (N_16839,N_15078,N_15452);
and U16840 (N_16840,N_15219,N_15782);
or U16841 (N_16841,N_15637,N_15695);
nand U16842 (N_16842,N_15094,N_15459);
nand U16843 (N_16843,N_15685,N_15457);
and U16844 (N_16844,N_15298,N_15565);
nand U16845 (N_16845,N_15675,N_15108);
nand U16846 (N_16846,N_15117,N_15212);
nand U16847 (N_16847,N_15722,N_15180);
nor U16848 (N_16848,N_15053,N_15693);
nand U16849 (N_16849,N_15623,N_15989);
nor U16850 (N_16850,N_15929,N_15469);
and U16851 (N_16851,N_15020,N_15615);
or U16852 (N_16852,N_15580,N_15722);
and U16853 (N_16853,N_15579,N_15622);
or U16854 (N_16854,N_15579,N_15187);
or U16855 (N_16855,N_15885,N_15386);
nor U16856 (N_16856,N_15634,N_15388);
nand U16857 (N_16857,N_15997,N_15522);
xnor U16858 (N_16858,N_15218,N_15727);
and U16859 (N_16859,N_15182,N_15824);
nand U16860 (N_16860,N_15712,N_15263);
xnor U16861 (N_16861,N_15155,N_15143);
xor U16862 (N_16862,N_15372,N_15119);
or U16863 (N_16863,N_15440,N_15239);
and U16864 (N_16864,N_15766,N_15068);
nand U16865 (N_16865,N_15733,N_15579);
nand U16866 (N_16866,N_15656,N_15111);
xor U16867 (N_16867,N_15641,N_15354);
and U16868 (N_16868,N_15158,N_15179);
or U16869 (N_16869,N_15840,N_15450);
nor U16870 (N_16870,N_15391,N_15808);
or U16871 (N_16871,N_15961,N_15501);
and U16872 (N_16872,N_15934,N_15241);
nor U16873 (N_16873,N_15145,N_15339);
xor U16874 (N_16874,N_15717,N_15768);
nor U16875 (N_16875,N_15977,N_15487);
or U16876 (N_16876,N_15597,N_15370);
or U16877 (N_16877,N_15594,N_15918);
nor U16878 (N_16878,N_15546,N_15949);
nor U16879 (N_16879,N_15766,N_15477);
or U16880 (N_16880,N_15798,N_15164);
xnor U16881 (N_16881,N_15825,N_15329);
nand U16882 (N_16882,N_15536,N_15711);
xnor U16883 (N_16883,N_15037,N_15940);
or U16884 (N_16884,N_15331,N_15313);
nor U16885 (N_16885,N_15517,N_15368);
xor U16886 (N_16886,N_15674,N_15520);
xor U16887 (N_16887,N_15993,N_15017);
xor U16888 (N_16888,N_15579,N_15486);
and U16889 (N_16889,N_15110,N_15355);
nor U16890 (N_16890,N_15411,N_15874);
or U16891 (N_16891,N_15822,N_15865);
nand U16892 (N_16892,N_15043,N_15856);
nand U16893 (N_16893,N_15198,N_15544);
xor U16894 (N_16894,N_15649,N_15230);
and U16895 (N_16895,N_15543,N_15971);
nand U16896 (N_16896,N_15136,N_15876);
and U16897 (N_16897,N_15352,N_15171);
xor U16898 (N_16898,N_15948,N_15385);
xnor U16899 (N_16899,N_15084,N_15630);
nor U16900 (N_16900,N_15664,N_15822);
or U16901 (N_16901,N_15902,N_15700);
and U16902 (N_16902,N_15766,N_15336);
and U16903 (N_16903,N_15695,N_15087);
nand U16904 (N_16904,N_15288,N_15963);
or U16905 (N_16905,N_15494,N_15358);
xnor U16906 (N_16906,N_15433,N_15725);
nand U16907 (N_16907,N_15644,N_15440);
and U16908 (N_16908,N_15617,N_15241);
xor U16909 (N_16909,N_15407,N_15939);
nand U16910 (N_16910,N_15467,N_15423);
nor U16911 (N_16911,N_15768,N_15636);
xnor U16912 (N_16912,N_15103,N_15002);
nor U16913 (N_16913,N_15595,N_15845);
nand U16914 (N_16914,N_15620,N_15561);
nor U16915 (N_16915,N_15079,N_15812);
and U16916 (N_16916,N_15000,N_15654);
nor U16917 (N_16917,N_15227,N_15278);
xnor U16918 (N_16918,N_15491,N_15609);
or U16919 (N_16919,N_15188,N_15818);
or U16920 (N_16920,N_15979,N_15351);
or U16921 (N_16921,N_15495,N_15191);
nand U16922 (N_16922,N_15816,N_15487);
nor U16923 (N_16923,N_15626,N_15940);
and U16924 (N_16924,N_15645,N_15601);
nor U16925 (N_16925,N_15323,N_15885);
or U16926 (N_16926,N_15722,N_15414);
nor U16927 (N_16927,N_15647,N_15191);
nand U16928 (N_16928,N_15631,N_15261);
or U16929 (N_16929,N_15805,N_15020);
nand U16930 (N_16930,N_15076,N_15124);
or U16931 (N_16931,N_15683,N_15596);
xnor U16932 (N_16932,N_15789,N_15026);
nor U16933 (N_16933,N_15834,N_15121);
nand U16934 (N_16934,N_15758,N_15706);
nand U16935 (N_16935,N_15771,N_15217);
nand U16936 (N_16936,N_15847,N_15064);
nand U16937 (N_16937,N_15103,N_15700);
or U16938 (N_16938,N_15278,N_15799);
nand U16939 (N_16939,N_15495,N_15091);
xnor U16940 (N_16940,N_15443,N_15566);
or U16941 (N_16941,N_15472,N_15848);
xnor U16942 (N_16942,N_15631,N_15879);
and U16943 (N_16943,N_15857,N_15621);
and U16944 (N_16944,N_15252,N_15642);
and U16945 (N_16945,N_15402,N_15799);
nor U16946 (N_16946,N_15508,N_15544);
and U16947 (N_16947,N_15753,N_15129);
xor U16948 (N_16948,N_15208,N_15410);
nand U16949 (N_16949,N_15303,N_15896);
nand U16950 (N_16950,N_15023,N_15143);
nor U16951 (N_16951,N_15271,N_15409);
xor U16952 (N_16952,N_15653,N_15428);
and U16953 (N_16953,N_15524,N_15613);
xnor U16954 (N_16954,N_15268,N_15638);
or U16955 (N_16955,N_15164,N_15269);
nor U16956 (N_16956,N_15575,N_15618);
nor U16957 (N_16957,N_15271,N_15515);
xnor U16958 (N_16958,N_15090,N_15367);
nor U16959 (N_16959,N_15630,N_15979);
xnor U16960 (N_16960,N_15580,N_15286);
nor U16961 (N_16961,N_15989,N_15054);
or U16962 (N_16962,N_15417,N_15171);
nand U16963 (N_16963,N_15389,N_15967);
xnor U16964 (N_16964,N_15828,N_15050);
and U16965 (N_16965,N_15714,N_15315);
nor U16966 (N_16966,N_15516,N_15961);
xnor U16967 (N_16967,N_15310,N_15010);
nand U16968 (N_16968,N_15057,N_15404);
nand U16969 (N_16969,N_15949,N_15076);
nor U16970 (N_16970,N_15501,N_15818);
and U16971 (N_16971,N_15553,N_15033);
xor U16972 (N_16972,N_15150,N_15288);
and U16973 (N_16973,N_15818,N_15460);
nand U16974 (N_16974,N_15240,N_15612);
nand U16975 (N_16975,N_15445,N_15620);
nor U16976 (N_16976,N_15422,N_15516);
nand U16977 (N_16977,N_15223,N_15828);
xor U16978 (N_16978,N_15590,N_15576);
xor U16979 (N_16979,N_15308,N_15797);
xnor U16980 (N_16980,N_15599,N_15154);
xnor U16981 (N_16981,N_15430,N_15647);
and U16982 (N_16982,N_15746,N_15800);
nor U16983 (N_16983,N_15041,N_15599);
and U16984 (N_16984,N_15254,N_15762);
nor U16985 (N_16985,N_15800,N_15252);
and U16986 (N_16986,N_15306,N_15846);
nor U16987 (N_16987,N_15247,N_15113);
or U16988 (N_16988,N_15088,N_15507);
nand U16989 (N_16989,N_15817,N_15752);
or U16990 (N_16990,N_15819,N_15368);
or U16991 (N_16991,N_15271,N_15697);
nor U16992 (N_16992,N_15367,N_15689);
nor U16993 (N_16993,N_15626,N_15355);
nor U16994 (N_16994,N_15914,N_15514);
and U16995 (N_16995,N_15013,N_15292);
or U16996 (N_16996,N_15458,N_15172);
and U16997 (N_16997,N_15329,N_15245);
and U16998 (N_16998,N_15803,N_15329);
xnor U16999 (N_16999,N_15775,N_15901);
xnor U17000 (N_17000,N_16840,N_16630);
or U17001 (N_17001,N_16599,N_16554);
or U17002 (N_17002,N_16883,N_16976);
nand U17003 (N_17003,N_16548,N_16658);
xor U17004 (N_17004,N_16953,N_16798);
nor U17005 (N_17005,N_16206,N_16593);
nor U17006 (N_17006,N_16961,N_16329);
nor U17007 (N_17007,N_16971,N_16861);
nand U17008 (N_17008,N_16233,N_16401);
nor U17009 (N_17009,N_16801,N_16078);
xor U17010 (N_17010,N_16140,N_16142);
nand U17011 (N_17011,N_16001,N_16046);
or U17012 (N_17012,N_16562,N_16956);
xor U17013 (N_17013,N_16287,N_16405);
nor U17014 (N_17014,N_16446,N_16717);
and U17015 (N_17015,N_16704,N_16478);
or U17016 (N_17016,N_16999,N_16937);
xor U17017 (N_17017,N_16396,N_16508);
and U17018 (N_17018,N_16458,N_16439);
xor U17019 (N_17019,N_16754,N_16687);
nand U17020 (N_17020,N_16064,N_16910);
nand U17021 (N_17021,N_16133,N_16387);
or U17022 (N_17022,N_16277,N_16180);
xnor U17023 (N_17023,N_16926,N_16870);
and U17024 (N_17024,N_16669,N_16829);
nand U17025 (N_17025,N_16194,N_16238);
and U17026 (N_17026,N_16952,N_16369);
nor U17027 (N_17027,N_16404,N_16311);
nand U17028 (N_17028,N_16815,N_16964);
and U17029 (N_17029,N_16573,N_16411);
nor U17030 (N_17030,N_16553,N_16093);
xor U17031 (N_17031,N_16675,N_16740);
and U17032 (N_17032,N_16294,N_16415);
xor U17033 (N_17033,N_16111,N_16723);
or U17034 (N_17034,N_16677,N_16544);
and U17035 (N_17035,N_16940,N_16278);
xnor U17036 (N_17036,N_16388,N_16853);
xor U17037 (N_17037,N_16533,N_16510);
or U17038 (N_17038,N_16598,N_16733);
xor U17039 (N_17039,N_16463,N_16392);
xnor U17040 (N_17040,N_16274,N_16184);
nor U17041 (N_17041,N_16412,N_16484);
and U17042 (N_17042,N_16907,N_16837);
nor U17043 (N_17043,N_16247,N_16930);
xnor U17044 (N_17044,N_16252,N_16582);
and U17045 (N_17045,N_16399,N_16110);
nor U17046 (N_17046,N_16128,N_16119);
and U17047 (N_17047,N_16254,N_16962);
nor U17048 (N_17048,N_16890,N_16153);
nor U17049 (N_17049,N_16877,N_16340);
xor U17050 (N_17050,N_16793,N_16958);
nand U17051 (N_17051,N_16509,N_16270);
or U17052 (N_17052,N_16359,N_16182);
nor U17053 (N_17053,N_16306,N_16646);
nor U17054 (N_17054,N_16413,N_16283);
or U17055 (N_17055,N_16747,N_16087);
nand U17056 (N_17056,N_16944,N_16059);
nand U17057 (N_17057,N_16679,N_16792);
nand U17058 (N_17058,N_16070,N_16539);
nand U17059 (N_17059,N_16227,N_16950);
xnor U17060 (N_17060,N_16858,N_16806);
xnor U17061 (N_17061,N_16874,N_16368);
nor U17062 (N_17062,N_16394,N_16529);
and U17063 (N_17063,N_16876,N_16315);
nand U17064 (N_17064,N_16805,N_16498);
and U17065 (N_17065,N_16807,N_16290);
or U17066 (N_17066,N_16225,N_16019);
or U17067 (N_17067,N_16260,N_16159);
xor U17068 (N_17068,N_16702,N_16796);
nor U17069 (N_17069,N_16844,N_16766);
nand U17070 (N_17070,N_16812,N_16645);
or U17071 (N_17071,N_16178,N_16370);
nand U17072 (N_17072,N_16731,N_16381);
or U17073 (N_17073,N_16467,N_16674);
nand U17074 (N_17074,N_16273,N_16165);
or U17075 (N_17075,N_16568,N_16209);
and U17076 (N_17076,N_16709,N_16830);
nand U17077 (N_17077,N_16557,N_16968);
nand U17078 (N_17078,N_16210,N_16347);
xor U17079 (N_17079,N_16694,N_16008);
or U17080 (N_17080,N_16822,N_16433);
nand U17081 (N_17081,N_16264,N_16288);
xor U17082 (N_17082,N_16664,N_16672);
or U17083 (N_17083,N_16085,N_16318);
nor U17084 (N_17084,N_16574,N_16231);
nand U17085 (N_17085,N_16915,N_16602);
xor U17086 (N_17086,N_16328,N_16158);
nand U17087 (N_17087,N_16698,N_16355);
or U17088 (N_17088,N_16567,N_16762);
nand U17089 (N_17089,N_16635,N_16163);
or U17090 (N_17090,N_16765,N_16846);
nor U17091 (N_17091,N_16025,N_16503);
nor U17092 (N_17092,N_16092,N_16989);
or U17093 (N_17093,N_16735,N_16454);
or U17094 (N_17094,N_16847,N_16098);
nor U17095 (N_17095,N_16734,N_16699);
or U17096 (N_17096,N_16432,N_16560);
nand U17097 (N_17097,N_16337,N_16443);
or U17098 (N_17098,N_16452,N_16591);
xor U17099 (N_17099,N_16515,N_16058);
nand U17100 (N_17100,N_16872,N_16052);
nor U17101 (N_17101,N_16549,N_16650);
or U17102 (N_17102,N_16230,N_16229);
nor U17103 (N_17103,N_16933,N_16938);
or U17104 (N_17104,N_16016,N_16050);
or U17105 (N_17105,N_16346,N_16295);
nand U17106 (N_17106,N_16045,N_16753);
xor U17107 (N_17107,N_16320,N_16339);
xor U17108 (N_17108,N_16258,N_16500);
nor U17109 (N_17109,N_16795,N_16176);
or U17110 (N_17110,N_16901,N_16151);
or U17111 (N_17111,N_16228,N_16168);
and U17112 (N_17112,N_16895,N_16586);
or U17113 (N_17113,N_16018,N_16980);
xor U17114 (N_17114,N_16639,N_16007);
nand U17115 (N_17115,N_16038,N_16365);
or U17116 (N_17116,N_16345,N_16362);
xnor U17117 (N_17117,N_16817,N_16714);
nand U17118 (N_17118,N_16905,N_16994);
or U17119 (N_17119,N_16564,N_16712);
xnor U17120 (N_17120,N_16730,N_16308);
nor U17121 (N_17121,N_16935,N_16809);
or U17122 (N_17122,N_16237,N_16426);
or U17123 (N_17123,N_16169,N_16957);
xor U17124 (N_17124,N_16073,N_16794);
or U17125 (N_17125,N_16450,N_16124);
and U17126 (N_17126,N_16029,N_16756);
and U17127 (N_17127,N_16610,N_16902);
nor U17128 (N_17128,N_16407,N_16843);
and U17129 (N_17129,N_16470,N_16845);
nor U17130 (N_17130,N_16114,N_16927);
nand U17131 (N_17131,N_16973,N_16688);
nand U17132 (N_17132,N_16545,N_16033);
nand U17133 (N_17133,N_16784,N_16848);
nand U17134 (N_17134,N_16918,N_16720);
xnor U17135 (N_17135,N_16267,N_16280);
nor U17136 (N_17136,N_16473,N_16623);
nand U17137 (N_17137,N_16965,N_16997);
or U17138 (N_17138,N_16697,N_16494);
or U17139 (N_17139,N_16268,N_16571);
nand U17140 (N_17140,N_16523,N_16010);
xor U17141 (N_17141,N_16285,N_16071);
nor U17142 (N_17142,N_16887,N_16827);
nand U17143 (N_17143,N_16036,N_16390);
xor U17144 (N_17144,N_16269,N_16350);
xnor U17145 (N_17145,N_16517,N_16035);
nand U17146 (N_17146,N_16682,N_16992);
nor U17147 (N_17147,N_16491,N_16116);
nand U17148 (N_17148,N_16441,N_16242);
nor U17149 (N_17149,N_16621,N_16057);
and U17150 (N_17150,N_16651,N_16929);
and U17151 (N_17151,N_16606,N_16696);
or U17152 (N_17152,N_16767,N_16167);
and U17153 (N_17153,N_16461,N_16305);
nand U17154 (N_17154,N_16455,N_16608);
and U17155 (N_17155,N_16779,N_16297);
and U17156 (N_17156,N_16501,N_16683);
or U17157 (N_17157,N_16084,N_16541);
nand U17158 (N_17158,N_16187,N_16185);
nand U17159 (N_17159,N_16946,N_16521);
and U17160 (N_17160,N_16898,N_16863);
and U17161 (N_17161,N_16963,N_16145);
nor U17162 (N_17162,N_16855,N_16575);
nor U17163 (N_17163,N_16813,N_16129);
or U17164 (N_17164,N_16922,N_16040);
nand U17165 (N_17165,N_16186,N_16743);
xor U17166 (N_17166,N_16425,N_16179);
nand U17167 (N_17167,N_16333,N_16917);
nand U17168 (N_17168,N_16527,N_16903);
nand U17169 (N_17169,N_16649,N_16978);
or U17170 (N_17170,N_16969,N_16559);
xor U17171 (N_17171,N_16459,N_16859);
and U17172 (N_17172,N_16246,N_16875);
nor U17173 (N_17173,N_16482,N_16244);
xor U17174 (N_17174,N_16594,N_16892);
nor U17175 (N_17175,N_16449,N_16495);
nor U17176 (N_17176,N_16291,N_16641);
and U17177 (N_17177,N_16109,N_16881);
and U17178 (N_17178,N_16834,N_16836);
xnor U17179 (N_17179,N_16744,N_16886);
nor U17180 (N_17180,N_16620,N_16919);
nor U17181 (N_17181,N_16466,N_16344);
nand U17182 (N_17182,N_16703,N_16864);
xnor U17183 (N_17183,N_16015,N_16204);
or U17184 (N_17184,N_16120,N_16437);
xor U17185 (N_17185,N_16076,N_16808);
nor U17186 (N_17186,N_16511,N_16048);
xor U17187 (N_17187,N_16155,N_16728);
nand U17188 (N_17188,N_16654,N_16257);
nor U17189 (N_17189,N_16445,N_16826);
nand U17190 (N_17190,N_16082,N_16906);
nor U17191 (N_17191,N_16923,N_16556);
or U17192 (N_17192,N_16122,N_16661);
xor U17193 (N_17193,N_16094,N_16190);
xor U17194 (N_17194,N_16716,N_16604);
or U17195 (N_17195,N_16148,N_16420);
xor U17196 (N_17196,N_16424,N_16970);
nand U17197 (N_17197,N_16692,N_16024);
nand U17198 (N_17198,N_16310,N_16841);
or U17199 (N_17199,N_16607,N_16115);
nor U17200 (N_17200,N_16732,N_16357);
xor U17201 (N_17201,N_16833,N_16665);
and U17202 (N_17202,N_16587,N_16982);
and U17203 (N_17203,N_16854,N_16324);
or U17204 (N_17204,N_16331,N_16090);
xnor U17205 (N_17205,N_16668,N_16781);
nand U17206 (N_17206,N_16410,N_16525);
or U17207 (N_17207,N_16197,N_16819);
nor U17208 (N_17208,N_16408,N_16660);
nor U17209 (N_17209,N_16232,N_16374);
nor U17210 (N_17210,N_16043,N_16343);
nor U17211 (N_17211,N_16802,N_16416);
nand U17212 (N_17212,N_16519,N_16107);
nor U17213 (N_17213,N_16528,N_16749);
or U17214 (N_17214,N_16212,N_16729);
and U17215 (N_17215,N_16266,N_16030);
nand U17216 (N_17216,N_16219,N_16351);
xnor U17217 (N_17217,N_16823,N_16403);
or U17218 (N_17218,N_16485,N_16220);
nor U17219 (N_17219,N_16986,N_16436);
nand U17220 (N_17220,N_16380,N_16972);
nor U17221 (N_17221,N_16341,N_16289);
xor U17222 (N_17222,N_16880,N_16656);
xnor U17223 (N_17223,N_16745,N_16601);
nand U17224 (N_17224,N_16298,N_16505);
xnor U17225 (N_17225,N_16195,N_16199);
nand U17226 (N_17226,N_16442,N_16975);
and U17227 (N_17227,N_16106,N_16398);
or U17228 (N_17228,N_16924,N_16504);
nand U17229 (N_17229,N_16263,N_16386);
nand U17230 (N_17230,N_16166,N_16695);
or U17231 (N_17231,N_16105,N_16780);
and U17232 (N_17232,N_16526,N_16021);
nand U17233 (N_17233,N_16502,N_16349);
xor U17234 (N_17234,N_16857,N_16047);
xor U17235 (N_17235,N_16261,N_16418);
and U17236 (N_17236,N_16925,N_16136);
or U17237 (N_17237,N_16967,N_16304);
nor U17238 (N_17238,N_16395,N_16002);
and U17239 (N_17239,N_16832,N_16787);
nand U17240 (N_17240,N_16617,N_16786);
nand U17241 (N_17241,N_16625,N_16026);
and U17242 (N_17242,N_16543,N_16170);
xnor U17243 (N_17243,N_16949,N_16321);
xnor U17244 (N_17244,N_16056,N_16160);
and U17245 (N_17245,N_16065,N_16516);
and U17246 (N_17246,N_16055,N_16474);
or U17247 (N_17247,N_16079,N_16979);
and U17248 (N_17248,N_16772,N_16137);
xnor U17249 (N_17249,N_16039,N_16987);
nand U17250 (N_17250,N_16372,N_16081);
nor U17251 (N_17251,N_16626,N_16685);
and U17252 (N_17252,N_16427,N_16518);
xor U17253 (N_17253,N_16913,N_16939);
or U17254 (N_17254,N_16123,N_16684);
nor U17255 (N_17255,N_16921,N_16431);
nand U17256 (N_17256,N_16768,N_16570);
or U17257 (N_17257,N_16173,N_16208);
xor U17258 (N_17258,N_16300,N_16118);
nand U17259 (N_17259,N_16095,N_16882);
and U17260 (N_17260,N_16681,N_16138);
and U17261 (N_17261,N_16271,N_16147);
nand U17262 (N_17262,N_16551,N_16746);
or U17263 (N_17263,N_16423,N_16154);
nor U17264 (N_17264,N_16430,N_16959);
and U17265 (N_17265,N_16755,N_16713);
or U17266 (N_17266,N_16108,N_16721);
and U17267 (N_17267,N_16904,N_16005);
nand U17268 (N_17268,N_16616,N_16996);
nand U17269 (N_17269,N_16552,N_16286);
nand U17270 (N_17270,N_16644,N_16149);
or U17271 (N_17271,N_16991,N_16215);
and U17272 (N_17272,N_16532,N_16497);
and U17273 (N_17273,N_16307,N_16448);
nand U17274 (N_17274,N_16619,N_16471);
nor U17275 (N_17275,N_16891,N_16314);
or U17276 (N_17276,N_16479,N_16800);
and U17277 (N_17277,N_16818,N_16476);
xnor U17278 (N_17278,N_16850,N_16330);
or U17279 (N_17279,N_16156,N_16657);
xnor U17280 (N_17280,N_16382,N_16977);
xor U17281 (N_17281,N_16336,N_16327);
nor U17282 (N_17282,N_16900,N_16783);
nor U17283 (N_17283,N_16579,N_16634);
or U17284 (N_17284,N_16565,N_16583);
xor U17285 (N_17285,N_16101,N_16096);
nor U17286 (N_17286,N_16871,N_16004);
and U17287 (N_17287,N_16259,N_16652);
nand U17288 (N_17288,N_16255,N_16014);
and U17289 (N_17289,N_16788,N_16605);
or U17290 (N_17290,N_16663,N_16947);
nand U17291 (N_17291,N_16748,N_16611);
nand U17292 (N_17292,N_16912,N_16993);
nand U17293 (N_17293,N_16711,N_16239);
or U17294 (N_17294,N_16360,N_16540);
nor U17295 (N_17295,N_16726,N_16332);
and U17296 (N_17296,N_16581,N_16974);
nand U17297 (N_17297,N_16642,N_16188);
xor U17298 (N_17298,N_16542,N_16032);
nor U17299 (N_17299,N_16217,N_16804);
xnor U17300 (N_17300,N_16421,N_16691);
nor U17301 (N_17301,N_16348,N_16810);
and U17302 (N_17302,N_16356,N_16856);
xnor U17303 (N_17303,N_16936,N_16865);
xor U17304 (N_17304,N_16177,N_16161);
nand U17305 (N_17305,N_16453,N_16104);
and U17306 (N_17306,N_16223,N_16839);
xor U17307 (N_17307,N_16707,N_16584);
nand U17308 (N_17308,N_16499,N_16488);
nor U17309 (N_17309,N_16908,N_16736);
and U17310 (N_17310,N_16376,N_16816);
nor U17311 (N_17311,N_16724,N_16867);
and U17312 (N_17312,N_16221,N_16130);
nand U17313 (N_17313,N_16613,N_16135);
xor U17314 (N_17314,N_16366,N_16911);
or U17315 (N_17315,N_16440,N_16477);
nand U17316 (N_17316,N_16031,N_16868);
nand U17317 (N_17317,N_16507,N_16690);
or U17318 (N_17318,N_16146,N_16060);
nand U17319 (N_17319,N_16292,N_16770);
xor U17320 (N_17320,N_16757,N_16378);
nand U17321 (N_17321,N_16889,N_16852);
and U17322 (N_17322,N_16742,N_16216);
nand U17323 (N_17323,N_16282,N_16981);
or U17324 (N_17324,N_16438,N_16434);
xnor U17325 (N_17325,N_16067,N_16132);
nand U17326 (N_17326,N_16546,N_16322);
and U17327 (N_17327,N_16667,N_16486);
nor U17328 (N_17328,N_16472,N_16866);
or U17329 (N_17329,N_16272,N_16066);
nand U17330 (N_17330,N_16671,N_16998);
nor U17331 (N_17331,N_16086,N_16647);
and U17332 (N_17332,N_16535,N_16000);
nand U17333 (N_17333,N_16522,N_16465);
nor U17334 (N_17334,N_16253,N_16489);
nand U17335 (N_17335,N_16088,N_16384);
xor U17336 (N_17336,N_16774,N_16791);
nor U17337 (N_17337,N_16612,N_16480);
and U17338 (N_17338,N_16831,N_16701);
and U17339 (N_17339,N_16638,N_16954);
nand U17340 (N_17340,N_16256,N_16323);
or U17341 (N_17341,N_16689,N_16706);
and U17342 (N_17342,N_16012,N_16849);
nand U17343 (N_17343,N_16966,N_16771);
nor U17344 (N_17344,N_16960,N_16763);
xnor U17345 (N_17345,N_16371,N_16838);
and U17346 (N_17346,N_16629,N_16775);
or U17347 (N_17347,N_16017,N_16633);
nor U17348 (N_17348,N_16537,N_16493);
or U17349 (N_17349,N_16335,N_16131);
xor U17350 (N_17350,N_16444,N_16006);
xnor U17351 (N_17351,N_16400,N_16592);
nor U17352 (N_17352,N_16985,N_16174);
nor U17353 (N_17353,N_16490,N_16631);
xor U17354 (N_17354,N_16761,N_16162);
or U17355 (N_17355,N_16879,N_16296);
xnor U17356 (N_17356,N_16203,N_16572);
nor U17357 (N_17357,N_16099,N_16191);
xnor U17358 (N_17358,N_16429,N_16597);
and U17359 (N_17359,N_16385,N_16074);
nand U17360 (N_17360,N_16091,N_16512);
nand U17361 (N_17361,N_16062,N_16799);
nand U17362 (N_17362,N_16023,N_16680);
xor U17363 (N_17363,N_16492,N_16192);
nor U17364 (N_17364,N_16250,N_16778);
xor U17365 (N_17365,N_16224,N_16334);
nand U17366 (N_17366,N_16725,N_16739);
xor U17367 (N_17367,N_16377,N_16069);
nor U17368 (N_17368,N_16075,N_16113);
nand U17369 (N_17369,N_16632,N_16715);
nor U17370 (N_17370,N_16103,N_16600);
and U17371 (N_17371,N_16097,N_16054);
and U17372 (N_17372,N_16083,N_16955);
or U17373 (N_17373,N_16279,N_16851);
nor U17374 (N_17374,N_16243,N_16041);
and U17375 (N_17375,N_16653,N_16811);
nand U17376 (N_17376,N_16496,N_16789);
nand U17377 (N_17377,N_16013,N_16759);
nor U17378 (N_17378,N_16211,N_16189);
or U17379 (N_17379,N_16234,N_16044);
nor U17380 (N_17380,N_16643,N_16988);
nor U17381 (N_17381,N_16589,N_16820);
nor U17382 (N_17382,N_16555,N_16201);
and U17383 (N_17383,N_16894,N_16205);
xnor U17384 (N_17384,N_16764,N_16457);
nor U17385 (N_17385,N_16481,N_16577);
or U17386 (N_17386,N_16063,N_16576);
or U17387 (N_17387,N_16899,N_16226);
nand U17388 (N_17388,N_16536,N_16708);
xor U17389 (N_17389,N_16878,N_16373);
nor U17390 (N_17390,N_16941,N_16468);
and U17391 (N_17391,N_16265,N_16100);
xnor U17392 (N_17392,N_16666,N_16181);
or U17393 (N_17393,N_16051,N_16750);
and U17394 (N_17394,N_16776,N_16121);
nor U17395 (N_17395,N_16700,N_16338);
or U17396 (N_17396,N_16718,N_16316);
and U17397 (N_17397,N_16309,N_16428);
and U17398 (N_17398,N_16785,N_16352);
xnor U17399 (N_17399,N_16686,N_16451);
or U17400 (N_17400,N_16245,N_16460);
nand U17401 (N_17401,N_16462,N_16172);
nand U17402 (N_17402,N_16578,N_16397);
or U17403 (N_17403,N_16609,N_16585);
nor U17404 (N_17404,N_16353,N_16896);
nor U17405 (N_17405,N_16627,N_16112);
xor U17406 (N_17406,N_16990,N_16034);
or U17407 (N_17407,N_16550,N_16475);
nor U17408 (N_17408,N_16530,N_16534);
and U17409 (N_17409,N_16928,N_16943);
and U17410 (N_17410,N_16821,N_16655);
or U17411 (N_17411,N_16751,N_16009);
nor U17412 (N_17412,N_16464,N_16752);
xor U17413 (N_17413,N_16828,N_16251);
or U17414 (N_17414,N_16628,N_16862);
or U17415 (N_17415,N_16175,N_16143);
nand U17416 (N_17416,N_16003,N_16236);
or U17417 (N_17417,N_16152,N_16603);
and U17418 (N_17418,N_16213,N_16367);
nand U17419 (N_17419,N_16790,N_16547);
xnor U17420 (N_17420,N_16769,N_16435);
xnor U17421 (N_17421,N_16402,N_16738);
nand U17422 (N_17422,N_16524,N_16916);
nand U17423 (N_17423,N_16342,N_16514);
nor U17424 (N_17424,N_16614,N_16299);
xor U17425 (N_17425,N_16760,N_16214);
nand U17426 (N_17426,N_16659,N_16117);
or U17427 (N_17427,N_16301,N_16080);
and U17428 (N_17428,N_16157,N_16102);
nor U17429 (N_17429,N_16814,N_16354);
xor U17430 (N_17430,N_16558,N_16673);
or U17431 (N_17431,N_16487,N_16984);
nor U17432 (N_17432,N_16202,N_16141);
nor U17433 (N_17433,N_16361,N_16207);
nor U17434 (N_17434,N_16676,N_16183);
nor U17435 (N_17435,N_16580,N_16563);
and U17436 (N_17436,N_16281,N_16825);
nand U17437 (N_17437,N_16596,N_16951);
or U17438 (N_17438,N_16406,N_16678);
and U17439 (N_17439,N_16358,N_16139);
xor U17440 (N_17440,N_16248,N_16920);
or U17441 (N_17441,N_16125,N_16293);
and U17442 (N_17442,N_16931,N_16782);
xor U17443 (N_17443,N_16670,N_16164);
xor U17444 (N_17444,N_16218,N_16417);
nand U17445 (N_17445,N_16319,N_16897);
nor U17446 (N_17446,N_16042,N_16196);
nor U17447 (N_17447,N_16758,N_16171);
and U17448 (N_17448,N_16945,N_16835);
and U17449 (N_17449,N_16727,N_16028);
nand U17450 (N_17450,N_16506,N_16303);
and U17451 (N_17451,N_16150,N_16262);
nand U17452 (N_17452,N_16302,N_16869);
xor U17453 (N_17453,N_16719,N_16636);
nor U17454 (N_17454,N_16595,N_16379);
nand U17455 (N_17455,N_16797,N_16077);
and U17456 (N_17456,N_16873,N_16312);
nor U17457 (N_17457,N_16020,N_16364);
nand U17458 (N_17458,N_16089,N_16027);
and U17459 (N_17459,N_16741,N_16590);
or U17460 (N_17460,N_16520,N_16934);
nor U17461 (N_17461,N_16235,N_16389);
and U17462 (N_17462,N_16914,N_16932);
nand U17463 (N_17463,N_16325,N_16313);
and U17464 (N_17464,N_16942,N_16422);
nand U17465 (N_17465,N_16284,N_16068);
or U17466 (N_17466,N_16588,N_16375);
nor U17467 (N_17467,N_16037,N_16363);
nor U17468 (N_17468,N_16126,N_16276);
or U17469 (N_17469,N_16693,N_16842);
and U17470 (N_17470,N_16569,N_16995);
and U17471 (N_17471,N_16884,N_16383);
and U17472 (N_17472,N_16409,N_16419);
or U17473 (N_17473,N_16011,N_16317);
and U17474 (N_17474,N_16648,N_16640);
and U17475 (N_17475,N_16072,N_16566);
or U17476 (N_17476,N_16561,N_16193);
nor U17477 (N_17477,N_16622,N_16022);
nand U17478 (N_17478,N_16948,N_16618);
or U17479 (N_17479,N_16722,N_16624);
nand U17480 (N_17480,N_16275,N_16637);
nor U17481 (N_17481,N_16061,N_16249);
or U17482 (N_17482,N_16134,N_16200);
xor U17483 (N_17483,N_16893,N_16483);
xnor U17484 (N_17484,N_16391,N_16538);
xor U17485 (N_17485,N_16127,N_16983);
nand U17486 (N_17486,N_16860,N_16513);
nand U17487 (N_17487,N_16773,N_16198);
nor U17488 (N_17488,N_16885,N_16777);
nand U17489 (N_17489,N_16824,N_16447);
nand U17490 (N_17490,N_16240,N_16326);
nand U17491 (N_17491,N_16393,N_16049);
nor U17492 (N_17492,N_16144,N_16615);
or U17493 (N_17493,N_16469,N_16705);
nand U17494 (N_17494,N_16456,N_16737);
nor U17495 (N_17495,N_16803,N_16662);
nor U17496 (N_17496,N_16909,N_16531);
or U17497 (N_17497,N_16414,N_16710);
nand U17498 (N_17498,N_16888,N_16222);
nand U17499 (N_17499,N_16053,N_16241);
nand U17500 (N_17500,N_16891,N_16414);
and U17501 (N_17501,N_16823,N_16748);
or U17502 (N_17502,N_16019,N_16817);
nand U17503 (N_17503,N_16093,N_16671);
nand U17504 (N_17504,N_16335,N_16641);
nand U17505 (N_17505,N_16050,N_16974);
xor U17506 (N_17506,N_16727,N_16358);
or U17507 (N_17507,N_16919,N_16037);
or U17508 (N_17508,N_16537,N_16713);
and U17509 (N_17509,N_16573,N_16704);
nand U17510 (N_17510,N_16637,N_16272);
nand U17511 (N_17511,N_16749,N_16901);
nor U17512 (N_17512,N_16467,N_16989);
xor U17513 (N_17513,N_16158,N_16743);
nand U17514 (N_17514,N_16858,N_16974);
and U17515 (N_17515,N_16597,N_16407);
nand U17516 (N_17516,N_16006,N_16406);
nand U17517 (N_17517,N_16065,N_16536);
xnor U17518 (N_17518,N_16309,N_16923);
nand U17519 (N_17519,N_16905,N_16619);
nor U17520 (N_17520,N_16186,N_16804);
and U17521 (N_17521,N_16272,N_16091);
xor U17522 (N_17522,N_16820,N_16359);
or U17523 (N_17523,N_16700,N_16047);
and U17524 (N_17524,N_16814,N_16038);
xnor U17525 (N_17525,N_16006,N_16576);
or U17526 (N_17526,N_16471,N_16514);
nor U17527 (N_17527,N_16716,N_16060);
and U17528 (N_17528,N_16519,N_16701);
or U17529 (N_17529,N_16836,N_16786);
nand U17530 (N_17530,N_16260,N_16651);
nor U17531 (N_17531,N_16402,N_16417);
xnor U17532 (N_17532,N_16918,N_16729);
or U17533 (N_17533,N_16078,N_16358);
xnor U17534 (N_17534,N_16857,N_16951);
nor U17535 (N_17535,N_16472,N_16996);
xor U17536 (N_17536,N_16633,N_16731);
and U17537 (N_17537,N_16079,N_16980);
and U17538 (N_17538,N_16957,N_16381);
xnor U17539 (N_17539,N_16572,N_16147);
nand U17540 (N_17540,N_16493,N_16029);
or U17541 (N_17541,N_16808,N_16321);
or U17542 (N_17542,N_16935,N_16323);
and U17543 (N_17543,N_16289,N_16559);
nor U17544 (N_17544,N_16160,N_16298);
xor U17545 (N_17545,N_16868,N_16367);
nand U17546 (N_17546,N_16483,N_16325);
nor U17547 (N_17547,N_16237,N_16840);
nor U17548 (N_17548,N_16291,N_16155);
nand U17549 (N_17549,N_16530,N_16500);
nor U17550 (N_17550,N_16334,N_16504);
nor U17551 (N_17551,N_16974,N_16838);
and U17552 (N_17552,N_16432,N_16356);
nand U17553 (N_17553,N_16509,N_16457);
nor U17554 (N_17554,N_16558,N_16344);
xor U17555 (N_17555,N_16095,N_16839);
nand U17556 (N_17556,N_16300,N_16163);
nand U17557 (N_17557,N_16115,N_16728);
xor U17558 (N_17558,N_16744,N_16268);
and U17559 (N_17559,N_16518,N_16315);
xor U17560 (N_17560,N_16317,N_16616);
xor U17561 (N_17561,N_16366,N_16886);
nand U17562 (N_17562,N_16026,N_16932);
xnor U17563 (N_17563,N_16753,N_16234);
and U17564 (N_17564,N_16603,N_16118);
xor U17565 (N_17565,N_16205,N_16942);
nand U17566 (N_17566,N_16624,N_16486);
and U17567 (N_17567,N_16262,N_16555);
and U17568 (N_17568,N_16558,N_16387);
xnor U17569 (N_17569,N_16745,N_16292);
and U17570 (N_17570,N_16040,N_16307);
and U17571 (N_17571,N_16836,N_16099);
and U17572 (N_17572,N_16350,N_16925);
nor U17573 (N_17573,N_16942,N_16945);
nor U17574 (N_17574,N_16148,N_16593);
and U17575 (N_17575,N_16502,N_16171);
or U17576 (N_17576,N_16910,N_16572);
or U17577 (N_17577,N_16062,N_16881);
xor U17578 (N_17578,N_16784,N_16993);
and U17579 (N_17579,N_16055,N_16270);
and U17580 (N_17580,N_16820,N_16008);
xor U17581 (N_17581,N_16427,N_16772);
nand U17582 (N_17582,N_16980,N_16734);
nor U17583 (N_17583,N_16821,N_16851);
or U17584 (N_17584,N_16135,N_16230);
and U17585 (N_17585,N_16189,N_16202);
and U17586 (N_17586,N_16265,N_16409);
and U17587 (N_17587,N_16093,N_16160);
and U17588 (N_17588,N_16132,N_16358);
and U17589 (N_17589,N_16407,N_16595);
and U17590 (N_17590,N_16073,N_16281);
and U17591 (N_17591,N_16573,N_16778);
xor U17592 (N_17592,N_16670,N_16786);
nor U17593 (N_17593,N_16575,N_16379);
xor U17594 (N_17594,N_16059,N_16463);
nor U17595 (N_17595,N_16347,N_16358);
and U17596 (N_17596,N_16182,N_16826);
xnor U17597 (N_17597,N_16738,N_16243);
and U17598 (N_17598,N_16176,N_16076);
and U17599 (N_17599,N_16776,N_16115);
and U17600 (N_17600,N_16923,N_16218);
and U17601 (N_17601,N_16444,N_16218);
or U17602 (N_17602,N_16739,N_16451);
xnor U17603 (N_17603,N_16687,N_16543);
nor U17604 (N_17604,N_16320,N_16483);
and U17605 (N_17605,N_16596,N_16180);
xor U17606 (N_17606,N_16275,N_16606);
xnor U17607 (N_17607,N_16073,N_16225);
xor U17608 (N_17608,N_16732,N_16755);
xor U17609 (N_17609,N_16404,N_16715);
xnor U17610 (N_17610,N_16695,N_16563);
or U17611 (N_17611,N_16812,N_16155);
nor U17612 (N_17612,N_16885,N_16196);
xnor U17613 (N_17613,N_16378,N_16422);
and U17614 (N_17614,N_16049,N_16503);
nor U17615 (N_17615,N_16194,N_16195);
nor U17616 (N_17616,N_16516,N_16774);
nor U17617 (N_17617,N_16390,N_16279);
or U17618 (N_17618,N_16514,N_16152);
or U17619 (N_17619,N_16733,N_16716);
nand U17620 (N_17620,N_16470,N_16394);
nor U17621 (N_17621,N_16329,N_16181);
xnor U17622 (N_17622,N_16986,N_16909);
nor U17623 (N_17623,N_16540,N_16350);
nor U17624 (N_17624,N_16627,N_16651);
xnor U17625 (N_17625,N_16188,N_16958);
xnor U17626 (N_17626,N_16163,N_16446);
nor U17627 (N_17627,N_16870,N_16307);
and U17628 (N_17628,N_16069,N_16342);
nand U17629 (N_17629,N_16593,N_16336);
nand U17630 (N_17630,N_16098,N_16237);
nor U17631 (N_17631,N_16757,N_16737);
or U17632 (N_17632,N_16016,N_16518);
or U17633 (N_17633,N_16794,N_16401);
or U17634 (N_17634,N_16470,N_16400);
nand U17635 (N_17635,N_16225,N_16221);
nand U17636 (N_17636,N_16042,N_16720);
and U17637 (N_17637,N_16829,N_16464);
or U17638 (N_17638,N_16043,N_16093);
and U17639 (N_17639,N_16819,N_16614);
or U17640 (N_17640,N_16197,N_16271);
nor U17641 (N_17641,N_16797,N_16384);
xor U17642 (N_17642,N_16191,N_16199);
and U17643 (N_17643,N_16775,N_16419);
nor U17644 (N_17644,N_16235,N_16126);
nor U17645 (N_17645,N_16083,N_16594);
and U17646 (N_17646,N_16644,N_16688);
nor U17647 (N_17647,N_16134,N_16097);
and U17648 (N_17648,N_16329,N_16317);
or U17649 (N_17649,N_16068,N_16519);
and U17650 (N_17650,N_16103,N_16299);
xor U17651 (N_17651,N_16761,N_16046);
nor U17652 (N_17652,N_16156,N_16533);
xor U17653 (N_17653,N_16389,N_16557);
xor U17654 (N_17654,N_16638,N_16771);
nand U17655 (N_17655,N_16243,N_16797);
or U17656 (N_17656,N_16145,N_16938);
nand U17657 (N_17657,N_16299,N_16483);
nand U17658 (N_17658,N_16736,N_16884);
or U17659 (N_17659,N_16469,N_16637);
or U17660 (N_17660,N_16990,N_16410);
xor U17661 (N_17661,N_16705,N_16959);
or U17662 (N_17662,N_16647,N_16558);
or U17663 (N_17663,N_16933,N_16169);
nand U17664 (N_17664,N_16706,N_16359);
or U17665 (N_17665,N_16839,N_16535);
or U17666 (N_17666,N_16734,N_16431);
nand U17667 (N_17667,N_16784,N_16681);
and U17668 (N_17668,N_16658,N_16876);
nand U17669 (N_17669,N_16092,N_16660);
or U17670 (N_17670,N_16245,N_16486);
xor U17671 (N_17671,N_16076,N_16072);
nand U17672 (N_17672,N_16914,N_16213);
xor U17673 (N_17673,N_16062,N_16469);
xnor U17674 (N_17674,N_16693,N_16502);
xnor U17675 (N_17675,N_16935,N_16808);
nor U17676 (N_17676,N_16414,N_16455);
nand U17677 (N_17677,N_16282,N_16499);
nor U17678 (N_17678,N_16108,N_16748);
nand U17679 (N_17679,N_16497,N_16242);
or U17680 (N_17680,N_16636,N_16642);
nor U17681 (N_17681,N_16623,N_16328);
nand U17682 (N_17682,N_16969,N_16070);
nor U17683 (N_17683,N_16730,N_16183);
and U17684 (N_17684,N_16953,N_16610);
or U17685 (N_17685,N_16686,N_16064);
and U17686 (N_17686,N_16134,N_16711);
nand U17687 (N_17687,N_16697,N_16336);
and U17688 (N_17688,N_16171,N_16163);
and U17689 (N_17689,N_16470,N_16926);
and U17690 (N_17690,N_16404,N_16806);
and U17691 (N_17691,N_16766,N_16480);
nand U17692 (N_17692,N_16880,N_16405);
or U17693 (N_17693,N_16089,N_16431);
xor U17694 (N_17694,N_16858,N_16345);
nand U17695 (N_17695,N_16540,N_16367);
nor U17696 (N_17696,N_16305,N_16517);
xor U17697 (N_17697,N_16175,N_16169);
nor U17698 (N_17698,N_16879,N_16812);
xor U17699 (N_17699,N_16922,N_16443);
nor U17700 (N_17700,N_16883,N_16820);
nand U17701 (N_17701,N_16016,N_16749);
nor U17702 (N_17702,N_16426,N_16657);
xor U17703 (N_17703,N_16517,N_16930);
and U17704 (N_17704,N_16813,N_16457);
xnor U17705 (N_17705,N_16596,N_16692);
and U17706 (N_17706,N_16084,N_16178);
and U17707 (N_17707,N_16059,N_16138);
xnor U17708 (N_17708,N_16806,N_16220);
or U17709 (N_17709,N_16347,N_16605);
nor U17710 (N_17710,N_16174,N_16411);
xor U17711 (N_17711,N_16977,N_16323);
nand U17712 (N_17712,N_16349,N_16298);
or U17713 (N_17713,N_16416,N_16470);
nor U17714 (N_17714,N_16742,N_16886);
nor U17715 (N_17715,N_16631,N_16287);
and U17716 (N_17716,N_16422,N_16865);
or U17717 (N_17717,N_16757,N_16235);
nor U17718 (N_17718,N_16918,N_16673);
and U17719 (N_17719,N_16143,N_16450);
and U17720 (N_17720,N_16618,N_16020);
nand U17721 (N_17721,N_16088,N_16398);
or U17722 (N_17722,N_16981,N_16119);
nor U17723 (N_17723,N_16322,N_16923);
and U17724 (N_17724,N_16558,N_16056);
and U17725 (N_17725,N_16171,N_16343);
nor U17726 (N_17726,N_16358,N_16034);
or U17727 (N_17727,N_16807,N_16216);
xnor U17728 (N_17728,N_16880,N_16008);
nor U17729 (N_17729,N_16898,N_16573);
and U17730 (N_17730,N_16972,N_16079);
or U17731 (N_17731,N_16007,N_16625);
nor U17732 (N_17732,N_16735,N_16523);
xnor U17733 (N_17733,N_16285,N_16450);
xor U17734 (N_17734,N_16444,N_16317);
nand U17735 (N_17735,N_16574,N_16964);
nor U17736 (N_17736,N_16813,N_16278);
nand U17737 (N_17737,N_16303,N_16062);
nor U17738 (N_17738,N_16399,N_16178);
and U17739 (N_17739,N_16604,N_16844);
and U17740 (N_17740,N_16423,N_16927);
nand U17741 (N_17741,N_16597,N_16368);
xor U17742 (N_17742,N_16785,N_16979);
nor U17743 (N_17743,N_16214,N_16791);
nand U17744 (N_17744,N_16167,N_16424);
xnor U17745 (N_17745,N_16476,N_16263);
nor U17746 (N_17746,N_16901,N_16838);
nor U17747 (N_17747,N_16547,N_16655);
and U17748 (N_17748,N_16196,N_16915);
and U17749 (N_17749,N_16996,N_16543);
or U17750 (N_17750,N_16923,N_16826);
or U17751 (N_17751,N_16977,N_16488);
nor U17752 (N_17752,N_16988,N_16723);
and U17753 (N_17753,N_16083,N_16730);
nand U17754 (N_17754,N_16504,N_16385);
xnor U17755 (N_17755,N_16964,N_16806);
nor U17756 (N_17756,N_16642,N_16805);
and U17757 (N_17757,N_16086,N_16121);
or U17758 (N_17758,N_16357,N_16888);
or U17759 (N_17759,N_16197,N_16837);
nand U17760 (N_17760,N_16306,N_16102);
or U17761 (N_17761,N_16591,N_16756);
and U17762 (N_17762,N_16279,N_16550);
nor U17763 (N_17763,N_16890,N_16201);
nor U17764 (N_17764,N_16350,N_16784);
xnor U17765 (N_17765,N_16646,N_16376);
nand U17766 (N_17766,N_16804,N_16409);
xnor U17767 (N_17767,N_16378,N_16067);
xor U17768 (N_17768,N_16586,N_16659);
and U17769 (N_17769,N_16339,N_16347);
nand U17770 (N_17770,N_16026,N_16495);
nand U17771 (N_17771,N_16119,N_16343);
or U17772 (N_17772,N_16187,N_16779);
xor U17773 (N_17773,N_16385,N_16583);
or U17774 (N_17774,N_16743,N_16049);
or U17775 (N_17775,N_16621,N_16130);
nand U17776 (N_17776,N_16676,N_16086);
nor U17777 (N_17777,N_16245,N_16947);
xor U17778 (N_17778,N_16801,N_16443);
xnor U17779 (N_17779,N_16642,N_16929);
and U17780 (N_17780,N_16794,N_16214);
nand U17781 (N_17781,N_16476,N_16945);
xnor U17782 (N_17782,N_16222,N_16395);
or U17783 (N_17783,N_16281,N_16734);
nand U17784 (N_17784,N_16831,N_16265);
nor U17785 (N_17785,N_16085,N_16493);
nand U17786 (N_17786,N_16276,N_16611);
nor U17787 (N_17787,N_16156,N_16329);
or U17788 (N_17788,N_16007,N_16060);
and U17789 (N_17789,N_16559,N_16956);
and U17790 (N_17790,N_16797,N_16496);
or U17791 (N_17791,N_16122,N_16774);
xor U17792 (N_17792,N_16101,N_16284);
and U17793 (N_17793,N_16043,N_16951);
or U17794 (N_17794,N_16545,N_16040);
nand U17795 (N_17795,N_16113,N_16915);
or U17796 (N_17796,N_16839,N_16200);
nor U17797 (N_17797,N_16904,N_16336);
xor U17798 (N_17798,N_16292,N_16056);
nand U17799 (N_17799,N_16560,N_16431);
xnor U17800 (N_17800,N_16977,N_16487);
and U17801 (N_17801,N_16036,N_16412);
nand U17802 (N_17802,N_16072,N_16947);
or U17803 (N_17803,N_16429,N_16605);
or U17804 (N_17804,N_16487,N_16999);
nor U17805 (N_17805,N_16432,N_16017);
and U17806 (N_17806,N_16158,N_16658);
and U17807 (N_17807,N_16287,N_16400);
nand U17808 (N_17808,N_16392,N_16845);
nor U17809 (N_17809,N_16430,N_16090);
nand U17810 (N_17810,N_16607,N_16267);
nand U17811 (N_17811,N_16398,N_16868);
xnor U17812 (N_17812,N_16964,N_16619);
and U17813 (N_17813,N_16002,N_16057);
and U17814 (N_17814,N_16647,N_16848);
nor U17815 (N_17815,N_16116,N_16123);
xnor U17816 (N_17816,N_16791,N_16635);
xor U17817 (N_17817,N_16472,N_16029);
nor U17818 (N_17818,N_16089,N_16140);
nor U17819 (N_17819,N_16667,N_16500);
or U17820 (N_17820,N_16776,N_16320);
and U17821 (N_17821,N_16365,N_16370);
and U17822 (N_17822,N_16969,N_16366);
or U17823 (N_17823,N_16890,N_16313);
and U17824 (N_17824,N_16626,N_16768);
and U17825 (N_17825,N_16169,N_16394);
or U17826 (N_17826,N_16934,N_16030);
and U17827 (N_17827,N_16912,N_16611);
xor U17828 (N_17828,N_16707,N_16037);
nor U17829 (N_17829,N_16315,N_16879);
and U17830 (N_17830,N_16637,N_16180);
nand U17831 (N_17831,N_16250,N_16515);
xnor U17832 (N_17832,N_16476,N_16607);
and U17833 (N_17833,N_16451,N_16933);
xor U17834 (N_17834,N_16204,N_16486);
nor U17835 (N_17835,N_16568,N_16752);
and U17836 (N_17836,N_16732,N_16122);
and U17837 (N_17837,N_16496,N_16170);
xor U17838 (N_17838,N_16504,N_16834);
nand U17839 (N_17839,N_16120,N_16701);
nand U17840 (N_17840,N_16599,N_16653);
xnor U17841 (N_17841,N_16858,N_16246);
and U17842 (N_17842,N_16522,N_16644);
nor U17843 (N_17843,N_16550,N_16564);
xnor U17844 (N_17844,N_16145,N_16307);
nand U17845 (N_17845,N_16874,N_16343);
xnor U17846 (N_17846,N_16339,N_16791);
nand U17847 (N_17847,N_16402,N_16497);
or U17848 (N_17848,N_16293,N_16421);
and U17849 (N_17849,N_16082,N_16895);
nand U17850 (N_17850,N_16354,N_16958);
nor U17851 (N_17851,N_16606,N_16965);
and U17852 (N_17852,N_16210,N_16266);
or U17853 (N_17853,N_16689,N_16941);
and U17854 (N_17854,N_16837,N_16684);
nor U17855 (N_17855,N_16896,N_16780);
nand U17856 (N_17856,N_16159,N_16829);
xor U17857 (N_17857,N_16646,N_16463);
nor U17858 (N_17858,N_16413,N_16684);
and U17859 (N_17859,N_16216,N_16798);
nor U17860 (N_17860,N_16874,N_16830);
xnor U17861 (N_17861,N_16202,N_16407);
and U17862 (N_17862,N_16537,N_16833);
nand U17863 (N_17863,N_16191,N_16251);
nor U17864 (N_17864,N_16524,N_16797);
nor U17865 (N_17865,N_16739,N_16185);
and U17866 (N_17866,N_16837,N_16240);
and U17867 (N_17867,N_16925,N_16969);
and U17868 (N_17868,N_16468,N_16721);
nand U17869 (N_17869,N_16399,N_16793);
nand U17870 (N_17870,N_16920,N_16158);
nor U17871 (N_17871,N_16287,N_16923);
nor U17872 (N_17872,N_16603,N_16726);
nor U17873 (N_17873,N_16749,N_16820);
nor U17874 (N_17874,N_16176,N_16769);
xnor U17875 (N_17875,N_16967,N_16031);
or U17876 (N_17876,N_16030,N_16033);
xor U17877 (N_17877,N_16271,N_16039);
xor U17878 (N_17878,N_16807,N_16543);
xnor U17879 (N_17879,N_16995,N_16253);
nand U17880 (N_17880,N_16298,N_16989);
xnor U17881 (N_17881,N_16888,N_16683);
and U17882 (N_17882,N_16977,N_16932);
xnor U17883 (N_17883,N_16900,N_16236);
or U17884 (N_17884,N_16928,N_16330);
nor U17885 (N_17885,N_16089,N_16462);
or U17886 (N_17886,N_16545,N_16839);
xor U17887 (N_17887,N_16942,N_16585);
nor U17888 (N_17888,N_16584,N_16750);
or U17889 (N_17889,N_16274,N_16135);
nand U17890 (N_17890,N_16119,N_16645);
xor U17891 (N_17891,N_16022,N_16547);
or U17892 (N_17892,N_16628,N_16824);
xor U17893 (N_17893,N_16850,N_16882);
and U17894 (N_17894,N_16796,N_16040);
and U17895 (N_17895,N_16017,N_16842);
or U17896 (N_17896,N_16213,N_16011);
or U17897 (N_17897,N_16655,N_16687);
nor U17898 (N_17898,N_16006,N_16960);
nand U17899 (N_17899,N_16481,N_16798);
xnor U17900 (N_17900,N_16875,N_16651);
or U17901 (N_17901,N_16521,N_16810);
and U17902 (N_17902,N_16306,N_16900);
and U17903 (N_17903,N_16581,N_16013);
xor U17904 (N_17904,N_16893,N_16719);
nor U17905 (N_17905,N_16090,N_16995);
or U17906 (N_17906,N_16478,N_16246);
or U17907 (N_17907,N_16628,N_16142);
and U17908 (N_17908,N_16019,N_16754);
xor U17909 (N_17909,N_16544,N_16766);
nor U17910 (N_17910,N_16324,N_16845);
and U17911 (N_17911,N_16281,N_16193);
and U17912 (N_17912,N_16673,N_16139);
and U17913 (N_17913,N_16616,N_16215);
nand U17914 (N_17914,N_16637,N_16172);
and U17915 (N_17915,N_16604,N_16636);
and U17916 (N_17916,N_16199,N_16543);
nand U17917 (N_17917,N_16479,N_16828);
or U17918 (N_17918,N_16916,N_16541);
nand U17919 (N_17919,N_16700,N_16276);
nand U17920 (N_17920,N_16681,N_16642);
nand U17921 (N_17921,N_16880,N_16312);
and U17922 (N_17922,N_16176,N_16809);
and U17923 (N_17923,N_16518,N_16103);
or U17924 (N_17924,N_16640,N_16179);
xnor U17925 (N_17925,N_16852,N_16372);
nor U17926 (N_17926,N_16125,N_16747);
or U17927 (N_17927,N_16362,N_16205);
xnor U17928 (N_17928,N_16888,N_16057);
or U17929 (N_17929,N_16704,N_16481);
xor U17930 (N_17930,N_16896,N_16491);
or U17931 (N_17931,N_16515,N_16554);
or U17932 (N_17932,N_16768,N_16656);
nor U17933 (N_17933,N_16629,N_16554);
xor U17934 (N_17934,N_16919,N_16926);
nand U17935 (N_17935,N_16906,N_16273);
nand U17936 (N_17936,N_16037,N_16961);
nor U17937 (N_17937,N_16661,N_16551);
and U17938 (N_17938,N_16930,N_16714);
nand U17939 (N_17939,N_16354,N_16443);
or U17940 (N_17940,N_16353,N_16984);
nor U17941 (N_17941,N_16855,N_16129);
or U17942 (N_17942,N_16450,N_16178);
nor U17943 (N_17943,N_16924,N_16797);
nand U17944 (N_17944,N_16854,N_16864);
xor U17945 (N_17945,N_16719,N_16086);
nand U17946 (N_17946,N_16560,N_16191);
xnor U17947 (N_17947,N_16334,N_16487);
nand U17948 (N_17948,N_16999,N_16988);
xnor U17949 (N_17949,N_16358,N_16272);
and U17950 (N_17950,N_16554,N_16149);
nand U17951 (N_17951,N_16963,N_16203);
or U17952 (N_17952,N_16120,N_16734);
and U17953 (N_17953,N_16144,N_16559);
or U17954 (N_17954,N_16891,N_16932);
nor U17955 (N_17955,N_16051,N_16280);
nand U17956 (N_17956,N_16259,N_16595);
and U17957 (N_17957,N_16474,N_16635);
nor U17958 (N_17958,N_16399,N_16850);
or U17959 (N_17959,N_16586,N_16554);
xnor U17960 (N_17960,N_16873,N_16755);
xor U17961 (N_17961,N_16038,N_16459);
nor U17962 (N_17962,N_16633,N_16924);
or U17963 (N_17963,N_16507,N_16750);
nand U17964 (N_17964,N_16380,N_16865);
nand U17965 (N_17965,N_16274,N_16183);
xnor U17966 (N_17966,N_16287,N_16134);
nor U17967 (N_17967,N_16864,N_16067);
xnor U17968 (N_17968,N_16876,N_16915);
and U17969 (N_17969,N_16318,N_16839);
and U17970 (N_17970,N_16503,N_16907);
and U17971 (N_17971,N_16043,N_16129);
or U17972 (N_17972,N_16688,N_16452);
nor U17973 (N_17973,N_16792,N_16848);
or U17974 (N_17974,N_16799,N_16222);
nor U17975 (N_17975,N_16541,N_16174);
and U17976 (N_17976,N_16840,N_16108);
and U17977 (N_17977,N_16020,N_16788);
xor U17978 (N_17978,N_16744,N_16680);
xor U17979 (N_17979,N_16782,N_16839);
nor U17980 (N_17980,N_16913,N_16551);
and U17981 (N_17981,N_16285,N_16657);
or U17982 (N_17982,N_16461,N_16244);
xnor U17983 (N_17983,N_16527,N_16035);
and U17984 (N_17984,N_16737,N_16351);
nand U17985 (N_17985,N_16009,N_16284);
or U17986 (N_17986,N_16661,N_16765);
nor U17987 (N_17987,N_16230,N_16269);
nand U17988 (N_17988,N_16064,N_16798);
and U17989 (N_17989,N_16465,N_16138);
and U17990 (N_17990,N_16943,N_16867);
xnor U17991 (N_17991,N_16337,N_16666);
xor U17992 (N_17992,N_16374,N_16286);
xnor U17993 (N_17993,N_16036,N_16739);
nor U17994 (N_17994,N_16617,N_16968);
or U17995 (N_17995,N_16108,N_16389);
or U17996 (N_17996,N_16611,N_16483);
nor U17997 (N_17997,N_16839,N_16701);
nand U17998 (N_17998,N_16986,N_16731);
xnor U17999 (N_17999,N_16870,N_16839);
or U18000 (N_18000,N_17872,N_17821);
or U18001 (N_18001,N_17622,N_17077);
nand U18002 (N_18002,N_17048,N_17595);
nor U18003 (N_18003,N_17024,N_17900);
xnor U18004 (N_18004,N_17800,N_17239);
xor U18005 (N_18005,N_17925,N_17798);
and U18006 (N_18006,N_17807,N_17736);
or U18007 (N_18007,N_17747,N_17316);
nor U18008 (N_18008,N_17149,N_17330);
nand U18009 (N_18009,N_17792,N_17573);
or U18010 (N_18010,N_17210,N_17170);
xor U18011 (N_18011,N_17655,N_17213);
nand U18012 (N_18012,N_17547,N_17556);
and U18013 (N_18013,N_17723,N_17388);
and U18014 (N_18014,N_17776,N_17649);
nand U18015 (N_18015,N_17587,N_17298);
nor U18016 (N_18016,N_17047,N_17322);
and U18017 (N_18017,N_17893,N_17232);
nand U18018 (N_18018,N_17916,N_17613);
or U18019 (N_18019,N_17257,N_17791);
nor U18020 (N_18020,N_17191,N_17721);
nor U18021 (N_18021,N_17460,N_17419);
xor U18022 (N_18022,N_17100,N_17690);
nand U18023 (N_18023,N_17069,N_17135);
or U18024 (N_18024,N_17007,N_17430);
nand U18025 (N_18025,N_17078,N_17778);
or U18026 (N_18026,N_17852,N_17718);
xnor U18027 (N_18027,N_17891,N_17114);
nor U18028 (N_18028,N_17770,N_17489);
nand U18029 (N_18029,N_17625,N_17981);
nor U18030 (N_18030,N_17096,N_17699);
or U18031 (N_18031,N_17890,N_17968);
xor U18032 (N_18032,N_17246,N_17766);
or U18033 (N_18033,N_17666,N_17409);
nor U18034 (N_18034,N_17739,N_17932);
or U18035 (N_18035,N_17612,N_17802);
xnor U18036 (N_18036,N_17695,N_17864);
nand U18037 (N_18037,N_17041,N_17976);
nand U18038 (N_18038,N_17299,N_17339);
and U18039 (N_18039,N_17089,N_17144);
or U18040 (N_18040,N_17860,N_17727);
xnor U18041 (N_18041,N_17532,N_17597);
nand U18042 (N_18042,N_17657,N_17518);
nor U18043 (N_18043,N_17970,N_17995);
or U18044 (N_18044,N_17407,N_17732);
or U18045 (N_18045,N_17901,N_17992);
and U18046 (N_18046,N_17468,N_17974);
xnor U18047 (N_18047,N_17383,N_17725);
nor U18048 (N_18048,N_17125,N_17618);
nor U18049 (N_18049,N_17762,N_17260);
xor U18050 (N_18050,N_17351,N_17504);
xor U18051 (N_18051,N_17331,N_17895);
or U18052 (N_18052,N_17334,N_17876);
and U18053 (N_18053,N_17865,N_17009);
nor U18054 (N_18054,N_17417,N_17245);
xor U18055 (N_18055,N_17352,N_17459);
nand U18056 (N_18056,N_17844,N_17400);
or U18057 (N_18057,N_17730,N_17101);
nor U18058 (N_18058,N_17643,N_17415);
nand U18059 (N_18059,N_17359,N_17190);
nor U18060 (N_18060,N_17584,N_17606);
nor U18061 (N_18061,N_17122,N_17814);
nor U18062 (N_18062,N_17054,N_17517);
nor U18063 (N_18063,N_17989,N_17343);
or U18064 (N_18064,N_17617,N_17534);
or U18065 (N_18065,N_17759,N_17332);
nand U18066 (N_18066,N_17464,N_17526);
nand U18067 (N_18067,N_17551,N_17710);
nand U18068 (N_18068,N_17471,N_17083);
xnor U18069 (N_18069,N_17010,N_17368);
or U18070 (N_18070,N_17060,N_17871);
and U18071 (N_18071,N_17071,N_17775);
and U18072 (N_18072,N_17544,N_17425);
nand U18073 (N_18073,N_17001,N_17877);
nor U18074 (N_18074,N_17495,N_17093);
xnor U18075 (N_18075,N_17307,N_17636);
nand U18076 (N_18076,N_17769,N_17683);
or U18077 (N_18077,N_17333,N_17022);
xor U18078 (N_18078,N_17528,N_17050);
nand U18079 (N_18079,N_17867,N_17401);
nor U18080 (N_18080,N_17261,N_17420);
nor U18081 (N_18081,N_17574,N_17212);
and U18082 (N_18082,N_17218,N_17930);
nor U18083 (N_18083,N_17475,N_17315);
or U18084 (N_18084,N_17196,N_17520);
or U18085 (N_18085,N_17529,N_17158);
and U18086 (N_18086,N_17822,N_17364);
nor U18087 (N_18087,N_17441,N_17107);
or U18088 (N_18088,N_17066,N_17427);
xor U18089 (N_18089,N_17361,N_17244);
nor U18090 (N_18090,N_17395,N_17972);
nand U18091 (N_18091,N_17758,N_17812);
nor U18092 (N_18092,N_17494,N_17987);
or U18093 (N_18093,N_17026,N_17805);
or U18094 (N_18094,N_17373,N_17575);
xor U18095 (N_18095,N_17192,N_17102);
and U18096 (N_18096,N_17500,N_17788);
and U18097 (N_18097,N_17080,N_17946);
xnor U18098 (N_18098,N_17278,N_17920);
nor U18099 (N_18099,N_17248,N_17328);
nand U18100 (N_18100,N_17275,N_17112);
xnor U18101 (N_18101,N_17304,N_17652);
nand U18102 (N_18102,N_17983,N_17028);
and U18103 (N_18103,N_17319,N_17450);
nor U18104 (N_18104,N_17085,N_17845);
xnor U18105 (N_18105,N_17883,N_17226);
and U18106 (N_18106,N_17340,N_17123);
nor U18107 (N_18107,N_17061,N_17169);
nor U18108 (N_18108,N_17011,N_17856);
or U18109 (N_18109,N_17961,N_17664);
nor U18110 (N_18110,N_17150,N_17729);
xnor U18111 (N_18111,N_17477,N_17111);
xnor U18112 (N_18112,N_17079,N_17233);
and U18113 (N_18113,N_17090,N_17252);
nand U18114 (N_18114,N_17672,N_17437);
nor U18115 (N_18115,N_17926,N_17851);
or U18116 (N_18116,N_17473,N_17733);
nor U18117 (N_18117,N_17586,N_17660);
xor U18118 (N_18118,N_17157,N_17750);
nand U18119 (N_18119,N_17859,N_17939);
nand U18120 (N_18120,N_17493,N_17627);
nand U18121 (N_18121,N_17549,N_17915);
xnor U18122 (N_18122,N_17300,N_17043);
and U18123 (N_18123,N_17366,N_17578);
nor U18124 (N_18124,N_17843,N_17168);
and U18125 (N_18125,N_17786,N_17285);
nor U18126 (N_18126,N_17941,N_17422);
and U18127 (N_18127,N_17760,N_17507);
nand U18128 (N_18128,N_17969,N_17155);
and U18129 (N_18129,N_17580,N_17693);
nand U18130 (N_18130,N_17662,N_17200);
or U18131 (N_18131,N_17142,N_17839);
and U18132 (N_18132,N_17403,N_17677);
and U18133 (N_18133,N_17673,N_17658);
or U18134 (N_18134,N_17378,N_17633);
and U18135 (N_18135,N_17910,N_17572);
and U18136 (N_18136,N_17632,N_17385);
or U18137 (N_18137,N_17335,N_17737);
xnor U18138 (N_18138,N_17589,N_17076);
and U18139 (N_18139,N_17596,N_17120);
xor U18140 (N_18140,N_17785,N_17097);
xnor U18141 (N_18141,N_17313,N_17803);
or U18142 (N_18142,N_17341,N_17914);
nand U18143 (N_18143,N_17291,N_17431);
or U18144 (N_18144,N_17065,N_17832);
and U18145 (N_18145,N_17620,N_17002);
or U18146 (N_18146,N_17286,N_17855);
xnor U18147 (N_18147,N_17697,N_17647);
nand U18148 (N_18148,N_17035,N_17881);
or U18149 (N_18149,N_17588,N_17524);
nand U18150 (N_18150,N_17453,N_17131);
nand U18151 (N_18151,N_17519,N_17472);
or U18152 (N_18152,N_17499,N_17264);
xor U18153 (N_18153,N_17134,N_17945);
and U18154 (N_18154,N_17449,N_17282);
nand U18155 (N_18155,N_17645,N_17167);
or U18156 (N_18156,N_17317,N_17163);
nor U18157 (N_18157,N_17590,N_17204);
or U18158 (N_18158,N_17787,N_17846);
nand U18159 (N_18159,N_17074,N_17225);
and U18160 (N_18160,N_17370,N_17292);
xnor U18161 (N_18161,N_17908,N_17109);
or U18162 (N_18162,N_17016,N_17326);
nand U18163 (N_18163,N_17042,N_17132);
nor U18164 (N_18164,N_17862,N_17903);
nand U18165 (N_18165,N_17682,N_17906);
and U18166 (N_18166,N_17641,N_17140);
xor U18167 (N_18167,N_17369,N_17501);
nor U18168 (N_18168,N_17462,N_17861);
or U18169 (N_18169,N_17646,N_17553);
xnor U18170 (N_18170,N_17734,N_17583);
or U18171 (N_18171,N_17034,N_17508);
and U18172 (N_18172,N_17187,N_17301);
and U18173 (N_18173,N_17470,N_17988);
and U18174 (N_18174,N_17238,N_17503);
nor U18175 (N_18175,N_17779,N_17355);
nand U18176 (N_18176,N_17029,N_17297);
and U18177 (N_18177,N_17929,N_17365);
and U18178 (N_18178,N_17208,N_17560);
nor U18179 (N_18179,N_17160,N_17311);
nand U18180 (N_18180,N_17241,N_17438);
nor U18181 (N_18181,N_17189,N_17923);
or U18182 (N_18182,N_17581,N_17234);
nor U18183 (N_18183,N_17153,N_17406);
xor U18184 (N_18184,N_17804,N_17527);
nor U18185 (N_18185,N_17994,N_17990);
nor U18186 (N_18186,N_17303,N_17325);
nand U18187 (N_18187,N_17548,N_17767);
nor U18188 (N_18188,N_17428,N_17561);
nor U18189 (N_18189,N_17492,N_17392);
or U18190 (N_18190,N_17505,N_17512);
nand U18191 (N_18191,N_17336,N_17985);
xnor U18192 (N_18192,N_17774,N_17975);
and U18193 (N_18193,N_17514,N_17147);
xnor U18194 (N_18194,N_17094,N_17713);
xnor U18195 (N_18195,N_17413,N_17748);
or U18196 (N_18196,N_17886,N_17691);
nand U18197 (N_18197,N_17999,N_17654);
and U18198 (N_18198,N_17411,N_17497);
nand U18199 (N_18199,N_17562,N_17262);
and U18200 (N_18200,N_17907,N_17878);
and U18201 (N_18201,N_17899,N_17863);
nor U18202 (N_18202,N_17360,N_17138);
or U18203 (N_18203,N_17688,N_17379);
and U18204 (N_18204,N_17110,N_17746);
nor U18205 (N_18205,N_17712,N_17484);
nand U18206 (N_18206,N_17224,N_17457);
xor U18207 (N_18207,N_17087,N_17623);
xnor U18208 (N_18208,N_17092,N_17571);
and U18209 (N_18209,N_17817,N_17887);
or U18210 (N_18210,N_17741,N_17454);
nand U18211 (N_18211,N_17870,N_17040);
and U18212 (N_18212,N_17965,N_17585);
nand U18213 (N_18213,N_17854,N_17253);
nor U18214 (N_18214,N_17435,N_17393);
xor U18215 (N_18215,N_17025,N_17130);
or U18216 (N_18216,N_17781,N_17771);
and U18217 (N_18217,N_17919,N_17136);
nor U18218 (N_18218,N_17940,N_17717);
and U18219 (N_18219,N_17884,N_17266);
xor U18220 (N_18220,N_17117,N_17354);
nand U18221 (N_18221,N_17320,N_17698);
nor U18222 (N_18222,N_17115,N_17820);
or U18223 (N_18223,N_17591,N_17310);
and U18224 (N_18224,N_17963,N_17535);
or U18225 (N_18225,N_17849,N_17386);
xnor U18226 (N_18226,N_17638,N_17219);
nand U18227 (N_18227,N_17498,N_17557);
or U18228 (N_18228,N_17273,N_17897);
xor U18229 (N_18229,N_17530,N_17600);
nor U18230 (N_18230,N_17391,N_17440);
and U18231 (N_18231,N_17314,N_17467);
and U18232 (N_18232,N_17161,N_17305);
nand U18233 (N_18233,N_17108,N_17235);
or U18234 (N_18234,N_17382,N_17159);
or U18235 (N_18235,N_17829,N_17541);
nand U18236 (N_18236,N_17601,N_17938);
and U18237 (N_18237,N_17162,N_17452);
or U18238 (N_18238,N_17644,N_17840);
nor U18239 (N_18239,N_17823,N_17836);
and U18240 (N_18240,N_17979,N_17566);
and U18241 (N_18241,N_17599,N_17631);
xor U18242 (N_18242,N_17439,N_17934);
nand U18243 (N_18243,N_17116,N_17198);
nor U18244 (N_18244,N_17004,N_17991);
nand U18245 (N_18245,N_17461,N_17309);
or U18246 (N_18246,N_17081,N_17554);
and U18247 (N_18247,N_17014,N_17259);
and U18248 (N_18248,N_17609,N_17782);
or U18249 (N_18249,N_17476,N_17790);
nand U18250 (N_18250,N_17608,N_17429);
or U18251 (N_18251,N_17605,N_17312);
nor U18252 (N_18252,N_17318,N_17230);
nor U18253 (N_18253,N_17742,N_17152);
or U18254 (N_18254,N_17088,N_17242);
and U18255 (N_18255,N_17577,N_17099);
nor U18256 (N_18256,N_17833,N_17017);
and U18257 (N_18257,N_17251,N_17174);
or U18258 (N_18258,N_17521,N_17780);
or U18259 (N_18259,N_17686,N_17815);
or U18260 (N_18260,N_17045,N_17416);
or U18261 (N_18261,N_17199,N_17396);
and U18262 (N_18262,N_17055,N_17062);
nor U18263 (N_18263,N_17761,N_17270);
nor U18264 (N_18264,N_17955,N_17793);
and U18265 (N_18265,N_17496,N_17084);
xnor U18266 (N_18266,N_17276,N_17598);
nor U18267 (N_18267,N_17447,N_17070);
nor U18268 (N_18268,N_17768,N_17442);
nor U18269 (N_18269,N_17129,N_17831);
xor U18270 (N_18270,N_17372,N_17349);
and U18271 (N_18271,N_17185,N_17082);
and U18272 (N_18272,N_17894,N_17448);
xnor U18273 (N_18273,N_17667,N_17203);
nor U18274 (N_18274,N_17105,N_17651);
nor U18275 (N_18275,N_17342,N_17885);
xor U18276 (N_18276,N_17072,N_17258);
and U18277 (N_18277,N_17896,N_17942);
nor U18278 (N_18278,N_17801,N_17426);
and U18279 (N_18279,N_17446,N_17921);
nor U18280 (N_18280,N_17295,N_17306);
nand U18281 (N_18281,N_17058,N_17735);
xor U18282 (N_18282,N_17794,N_17656);
and U18283 (N_18283,N_17869,N_17337);
nor U18284 (N_18284,N_17931,N_17594);
and U18285 (N_18285,N_17329,N_17882);
and U18286 (N_18286,N_17952,N_17179);
or U18287 (N_18287,N_17231,N_17515);
nand U18288 (N_18288,N_17971,N_17949);
nor U18289 (N_18289,N_17338,N_17348);
or U18290 (N_18290,N_17480,N_17394);
xor U18291 (N_18291,N_17687,N_17380);
nand U18292 (N_18292,N_17937,N_17502);
nand U18293 (N_18293,N_17709,N_17175);
nand U18294 (N_18294,N_17513,N_17280);
nor U18295 (N_18295,N_17810,N_17182);
or U18296 (N_18296,N_17986,N_17956);
xnor U18297 (N_18297,N_17516,N_17640);
or U18298 (N_18298,N_17240,N_17954);
and U18299 (N_18299,N_17997,N_17127);
nor U18300 (N_18300,N_17121,N_17511);
xnor U18301 (N_18301,N_17487,N_17834);
xor U18302 (N_18302,N_17950,N_17145);
xor U18303 (N_18303,N_17694,N_17816);
xnor U18304 (N_18304,N_17616,N_17888);
or U18305 (N_18305,N_17183,N_17933);
xnor U18306 (N_18306,N_17249,N_17740);
xnor U18307 (N_18307,N_17113,N_17809);
or U18308 (N_18308,N_17481,N_17284);
or U18309 (N_18309,N_17255,N_17021);
or U18310 (N_18310,N_17243,N_17828);
and U18311 (N_18311,N_17165,N_17018);
xnor U18312 (N_18312,N_17263,N_17008);
or U18313 (N_18313,N_17023,N_17973);
and U18314 (N_18314,N_17483,N_17051);
or U18315 (N_18315,N_17716,N_17724);
nand U18316 (N_18316,N_17281,N_17172);
xor U18317 (N_18317,N_17924,N_17287);
xor U18318 (N_18318,N_17668,N_17764);
nand U18319 (N_18319,N_17387,N_17046);
xor U18320 (N_18320,N_17294,N_17247);
or U18321 (N_18321,N_17777,N_17648);
nor U18322 (N_18322,N_17271,N_17091);
nand U18323 (N_18323,N_17962,N_17033);
xor U18324 (N_18324,N_17133,N_17918);
xnor U18325 (N_18325,N_17818,N_17277);
xnor U18326 (N_18326,N_17993,N_17700);
or U18327 (N_18327,N_17958,N_17796);
nor U18328 (N_18328,N_17674,N_17509);
nand U18329 (N_18329,N_17565,N_17789);
nand U18330 (N_18330,N_17957,N_17478);
nand U18331 (N_18331,N_17059,N_17685);
xor U18332 (N_18332,N_17542,N_17948);
nor U18333 (N_18333,N_17754,N_17669);
nor U18334 (N_18334,N_17808,N_17289);
nor U18335 (N_18335,N_17848,N_17490);
and U18336 (N_18336,N_17722,N_17207);
and U18337 (N_18337,N_17098,N_17671);
nor U18338 (N_18338,N_17784,N_17272);
nor U18339 (N_18339,N_17569,N_17642);
and U18340 (N_18340,N_17902,N_17268);
xnor U18341 (N_18341,N_17592,N_17537);
xnor U18342 (N_18342,N_17593,N_17434);
nand U18343 (N_18343,N_17466,N_17824);
or U18344 (N_18344,N_17912,N_17491);
nand U18345 (N_18345,N_17838,N_17356);
xor U18346 (N_18346,N_17892,N_17728);
and U18347 (N_18347,N_17039,N_17486);
nand U18348 (N_18348,N_17719,N_17104);
and U18349 (N_18349,N_17536,N_17563);
and U18350 (N_18350,N_17012,N_17783);
and U18351 (N_18351,N_17753,N_17559);
nand U18352 (N_18352,N_17038,N_17659);
and U18353 (N_18353,N_17639,N_17205);
and U18354 (N_18354,N_17119,N_17015);
or U18355 (N_18355,N_17164,N_17269);
or U18356 (N_18356,N_17543,N_17423);
nand U18357 (N_18357,N_17607,N_17980);
or U18358 (N_18358,N_17582,N_17745);
or U18359 (N_18359,N_17917,N_17602);
nand U18360 (N_18360,N_17680,N_17692);
and U18361 (N_18361,N_17708,N_17755);
or U18362 (N_18362,N_17217,N_17103);
and U18363 (N_18363,N_17555,N_17184);
and U18364 (N_18364,N_17880,N_17397);
and U18365 (N_18365,N_17445,N_17194);
xor U18366 (N_18366,N_17837,N_17367);
nor U18367 (N_18367,N_17797,N_17650);
and U18368 (N_18368,N_17953,N_17178);
nand U18369 (N_18369,N_17951,N_17482);
xor U18370 (N_18370,N_17402,N_17675);
and U18371 (N_18371,N_17049,N_17064);
nor U18372 (N_18372,N_17321,N_17375);
nand U18373 (N_18373,N_17324,N_17531);
nor U18374 (N_18374,N_17567,N_17552);
nor U18375 (N_18375,N_17229,N_17538);
xnor U18376 (N_18376,N_17670,N_17209);
xnor U18377 (N_18377,N_17978,N_17384);
and U18378 (N_18378,N_17715,N_17465);
and U18379 (N_18379,N_17634,N_17889);
nor U18380 (N_18380,N_17635,N_17053);
nand U18381 (N_18381,N_17031,N_17546);
xnor U18382 (N_18382,N_17873,N_17463);
or U18383 (N_18383,N_17928,N_17180);
nand U18384 (N_18384,N_17827,N_17738);
or U18385 (N_18385,N_17381,N_17911);
nand U18386 (N_18386,N_17436,N_17626);
xor U18387 (N_18387,N_17705,N_17603);
nand U18388 (N_18388,N_17533,N_17410);
nand U18389 (N_18389,N_17086,N_17485);
nand U18390 (N_18390,N_17228,N_17451);
nand U18391 (N_18391,N_17960,N_17327);
or U18392 (N_18392,N_17433,N_17944);
nor U18393 (N_18393,N_17702,N_17371);
xor U18394 (N_18394,N_17663,N_17019);
nor U18395 (N_18395,N_17003,N_17274);
nor U18396 (N_18396,N_17146,N_17811);
and U18397 (N_18397,N_17000,N_17795);
nor U18398 (N_18398,N_17898,N_17703);
or U18399 (N_18399,N_17095,N_17414);
and U18400 (N_18400,N_17568,N_17236);
xor U18401 (N_18401,N_17220,N_17696);
xnor U18402 (N_18402,N_17570,N_17075);
or U18403 (N_18403,N_17267,N_17037);
nor U18404 (N_18404,N_17353,N_17265);
or U18405 (N_18405,N_17922,N_17128);
or U18406 (N_18406,N_17825,N_17510);
xnor U18407 (N_18407,N_17346,N_17357);
or U18408 (N_18408,N_17558,N_17154);
nor U18409 (N_18409,N_17399,N_17936);
xor U18410 (N_18410,N_17964,N_17506);
nand U18411 (N_18411,N_17068,N_17676);
and U18412 (N_18412,N_17756,N_17539);
nand U18413 (N_18413,N_17615,N_17689);
nor U18414 (N_18414,N_17665,N_17629);
nand U18415 (N_18415,N_17181,N_17614);
nor U18416 (N_18416,N_17679,N_17847);
nor U18417 (N_18417,N_17830,N_17412);
nor U18418 (N_18418,N_17904,N_17176);
nand U18419 (N_18419,N_17773,N_17148);
or U18420 (N_18420,N_17678,N_17522);
xor U18421 (N_18421,N_17935,N_17456);
or U18422 (N_18422,N_17604,N_17290);
xnor U18423 (N_18423,N_17661,N_17027);
xnor U18424 (N_18424,N_17905,N_17743);
nor U18425 (N_18425,N_17874,N_17850);
or U18426 (N_18426,N_17376,N_17799);
nor U18427 (N_18427,N_17044,N_17757);
nor U18428 (N_18428,N_17171,N_17458);
or U18429 (N_18429,N_17443,N_17813);
nor U18430 (N_18430,N_17432,N_17195);
or U18431 (N_18431,N_17474,N_17749);
and U18432 (N_18432,N_17706,N_17405);
and U18433 (N_18433,N_17841,N_17624);
nor U18434 (N_18434,N_17193,N_17374);
nand U18435 (N_18435,N_17030,N_17227);
and U18436 (N_18436,N_17222,N_17323);
or U18437 (N_18437,N_17424,N_17982);
and U18438 (N_18438,N_17469,N_17067);
or U18439 (N_18439,N_17576,N_17523);
xor U18440 (N_18440,N_17720,N_17826);
or U18441 (N_18441,N_17868,N_17765);
xnor U18442 (N_18442,N_17063,N_17488);
and U18443 (N_18443,N_17345,N_17350);
and U18444 (N_18444,N_17681,N_17610);
and U18445 (N_18445,N_17137,N_17126);
and U18446 (N_18446,N_17875,N_17418);
nand U18447 (N_18447,N_17927,N_17714);
xnor U18448 (N_18448,N_17106,N_17250);
nor U18449 (N_18449,N_17966,N_17835);
xnor U18450 (N_18450,N_17579,N_17806);
or U18451 (N_18451,N_17857,N_17545);
and U18452 (N_18452,N_17752,N_17052);
nor U18453 (N_18453,N_17173,N_17216);
nor U18454 (N_18454,N_17221,N_17637);
xor U18455 (N_18455,N_17197,N_17166);
nor U18456 (N_18456,N_17223,N_17621);
and U18457 (N_18457,N_17279,N_17684);
nor U18458 (N_18458,N_17005,N_17967);
xor U18459 (N_18459,N_17984,N_17141);
or U18460 (N_18460,N_17237,N_17996);
or U18461 (N_18461,N_17842,N_17751);
or U18462 (N_18462,N_17308,N_17288);
and U18463 (N_18463,N_17959,N_17214);
and U18464 (N_18464,N_17444,N_17977);
xnor U18465 (N_18465,N_17362,N_17377);
nor U18466 (N_18466,N_17711,N_17611);
and U18467 (N_18467,N_17143,N_17408);
and U18468 (N_18468,N_17731,N_17879);
nand U18469 (N_18469,N_17525,N_17866);
or U18470 (N_18470,N_17455,N_17177);
or U18471 (N_18471,N_17479,N_17032);
nand U18472 (N_18472,N_17256,N_17653);
or U18473 (N_18473,N_17701,N_17283);
nor U18474 (N_18474,N_17302,N_17540);
nor U18475 (N_18475,N_17772,N_17726);
nand U18476 (N_18476,N_17909,N_17215);
xor U18477 (N_18477,N_17628,N_17202);
nor U18478 (N_18478,N_17943,N_17390);
or U18479 (N_18479,N_17998,N_17550);
and U18480 (N_18480,N_17186,N_17254);
nand U18481 (N_18481,N_17358,N_17421);
or U18482 (N_18482,N_17057,N_17201);
nand U18483 (N_18483,N_17296,N_17744);
or U18484 (N_18484,N_17389,N_17564);
and U18485 (N_18485,N_17020,N_17619);
nand U18486 (N_18486,N_17704,N_17763);
and U18487 (N_18487,N_17206,N_17398);
and U18488 (N_18488,N_17947,N_17819);
nor U18489 (N_18489,N_17913,N_17006);
nand U18490 (N_18490,N_17156,N_17124);
and U18491 (N_18491,N_17211,N_17188);
and U18492 (N_18492,N_17404,N_17036);
nor U18493 (N_18493,N_17630,N_17363);
nor U18494 (N_18494,N_17293,N_17013);
or U18495 (N_18495,N_17056,N_17707);
nor U18496 (N_18496,N_17347,N_17151);
nand U18497 (N_18497,N_17853,N_17858);
nor U18498 (N_18498,N_17139,N_17344);
nand U18499 (N_18499,N_17073,N_17118);
and U18500 (N_18500,N_17330,N_17132);
or U18501 (N_18501,N_17858,N_17397);
nor U18502 (N_18502,N_17882,N_17754);
nor U18503 (N_18503,N_17947,N_17130);
and U18504 (N_18504,N_17823,N_17484);
xnor U18505 (N_18505,N_17261,N_17421);
nor U18506 (N_18506,N_17556,N_17095);
nor U18507 (N_18507,N_17643,N_17180);
and U18508 (N_18508,N_17635,N_17831);
nor U18509 (N_18509,N_17626,N_17908);
and U18510 (N_18510,N_17133,N_17775);
nand U18511 (N_18511,N_17109,N_17042);
nand U18512 (N_18512,N_17852,N_17445);
nand U18513 (N_18513,N_17006,N_17111);
or U18514 (N_18514,N_17547,N_17870);
or U18515 (N_18515,N_17828,N_17804);
nand U18516 (N_18516,N_17846,N_17875);
nor U18517 (N_18517,N_17237,N_17491);
and U18518 (N_18518,N_17822,N_17012);
and U18519 (N_18519,N_17313,N_17466);
nand U18520 (N_18520,N_17823,N_17979);
and U18521 (N_18521,N_17798,N_17945);
or U18522 (N_18522,N_17413,N_17312);
and U18523 (N_18523,N_17830,N_17648);
xnor U18524 (N_18524,N_17886,N_17582);
nor U18525 (N_18525,N_17211,N_17366);
or U18526 (N_18526,N_17404,N_17180);
or U18527 (N_18527,N_17190,N_17045);
xor U18528 (N_18528,N_17131,N_17591);
xor U18529 (N_18529,N_17077,N_17665);
xor U18530 (N_18530,N_17143,N_17260);
or U18531 (N_18531,N_17623,N_17422);
xnor U18532 (N_18532,N_17913,N_17360);
or U18533 (N_18533,N_17947,N_17418);
xor U18534 (N_18534,N_17250,N_17678);
or U18535 (N_18535,N_17723,N_17027);
nand U18536 (N_18536,N_17860,N_17571);
xor U18537 (N_18537,N_17612,N_17479);
or U18538 (N_18538,N_17493,N_17656);
and U18539 (N_18539,N_17477,N_17371);
nor U18540 (N_18540,N_17669,N_17212);
and U18541 (N_18541,N_17374,N_17710);
or U18542 (N_18542,N_17894,N_17722);
and U18543 (N_18543,N_17279,N_17038);
and U18544 (N_18544,N_17621,N_17327);
nand U18545 (N_18545,N_17115,N_17156);
xnor U18546 (N_18546,N_17004,N_17147);
and U18547 (N_18547,N_17828,N_17470);
nor U18548 (N_18548,N_17203,N_17176);
nor U18549 (N_18549,N_17962,N_17674);
or U18550 (N_18550,N_17143,N_17469);
and U18551 (N_18551,N_17292,N_17567);
or U18552 (N_18552,N_17898,N_17409);
or U18553 (N_18553,N_17084,N_17716);
nand U18554 (N_18554,N_17164,N_17442);
nor U18555 (N_18555,N_17083,N_17711);
nand U18556 (N_18556,N_17909,N_17163);
xnor U18557 (N_18557,N_17924,N_17867);
or U18558 (N_18558,N_17114,N_17591);
xor U18559 (N_18559,N_17443,N_17252);
nor U18560 (N_18560,N_17399,N_17362);
xnor U18561 (N_18561,N_17556,N_17001);
xor U18562 (N_18562,N_17666,N_17004);
nand U18563 (N_18563,N_17859,N_17118);
nand U18564 (N_18564,N_17371,N_17063);
nor U18565 (N_18565,N_17502,N_17192);
nor U18566 (N_18566,N_17429,N_17964);
nor U18567 (N_18567,N_17694,N_17541);
nand U18568 (N_18568,N_17580,N_17348);
nor U18569 (N_18569,N_17579,N_17595);
xor U18570 (N_18570,N_17305,N_17951);
nor U18571 (N_18571,N_17578,N_17983);
nand U18572 (N_18572,N_17847,N_17423);
or U18573 (N_18573,N_17684,N_17581);
nand U18574 (N_18574,N_17927,N_17844);
or U18575 (N_18575,N_17490,N_17429);
xnor U18576 (N_18576,N_17877,N_17767);
nor U18577 (N_18577,N_17465,N_17606);
xnor U18578 (N_18578,N_17338,N_17257);
nor U18579 (N_18579,N_17275,N_17624);
nor U18580 (N_18580,N_17539,N_17810);
nand U18581 (N_18581,N_17061,N_17059);
nand U18582 (N_18582,N_17732,N_17150);
xor U18583 (N_18583,N_17003,N_17051);
xnor U18584 (N_18584,N_17413,N_17540);
or U18585 (N_18585,N_17119,N_17133);
nand U18586 (N_18586,N_17173,N_17205);
nor U18587 (N_18587,N_17910,N_17612);
nor U18588 (N_18588,N_17751,N_17056);
and U18589 (N_18589,N_17410,N_17347);
nand U18590 (N_18590,N_17616,N_17678);
and U18591 (N_18591,N_17599,N_17603);
nand U18592 (N_18592,N_17646,N_17958);
nand U18593 (N_18593,N_17814,N_17892);
and U18594 (N_18594,N_17306,N_17479);
nor U18595 (N_18595,N_17691,N_17512);
and U18596 (N_18596,N_17698,N_17901);
nand U18597 (N_18597,N_17202,N_17899);
xnor U18598 (N_18598,N_17991,N_17404);
xor U18599 (N_18599,N_17221,N_17133);
or U18600 (N_18600,N_17055,N_17779);
nand U18601 (N_18601,N_17098,N_17521);
and U18602 (N_18602,N_17917,N_17042);
or U18603 (N_18603,N_17532,N_17456);
or U18604 (N_18604,N_17895,N_17936);
and U18605 (N_18605,N_17123,N_17789);
nand U18606 (N_18606,N_17903,N_17101);
and U18607 (N_18607,N_17314,N_17206);
xnor U18608 (N_18608,N_17386,N_17214);
nand U18609 (N_18609,N_17981,N_17929);
xor U18610 (N_18610,N_17702,N_17378);
or U18611 (N_18611,N_17233,N_17831);
and U18612 (N_18612,N_17601,N_17995);
nand U18613 (N_18613,N_17385,N_17949);
or U18614 (N_18614,N_17317,N_17329);
nand U18615 (N_18615,N_17196,N_17086);
xor U18616 (N_18616,N_17828,N_17087);
xnor U18617 (N_18617,N_17117,N_17581);
nor U18618 (N_18618,N_17622,N_17554);
and U18619 (N_18619,N_17053,N_17274);
and U18620 (N_18620,N_17860,N_17105);
nand U18621 (N_18621,N_17277,N_17279);
nand U18622 (N_18622,N_17690,N_17549);
nand U18623 (N_18623,N_17752,N_17009);
xnor U18624 (N_18624,N_17296,N_17785);
or U18625 (N_18625,N_17471,N_17551);
and U18626 (N_18626,N_17959,N_17775);
xor U18627 (N_18627,N_17634,N_17613);
and U18628 (N_18628,N_17189,N_17386);
nor U18629 (N_18629,N_17393,N_17264);
nor U18630 (N_18630,N_17723,N_17925);
nor U18631 (N_18631,N_17400,N_17716);
and U18632 (N_18632,N_17555,N_17598);
nand U18633 (N_18633,N_17347,N_17419);
and U18634 (N_18634,N_17652,N_17840);
and U18635 (N_18635,N_17432,N_17241);
nor U18636 (N_18636,N_17672,N_17310);
nor U18637 (N_18637,N_17811,N_17971);
nor U18638 (N_18638,N_17827,N_17683);
nand U18639 (N_18639,N_17662,N_17498);
xnor U18640 (N_18640,N_17020,N_17573);
and U18641 (N_18641,N_17361,N_17052);
xor U18642 (N_18642,N_17293,N_17963);
nand U18643 (N_18643,N_17630,N_17962);
and U18644 (N_18644,N_17826,N_17971);
nor U18645 (N_18645,N_17547,N_17822);
or U18646 (N_18646,N_17359,N_17891);
and U18647 (N_18647,N_17065,N_17934);
nor U18648 (N_18648,N_17160,N_17458);
xor U18649 (N_18649,N_17654,N_17250);
or U18650 (N_18650,N_17443,N_17487);
xor U18651 (N_18651,N_17474,N_17988);
nor U18652 (N_18652,N_17208,N_17513);
xor U18653 (N_18653,N_17253,N_17628);
or U18654 (N_18654,N_17644,N_17011);
xor U18655 (N_18655,N_17877,N_17385);
or U18656 (N_18656,N_17941,N_17450);
xnor U18657 (N_18657,N_17290,N_17935);
and U18658 (N_18658,N_17435,N_17970);
nor U18659 (N_18659,N_17242,N_17988);
nand U18660 (N_18660,N_17532,N_17047);
xnor U18661 (N_18661,N_17317,N_17745);
xnor U18662 (N_18662,N_17850,N_17096);
or U18663 (N_18663,N_17669,N_17947);
or U18664 (N_18664,N_17129,N_17455);
xor U18665 (N_18665,N_17091,N_17584);
or U18666 (N_18666,N_17974,N_17146);
nand U18667 (N_18667,N_17000,N_17598);
nor U18668 (N_18668,N_17324,N_17736);
or U18669 (N_18669,N_17363,N_17155);
or U18670 (N_18670,N_17233,N_17957);
or U18671 (N_18671,N_17640,N_17780);
and U18672 (N_18672,N_17514,N_17712);
or U18673 (N_18673,N_17263,N_17889);
or U18674 (N_18674,N_17769,N_17717);
xor U18675 (N_18675,N_17400,N_17917);
or U18676 (N_18676,N_17965,N_17666);
nor U18677 (N_18677,N_17453,N_17442);
and U18678 (N_18678,N_17379,N_17616);
xor U18679 (N_18679,N_17624,N_17144);
and U18680 (N_18680,N_17923,N_17917);
or U18681 (N_18681,N_17081,N_17665);
nor U18682 (N_18682,N_17561,N_17443);
and U18683 (N_18683,N_17457,N_17653);
and U18684 (N_18684,N_17560,N_17412);
nand U18685 (N_18685,N_17577,N_17695);
nor U18686 (N_18686,N_17298,N_17966);
and U18687 (N_18687,N_17885,N_17266);
nor U18688 (N_18688,N_17398,N_17583);
nand U18689 (N_18689,N_17850,N_17610);
nor U18690 (N_18690,N_17654,N_17070);
xor U18691 (N_18691,N_17323,N_17766);
xnor U18692 (N_18692,N_17910,N_17604);
and U18693 (N_18693,N_17792,N_17628);
and U18694 (N_18694,N_17060,N_17804);
nor U18695 (N_18695,N_17019,N_17083);
and U18696 (N_18696,N_17146,N_17409);
xnor U18697 (N_18697,N_17737,N_17866);
and U18698 (N_18698,N_17976,N_17249);
and U18699 (N_18699,N_17814,N_17186);
or U18700 (N_18700,N_17316,N_17932);
xor U18701 (N_18701,N_17864,N_17593);
xor U18702 (N_18702,N_17050,N_17132);
nor U18703 (N_18703,N_17415,N_17895);
and U18704 (N_18704,N_17785,N_17420);
or U18705 (N_18705,N_17844,N_17155);
nor U18706 (N_18706,N_17427,N_17705);
or U18707 (N_18707,N_17877,N_17860);
xnor U18708 (N_18708,N_17303,N_17202);
nand U18709 (N_18709,N_17416,N_17984);
xor U18710 (N_18710,N_17608,N_17024);
and U18711 (N_18711,N_17169,N_17803);
and U18712 (N_18712,N_17606,N_17353);
and U18713 (N_18713,N_17373,N_17226);
xor U18714 (N_18714,N_17578,N_17268);
nor U18715 (N_18715,N_17993,N_17552);
and U18716 (N_18716,N_17245,N_17037);
or U18717 (N_18717,N_17861,N_17343);
nand U18718 (N_18718,N_17400,N_17824);
xor U18719 (N_18719,N_17996,N_17442);
nand U18720 (N_18720,N_17694,N_17844);
nand U18721 (N_18721,N_17775,N_17735);
and U18722 (N_18722,N_17531,N_17779);
nand U18723 (N_18723,N_17969,N_17284);
nand U18724 (N_18724,N_17616,N_17046);
or U18725 (N_18725,N_17438,N_17407);
nor U18726 (N_18726,N_17796,N_17478);
or U18727 (N_18727,N_17775,N_17809);
and U18728 (N_18728,N_17994,N_17629);
xnor U18729 (N_18729,N_17988,N_17219);
xnor U18730 (N_18730,N_17571,N_17603);
and U18731 (N_18731,N_17065,N_17058);
or U18732 (N_18732,N_17728,N_17258);
or U18733 (N_18733,N_17047,N_17319);
nand U18734 (N_18734,N_17966,N_17635);
nand U18735 (N_18735,N_17834,N_17898);
nor U18736 (N_18736,N_17090,N_17357);
xor U18737 (N_18737,N_17918,N_17207);
xor U18738 (N_18738,N_17260,N_17836);
nand U18739 (N_18739,N_17896,N_17495);
or U18740 (N_18740,N_17141,N_17920);
nor U18741 (N_18741,N_17946,N_17132);
and U18742 (N_18742,N_17491,N_17090);
and U18743 (N_18743,N_17730,N_17327);
nor U18744 (N_18744,N_17649,N_17195);
and U18745 (N_18745,N_17832,N_17887);
nor U18746 (N_18746,N_17319,N_17119);
xnor U18747 (N_18747,N_17700,N_17019);
nor U18748 (N_18748,N_17058,N_17010);
nor U18749 (N_18749,N_17883,N_17125);
or U18750 (N_18750,N_17224,N_17647);
or U18751 (N_18751,N_17755,N_17226);
xnor U18752 (N_18752,N_17970,N_17437);
xor U18753 (N_18753,N_17646,N_17001);
xnor U18754 (N_18754,N_17801,N_17230);
and U18755 (N_18755,N_17104,N_17399);
xor U18756 (N_18756,N_17723,N_17198);
nand U18757 (N_18757,N_17914,N_17540);
nand U18758 (N_18758,N_17467,N_17291);
or U18759 (N_18759,N_17481,N_17742);
and U18760 (N_18760,N_17227,N_17043);
and U18761 (N_18761,N_17236,N_17157);
nor U18762 (N_18762,N_17938,N_17897);
or U18763 (N_18763,N_17707,N_17532);
nor U18764 (N_18764,N_17180,N_17366);
or U18765 (N_18765,N_17066,N_17396);
xor U18766 (N_18766,N_17643,N_17759);
nor U18767 (N_18767,N_17811,N_17965);
or U18768 (N_18768,N_17455,N_17166);
nand U18769 (N_18769,N_17446,N_17475);
nor U18770 (N_18770,N_17190,N_17702);
nand U18771 (N_18771,N_17626,N_17510);
xor U18772 (N_18772,N_17437,N_17032);
or U18773 (N_18773,N_17394,N_17309);
nand U18774 (N_18774,N_17548,N_17036);
and U18775 (N_18775,N_17057,N_17981);
xor U18776 (N_18776,N_17630,N_17407);
or U18777 (N_18777,N_17790,N_17893);
or U18778 (N_18778,N_17921,N_17641);
nand U18779 (N_18779,N_17768,N_17483);
nor U18780 (N_18780,N_17673,N_17452);
nor U18781 (N_18781,N_17325,N_17785);
nand U18782 (N_18782,N_17149,N_17371);
or U18783 (N_18783,N_17178,N_17477);
and U18784 (N_18784,N_17347,N_17082);
xor U18785 (N_18785,N_17603,N_17978);
xnor U18786 (N_18786,N_17387,N_17622);
xnor U18787 (N_18787,N_17129,N_17777);
and U18788 (N_18788,N_17851,N_17027);
xor U18789 (N_18789,N_17990,N_17636);
nand U18790 (N_18790,N_17781,N_17420);
nand U18791 (N_18791,N_17782,N_17668);
and U18792 (N_18792,N_17179,N_17754);
nand U18793 (N_18793,N_17841,N_17346);
or U18794 (N_18794,N_17221,N_17792);
nor U18795 (N_18795,N_17049,N_17897);
nand U18796 (N_18796,N_17329,N_17363);
nand U18797 (N_18797,N_17842,N_17256);
and U18798 (N_18798,N_17802,N_17226);
or U18799 (N_18799,N_17182,N_17208);
or U18800 (N_18800,N_17389,N_17912);
and U18801 (N_18801,N_17630,N_17242);
nor U18802 (N_18802,N_17134,N_17007);
or U18803 (N_18803,N_17076,N_17020);
nand U18804 (N_18804,N_17406,N_17983);
nand U18805 (N_18805,N_17864,N_17738);
or U18806 (N_18806,N_17415,N_17126);
nor U18807 (N_18807,N_17219,N_17797);
nand U18808 (N_18808,N_17112,N_17445);
xnor U18809 (N_18809,N_17567,N_17667);
nor U18810 (N_18810,N_17284,N_17837);
xnor U18811 (N_18811,N_17757,N_17068);
or U18812 (N_18812,N_17118,N_17628);
and U18813 (N_18813,N_17867,N_17088);
or U18814 (N_18814,N_17570,N_17129);
xor U18815 (N_18815,N_17699,N_17249);
xor U18816 (N_18816,N_17271,N_17001);
xnor U18817 (N_18817,N_17953,N_17322);
or U18818 (N_18818,N_17789,N_17219);
nor U18819 (N_18819,N_17862,N_17634);
xnor U18820 (N_18820,N_17490,N_17596);
nand U18821 (N_18821,N_17044,N_17482);
nor U18822 (N_18822,N_17477,N_17928);
and U18823 (N_18823,N_17582,N_17180);
nor U18824 (N_18824,N_17376,N_17453);
nand U18825 (N_18825,N_17560,N_17571);
nand U18826 (N_18826,N_17627,N_17948);
and U18827 (N_18827,N_17871,N_17370);
and U18828 (N_18828,N_17620,N_17387);
nor U18829 (N_18829,N_17624,N_17505);
nand U18830 (N_18830,N_17063,N_17813);
nand U18831 (N_18831,N_17996,N_17739);
xor U18832 (N_18832,N_17706,N_17769);
xor U18833 (N_18833,N_17898,N_17830);
and U18834 (N_18834,N_17992,N_17927);
nand U18835 (N_18835,N_17878,N_17495);
or U18836 (N_18836,N_17429,N_17335);
and U18837 (N_18837,N_17372,N_17330);
and U18838 (N_18838,N_17168,N_17349);
nand U18839 (N_18839,N_17672,N_17580);
or U18840 (N_18840,N_17753,N_17016);
or U18841 (N_18841,N_17462,N_17472);
nor U18842 (N_18842,N_17661,N_17778);
nand U18843 (N_18843,N_17444,N_17187);
nor U18844 (N_18844,N_17846,N_17465);
nor U18845 (N_18845,N_17966,N_17329);
nor U18846 (N_18846,N_17196,N_17307);
or U18847 (N_18847,N_17235,N_17067);
and U18848 (N_18848,N_17757,N_17486);
nand U18849 (N_18849,N_17473,N_17303);
or U18850 (N_18850,N_17013,N_17388);
nor U18851 (N_18851,N_17586,N_17965);
xnor U18852 (N_18852,N_17601,N_17749);
nor U18853 (N_18853,N_17786,N_17653);
xnor U18854 (N_18854,N_17646,N_17934);
xor U18855 (N_18855,N_17931,N_17402);
or U18856 (N_18856,N_17094,N_17655);
or U18857 (N_18857,N_17894,N_17846);
or U18858 (N_18858,N_17921,N_17883);
or U18859 (N_18859,N_17612,N_17477);
and U18860 (N_18860,N_17664,N_17376);
xnor U18861 (N_18861,N_17033,N_17072);
nand U18862 (N_18862,N_17809,N_17579);
and U18863 (N_18863,N_17049,N_17809);
xor U18864 (N_18864,N_17892,N_17210);
and U18865 (N_18865,N_17341,N_17717);
nor U18866 (N_18866,N_17004,N_17327);
and U18867 (N_18867,N_17485,N_17742);
nor U18868 (N_18868,N_17416,N_17993);
nand U18869 (N_18869,N_17828,N_17630);
nand U18870 (N_18870,N_17698,N_17541);
xnor U18871 (N_18871,N_17541,N_17451);
xor U18872 (N_18872,N_17693,N_17240);
xnor U18873 (N_18873,N_17249,N_17708);
nor U18874 (N_18874,N_17621,N_17782);
xnor U18875 (N_18875,N_17604,N_17801);
xor U18876 (N_18876,N_17294,N_17840);
nand U18877 (N_18877,N_17687,N_17164);
and U18878 (N_18878,N_17750,N_17253);
and U18879 (N_18879,N_17836,N_17955);
or U18880 (N_18880,N_17561,N_17981);
or U18881 (N_18881,N_17368,N_17683);
or U18882 (N_18882,N_17575,N_17352);
nand U18883 (N_18883,N_17269,N_17394);
and U18884 (N_18884,N_17372,N_17146);
nor U18885 (N_18885,N_17513,N_17305);
nand U18886 (N_18886,N_17899,N_17550);
or U18887 (N_18887,N_17732,N_17179);
or U18888 (N_18888,N_17847,N_17805);
or U18889 (N_18889,N_17260,N_17434);
xnor U18890 (N_18890,N_17505,N_17911);
or U18891 (N_18891,N_17854,N_17848);
and U18892 (N_18892,N_17931,N_17898);
and U18893 (N_18893,N_17492,N_17487);
and U18894 (N_18894,N_17431,N_17429);
or U18895 (N_18895,N_17818,N_17997);
nor U18896 (N_18896,N_17496,N_17677);
nor U18897 (N_18897,N_17570,N_17178);
or U18898 (N_18898,N_17503,N_17583);
and U18899 (N_18899,N_17940,N_17809);
nand U18900 (N_18900,N_17123,N_17809);
and U18901 (N_18901,N_17190,N_17895);
nor U18902 (N_18902,N_17645,N_17041);
xor U18903 (N_18903,N_17186,N_17219);
xnor U18904 (N_18904,N_17295,N_17855);
nor U18905 (N_18905,N_17157,N_17507);
or U18906 (N_18906,N_17688,N_17959);
nand U18907 (N_18907,N_17700,N_17434);
nand U18908 (N_18908,N_17244,N_17528);
or U18909 (N_18909,N_17762,N_17207);
nor U18910 (N_18910,N_17194,N_17413);
or U18911 (N_18911,N_17522,N_17195);
and U18912 (N_18912,N_17918,N_17908);
nand U18913 (N_18913,N_17402,N_17194);
nor U18914 (N_18914,N_17234,N_17073);
xor U18915 (N_18915,N_17244,N_17933);
or U18916 (N_18916,N_17639,N_17273);
nand U18917 (N_18917,N_17450,N_17052);
nand U18918 (N_18918,N_17740,N_17815);
nand U18919 (N_18919,N_17924,N_17641);
and U18920 (N_18920,N_17285,N_17514);
nand U18921 (N_18921,N_17562,N_17823);
or U18922 (N_18922,N_17596,N_17532);
xor U18923 (N_18923,N_17805,N_17446);
or U18924 (N_18924,N_17712,N_17351);
nand U18925 (N_18925,N_17118,N_17485);
or U18926 (N_18926,N_17309,N_17005);
nand U18927 (N_18927,N_17975,N_17868);
nor U18928 (N_18928,N_17897,N_17334);
and U18929 (N_18929,N_17160,N_17757);
nor U18930 (N_18930,N_17274,N_17903);
and U18931 (N_18931,N_17632,N_17492);
nand U18932 (N_18932,N_17826,N_17571);
nand U18933 (N_18933,N_17718,N_17152);
xnor U18934 (N_18934,N_17403,N_17299);
or U18935 (N_18935,N_17603,N_17644);
nor U18936 (N_18936,N_17858,N_17154);
or U18937 (N_18937,N_17007,N_17947);
nand U18938 (N_18938,N_17980,N_17349);
nand U18939 (N_18939,N_17766,N_17673);
or U18940 (N_18940,N_17054,N_17275);
nor U18941 (N_18941,N_17023,N_17327);
or U18942 (N_18942,N_17912,N_17460);
or U18943 (N_18943,N_17594,N_17415);
nor U18944 (N_18944,N_17157,N_17464);
and U18945 (N_18945,N_17019,N_17236);
xor U18946 (N_18946,N_17411,N_17664);
nand U18947 (N_18947,N_17888,N_17270);
and U18948 (N_18948,N_17715,N_17056);
or U18949 (N_18949,N_17357,N_17420);
or U18950 (N_18950,N_17455,N_17291);
nor U18951 (N_18951,N_17922,N_17657);
nor U18952 (N_18952,N_17642,N_17200);
nand U18953 (N_18953,N_17219,N_17248);
nand U18954 (N_18954,N_17214,N_17082);
or U18955 (N_18955,N_17063,N_17735);
and U18956 (N_18956,N_17572,N_17114);
and U18957 (N_18957,N_17803,N_17178);
xnor U18958 (N_18958,N_17142,N_17326);
or U18959 (N_18959,N_17562,N_17148);
nor U18960 (N_18960,N_17821,N_17026);
or U18961 (N_18961,N_17779,N_17925);
nor U18962 (N_18962,N_17548,N_17613);
xnor U18963 (N_18963,N_17917,N_17382);
nor U18964 (N_18964,N_17788,N_17851);
and U18965 (N_18965,N_17770,N_17613);
nor U18966 (N_18966,N_17753,N_17950);
nand U18967 (N_18967,N_17113,N_17306);
nand U18968 (N_18968,N_17497,N_17199);
or U18969 (N_18969,N_17105,N_17086);
nor U18970 (N_18970,N_17917,N_17432);
and U18971 (N_18971,N_17346,N_17273);
nor U18972 (N_18972,N_17489,N_17989);
nor U18973 (N_18973,N_17408,N_17506);
and U18974 (N_18974,N_17842,N_17171);
or U18975 (N_18975,N_17609,N_17887);
or U18976 (N_18976,N_17644,N_17107);
xor U18977 (N_18977,N_17688,N_17790);
nand U18978 (N_18978,N_17811,N_17891);
nand U18979 (N_18979,N_17842,N_17362);
and U18980 (N_18980,N_17153,N_17173);
xor U18981 (N_18981,N_17547,N_17656);
xor U18982 (N_18982,N_17437,N_17270);
or U18983 (N_18983,N_17019,N_17696);
or U18984 (N_18984,N_17546,N_17271);
nor U18985 (N_18985,N_17325,N_17546);
nor U18986 (N_18986,N_17747,N_17410);
nand U18987 (N_18987,N_17888,N_17853);
nand U18988 (N_18988,N_17323,N_17996);
nand U18989 (N_18989,N_17617,N_17374);
nand U18990 (N_18990,N_17397,N_17654);
nand U18991 (N_18991,N_17336,N_17831);
nand U18992 (N_18992,N_17542,N_17665);
or U18993 (N_18993,N_17338,N_17708);
and U18994 (N_18994,N_17697,N_17000);
or U18995 (N_18995,N_17274,N_17560);
nand U18996 (N_18996,N_17263,N_17386);
xnor U18997 (N_18997,N_17256,N_17765);
nor U18998 (N_18998,N_17051,N_17387);
and U18999 (N_18999,N_17063,N_17539);
nand U19000 (N_19000,N_18553,N_18410);
and U19001 (N_19001,N_18531,N_18470);
xnor U19002 (N_19002,N_18827,N_18172);
nand U19003 (N_19003,N_18722,N_18919);
or U19004 (N_19004,N_18670,N_18492);
nor U19005 (N_19005,N_18023,N_18207);
nand U19006 (N_19006,N_18366,N_18467);
nand U19007 (N_19007,N_18689,N_18121);
xnor U19008 (N_19008,N_18376,N_18144);
and U19009 (N_19009,N_18063,N_18259);
nor U19010 (N_19010,N_18558,N_18715);
xnor U19011 (N_19011,N_18234,N_18385);
or U19012 (N_19012,N_18167,N_18658);
nand U19013 (N_19013,N_18671,N_18639);
nor U19014 (N_19014,N_18749,N_18915);
nand U19015 (N_19015,N_18101,N_18058);
or U19016 (N_19016,N_18816,N_18344);
nand U19017 (N_19017,N_18662,N_18434);
or U19018 (N_19018,N_18171,N_18659);
or U19019 (N_19019,N_18198,N_18609);
and U19020 (N_19020,N_18189,N_18582);
nand U19021 (N_19021,N_18059,N_18599);
nand U19022 (N_19022,N_18980,N_18907);
nand U19023 (N_19023,N_18991,N_18603);
nand U19024 (N_19024,N_18035,N_18415);
xnor U19025 (N_19025,N_18301,N_18889);
xnor U19026 (N_19026,N_18850,N_18329);
nand U19027 (N_19027,N_18038,N_18868);
and U19028 (N_19028,N_18217,N_18967);
xor U19029 (N_19029,N_18946,N_18491);
or U19030 (N_19030,N_18740,N_18400);
nand U19031 (N_19031,N_18709,N_18387);
nand U19032 (N_19032,N_18534,N_18176);
nor U19033 (N_19033,N_18962,N_18828);
xnor U19034 (N_19034,N_18285,N_18799);
and U19035 (N_19035,N_18651,N_18287);
nand U19036 (N_19036,N_18205,N_18897);
and U19037 (N_19037,N_18909,N_18421);
nand U19038 (N_19038,N_18583,N_18815);
and U19039 (N_19039,N_18142,N_18641);
nand U19040 (N_19040,N_18638,N_18890);
nand U19041 (N_19041,N_18832,N_18835);
xnor U19042 (N_19042,N_18841,N_18258);
or U19043 (N_19043,N_18923,N_18982);
nand U19044 (N_19044,N_18625,N_18314);
and U19045 (N_19045,N_18149,N_18621);
nor U19046 (N_19046,N_18587,N_18634);
nand U19047 (N_19047,N_18054,N_18053);
or U19048 (N_19048,N_18728,N_18163);
xnor U19049 (N_19049,N_18644,N_18336);
nor U19050 (N_19050,N_18877,N_18466);
nand U19051 (N_19051,N_18147,N_18377);
or U19052 (N_19052,N_18955,N_18575);
and U19053 (N_19053,N_18392,N_18484);
nor U19054 (N_19054,N_18527,N_18576);
or U19055 (N_19055,N_18795,N_18848);
xor U19056 (N_19056,N_18508,N_18204);
or U19057 (N_19057,N_18711,N_18006);
nand U19058 (N_19058,N_18928,N_18373);
nand U19059 (N_19059,N_18419,N_18283);
nor U19060 (N_19060,N_18705,N_18566);
nand U19061 (N_19061,N_18241,N_18218);
nand U19062 (N_19062,N_18028,N_18153);
nor U19063 (N_19063,N_18905,N_18326);
nor U19064 (N_19064,N_18118,N_18924);
nor U19065 (N_19065,N_18290,N_18618);
and U19066 (N_19066,N_18046,N_18507);
nor U19067 (N_19067,N_18297,N_18268);
nor U19068 (N_19068,N_18655,N_18519);
nand U19069 (N_19069,N_18833,N_18528);
nand U19070 (N_19070,N_18560,N_18341);
xor U19071 (N_19071,N_18102,N_18254);
nor U19072 (N_19072,N_18381,N_18648);
and U19073 (N_19073,N_18800,N_18733);
or U19074 (N_19074,N_18807,N_18572);
or U19075 (N_19075,N_18245,N_18224);
nor U19076 (N_19076,N_18347,N_18904);
and U19077 (N_19077,N_18994,N_18664);
xor U19078 (N_19078,N_18156,N_18953);
and U19079 (N_19079,N_18562,N_18013);
xnor U19080 (N_19080,N_18629,N_18674);
xnor U19081 (N_19081,N_18386,N_18422);
nand U19082 (N_19082,N_18371,N_18251);
nand U19083 (N_19083,N_18200,N_18650);
xor U19084 (N_19084,N_18922,N_18324);
xor U19085 (N_19085,N_18214,N_18108);
nand U19086 (N_19086,N_18201,N_18631);
and U19087 (N_19087,N_18256,N_18615);
or U19088 (N_19088,N_18601,N_18524);
xnor U19089 (N_19089,N_18313,N_18762);
xnor U19090 (N_19090,N_18143,N_18380);
or U19091 (N_19091,N_18180,N_18864);
nand U19092 (N_19092,N_18315,N_18413);
nor U19093 (N_19093,N_18279,N_18170);
nor U19094 (N_19094,N_18623,N_18015);
nand U19095 (N_19095,N_18744,N_18420);
or U19096 (N_19096,N_18875,N_18520);
or U19097 (N_19097,N_18497,N_18260);
and U19098 (N_19098,N_18117,N_18593);
nor U19099 (N_19099,N_18209,N_18049);
nor U19100 (N_19100,N_18363,N_18032);
xor U19101 (N_19101,N_18022,N_18624);
or U19102 (N_19102,N_18019,N_18505);
nor U19103 (N_19103,N_18783,N_18756);
and U19104 (N_19104,N_18383,N_18225);
nand U19105 (N_19105,N_18050,N_18277);
xnor U19106 (N_19106,N_18565,N_18970);
nand U19107 (N_19107,N_18514,N_18140);
or U19108 (N_19108,N_18839,N_18359);
xnor U19109 (N_19109,N_18809,N_18012);
xor U19110 (N_19110,N_18773,N_18455);
and U19111 (N_19111,N_18448,N_18779);
xor U19112 (N_19112,N_18228,N_18107);
nand U19113 (N_19113,N_18643,N_18401);
and U19114 (N_19114,N_18169,N_18369);
nand U19115 (N_19115,N_18766,N_18957);
and U19116 (N_19116,N_18340,N_18210);
or U19117 (N_19117,N_18939,N_18826);
or U19118 (N_19118,N_18811,N_18498);
or U19119 (N_19119,N_18495,N_18921);
nand U19120 (N_19120,N_18737,N_18517);
nand U19121 (N_19121,N_18777,N_18960);
nand U19122 (N_19122,N_18403,N_18468);
xnor U19123 (N_19123,N_18358,N_18139);
and U19124 (N_19124,N_18231,N_18262);
and U19125 (N_19125,N_18999,N_18034);
nor U19126 (N_19126,N_18918,N_18304);
or U19127 (N_19127,N_18067,N_18077);
and U19128 (N_19128,N_18001,N_18317);
and U19129 (N_19129,N_18652,N_18769);
or U19130 (N_19130,N_18956,N_18852);
and U19131 (N_19131,N_18567,N_18441);
and U19132 (N_19132,N_18122,N_18454);
and U19133 (N_19133,N_18099,N_18129);
xnor U19134 (N_19134,N_18197,N_18296);
and U19135 (N_19135,N_18612,N_18637);
nor U19136 (N_19136,N_18405,N_18246);
or U19137 (N_19137,N_18742,N_18299);
nand U19138 (N_19138,N_18354,N_18069);
or U19139 (N_19139,N_18713,N_18798);
or U19140 (N_19140,N_18808,N_18981);
nor U19141 (N_19141,N_18282,N_18834);
or U19142 (N_19142,N_18327,N_18851);
and U19143 (N_19143,N_18926,N_18735);
nor U19144 (N_19144,N_18330,N_18307);
xor U19145 (N_19145,N_18060,N_18025);
and U19146 (N_19146,N_18474,N_18398);
nor U19147 (N_19147,N_18791,N_18866);
and U19148 (N_19148,N_18916,N_18555);
and U19149 (N_19149,N_18554,N_18719);
xor U19150 (N_19150,N_18708,N_18684);
nor U19151 (N_19151,N_18765,N_18220);
nor U19152 (N_19152,N_18760,N_18596);
nor U19153 (N_19153,N_18408,N_18630);
nor U19154 (N_19154,N_18985,N_18842);
xor U19155 (N_19155,N_18346,N_18362);
or U19156 (N_19156,N_18082,N_18993);
xnor U19157 (N_19157,N_18654,N_18334);
or U19158 (N_19158,N_18098,N_18349);
and U19159 (N_19159,N_18511,N_18230);
or U19160 (N_19160,N_18306,N_18192);
nor U19161 (N_19161,N_18640,N_18071);
or U19162 (N_19162,N_18887,N_18772);
nor U19163 (N_19163,N_18364,N_18821);
xnor U19164 (N_19164,N_18064,N_18087);
nand U19165 (N_19165,N_18343,N_18845);
xnor U19166 (N_19166,N_18292,N_18097);
and U19167 (N_19167,N_18316,N_18780);
and U19168 (N_19168,N_18091,N_18607);
and U19169 (N_19169,N_18273,N_18042);
nand U19170 (N_19170,N_18095,N_18490);
and U19171 (N_19171,N_18571,N_18754);
and U19172 (N_19172,N_18423,N_18679);
nand U19173 (N_19173,N_18242,N_18523);
xor U19174 (N_19174,N_18130,N_18206);
nor U19175 (N_19175,N_18110,N_18280);
and U19176 (N_19176,N_18062,N_18456);
or U19177 (N_19177,N_18017,N_18240);
nand U19178 (N_19178,N_18266,N_18646);
nor U19179 (N_19179,N_18885,N_18504);
xor U19180 (N_19180,N_18177,N_18243);
nand U19181 (N_19181,N_18076,N_18849);
and U19182 (N_19182,N_18115,N_18547);
nor U19183 (N_19183,N_18509,N_18159);
nand U19184 (N_19184,N_18004,N_18407);
xor U19185 (N_19185,N_18861,N_18016);
nor U19186 (N_19186,N_18721,N_18611);
nor U19187 (N_19187,N_18181,N_18103);
and U19188 (N_19188,N_18033,N_18114);
nand U19189 (N_19189,N_18537,N_18899);
xor U19190 (N_19190,N_18429,N_18965);
nand U19191 (N_19191,N_18574,N_18440);
nor U19192 (N_19192,N_18310,N_18753);
xor U19193 (N_19193,N_18320,N_18188);
nor U19194 (N_19194,N_18901,N_18356);
or U19195 (N_19195,N_18426,N_18461);
nor U19196 (N_19196,N_18856,N_18548);
nand U19197 (N_19197,N_18862,N_18948);
or U19198 (N_19198,N_18613,N_18913);
and U19199 (N_19199,N_18578,N_18424);
or U19200 (N_19200,N_18409,N_18880);
nor U19201 (N_19201,N_18269,N_18941);
nor U19202 (N_19202,N_18820,N_18223);
nand U19203 (N_19203,N_18487,N_18831);
xor U19204 (N_19204,N_18529,N_18335);
nor U19205 (N_19205,N_18394,N_18871);
and U19206 (N_19206,N_18009,N_18372);
nor U19207 (N_19207,N_18930,N_18714);
nor U19208 (N_19208,N_18227,N_18074);
and U19209 (N_19209,N_18645,N_18594);
nand U19210 (N_19210,N_18723,N_18622);
or U19211 (N_19211,N_18318,N_18168);
xnor U19212 (N_19212,N_18044,N_18175);
and U19213 (N_19213,N_18183,N_18971);
and U19214 (N_19214,N_18378,N_18616);
or U19215 (N_19215,N_18263,N_18453);
nor U19216 (N_19216,N_18473,N_18226);
xnor U19217 (N_19217,N_18472,N_18801);
xnor U19218 (N_19218,N_18295,N_18996);
xnor U19219 (N_19219,N_18480,N_18912);
xor U19220 (N_19220,N_18432,N_18278);
or U19221 (N_19221,N_18478,N_18949);
or U19222 (N_19222,N_18312,N_18061);
nand U19223 (N_19223,N_18402,N_18886);
nor U19224 (N_19224,N_18112,N_18134);
and U19225 (N_19225,N_18669,N_18399);
nand U19226 (N_19226,N_18741,N_18846);
nand U19227 (N_19227,N_18556,N_18244);
or U19228 (N_19228,N_18893,N_18272);
xnor U19229 (N_19229,N_18152,N_18286);
or U19230 (N_19230,N_18443,N_18293);
nor U19231 (N_19231,N_18573,N_18840);
or U19232 (N_19232,N_18406,N_18736);
or U19233 (N_19233,N_18759,N_18825);
xnor U19234 (N_19234,N_18768,N_18917);
nand U19235 (N_19235,N_18961,N_18717);
and U19236 (N_19236,N_18521,N_18788);
and U19237 (N_19237,N_18822,N_18512);
nor U19238 (N_19238,N_18173,N_18663);
and U19239 (N_19239,N_18450,N_18345);
nor U19240 (N_19240,N_18361,N_18396);
nand U19241 (N_19241,N_18716,N_18983);
xor U19242 (N_19242,N_18681,N_18271);
xor U19243 (N_19243,N_18703,N_18465);
nor U19244 (N_19244,N_18043,N_18235);
or U19245 (N_19245,N_18133,N_18039);
nand U19246 (N_19246,N_18353,N_18388);
nor U19247 (N_19247,N_18692,N_18563);
or U19248 (N_19248,N_18416,N_18927);
xor U19249 (N_19249,N_18530,N_18804);
or U19250 (N_19250,N_18427,N_18270);
nor U19251 (N_19251,N_18264,N_18365);
and U19252 (N_19252,N_18789,N_18552);
xnor U19253 (N_19253,N_18124,N_18430);
nand U19254 (N_19254,N_18193,N_18963);
xnor U19255 (N_19255,N_18221,N_18029);
or U19256 (N_19256,N_18449,N_18704);
nand U19257 (N_19257,N_18105,N_18414);
xnor U19258 (N_19258,N_18649,N_18642);
or U19259 (N_19259,N_18933,N_18489);
nor U19260 (N_19260,N_18729,N_18357);
xnor U19261 (N_19261,N_18151,N_18431);
and U19262 (N_19262,N_18544,N_18675);
nor U19263 (N_19263,N_18802,N_18984);
or U19264 (N_19264,N_18632,N_18844);
and U19265 (N_19265,N_18874,N_18628);
xor U19266 (N_19266,N_18477,N_18191);
and U19267 (N_19267,N_18745,N_18819);
nor U19268 (N_19268,N_18732,N_18428);
nor U19269 (N_19269,N_18796,N_18202);
xnor U19270 (N_19270,N_18458,N_18954);
or U19271 (N_19271,N_18265,N_18792);
nor U19272 (N_19272,N_18724,N_18350);
nand U19273 (N_19273,N_18008,N_18602);
xnor U19274 (N_19274,N_18352,N_18031);
nor U19275 (N_19275,N_18561,N_18898);
nor U19276 (N_19276,N_18382,N_18138);
nand U19277 (N_19277,N_18738,N_18481);
xnor U19278 (N_19278,N_18667,N_18284);
or U19279 (N_19279,N_18355,N_18950);
or U19280 (N_19280,N_18123,N_18486);
nand U19281 (N_19281,N_18813,N_18485);
nor U19282 (N_19282,N_18065,N_18469);
or U19283 (N_19283,N_18761,N_18219);
or U19284 (N_19284,N_18476,N_18447);
nand U19285 (N_19285,N_18784,N_18750);
xor U19286 (N_19286,N_18688,N_18814);
nand U19287 (N_19287,N_18992,N_18920);
and U19288 (N_19288,N_18236,N_18974);
or U19289 (N_19289,N_18113,N_18146);
nor U19290 (N_19290,N_18579,N_18445);
nor U19291 (N_19291,N_18883,N_18942);
or U19292 (N_19292,N_18678,N_18627);
nand U19293 (N_19293,N_18620,N_18309);
xor U19294 (N_19294,N_18444,N_18906);
nand U19295 (N_19295,N_18559,N_18374);
nand U19296 (N_19296,N_18178,N_18018);
nor U19297 (N_19297,N_18185,N_18947);
nor U19298 (N_19298,N_18683,N_18702);
nor U19299 (N_19299,N_18212,N_18094);
or U19300 (N_19300,N_18536,N_18002);
nor U19301 (N_19301,N_18075,N_18569);
nor U19302 (N_19302,N_18057,N_18047);
nor U19303 (N_19303,N_18752,N_18125);
nor U19304 (N_19304,N_18328,N_18155);
nor U19305 (N_19305,N_18148,N_18005);
xnor U19306 (N_19306,N_18267,N_18194);
or U19307 (N_19307,N_18793,N_18546);
nand U19308 (N_19308,N_18882,N_18586);
xor U19309 (N_19309,N_18437,N_18545);
xnor U19310 (N_19310,N_18966,N_18687);
nor U19311 (N_19311,N_18010,N_18515);
nor U19312 (N_19312,N_18164,N_18847);
nor U19313 (N_19313,N_18810,N_18119);
and U19314 (N_19314,N_18084,N_18302);
xnor U19315 (N_19315,N_18782,N_18690);
xor U19316 (N_19316,N_18348,N_18676);
nand U19317 (N_19317,N_18248,N_18542);
and U19318 (N_19318,N_18462,N_18109);
nand U19319 (N_19319,N_18647,N_18510);
nor U19320 (N_19320,N_18900,N_18250);
nand U19321 (N_19321,N_18686,N_18958);
xnor U19322 (N_19322,N_18770,N_18935);
nor U19323 (N_19323,N_18786,N_18911);
and U19324 (N_19324,N_18199,N_18925);
or U19325 (N_19325,N_18308,N_18239);
or U19326 (N_19326,N_18584,N_18021);
nand U19327 (N_19327,N_18817,N_18591);
and U19328 (N_19328,N_18275,N_18829);
nor U19329 (N_19329,N_18493,N_18577);
xor U19330 (N_19330,N_18617,N_18072);
nand U19331 (N_19331,N_18812,N_18331);
or U19332 (N_19332,N_18636,N_18179);
nor U19333 (N_19333,N_18066,N_18778);
nand U19334 (N_19334,N_18860,N_18425);
nand U19335 (N_19335,N_18037,N_18055);
xor U19336 (N_19336,N_18951,N_18739);
xnor U19337 (N_19337,N_18274,N_18865);
nor U19338 (N_19338,N_18261,N_18150);
xor U19339 (N_19339,N_18891,N_18499);
xnor U19340 (N_19340,N_18333,N_18090);
nor U19341 (N_19341,N_18763,N_18294);
nand U19342 (N_19342,N_18525,N_18694);
nand U19343 (N_19343,N_18116,N_18978);
xor U19344 (N_19344,N_18325,N_18203);
and U19345 (N_19345,N_18903,N_18764);
and U19346 (N_19346,N_18024,N_18370);
nand U19347 (N_19347,N_18995,N_18502);
nand U19348 (N_19348,N_18154,N_18937);
xor U19349 (N_19349,N_18549,N_18797);
nor U19350 (N_19350,N_18668,N_18869);
and U19351 (N_19351,N_18597,N_18237);
nor U19352 (N_19352,N_18040,N_18700);
or U19353 (N_19353,N_18391,N_18619);
nand U19354 (N_19354,N_18712,N_18830);
and U19355 (N_19355,N_18106,N_18775);
or U19356 (N_19356,N_18186,N_18696);
nor U19357 (N_19357,N_18080,N_18589);
nor U19358 (N_19358,N_18252,N_18337);
xnor U19359 (N_19359,N_18677,N_18007);
or U19360 (N_19360,N_18691,N_18442);
nor U19361 (N_19361,N_18436,N_18936);
xnor U19362 (N_19362,N_18969,N_18513);
nor U19363 (N_19363,N_18052,N_18902);
nand U19364 (N_19364,N_18706,N_18141);
nor U19365 (N_19365,N_18934,N_18837);
xnor U19366 (N_19366,N_18757,N_18539);
or U19367 (N_19367,N_18661,N_18516);
xnor U19368 (N_19368,N_18247,N_18710);
xnor U19369 (N_19369,N_18070,N_18073);
or U19370 (N_19370,N_18463,N_18853);
nand U19371 (N_19371,N_18404,N_18501);
xnor U19372 (N_19372,N_18608,N_18718);
xnor U19373 (N_19373,N_18867,N_18276);
nor U19374 (N_19374,N_18990,N_18459);
and U19375 (N_19375,N_18541,N_18311);
nor U19376 (N_19376,N_18944,N_18518);
or U19377 (N_19377,N_18666,N_18976);
or U19378 (N_19378,N_18879,N_18592);
xnor U19379 (N_19379,N_18111,N_18446);
nor U19380 (N_19380,N_18471,N_18503);
or U19381 (N_19381,N_18083,N_18673);
xor U19382 (N_19382,N_18393,N_18943);
nand U19383 (N_19383,N_18532,N_18166);
and U19384 (N_19384,N_18838,N_18368);
nor U19385 (N_19385,N_18137,N_18892);
and U19386 (N_19386,N_18973,N_18748);
nor U19387 (N_19387,N_18526,N_18595);
xor U19388 (N_19388,N_18606,N_18635);
and U19389 (N_19389,N_18794,N_18127);
nand U19390 (N_19390,N_18417,N_18945);
xor U19391 (N_19391,N_18190,N_18418);
nor U19392 (N_19392,N_18633,N_18390);
and U19393 (N_19393,N_18751,N_18338);
nand U19394 (N_19394,N_18580,N_18216);
and U19395 (N_19395,N_18896,N_18100);
xor U19396 (N_19396,N_18698,N_18438);
and U19397 (N_19397,N_18535,N_18972);
nand U19398 (N_19398,N_18249,N_18196);
xor U19399 (N_19399,N_18026,N_18457);
xor U19400 (N_19400,N_18027,N_18379);
xor U19401 (N_19401,N_18452,N_18680);
or U19402 (N_19402,N_18790,N_18747);
or U19403 (N_19403,N_18165,N_18836);
nor U19404 (N_19404,N_18894,N_18540);
and U19405 (N_19405,N_18672,N_18051);
xor U19406 (N_19406,N_18588,N_18858);
or U19407 (N_19407,N_18045,N_18538);
and U19408 (N_19408,N_18030,N_18884);
xnor U19409 (N_19409,N_18360,N_18494);
nand U19410 (N_19410,N_18433,N_18411);
nand U19411 (N_19411,N_18078,N_18451);
xor U19412 (N_19412,N_18222,N_18182);
nor U19413 (N_19413,N_18755,N_18255);
xor U19414 (N_19414,N_18758,N_18598);
and U19415 (N_19415,N_18288,N_18701);
xor U19416 (N_19416,N_18987,N_18727);
nor U19417 (N_19417,N_18910,N_18162);
nor U19418 (N_19418,N_18351,N_18774);
xor U19419 (N_19419,N_18693,N_18726);
nor U19420 (N_19420,N_18781,N_18843);
or U19421 (N_19421,N_18367,N_18435);
xor U19422 (N_19422,N_18305,N_18776);
nor U19423 (N_19423,N_18384,N_18551);
nor U19424 (N_19424,N_18048,N_18460);
xor U19425 (N_19425,N_18041,N_18656);
or U19426 (N_19426,N_18986,N_18895);
nand U19427 (N_19427,N_18291,N_18931);
and U19428 (N_19428,N_18093,N_18975);
or U19429 (N_19429,N_18730,N_18158);
nand U19430 (N_19430,N_18605,N_18522);
or U19431 (N_19431,N_18854,N_18298);
or U19432 (N_19432,N_18233,N_18475);
xor U19433 (N_19433,N_18585,N_18707);
xnor U19434 (N_19434,N_18823,N_18136);
and U19435 (N_19435,N_18321,N_18743);
or U19436 (N_19436,N_18626,N_18003);
xor U19437 (N_19437,N_18581,N_18322);
xnor U19438 (N_19438,N_18998,N_18940);
nand U19439 (N_19439,N_18653,N_18731);
or U19440 (N_19440,N_18479,N_18303);
xnor U19441 (N_19441,N_18787,N_18085);
xor U19442 (N_19442,N_18697,N_18104);
nand U19443 (N_19443,N_18397,N_18281);
nand U19444 (N_19444,N_18908,N_18988);
xor U19445 (N_19445,N_18564,N_18253);
and U19446 (N_19446,N_18208,N_18855);
and U19447 (N_19447,N_18873,N_18187);
and U19448 (N_19448,N_18570,N_18682);
xor U19449 (N_19449,N_18859,N_18720);
nor U19450 (N_19450,N_18543,N_18699);
and U19451 (N_19451,N_18665,N_18300);
or U19452 (N_19452,N_18211,N_18323);
nor U19453 (N_19453,N_18257,N_18959);
nor U19454 (N_19454,N_18590,N_18160);
nand U19455 (N_19455,N_18550,N_18332);
and U19456 (N_19456,N_18932,N_18857);
nand U19457 (N_19457,N_18213,N_18036);
xor U19458 (N_19458,N_18870,N_18568);
and U19459 (N_19459,N_18600,N_18238);
xnor U19460 (N_19460,N_18824,N_18120);
nor U19461 (N_19461,N_18506,N_18929);
xnor U19462 (N_19462,N_18079,N_18614);
xnor U19463 (N_19463,N_18339,N_18135);
nand U19464 (N_19464,N_18734,N_18092);
and U19465 (N_19465,N_18088,N_18000);
and U19466 (N_19466,N_18086,N_18145);
nor U19467 (N_19467,N_18157,N_18968);
and U19468 (N_19468,N_18412,N_18232);
nor U19469 (N_19469,N_18806,N_18174);
and U19470 (N_19470,N_18771,N_18089);
and U19471 (N_19471,N_18488,N_18014);
or U19472 (N_19472,N_18805,N_18500);
and U19473 (N_19473,N_18767,N_18319);
nand U19474 (N_19474,N_18184,N_18660);
or U19475 (N_19475,N_18725,N_18126);
or U19476 (N_19476,N_18375,N_18482);
and U19477 (N_19477,N_18964,N_18557);
nor U19478 (N_19478,N_18161,N_18464);
xnor U19479 (N_19479,N_18439,N_18289);
nor U19480 (N_19480,N_18068,N_18389);
nor U19481 (N_19481,N_18610,N_18888);
or U19482 (N_19482,N_18483,N_18128);
xnor U19483 (N_19483,N_18803,N_18785);
nand U19484 (N_19484,N_18395,N_18979);
xor U19485 (N_19485,N_18881,N_18011);
or U19486 (N_19486,N_18878,N_18872);
and U19487 (N_19487,N_18342,N_18056);
nor U19488 (N_19488,N_18496,N_18695);
or U19489 (N_19489,N_18215,N_18818);
or U19490 (N_19490,N_18914,N_18604);
nand U19491 (N_19491,N_18132,N_18685);
and U19492 (N_19492,N_18533,N_18989);
nor U19493 (N_19493,N_18081,N_18952);
or U19494 (N_19494,N_18876,N_18131);
nor U19495 (N_19495,N_18020,N_18977);
nand U19496 (N_19496,N_18195,N_18657);
xor U19497 (N_19497,N_18863,N_18938);
and U19498 (N_19498,N_18096,N_18229);
or U19499 (N_19499,N_18997,N_18746);
xnor U19500 (N_19500,N_18951,N_18877);
or U19501 (N_19501,N_18501,N_18064);
and U19502 (N_19502,N_18982,N_18867);
nand U19503 (N_19503,N_18289,N_18994);
or U19504 (N_19504,N_18431,N_18073);
xor U19505 (N_19505,N_18379,N_18131);
and U19506 (N_19506,N_18205,N_18715);
or U19507 (N_19507,N_18400,N_18714);
xor U19508 (N_19508,N_18167,N_18244);
nor U19509 (N_19509,N_18857,N_18406);
xor U19510 (N_19510,N_18091,N_18708);
nor U19511 (N_19511,N_18302,N_18243);
nor U19512 (N_19512,N_18034,N_18582);
or U19513 (N_19513,N_18798,N_18013);
xnor U19514 (N_19514,N_18982,N_18598);
xor U19515 (N_19515,N_18483,N_18809);
nor U19516 (N_19516,N_18023,N_18977);
nor U19517 (N_19517,N_18675,N_18094);
xor U19518 (N_19518,N_18449,N_18347);
nor U19519 (N_19519,N_18223,N_18504);
nand U19520 (N_19520,N_18887,N_18850);
and U19521 (N_19521,N_18235,N_18742);
nand U19522 (N_19522,N_18954,N_18851);
nand U19523 (N_19523,N_18902,N_18513);
xor U19524 (N_19524,N_18591,N_18807);
or U19525 (N_19525,N_18493,N_18641);
nand U19526 (N_19526,N_18371,N_18906);
nor U19527 (N_19527,N_18940,N_18008);
or U19528 (N_19528,N_18362,N_18708);
nand U19529 (N_19529,N_18105,N_18532);
xnor U19530 (N_19530,N_18241,N_18024);
nand U19531 (N_19531,N_18071,N_18814);
xor U19532 (N_19532,N_18278,N_18428);
nor U19533 (N_19533,N_18566,N_18804);
and U19534 (N_19534,N_18846,N_18585);
nand U19535 (N_19535,N_18542,N_18899);
and U19536 (N_19536,N_18278,N_18852);
nor U19537 (N_19537,N_18658,N_18813);
xor U19538 (N_19538,N_18136,N_18787);
or U19539 (N_19539,N_18698,N_18977);
xor U19540 (N_19540,N_18734,N_18345);
or U19541 (N_19541,N_18287,N_18291);
nor U19542 (N_19542,N_18239,N_18193);
nor U19543 (N_19543,N_18816,N_18078);
or U19544 (N_19544,N_18332,N_18544);
or U19545 (N_19545,N_18908,N_18675);
or U19546 (N_19546,N_18904,N_18558);
nor U19547 (N_19547,N_18969,N_18468);
and U19548 (N_19548,N_18623,N_18566);
and U19549 (N_19549,N_18277,N_18771);
nor U19550 (N_19550,N_18094,N_18075);
nor U19551 (N_19551,N_18807,N_18731);
and U19552 (N_19552,N_18107,N_18278);
xnor U19553 (N_19553,N_18019,N_18194);
xor U19554 (N_19554,N_18099,N_18745);
or U19555 (N_19555,N_18957,N_18893);
and U19556 (N_19556,N_18435,N_18487);
and U19557 (N_19557,N_18152,N_18012);
and U19558 (N_19558,N_18612,N_18743);
xnor U19559 (N_19559,N_18424,N_18392);
or U19560 (N_19560,N_18518,N_18832);
and U19561 (N_19561,N_18031,N_18653);
and U19562 (N_19562,N_18425,N_18877);
and U19563 (N_19563,N_18702,N_18460);
and U19564 (N_19564,N_18140,N_18693);
xor U19565 (N_19565,N_18467,N_18626);
nand U19566 (N_19566,N_18419,N_18858);
nand U19567 (N_19567,N_18318,N_18015);
xor U19568 (N_19568,N_18022,N_18289);
xor U19569 (N_19569,N_18449,N_18888);
or U19570 (N_19570,N_18475,N_18198);
nor U19571 (N_19571,N_18057,N_18426);
nor U19572 (N_19572,N_18516,N_18909);
or U19573 (N_19573,N_18746,N_18948);
and U19574 (N_19574,N_18491,N_18505);
nor U19575 (N_19575,N_18721,N_18606);
nor U19576 (N_19576,N_18768,N_18311);
and U19577 (N_19577,N_18467,N_18844);
or U19578 (N_19578,N_18100,N_18674);
and U19579 (N_19579,N_18546,N_18836);
xor U19580 (N_19580,N_18209,N_18328);
and U19581 (N_19581,N_18320,N_18207);
or U19582 (N_19582,N_18328,N_18299);
xnor U19583 (N_19583,N_18905,N_18353);
nor U19584 (N_19584,N_18945,N_18333);
nand U19585 (N_19585,N_18043,N_18349);
or U19586 (N_19586,N_18020,N_18798);
or U19587 (N_19587,N_18543,N_18294);
nor U19588 (N_19588,N_18672,N_18349);
nor U19589 (N_19589,N_18909,N_18374);
nor U19590 (N_19590,N_18220,N_18958);
xor U19591 (N_19591,N_18866,N_18043);
xor U19592 (N_19592,N_18790,N_18875);
xnor U19593 (N_19593,N_18920,N_18394);
or U19594 (N_19594,N_18125,N_18587);
or U19595 (N_19595,N_18147,N_18160);
xor U19596 (N_19596,N_18183,N_18586);
xnor U19597 (N_19597,N_18996,N_18536);
nand U19598 (N_19598,N_18794,N_18758);
nor U19599 (N_19599,N_18360,N_18684);
or U19600 (N_19600,N_18933,N_18873);
and U19601 (N_19601,N_18307,N_18720);
or U19602 (N_19602,N_18585,N_18499);
nor U19603 (N_19603,N_18355,N_18788);
xnor U19604 (N_19604,N_18265,N_18370);
xnor U19605 (N_19605,N_18389,N_18742);
nand U19606 (N_19606,N_18999,N_18613);
nor U19607 (N_19607,N_18941,N_18920);
and U19608 (N_19608,N_18060,N_18040);
nor U19609 (N_19609,N_18010,N_18617);
and U19610 (N_19610,N_18214,N_18241);
or U19611 (N_19611,N_18321,N_18796);
and U19612 (N_19612,N_18623,N_18568);
nor U19613 (N_19613,N_18862,N_18684);
or U19614 (N_19614,N_18928,N_18762);
xor U19615 (N_19615,N_18229,N_18286);
or U19616 (N_19616,N_18642,N_18341);
or U19617 (N_19617,N_18052,N_18107);
or U19618 (N_19618,N_18002,N_18915);
nand U19619 (N_19619,N_18348,N_18751);
nor U19620 (N_19620,N_18070,N_18978);
or U19621 (N_19621,N_18601,N_18373);
nand U19622 (N_19622,N_18655,N_18573);
nor U19623 (N_19623,N_18637,N_18883);
xor U19624 (N_19624,N_18273,N_18691);
or U19625 (N_19625,N_18297,N_18547);
or U19626 (N_19626,N_18793,N_18801);
nor U19627 (N_19627,N_18385,N_18832);
nor U19628 (N_19628,N_18598,N_18640);
nand U19629 (N_19629,N_18840,N_18982);
nor U19630 (N_19630,N_18825,N_18289);
nand U19631 (N_19631,N_18491,N_18391);
nand U19632 (N_19632,N_18646,N_18154);
nor U19633 (N_19633,N_18005,N_18067);
nand U19634 (N_19634,N_18644,N_18263);
and U19635 (N_19635,N_18621,N_18311);
and U19636 (N_19636,N_18510,N_18174);
nand U19637 (N_19637,N_18042,N_18016);
or U19638 (N_19638,N_18483,N_18374);
or U19639 (N_19639,N_18320,N_18278);
and U19640 (N_19640,N_18051,N_18761);
nand U19641 (N_19641,N_18037,N_18283);
or U19642 (N_19642,N_18239,N_18071);
xor U19643 (N_19643,N_18666,N_18877);
or U19644 (N_19644,N_18315,N_18699);
nor U19645 (N_19645,N_18739,N_18975);
xor U19646 (N_19646,N_18413,N_18757);
and U19647 (N_19647,N_18381,N_18965);
xnor U19648 (N_19648,N_18928,N_18455);
nand U19649 (N_19649,N_18345,N_18481);
nor U19650 (N_19650,N_18686,N_18533);
and U19651 (N_19651,N_18488,N_18465);
xor U19652 (N_19652,N_18888,N_18131);
or U19653 (N_19653,N_18416,N_18919);
nor U19654 (N_19654,N_18896,N_18591);
nand U19655 (N_19655,N_18917,N_18204);
nand U19656 (N_19656,N_18242,N_18534);
and U19657 (N_19657,N_18923,N_18678);
and U19658 (N_19658,N_18940,N_18405);
nand U19659 (N_19659,N_18608,N_18272);
and U19660 (N_19660,N_18549,N_18361);
and U19661 (N_19661,N_18272,N_18160);
or U19662 (N_19662,N_18855,N_18760);
and U19663 (N_19663,N_18294,N_18683);
xnor U19664 (N_19664,N_18951,N_18442);
nor U19665 (N_19665,N_18167,N_18653);
nor U19666 (N_19666,N_18008,N_18499);
nand U19667 (N_19667,N_18880,N_18323);
nor U19668 (N_19668,N_18296,N_18792);
xor U19669 (N_19669,N_18272,N_18715);
nor U19670 (N_19670,N_18568,N_18036);
xor U19671 (N_19671,N_18092,N_18592);
and U19672 (N_19672,N_18293,N_18861);
and U19673 (N_19673,N_18193,N_18103);
and U19674 (N_19674,N_18308,N_18567);
and U19675 (N_19675,N_18353,N_18105);
or U19676 (N_19676,N_18197,N_18225);
nor U19677 (N_19677,N_18041,N_18403);
nand U19678 (N_19678,N_18507,N_18288);
or U19679 (N_19679,N_18828,N_18468);
and U19680 (N_19680,N_18715,N_18198);
nor U19681 (N_19681,N_18516,N_18523);
or U19682 (N_19682,N_18806,N_18388);
xor U19683 (N_19683,N_18066,N_18099);
nor U19684 (N_19684,N_18294,N_18610);
nor U19685 (N_19685,N_18441,N_18641);
or U19686 (N_19686,N_18445,N_18035);
xnor U19687 (N_19687,N_18206,N_18714);
and U19688 (N_19688,N_18116,N_18107);
nor U19689 (N_19689,N_18679,N_18388);
nor U19690 (N_19690,N_18898,N_18168);
or U19691 (N_19691,N_18507,N_18932);
and U19692 (N_19692,N_18811,N_18592);
or U19693 (N_19693,N_18377,N_18576);
nor U19694 (N_19694,N_18367,N_18561);
nand U19695 (N_19695,N_18077,N_18159);
or U19696 (N_19696,N_18712,N_18374);
and U19697 (N_19697,N_18066,N_18952);
xor U19698 (N_19698,N_18854,N_18719);
xor U19699 (N_19699,N_18830,N_18966);
and U19700 (N_19700,N_18707,N_18956);
xnor U19701 (N_19701,N_18851,N_18045);
or U19702 (N_19702,N_18074,N_18815);
xnor U19703 (N_19703,N_18556,N_18958);
xnor U19704 (N_19704,N_18286,N_18085);
or U19705 (N_19705,N_18497,N_18482);
nand U19706 (N_19706,N_18493,N_18632);
nor U19707 (N_19707,N_18328,N_18898);
xnor U19708 (N_19708,N_18059,N_18243);
and U19709 (N_19709,N_18922,N_18441);
or U19710 (N_19710,N_18486,N_18502);
and U19711 (N_19711,N_18013,N_18643);
nand U19712 (N_19712,N_18976,N_18002);
nand U19713 (N_19713,N_18924,N_18779);
and U19714 (N_19714,N_18370,N_18895);
and U19715 (N_19715,N_18196,N_18872);
or U19716 (N_19716,N_18834,N_18456);
and U19717 (N_19717,N_18204,N_18127);
xnor U19718 (N_19718,N_18159,N_18974);
nand U19719 (N_19719,N_18959,N_18936);
xnor U19720 (N_19720,N_18532,N_18203);
nor U19721 (N_19721,N_18726,N_18552);
or U19722 (N_19722,N_18484,N_18470);
nor U19723 (N_19723,N_18710,N_18626);
xnor U19724 (N_19724,N_18134,N_18728);
nor U19725 (N_19725,N_18872,N_18611);
nand U19726 (N_19726,N_18160,N_18545);
nand U19727 (N_19727,N_18804,N_18849);
xor U19728 (N_19728,N_18066,N_18397);
nand U19729 (N_19729,N_18249,N_18902);
xnor U19730 (N_19730,N_18157,N_18805);
nor U19731 (N_19731,N_18001,N_18764);
xnor U19732 (N_19732,N_18063,N_18078);
and U19733 (N_19733,N_18646,N_18109);
nand U19734 (N_19734,N_18032,N_18624);
nand U19735 (N_19735,N_18997,N_18315);
and U19736 (N_19736,N_18961,N_18550);
and U19737 (N_19737,N_18328,N_18249);
nand U19738 (N_19738,N_18560,N_18111);
or U19739 (N_19739,N_18837,N_18101);
and U19740 (N_19740,N_18969,N_18176);
xor U19741 (N_19741,N_18857,N_18970);
or U19742 (N_19742,N_18427,N_18118);
nand U19743 (N_19743,N_18711,N_18617);
or U19744 (N_19744,N_18601,N_18441);
and U19745 (N_19745,N_18154,N_18308);
and U19746 (N_19746,N_18388,N_18449);
nor U19747 (N_19747,N_18172,N_18865);
xor U19748 (N_19748,N_18635,N_18276);
nand U19749 (N_19749,N_18110,N_18747);
or U19750 (N_19750,N_18758,N_18337);
xor U19751 (N_19751,N_18097,N_18805);
and U19752 (N_19752,N_18752,N_18004);
nor U19753 (N_19753,N_18480,N_18676);
xor U19754 (N_19754,N_18123,N_18408);
xnor U19755 (N_19755,N_18975,N_18579);
or U19756 (N_19756,N_18962,N_18156);
nand U19757 (N_19757,N_18782,N_18364);
xor U19758 (N_19758,N_18300,N_18010);
nor U19759 (N_19759,N_18773,N_18652);
xor U19760 (N_19760,N_18897,N_18636);
and U19761 (N_19761,N_18290,N_18393);
nor U19762 (N_19762,N_18842,N_18681);
nand U19763 (N_19763,N_18823,N_18455);
xnor U19764 (N_19764,N_18897,N_18604);
or U19765 (N_19765,N_18609,N_18244);
and U19766 (N_19766,N_18605,N_18501);
or U19767 (N_19767,N_18401,N_18611);
nor U19768 (N_19768,N_18664,N_18627);
nor U19769 (N_19769,N_18751,N_18163);
nor U19770 (N_19770,N_18239,N_18904);
xnor U19771 (N_19771,N_18326,N_18239);
xor U19772 (N_19772,N_18401,N_18395);
nor U19773 (N_19773,N_18337,N_18699);
xnor U19774 (N_19774,N_18523,N_18352);
or U19775 (N_19775,N_18716,N_18763);
xor U19776 (N_19776,N_18276,N_18565);
xnor U19777 (N_19777,N_18362,N_18705);
nand U19778 (N_19778,N_18538,N_18403);
and U19779 (N_19779,N_18457,N_18285);
nor U19780 (N_19780,N_18638,N_18434);
or U19781 (N_19781,N_18673,N_18552);
and U19782 (N_19782,N_18180,N_18379);
xor U19783 (N_19783,N_18609,N_18262);
nor U19784 (N_19784,N_18582,N_18553);
or U19785 (N_19785,N_18773,N_18311);
nor U19786 (N_19786,N_18437,N_18491);
or U19787 (N_19787,N_18989,N_18763);
nor U19788 (N_19788,N_18280,N_18207);
nand U19789 (N_19789,N_18195,N_18399);
nor U19790 (N_19790,N_18182,N_18611);
nor U19791 (N_19791,N_18256,N_18130);
nor U19792 (N_19792,N_18605,N_18979);
and U19793 (N_19793,N_18786,N_18186);
nand U19794 (N_19794,N_18044,N_18599);
xor U19795 (N_19795,N_18238,N_18939);
and U19796 (N_19796,N_18629,N_18120);
xnor U19797 (N_19797,N_18798,N_18585);
nand U19798 (N_19798,N_18391,N_18772);
and U19799 (N_19799,N_18812,N_18769);
nor U19800 (N_19800,N_18815,N_18202);
or U19801 (N_19801,N_18813,N_18099);
xnor U19802 (N_19802,N_18082,N_18862);
xnor U19803 (N_19803,N_18402,N_18725);
nor U19804 (N_19804,N_18960,N_18374);
and U19805 (N_19805,N_18071,N_18403);
nor U19806 (N_19806,N_18951,N_18188);
nand U19807 (N_19807,N_18465,N_18919);
nor U19808 (N_19808,N_18539,N_18032);
xnor U19809 (N_19809,N_18165,N_18720);
nand U19810 (N_19810,N_18374,N_18789);
nor U19811 (N_19811,N_18774,N_18392);
or U19812 (N_19812,N_18392,N_18852);
and U19813 (N_19813,N_18748,N_18024);
nand U19814 (N_19814,N_18462,N_18438);
nand U19815 (N_19815,N_18691,N_18284);
or U19816 (N_19816,N_18028,N_18118);
nand U19817 (N_19817,N_18297,N_18773);
or U19818 (N_19818,N_18368,N_18668);
nand U19819 (N_19819,N_18307,N_18812);
nand U19820 (N_19820,N_18467,N_18755);
nor U19821 (N_19821,N_18189,N_18747);
xnor U19822 (N_19822,N_18710,N_18515);
and U19823 (N_19823,N_18042,N_18003);
nand U19824 (N_19824,N_18661,N_18345);
and U19825 (N_19825,N_18330,N_18611);
xnor U19826 (N_19826,N_18217,N_18577);
and U19827 (N_19827,N_18195,N_18946);
xnor U19828 (N_19828,N_18159,N_18950);
or U19829 (N_19829,N_18045,N_18516);
and U19830 (N_19830,N_18773,N_18783);
and U19831 (N_19831,N_18846,N_18597);
and U19832 (N_19832,N_18161,N_18629);
and U19833 (N_19833,N_18758,N_18963);
or U19834 (N_19834,N_18683,N_18309);
or U19835 (N_19835,N_18295,N_18596);
nand U19836 (N_19836,N_18489,N_18172);
and U19837 (N_19837,N_18628,N_18815);
nand U19838 (N_19838,N_18281,N_18137);
and U19839 (N_19839,N_18163,N_18772);
xnor U19840 (N_19840,N_18816,N_18792);
nand U19841 (N_19841,N_18032,N_18140);
nor U19842 (N_19842,N_18797,N_18847);
nor U19843 (N_19843,N_18655,N_18538);
xnor U19844 (N_19844,N_18257,N_18220);
and U19845 (N_19845,N_18244,N_18298);
and U19846 (N_19846,N_18511,N_18971);
nand U19847 (N_19847,N_18130,N_18236);
or U19848 (N_19848,N_18150,N_18232);
nor U19849 (N_19849,N_18833,N_18942);
and U19850 (N_19850,N_18854,N_18065);
xor U19851 (N_19851,N_18097,N_18449);
and U19852 (N_19852,N_18057,N_18889);
xnor U19853 (N_19853,N_18603,N_18212);
and U19854 (N_19854,N_18939,N_18662);
or U19855 (N_19855,N_18954,N_18104);
nand U19856 (N_19856,N_18938,N_18455);
or U19857 (N_19857,N_18444,N_18655);
and U19858 (N_19858,N_18350,N_18118);
and U19859 (N_19859,N_18672,N_18590);
nand U19860 (N_19860,N_18403,N_18803);
nor U19861 (N_19861,N_18803,N_18932);
nor U19862 (N_19862,N_18829,N_18037);
nand U19863 (N_19863,N_18701,N_18426);
xnor U19864 (N_19864,N_18539,N_18303);
and U19865 (N_19865,N_18976,N_18956);
nand U19866 (N_19866,N_18440,N_18981);
xnor U19867 (N_19867,N_18538,N_18457);
nor U19868 (N_19868,N_18534,N_18444);
nand U19869 (N_19869,N_18107,N_18884);
and U19870 (N_19870,N_18002,N_18040);
nor U19871 (N_19871,N_18968,N_18278);
and U19872 (N_19872,N_18548,N_18641);
nor U19873 (N_19873,N_18223,N_18740);
nor U19874 (N_19874,N_18800,N_18288);
and U19875 (N_19875,N_18600,N_18427);
nor U19876 (N_19876,N_18403,N_18440);
nand U19877 (N_19877,N_18922,N_18301);
nand U19878 (N_19878,N_18259,N_18395);
nor U19879 (N_19879,N_18455,N_18211);
nand U19880 (N_19880,N_18858,N_18964);
and U19881 (N_19881,N_18725,N_18976);
and U19882 (N_19882,N_18093,N_18709);
nor U19883 (N_19883,N_18544,N_18539);
nor U19884 (N_19884,N_18890,N_18540);
or U19885 (N_19885,N_18218,N_18422);
and U19886 (N_19886,N_18400,N_18127);
or U19887 (N_19887,N_18891,N_18906);
nand U19888 (N_19888,N_18180,N_18423);
and U19889 (N_19889,N_18097,N_18249);
nor U19890 (N_19890,N_18237,N_18277);
or U19891 (N_19891,N_18799,N_18360);
xor U19892 (N_19892,N_18376,N_18363);
and U19893 (N_19893,N_18622,N_18394);
or U19894 (N_19894,N_18935,N_18364);
or U19895 (N_19895,N_18632,N_18849);
nor U19896 (N_19896,N_18482,N_18835);
or U19897 (N_19897,N_18365,N_18487);
xnor U19898 (N_19898,N_18874,N_18541);
xor U19899 (N_19899,N_18374,N_18770);
nor U19900 (N_19900,N_18269,N_18044);
nor U19901 (N_19901,N_18695,N_18619);
nor U19902 (N_19902,N_18837,N_18294);
xor U19903 (N_19903,N_18299,N_18419);
nand U19904 (N_19904,N_18861,N_18801);
nor U19905 (N_19905,N_18288,N_18918);
and U19906 (N_19906,N_18848,N_18833);
nor U19907 (N_19907,N_18519,N_18017);
or U19908 (N_19908,N_18822,N_18376);
nand U19909 (N_19909,N_18587,N_18833);
nand U19910 (N_19910,N_18347,N_18158);
xor U19911 (N_19911,N_18606,N_18396);
xnor U19912 (N_19912,N_18960,N_18187);
nor U19913 (N_19913,N_18065,N_18434);
or U19914 (N_19914,N_18939,N_18682);
xor U19915 (N_19915,N_18176,N_18701);
xnor U19916 (N_19916,N_18084,N_18649);
nand U19917 (N_19917,N_18239,N_18657);
and U19918 (N_19918,N_18286,N_18646);
and U19919 (N_19919,N_18179,N_18735);
and U19920 (N_19920,N_18808,N_18649);
xnor U19921 (N_19921,N_18202,N_18086);
xnor U19922 (N_19922,N_18984,N_18644);
xnor U19923 (N_19923,N_18502,N_18619);
and U19924 (N_19924,N_18571,N_18394);
or U19925 (N_19925,N_18697,N_18550);
nand U19926 (N_19926,N_18415,N_18457);
xor U19927 (N_19927,N_18561,N_18858);
or U19928 (N_19928,N_18231,N_18536);
nor U19929 (N_19929,N_18999,N_18593);
nor U19930 (N_19930,N_18776,N_18386);
xnor U19931 (N_19931,N_18289,N_18193);
or U19932 (N_19932,N_18083,N_18659);
and U19933 (N_19933,N_18898,N_18025);
and U19934 (N_19934,N_18052,N_18177);
nand U19935 (N_19935,N_18659,N_18618);
and U19936 (N_19936,N_18281,N_18441);
xor U19937 (N_19937,N_18349,N_18920);
nor U19938 (N_19938,N_18927,N_18114);
or U19939 (N_19939,N_18627,N_18436);
xnor U19940 (N_19940,N_18371,N_18257);
nor U19941 (N_19941,N_18011,N_18046);
nor U19942 (N_19942,N_18299,N_18828);
and U19943 (N_19943,N_18031,N_18459);
nor U19944 (N_19944,N_18250,N_18458);
xor U19945 (N_19945,N_18823,N_18044);
or U19946 (N_19946,N_18263,N_18214);
or U19947 (N_19947,N_18539,N_18733);
xor U19948 (N_19948,N_18369,N_18812);
nor U19949 (N_19949,N_18302,N_18265);
and U19950 (N_19950,N_18190,N_18905);
and U19951 (N_19951,N_18090,N_18614);
and U19952 (N_19952,N_18732,N_18383);
nand U19953 (N_19953,N_18604,N_18582);
or U19954 (N_19954,N_18721,N_18684);
nand U19955 (N_19955,N_18139,N_18928);
nor U19956 (N_19956,N_18341,N_18570);
and U19957 (N_19957,N_18010,N_18086);
nand U19958 (N_19958,N_18435,N_18586);
nand U19959 (N_19959,N_18062,N_18449);
nand U19960 (N_19960,N_18821,N_18076);
xor U19961 (N_19961,N_18841,N_18604);
xor U19962 (N_19962,N_18201,N_18334);
and U19963 (N_19963,N_18259,N_18543);
or U19964 (N_19964,N_18115,N_18023);
or U19965 (N_19965,N_18733,N_18167);
nor U19966 (N_19966,N_18240,N_18104);
xnor U19967 (N_19967,N_18666,N_18518);
or U19968 (N_19968,N_18377,N_18696);
nor U19969 (N_19969,N_18896,N_18673);
nor U19970 (N_19970,N_18622,N_18582);
nand U19971 (N_19971,N_18217,N_18267);
or U19972 (N_19972,N_18768,N_18726);
and U19973 (N_19973,N_18090,N_18684);
nor U19974 (N_19974,N_18471,N_18073);
xor U19975 (N_19975,N_18138,N_18049);
or U19976 (N_19976,N_18811,N_18486);
xnor U19977 (N_19977,N_18081,N_18442);
nor U19978 (N_19978,N_18233,N_18133);
or U19979 (N_19979,N_18895,N_18896);
and U19980 (N_19980,N_18018,N_18583);
xor U19981 (N_19981,N_18344,N_18380);
nor U19982 (N_19982,N_18027,N_18778);
xor U19983 (N_19983,N_18184,N_18761);
and U19984 (N_19984,N_18642,N_18501);
or U19985 (N_19985,N_18313,N_18290);
xor U19986 (N_19986,N_18812,N_18521);
xnor U19987 (N_19987,N_18211,N_18847);
nor U19988 (N_19988,N_18437,N_18867);
and U19989 (N_19989,N_18428,N_18042);
and U19990 (N_19990,N_18446,N_18523);
nand U19991 (N_19991,N_18878,N_18277);
nor U19992 (N_19992,N_18437,N_18727);
and U19993 (N_19993,N_18587,N_18547);
or U19994 (N_19994,N_18250,N_18185);
nor U19995 (N_19995,N_18241,N_18817);
and U19996 (N_19996,N_18672,N_18538);
and U19997 (N_19997,N_18728,N_18392);
and U19998 (N_19998,N_18953,N_18286);
and U19999 (N_19999,N_18535,N_18082);
or U20000 (N_20000,N_19430,N_19740);
or U20001 (N_20001,N_19285,N_19220);
or U20002 (N_20002,N_19025,N_19247);
nor U20003 (N_20003,N_19949,N_19443);
nand U20004 (N_20004,N_19355,N_19624);
nand U20005 (N_20005,N_19792,N_19561);
nor U20006 (N_20006,N_19992,N_19349);
and U20007 (N_20007,N_19032,N_19238);
or U20008 (N_20008,N_19447,N_19436);
and U20009 (N_20009,N_19791,N_19028);
xor U20010 (N_20010,N_19834,N_19172);
and U20011 (N_20011,N_19521,N_19118);
and U20012 (N_20012,N_19309,N_19694);
xor U20013 (N_20013,N_19876,N_19395);
nand U20014 (N_20014,N_19124,N_19906);
and U20015 (N_20015,N_19986,N_19319);
nand U20016 (N_20016,N_19228,N_19940);
xor U20017 (N_20017,N_19081,N_19122);
and U20018 (N_20018,N_19932,N_19979);
nand U20019 (N_20019,N_19221,N_19223);
xnor U20020 (N_20020,N_19674,N_19704);
or U20021 (N_20021,N_19788,N_19782);
nand U20022 (N_20022,N_19564,N_19554);
xnor U20023 (N_20023,N_19604,N_19277);
xor U20024 (N_20024,N_19423,N_19983);
nor U20025 (N_20025,N_19398,N_19669);
or U20026 (N_20026,N_19354,N_19506);
and U20027 (N_20027,N_19017,N_19548);
or U20028 (N_20028,N_19311,N_19848);
nor U20029 (N_20029,N_19636,N_19997);
or U20030 (N_20030,N_19497,N_19568);
and U20031 (N_20031,N_19350,N_19952);
xor U20032 (N_20032,N_19996,N_19900);
and U20033 (N_20033,N_19327,N_19258);
nand U20034 (N_20034,N_19377,N_19212);
nand U20035 (N_20035,N_19918,N_19606);
nand U20036 (N_20036,N_19840,N_19888);
xnor U20037 (N_20037,N_19255,N_19382);
and U20038 (N_20038,N_19965,N_19747);
nor U20039 (N_20039,N_19441,N_19597);
and U20040 (N_20040,N_19093,N_19544);
or U20041 (N_20041,N_19562,N_19806);
nand U20042 (N_20042,N_19077,N_19558);
nor U20043 (N_20043,N_19330,N_19390);
nor U20044 (N_20044,N_19938,N_19642);
nor U20045 (N_20045,N_19268,N_19131);
nand U20046 (N_20046,N_19383,N_19452);
and U20047 (N_20047,N_19407,N_19508);
nor U20048 (N_20048,N_19162,N_19372);
nor U20049 (N_20049,N_19192,N_19088);
xnor U20050 (N_20050,N_19978,N_19967);
or U20051 (N_20051,N_19920,N_19789);
nor U20052 (N_20052,N_19805,N_19307);
or U20053 (N_20053,N_19030,N_19526);
nand U20054 (N_20054,N_19408,N_19942);
nand U20055 (N_20055,N_19075,N_19535);
and U20056 (N_20056,N_19478,N_19274);
nor U20057 (N_20057,N_19374,N_19150);
nand U20058 (N_20058,N_19240,N_19061);
nand U20059 (N_20059,N_19721,N_19546);
nor U20060 (N_20060,N_19011,N_19995);
nor U20061 (N_20061,N_19640,N_19998);
and U20062 (N_20062,N_19246,N_19818);
nand U20063 (N_20063,N_19830,N_19187);
nor U20064 (N_20064,N_19801,N_19727);
nand U20065 (N_20065,N_19076,N_19643);
xnor U20066 (N_20066,N_19144,N_19052);
or U20067 (N_20067,N_19582,N_19173);
or U20068 (N_20068,N_19631,N_19917);
nor U20069 (N_20069,N_19778,N_19074);
and U20070 (N_20070,N_19632,N_19233);
or U20071 (N_20071,N_19001,N_19894);
xnor U20072 (N_20072,N_19874,N_19990);
nand U20073 (N_20073,N_19413,N_19189);
nand U20074 (N_20074,N_19931,N_19108);
and U20075 (N_20075,N_19344,N_19007);
nand U20076 (N_20076,N_19112,N_19299);
nand U20077 (N_20077,N_19819,N_19677);
nor U20078 (N_20078,N_19097,N_19483);
nand U20079 (N_20079,N_19324,N_19200);
nor U20080 (N_20080,N_19058,N_19620);
or U20081 (N_20081,N_19461,N_19852);
nor U20082 (N_20082,N_19293,N_19456);
or U20083 (N_20083,N_19595,N_19831);
xor U20084 (N_20084,N_19132,N_19099);
nand U20085 (N_20085,N_19439,N_19589);
nand U20086 (N_20086,N_19066,N_19466);
and U20087 (N_20087,N_19947,N_19684);
nor U20088 (N_20088,N_19808,N_19579);
xor U20089 (N_20089,N_19550,N_19667);
or U20090 (N_20090,N_19446,N_19871);
and U20091 (N_20091,N_19037,N_19518);
nor U20092 (N_20092,N_19083,N_19839);
or U20093 (N_20093,N_19264,N_19208);
and U20094 (N_20094,N_19257,N_19096);
or U20095 (N_20095,N_19085,N_19087);
xor U20096 (N_20096,N_19485,N_19051);
nor U20097 (N_20097,N_19270,N_19272);
or U20098 (N_20098,N_19673,N_19714);
and U20099 (N_20099,N_19232,N_19929);
xnor U20100 (N_20100,N_19154,N_19729);
or U20101 (N_20101,N_19474,N_19498);
or U20102 (N_20102,N_19351,N_19322);
and U20103 (N_20103,N_19204,N_19610);
nand U20104 (N_20104,N_19142,N_19072);
and U20105 (N_20105,N_19889,N_19502);
and U20106 (N_20106,N_19475,N_19434);
or U20107 (N_20107,N_19013,N_19703);
or U20108 (N_20108,N_19754,N_19892);
or U20109 (N_20109,N_19445,N_19868);
nand U20110 (N_20110,N_19024,N_19411);
nor U20111 (N_20111,N_19707,N_19713);
or U20112 (N_20112,N_19731,N_19572);
or U20113 (N_20113,N_19607,N_19010);
xor U20114 (N_20114,N_19281,N_19545);
and U20115 (N_20115,N_19301,N_19416);
nand U20116 (N_20116,N_19450,N_19205);
and U20117 (N_20117,N_19811,N_19318);
or U20118 (N_20118,N_19662,N_19380);
nor U20119 (N_20119,N_19050,N_19251);
nor U20120 (N_20120,N_19280,N_19214);
and U20121 (N_20121,N_19883,N_19089);
xnor U20122 (N_20122,N_19019,N_19463);
nand U20123 (N_20123,N_19578,N_19537);
or U20124 (N_20124,N_19580,N_19215);
xor U20125 (N_20125,N_19143,N_19614);
nand U20126 (N_20126,N_19903,N_19798);
nor U20127 (N_20127,N_19298,N_19807);
and U20128 (N_20128,N_19827,N_19339);
nor U20129 (N_20129,N_19417,N_19273);
and U20130 (N_20130,N_19371,N_19147);
nand U20131 (N_20131,N_19628,N_19209);
or U20132 (N_20132,N_19263,N_19911);
nor U20133 (N_20133,N_19760,N_19464);
xnor U20134 (N_20134,N_19676,N_19974);
nand U20135 (N_20135,N_19259,N_19287);
nand U20136 (N_20136,N_19551,N_19936);
nor U20137 (N_20137,N_19762,N_19338);
and U20138 (N_20138,N_19513,N_19717);
nor U20139 (N_20139,N_19822,N_19552);
nor U20140 (N_20140,N_19419,N_19886);
nor U20141 (N_20141,N_19457,N_19119);
xnor U20142 (N_20142,N_19418,N_19412);
xnor U20143 (N_20143,N_19756,N_19896);
nor U20144 (N_20144,N_19786,N_19031);
and U20145 (N_20145,N_19183,N_19718);
xnor U20146 (N_20146,N_19970,N_19869);
nor U20147 (N_20147,N_19235,N_19193);
xnor U20148 (N_20148,N_19462,N_19658);
xnor U20149 (N_20149,N_19977,N_19388);
nand U20150 (N_20150,N_19916,N_19337);
or U20151 (N_20151,N_19837,N_19184);
and U20152 (N_20152,N_19661,N_19780);
and U20153 (N_20153,N_19591,N_19878);
or U20154 (N_20154,N_19531,N_19895);
and U20155 (N_20155,N_19176,N_19117);
and U20156 (N_20156,N_19091,N_19328);
or U20157 (N_20157,N_19167,N_19006);
nand U20158 (N_20158,N_19752,N_19841);
nor U20159 (N_20159,N_19758,N_19104);
and U20160 (N_20160,N_19479,N_19647);
and U20161 (N_20161,N_19206,N_19467);
nor U20162 (N_20162,N_19700,N_19465);
nand U20163 (N_20163,N_19080,N_19849);
nor U20164 (N_20164,N_19799,N_19512);
nor U20165 (N_20165,N_19429,N_19295);
or U20166 (N_20166,N_19079,N_19260);
nand U20167 (N_20167,N_19415,N_19427);
xnor U20168 (N_20168,N_19044,N_19120);
nand U20169 (N_20169,N_19660,N_19757);
xor U20170 (N_20170,N_19618,N_19809);
and U20171 (N_20171,N_19766,N_19516);
or U20172 (N_20172,N_19431,N_19765);
nand U20173 (N_20173,N_19034,N_19015);
nand U20174 (N_20174,N_19616,N_19627);
nor U20175 (N_20175,N_19770,N_19370);
and U20176 (N_20176,N_19468,N_19865);
and U20177 (N_20177,N_19243,N_19541);
or U20178 (N_20178,N_19279,N_19697);
and U20179 (N_20179,N_19369,N_19347);
nor U20180 (N_20180,N_19596,N_19510);
nor U20181 (N_20181,N_19123,N_19067);
nand U20182 (N_20182,N_19743,N_19316);
nand U20183 (N_20183,N_19891,N_19585);
xnor U20184 (N_20184,N_19432,N_19321);
xor U20185 (N_20185,N_19082,N_19353);
nand U20186 (N_20186,N_19605,N_19068);
xor U20187 (N_20187,N_19682,N_19018);
nor U20188 (N_20188,N_19042,N_19857);
or U20189 (N_20189,N_19484,N_19248);
and U20190 (N_20190,N_19725,N_19414);
or U20191 (N_20191,N_19146,N_19609);
and U20192 (N_20192,N_19135,N_19543);
or U20193 (N_20193,N_19312,N_19515);
xnor U20194 (N_20194,N_19329,N_19164);
nor U20195 (N_20195,N_19879,N_19185);
xor U20196 (N_20196,N_19125,N_19884);
xnor U20197 (N_20197,N_19138,N_19368);
or U20198 (N_20198,N_19856,N_19656);
xnor U20199 (N_20199,N_19955,N_19245);
nor U20200 (N_20200,N_19927,N_19492);
and U20201 (N_20201,N_19045,N_19675);
or U20202 (N_20202,N_19207,N_19824);
or U20203 (N_20203,N_19180,N_19004);
or U20204 (N_20204,N_19800,N_19750);
nor U20205 (N_20205,N_19113,N_19406);
nand U20206 (N_20206,N_19576,N_19379);
nand U20207 (N_20207,N_19644,N_19386);
nand U20208 (N_20208,N_19962,N_19313);
nor U20209 (N_20209,N_19863,N_19570);
or U20210 (N_20210,N_19236,N_19823);
or U20211 (N_20211,N_19688,N_19654);
xor U20212 (N_20212,N_19873,N_19401);
xnor U20213 (N_20213,N_19198,N_19393);
or U20214 (N_20214,N_19128,N_19016);
and U20215 (N_20215,N_19336,N_19744);
xor U20216 (N_20216,N_19389,N_19957);
or U20217 (N_20217,N_19496,N_19709);
or U20218 (N_20218,N_19772,N_19608);
or U20219 (N_20219,N_19774,N_19925);
or U20220 (N_20220,N_19861,N_19821);
nor U20221 (N_20221,N_19685,N_19095);
and U20222 (N_20222,N_19064,N_19086);
nor U20223 (N_20223,N_19733,N_19972);
and U20224 (N_20224,N_19194,N_19375);
nand U20225 (N_20225,N_19812,N_19795);
or U20226 (N_20226,N_19509,N_19532);
xnor U20227 (N_20227,N_19899,N_19262);
or U20228 (N_20228,N_19078,N_19043);
or U20229 (N_20229,N_19569,N_19603);
xor U20230 (N_20230,N_19790,N_19993);
nor U20231 (N_20231,N_19420,N_19858);
xnor U20232 (N_20232,N_19216,N_19424);
or U20233 (N_20233,N_19964,N_19875);
xnor U20234 (N_20234,N_19060,N_19810);
or U20235 (N_20235,N_19181,N_19951);
xnor U20236 (N_20236,N_19842,N_19168);
and U20237 (N_20237,N_19622,N_19003);
xor U20238 (N_20238,N_19557,N_19469);
and U20239 (N_20239,N_19559,N_19470);
xnor U20240 (N_20240,N_19308,N_19035);
and U20241 (N_20241,N_19290,N_19499);
nand U20242 (N_20242,N_19706,N_19009);
xor U20243 (N_20243,N_19738,N_19110);
and U20244 (N_20244,N_19048,N_19663);
nand U20245 (N_20245,N_19981,N_19956);
or U20246 (N_20246,N_19057,N_19224);
nor U20247 (N_20247,N_19053,N_19271);
xor U20248 (N_20248,N_19503,N_19973);
or U20249 (N_20249,N_19571,N_19156);
or U20250 (N_20250,N_19681,N_19333);
xor U20251 (N_20251,N_19442,N_19332);
or U20252 (N_20252,N_19672,N_19635);
nor U20253 (N_20253,N_19493,N_19140);
xnor U20254 (N_20254,N_19930,N_19149);
nor U20255 (N_20255,N_19405,N_19989);
and U20256 (N_20256,N_19239,N_19202);
xor U20257 (N_20257,N_19433,N_19828);
nand U20258 (N_20258,N_19387,N_19103);
xnor U20259 (N_20259,N_19400,N_19749);
and U20260 (N_20260,N_19779,N_19267);
xnor U20261 (N_20261,N_19802,N_19555);
nor U20262 (N_20262,N_19547,N_19489);
nand U20263 (N_20263,N_19437,N_19381);
xor U20264 (N_20264,N_19678,N_19665);
and U20265 (N_20265,N_19907,N_19121);
or U20266 (N_20266,N_19577,N_19645);
nand U20267 (N_20267,N_19594,N_19623);
nand U20268 (N_20268,N_19190,N_19567);
nor U20269 (N_20269,N_19860,N_19084);
xor U20270 (N_20270,N_19928,N_19314);
and U20271 (N_20271,N_19683,N_19519);
nand U20272 (N_20272,N_19611,N_19944);
nor U20273 (N_20273,N_19305,N_19453);
nand U20274 (N_20274,N_19679,N_19961);
nor U20275 (N_20275,N_19670,N_19012);
xor U20276 (N_20276,N_19127,N_19363);
or U20277 (N_20277,N_19912,N_19999);
nor U20278 (N_20278,N_19399,N_19935);
nor U20279 (N_20279,N_19708,N_19639);
xor U20280 (N_20280,N_19748,N_19094);
nor U20281 (N_20281,N_19473,N_19225);
xor U20282 (N_20282,N_19793,N_19817);
nand U20283 (N_20283,N_19695,N_19111);
nand U20284 (N_20284,N_19211,N_19556);
and U20285 (N_20285,N_19573,N_19870);
and U20286 (N_20286,N_19219,N_19195);
nor U20287 (N_20287,N_19540,N_19887);
nor U20288 (N_20288,N_19833,N_19459);
and U20289 (N_20289,N_19291,N_19230);
nand U20290 (N_20290,N_19227,N_19534);
xor U20291 (N_20291,N_19777,N_19361);
nand U20292 (N_20292,N_19056,N_19002);
xnor U20293 (N_20293,N_19449,N_19910);
xor U20294 (N_20294,N_19836,N_19813);
and U20295 (N_20295,N_19711,N_19784);
or U20296 (N_20296,N_19523,N_19101);
and U20297 (N_20297,N_19862,N_19692);
and U20298 (N_20298,N_19880,N_19397);
or U20299 (N_20299,N_19844,N_19289);
nand U20300 (N_20300,N_19601,N_19297);
nand U20301 (N_20301,N_19574,N_19008);
or U20302 (N_20302,N_19092,N_19536);
nor U20303 (N_20303,N_19356,N_19719);
xor U20304 (N_20304,N_19488,N_19746);
xor U20305 (N_20305,N_19693,N_19376);
xnor U20306 (N_20306,N_19460,N_19587);
xnor U20307 (N_20307,N_19520,N_19481);
and U20308 (N_20308,N_19155,N_19373);
nand U20309 (N_20309,N_19775,N_19764);
nor U20310 (N_20310,N_19166,N_19507);
and U20311 (N_20311,N_19710,N_19438);
or U20312 (N_20312,N_19838,N_19161);
or U20313 (N_20313,N_19022,N_19751);
xor U20314 (N_20314,N_19549,N_19539);
nor U20315 (N_20315,N_19741,N_19114);
or U20316 (N_20316,N_19410,N_19486);
nor U20317 (N_20317,N_19511,N_19637);
or U20318 (N_20318,N_19106,N_19901);
or U20319 (N_20319,N_19040,N_19340);
nor U20320 (N_20320,N_19046,N_19855);
xnor U20321 (N_20321,N_19626,N_19435);
and U20322 (N_20322,N_19222,N_19881);
or U20323 (N_20323,N_19612,N_19027);
xnor U20324 (N_20324,N_19179,N_19480);
xor U20325 (N_20325,N_19794,N_19458);
nand U20326 (N_20326,N_19186,N_19864);
or U20327 (N_20327,N_19409,N_19755);
xor U20328 (N_20328,N_19249,N_19139);
or U20329 (N_20329,N_19565,N_19563);
xor U20330 (N_20330,N_19256,N_19177);
nand U20331 (N_20331,N_19734,N_19958);
nand U20332 (N_20332,N_19334,N_19945);
and U20333 (N_20333,N_19722,N_19275);
nand U20334 (N_20334,N_19199,N_19505);
nand U20335 (N_20335,N_19394,N_19843);
nor U20336 (N_20336,N_19472,N_19196);
nor U20337 (N_20337,N_19145,N_19129);
or U20338 (N_20338,N_19987,N_19953);
nand U20339 (N_20339,N_19923,N_19362);
or U20340 (N_20340,N_19615,N_19702);
nor U20341 (N_20341,N_19638,N_19698);
or U20342 (N_20342,N_19882,N_19763);
xor U20343 (N_20343,N_19317,N_19598);
and U20344 (N_20344,N_19524,N_19921);
and U20345 (N_20345,N_19422,N_19530);
xnor U20346 (N_20346,N_19366,N_19933);
xor U20347 (N_20347,N_19490,N_19872);
nand U20348 (N_20348,N_19231,N_19845);
nor U20349 (N_20349,N_19165,N_19253);
and U20350 (N_20350,N_19304,N_19278);
or U20351 (N_20351,N_19100,N_19252);
or U20352 (N_20352,N_19266,N_19360);
nand U20353 (N_20353,N_19835,N_19847);
or U20354 (N_20354,N_19197,N_19527);
or U20355 (N_20355,N_19343,N_19866);
or U20356 (N_20356,N_19021,N_19671);
or U20357 (N_20357,N_19217,N_19629);
nor U20358 (N_20358,N_19384,N_19716);
and U20359 (N_20359,N_19396,N_19724);
nand U20360 (N_20360,N_19153,N_19768);
nand U20361 (N_20361,N_19890,N_19804);
xnor U20362 (N_20362,N_19500,N_19728);
xor U20363 (N_20363,N_19403,N_19310);
and U20364 (N_20364,N_19630,N_19471);
xor U20365 (N_20365,N_19991,N_19054);
nor U20366 (N_20366,N_19593,N_19980);
and U20367 (N_20367,N_19924,N_19657);
nand U20368 (N_20368,N_19915,N_19325);
nand U20369 (N_20369,N_19542,N_19946);
or U20370 (N_20370,N_19038,N_19158);
and U20371 (N_20371,N_19528,N_19617);
and U20372 (N_20372,N_19976,N_19136);
or U20373 (N_20373,N_19680,N_19583);
nand U20374 (N_20374,N_19689,N_19908);
and U20375 (N_20375,N_19323,N_19282);
nand U20376 (N_20376,N_19276,N_19994);
or U20377 (N_20377,N_19047,N_19364);
nor U20378 (N_20378,N_19742,N_19444);
xor U20379 (N_20379,N_19699,N_19402);
nand U20380 (N_20380,N_19820,N_19306);
nor U20381 (N_20381,N_19455,N_19062);
and U20382 (N_20382,N_19071,N_19041);
or U20383 (N_20383,N_19476,N_19592);
and U20384 (N_20384,N_19226,N_19352);
and U20385 (N_20385,N_19115,N_19055);
xor U20386 (N_20386,N_19283,N_19781);
nor U20387 (N_20387,N_19948,N_19909);
xnor U20388 (N_20388,N_19581,N_19826);
and U20389 (N_20389,N_19234,N_19504);
nand U20390 (N_20390,N_19602,N_19613);
xnor U20391 (N_20391,N_19664,N_19169);
and U20392 (N_20392,N_19898,N_19367);
nor U20393 (N_20393,N_19959,N_19982);
nor U20394 (N_20394,N_19715,N_19553);
nor U20395 (N_20395,N_19098,N_19296);
nand U20396 (N_20396,N_19803,N_19648);
nand U20397 (N_20397,N_19365,N_19600);
and U20398 (N_20398,N_19421,N_19939);
and U20399 (N_20399,N_19178,N_19175);
and U20400 (N_20400,N_19913,N_19392);
or U20401 (N_20401,N_19269,N_19157);
nand U20402 (N_20402,N_19163,N_19482);
and U20403 (N_20403,N_19853,N_19065);
xnor U20404 (N_20404,N_19130,N_19914);
or U20405 (N_20405,N_19854,N_19425);
xnor U20406 (N_20406,N_19171,N_19491);
and U20407 (N_20407,N_19391,N_19102);
nand U20408 (N_20408,N_19797,N_19753);
xor U20409 (N_20409,N_19937,N_19825);
nor U20410 (N_20410,N_19023,N_19730);
nor U20411 (N_20411,N_19776,N_19292);
and U20412 (N_20412,N_19877,N_19090);
and U20413 (N_20413,N_19904,N_19960);
xnor U20414 (N_20414,N_19922,N_19487);
and U20415 (N_20415,N_19341,N_19653);
xor U20416 (N_20416,N_19621,N_19655);
nor U20417 (N_20417,N_19326,N_19969);
nor U20418 (N_20418,N_19448,N_19033);
xor U20419 (N_20419,N_19796,N_19566);
or U20420 (N_20420,N_19735,N_19160);
xor U20421 (N_20421,N_19315,N_19346);
nor U20422 (N_20422,N_19723,N_19651);
or U20423 (N_20423,N_19771,N_19404);
or U20424 (N_20424,N_19966,N_19934);
and U20425 (N_20425,N_19288,N_19885);
or U20426 (N_20426,N_19634,N_19737);
nor U20427 (N_20427,N_19451,N_19893);
and U20428 (N_20428,N_19494,N_19850);
nor U20429 (N_20429,N_19345,N_19059);
and U20430 (N_20430,N_19649,N_19652);
and U20431 (N_20431,N_19529,N_19303);
xnor U20432 (N_20432,N_19668,N_19440);
xor U20433 (N_20433,N_19761,N_19696);
nor U20434 (N_20434,N_19701,N_19666);
nand U20435 (N_20435,N_19968,N_19029);
or U20436 (N_20436,N_19941,N_19633);
nor U20437 (N_20437,N_19000,N_19203);
nand U20438 (N_20438,N_19152,N_19182);
nand U20439 (N_20439,N_19590,N_19141);
nor U20440 (N_20440,N_19357,N_19174);
xor U20441 (N_20441,N_19428,N_19584);
nor U20442 (N_20442,N_19359,N_19829);
or U20443 (N_20443,N_19241,N_19134);
nand U20444 (N_20444,N_19650,N_19063);
nand U20445 (N_20445,N_19816,N_19105);
xor U20446 (N_20446,N_19641,N_19599);
and U20447 (N_20447,N_19244,N_19984);
or U20448 (N_20448,N_19963,N_19213);
or U20449 (N_20449,N_19191,N_19905);
or U20450 (N_20450,N_19646,N_19320);
or U20451 (N_20451,N_19039,N_19342);
and U20452 (N_20452,N_19107,N_19358);
or U20453 (N_20453,N_19815,N_19294);
nand U20454 (N_20454,N_19170,N_19335);
and U20455 (N_20455,N_19284,N_19302);
nand U20456 (N_20456,N_19148,N_19210);
or U20457 (N_20457,N_19514,N_19159);
or U20458 (N_20458,N_19787,N_19036);
and U20459 (N_20459,N_19261,N_19736);
and U20460 (N_20460,N_19188,N_19070);
xnor U20461 (N_20461,N_19785,N_19732);
nand U20462 (N_20462,N_19495,N_19348);
nand U20463 (N_20463,N_19686,N_19851);
nand U20464 (N_20464,N_19926,N_19151);
xnor U20465 (N_20465,N_19229,N_19739);
or U20466 (N_20466,N_19902,N_19250);
nand U20467 (N_20467,N_19560,N_19586);
and U20468 (N_20468,N_19218,N_19687);
and U20469 (N_20469,N_19109,N_19659);
or U20470 (N_20470,N_19454,N_19767);
and U20471 (N_20471,N_19759,N_19477);
xnor U20472 (N_20472,N_19378,N_19588);
xnor U20473 (N_20473,N_19265,N_19691);
xnor U20474 (N_20474,N_19049,N_19426);
nor U20475 (N_20475,N_19954,N_19773);
nor U20476 (N_20476,N_19126,N_19745);
nor U20477 (N_20477,N_19705,N_19867);
nor U20478 (N_20478,N_19919,N_19517);
xnor U20479 (N_20479,N_19300,N_19575);
and U20480 (N_20480,N_19988,N_19069);
nor U20481 (N_20481,N_19690,N_19625);
nor U20482 (N_20482,N_19237,N_19975);
nor U20483 (N_20483,N_19026,N_19769);
nor U20484 (N_20484,N_19859,N_19137);
xor U20485 (N_20485,N_19897,N_19286);
or U20486 (N_20486,N_19385,N_19254);
nand U20487 (N_20487,N_19943,N_19201);
xnor U20488 (N_20488,N_19005,N_19014);
nand U20489 (N_20489,N_19832,N_19846);
xor U20490 (N_20490,N_19522,N_19020);
xnor U20491 (N_20491,N_19533,N_19538);
or U20492 (N_20492,N_19720,N_19971);
or U20493 (N_20493,N_19073,N_19950);
xnor U20494 (N_20494,N_19783,N_19619);
nand U20495 (N_20495,N_19712,N_19726);
or U20496 (N_20496,N_19242,N_19814);
and U20497 (N_20497,N_19331,N_19116);
xor U20498 (N_20498,N_19501,N_19525);
nor U20499 (N_20499,N_19985,N_19133);
xnor U20500 (N_20500,N_19005,N_19241);
nor U20501 (N_20501,N_19801,N_19624);
nand U20502 (N_20502,N_19104,N_19112);
xnor U20503 (N_20503,N_19515,N_19144);
or U20504 (N_20504,N_19202,N_19107);
or U20505 (N_20505,N_19270,N_19474);
or U20506 (N_20506,N_19938,N_19593);
and U20507 (N_20507,N_19464,N_19369);
xnor U20508 (N_20508,N_19025,N_19630);
xor U20509 (N_20509,N_19444,N_19090);
nand U20510 (N_20510,N_19994,N_19821);
or U20511 (N_20511,N_19684,N_19152);
xor U20512 (N_20512,N_19318,N_19477);
or U20513 (N_20513,N_19851,N_19534);
xnor U20514 (N_20514,N_19251,N_19519);
xor U20515 (N_20515,N_19975,N_19179);
nand U20516 (N_20516,N_19302,N_19522);
or U20517 (N_20517,N_19513,N_19064);
nand U20518 (N_20518,N_19279,N_19521);
xor U20519 (N_20519,N_19728,N_19230);
nand U20520 (N_20520,N_19594,N_19428);
and U20521 (N_20521,N_19728,N_19534);
and U20522 (N_20522,N_19156,N_19699);
xnor U20523 (N_20523,N_19687,N_19431);
or U20524 (N_20524,N_19736,N_19815);
nor U20525 (N_20525,N_19425,N_19887);
nand U20526 (N_20526,N_19274,N_19308);
nand U20527 (N_20527,N_19113,N_19520);
nor U20528 (N_20528,N_19499,N_19143);
xnor U20529 (N_20529,N_19757,N_19845);
nor U20530 (N_20530,N_19620,N_19542);
nor U20531 (N_20531,N_19825,N_19151);
xor U20532 (N_20532,N_19929,N_19577);
or U20533 (N_20533,N_19589,N_19116);
nor U20534 (N_20534,N_19077,N_19334);
nor U20535 (N_20535,N_19827,N_19643);
nor U20536 (N_20536,N_19028,N_19634);
nor U20537 (N_20537,N_19549,N_19134);
nor U20538 (N_20538,N_19130,N_19570);
and U20539 (N_20539,N_19246,N_19465);
or U20540 (N_20540,N_19679,N_19477);
xor U20541 (N_20541,N_19902,N_19697);
xnor U20542 (N_20542,N_19379,N_19706);
and U20543 (N_20543,N_19018,N_19893);
or U20544 (N_20544,N_19193,N_19262);
or U20545 (N_20545,N_19971,N_19091);
nand U20546 (N_20546,N_19149,N_19341);
or U20547 (N_20547,N_19720,N_19309);
and U20548 (N_20548,N_19643,N_19885);
xor U20549 (N_20549,N_19229,N_19688);
or U20550 (N_20550,N_19964,N_19580);
nor U20551 (N_20551,N_19603,N_19662);
and U20552 (N_20552,N_19738,N_19073);
or U20553 (N_20553,N_19548,N_19755);
nand U20554 (N_20554,N_19205,N_19883);
xor U20555 (N_20555,N_19480,N_19148);
xnor U20556 (N_20556,N_19372,N_19961);
and U20557 (N_20557,N_19264,N_19923);
and U20558 (N_20558,N_19529,N_19098);
or U20559 (N_20559,N_19596,N_19518);
and U20560 (N_20560,N_19230,N_19465);
nand U20561 (N_20561,N_19275,N_19884);
or U20562 (N_20562,N_19593,N_19164);
nor U20563 (N_20563,N_19358,N_19128);
or U20564 (N_20564,N_19920,N_19740);
xor U20565 (N_20565,N_19253,N_19759);
and U20566 (N_20566,N_19541,N_19108);
nand U20567 (N_20567,N_19752,N_19319);
nor U20568 (N_20568,N_19680,N_19620);
nand U20569 (N_20569,N_19715,N_19519);
and U20570 (N_20570,N_19903,N_19596);
xor U20571 (N_20571,N_19473,N_19802);
nand U20572 (N_20572,N_19005,N_19372);
xnor U20573 (N_20573,N_19857,N_19024);
xor U20574 (N_20574,N_19775,N_19956);
xor U20575 (N_20575,N_19344,N_19695);
nor U20576 (N_20576,N_19376,N_19559);
xor U20577 (N_20577,N_19667,N_19716);
and U20578 (N_20578,N_19457,N_19065);
nand U20579 (N_20579,N_19431,N_19157);
xor U20580 (N_20580,N_19546,N_19292);
or U20581 (N_20581,N_19178,N_19025);
xor U20582 (N_20582,N_19374,N_19071);
xor U20583 (N_20583,N_19236,N_19442);
nand U20584 (N_20584,N_19325,N_19863);
xnor U20585 (N_20585,N_19832,N_19330);
and U20586 (N_20586,N_19479,N_19043);
or U20587 (N_20587,N_19906,N_19013);
or U20588 (N_20588,N_19338,N_19741);
or U20589 (N_20589,N_19322,N_19407);
nand U20590 (N_20590,N_19978,N_19412);
xor U20591 (N_20591,N_19771,N_19209);
nor U20592 (N_20592,N_19995,N_19237);
and U20593 (N_20593,N_19591,N_19047);
nand U20594 (N_20594,N_19110,N_19928);
nor U20595 (N_20595,N_19685,N_19532);
xnor U20596 (N_20596,N_19359,N_19646);
nor U20597 (N_20597,N_19817,N_19314);
nand U20598 (N_20598,N_19121,N_19633);
nor U20599 (N_20599,N_19613,N_19868);
nand U20600 (N_20600,N_19582,N_19317);
and U20601 (N_20601,N_19770,N_19322);
xnor U20602 (N_20602,N_19259,N_19227);
or U20603 (N_20603,N_19766,N_19786);
xor U20604 (N_20604,N_19966,N_19177);
nand U20605 (N_20605,N_19568,N_19796);
and U20606 (N_20606,N_19941,N_19659);
or U20607 (N_20607,N_19789,N_19337);
and U20608 (N_20608,N_19942,N_19913);
or U20609 (N_20609,N_19430,N_19443);
nand U20610 (N_20610,N_19276,N_19851);
xnor U20611 (N_20611,N_19916,N_19192);
nor U20612 (N_20612,N_19074,N_19002);
nor U20613 (N_20613,N_19325,N_19505);
nor U20614 (N_20614,N_19886,N_19577);
nand U20615 (N_20615,N_19842,N_19407);
nor U20616 (N_20616,N_19322,N_19766);
nand U20617 (N_20617,N_19506,N_19232);
xor U20618 (N_20618,N_19065,N_19942);
and U20619 (N_20619,N_19151,N_19930);
or U20620 (N_20620,N_19410,N_19405);
nand U20621 (N_20621,N_19811,N_19164);
nand U20622 (N_20622,N_19459,N_19900);
xnor U20623 (N_20623,N_19285,N_19463);
and U20624 (N_20624,N_19817,N_19171);
xor U20625 (N_20625,N_19909,N_19207);
nor U20626 (N_20626,N_19243,N_19221);
xor U20627 (N_20627,N_19740,N_19463);
or U20628 (N_20628,N_19856,N_19834);
nand U20629 (N_20629,N_19965,N_19316);
nor U20630 (N_20630,N_19044,N_19399);
and U20631 (N_20631,N_19805,N_19210);
and U20632 (N_20632,N_19339,N_19992);
xnor U20633 (N_20633,N_19811,N_19010);
nand U20634 (N_20634,N_19291,N_19114);
xor U20635 (N_20635,N_19817,N_19450);
nand U20636 (N_20636,N_19587,N_19316);
and U20637 (N_20637,N_19036,N_19708);
xor U20638 (N_20638,N_19859,N_19634);
xor U20639 (N_20639,N_19779,N_19585);
or U20640 (N_20640,N_19081,N_19682);
and U20641 (N_20641,N_19937,N_19358);
xnor U20642 (N_20642,N_19421,N_19637);
or U20643 (N_20643,N_19496,N_19030);
nand U20644 (N_20644,N_19511,N_19097);
or U20645 (N_20645,N_19893,N_19028);
or U20646 (N_20646,N_19052,N_19365);
or U20647 (N_20647,N_19003,N_19771);
nor U20648 (N_20648,N_19754,N_19889);
or U20649 (N_20649,N_19896,N_19025);
xor U20650 (N_20650,N_19227,N_19030);
nor U20651 (N_20651,N_19363,N_19301);
xnor U20652 (N_20652,N_19506,N_19068);
or U20653 (N_20653,N_19723,N_19571);
nand U20654 (N_20654,N_19154,N_19886);
or U20655 (N_20655,N_19094,N_19469);
and U20656 (N_20656,N_19661,N_19328);
and U20657 (N_20657,N_19061,N_19106);
or U20658 (N_20658,N_19212,N_19420);
xnor U20659 (N_20659,N_19701,N_19814);
xor U20660 (N_20660,N_19573,N_19550);
or U20661 (N_20661,N_19038,N_19322);
or U20662 (N_20662,N_19931,N_19362);
nor U20663 (N_20663,N_19399,N_19914);
and U20664 (N_20664,N_19076,N_19904);
nand U20665 (N_20665,N_19722,N_19224);
xor U20666 (N_20666,N_19753,N_19357);
nand U20667 (N_20667,N_19607,N_19309);
nand U20668 (N_20668,N_19832,N_19335);
nor U20669 (N_20669,N_19629,N_19787);
nor U20670 (N_20670,N_19641,N_19739);
nand U20671 (N_20671,N_19467,N_19870);
and U20672 (N_20672,N_19711,N_19181);
nand U20673 (N_20673,N_19445,N_19496);
nand U20674 (N_20674,N_19771,N_19742);
and U20675 (N_20675,N_19148,N_19734);
nand U20676 (N_20676,N_19723,N_19008);
or U20677 (N_20677,N_19858,N_19677);
or U20678 (N_20678,N_19911,N_19462);
nor U20679 (N_20679,N_19428,N_19492);
or U20680 (N_20680,N_19244,N_19938);
nor U20681 (N_20681,N_19180,N_19786);
nor U20682 (N_20682,N_19684,N_19974);
xnor U20683 (N_20683,N_19205,N_19322);
xor U20684 (N_20684,N_19924,N_19329);
xnor U20685 (N_20685,N_19332,N_19790);
xnor U20686 (N_20686,N_19927,N_19126);
nand U20687 (N_20687,N_19454,N_19943);
xor U20688 (N_20688,N_19734,N_19545);
or U20689 (N_20689,N_19884,N_19971);
and U20690 (N_20690,N_19241,N_19677);
and U20691 (N_20691,N_19061,N_19608);
or U20692 (N_20692,N_19249,N_19043);
nor U20693 (N_20693,N_19463,N_19716);
and U20694 (N_20694,N_19377,N_19987);
xor U20695 (N_20695,N_19135,N_19568);
or U20696 (N_20696,N_19976,N_19886);
and U20697 (N_20697,N_19607,N_19800);
or U20698 (N_20698,N_19373,N_19322);
xnor U20699 (N_20699,N_19309,N_19534);
xor U20700 (N_20700,N_19005,N_19837);
and U20701 (N_20701,N_19499,N_19370);
and U20702 (N_20702,N_19281,N_19149);
xor U20703 (N_20703,N_19182,N_19121);
or U20704 (N_20704,N_19213,N_19833);
or U20705 (N_20705,N_19328,N_19992);
and U20706 (N_20706,N_19901,N_19730);
or U20707 (N_20707,N_19913,N_19728);
nor U20708 (N_20708,N_19438,N_19563);
and U20709 (N_20709,N_19858,N_19154);
nor U20710 (N_20710,N_19438,N_19562);
nor U20711 (N_20711,N_19443,N_19615);
nor U20712 (N_20712,N_19778,N_19216);
or U20713 (N_20713,N_19862,N_19477);
or U20714 (N_20714,N_19934,N_19917);
nand U20715 (N_20715,N_19640,N_19909);
and U20716 (N_20716,N_19129,N_19533);
and U20717 (N_20717,N_19385,N_19046);
nor U20718 (N_20718,N_19963,N_19813);
xor U20719 (N_20719,N_19259,N_19057);
and U20720 (N_20720,N_19720,N_19700);
and U20721 (N_20721,N_19179,N_19665);
xnor U20722 (N_20722,N_19336,N_19955);
nor U20723 (N_20723,N_19198,N_19104);
and U20724 (N_20724,N_19496,N_19256);
nand U20725 (N_20725,N_19485,N_19792);
xor U20726 (N_20726,N_19879,N_19248);
xor U20727 (N_20727,N_19599,N_19094);
nor U20728 (N_20728,N_19880,N_19568);
and U20729 (N_20729,N_19641,N_19753);
nand U20730 (N_20730,N_19634,N_19147);
and U20731 (N_20731,N_19456,N_19011);
and U20732 (N_20732,N_19358,N_19625);
xnor U20733 (N_20733,N_19986,N_19027);
and U20734 (N_20734,N_19933,N_19314);
xnor U20735 (N_20735,N_19300,N_19005);
or U20736 (N_20736,N_19001,N_19554);
nand U20737 (N_20737,N_19086,N_19248);
and U20738 (N_20738,N_19574,N_19456);
nor U20739 (N_20739,N_19482,N_19962);
or U20740 (N_20740,N_19160,N_19220);
and U20741 (N_20741,N_19948,N_19816);
or U20742 (N_20742,N_19647,N_19589);
nand U20743 (N_20743,N_19521,N_19544);
nand U20744 (N_20744,N_19614,N_19621);
nor U20745 (N_20745,N_19646,N_19594);
or U20746 (N_20746,N_19856,N_19476);
or U20747 (N_20747,N_19698,N_19364);
or U20748 (N_20748,N_19317,N_19305);
xor U20749 (N_20749,N_19476,N_19905);
or U20750 (N_20750,N_19206,N_19716);
nor U20751 (N_20751,N_19912,N_19441);
or U20752 (N_20752,N_19132,N_19758);
nor U20753 (N_20753,N_19327,N_19510);
and U20754 (N_20754,N_19828,N_19341);
or U20755 (N_20755,N_19941,N_19427);
or U20756 (N_20756,N_19533,N_19006);
nand U20757 (N_20757,N_19486,N_19322);
nor U20758 (N_20758,N_19415,N_19309);
nand U20759 (N_20759,N_19052,N_19371);
nor U20760 (N_20760,N_19605,N_19542);
xnor U20761 (N_20761,N_19755,N_19950);
xor U20762 (N_20762,N_19096,N_19101);
nand U20763 (N_20763,N_19112,N_19317);
or U20764 (N_20764,N_19085,N_19349);
and U20765 (N_20765,N_19128,N_19498);
nand U20766 (N_20766,N_19690,N_19181);
nor U20767 (N_20767,N_19933,N_19908);
xor U20768 (N_20768,N_19594,N_19941);
nand U20769 (N_20769,N_19363,N_19550);
xor U20770 (N_20770,N_19516,N_19367);
xor U20771 (N_20771,N_19870,N_19734);
or U20772 (N_20772,N_19759,N_19594);
and U20773 (N_20773,N_19098,N_19031);
nor U20774 (N_20774,N_19139,N_19587);
nand U20775 (N_20775,N_19370,N_19139);
and U20776 (N_20776,N_19480,N_19802);
nand U20777 (N_20777,N_19332,N_19181);
nor U20778 (N_20778,N_19481,N_19204);
nand U20779 (N_20779,N_19343,N_19256);
xnor U20780 (N_20780,N_19000,N_19049);
nor U20781 (N_20781,N_19872,N_19917);
xnor U20782 (N_20782,N_19158,N_19049);
nor U20783 (N_20783,N_19084,N_19432);
and U20784 (N_20784,N_19877,N_19064);
or U20785 (N_20785,N_19258,N_19025);
and U20786 (N_20786,N_19386,N_19789);
or U20787 (N_20787,N_19466,N_19344);
or U20788 (N_20788,N_19677,N_19896);
xnor U20789 (N_20789,N_19158,N_19869);
nor U20790 (N_20790,N_19230,N_19666);
xnor U20791 (N_20791,N_19747,N_19873);
xor U20792 (N_20792,N_19350,N_19771);
nor U20793 (N_20793,N_19853,N_19409);
xnor U20794 (N_20794,N_19823,N_19674);
nand U20795 (N_20795,N_19761,N_19934);
nor U20796 (N_20796,N_19059,N_19667);
xor U20797 (N_20797,N_19510,N_19300);
nand U20798 (N_20798,N_19451,N_19467);
xnor U20799 (N_20799,N_19830,N_19447);
nor U20800 (N_20800,N_19053,N_19096);
xor U20801 (N_20801,N_19036,N_19032);
or U20802 (N_20802,N_19058,N_19196);
or U20803 (N_20803,N_19152,N_19776);
nand U20804 (N_20804,N_19420,N_19556);
and U20805 (N_20805,N_19714,N_19166);
or U20806 (N_20806,N_19763,N_19106);
and U20807 (N_20807,N_19884,N_19309);
xnor U20808 (N_20808,N_19203,N_19241);
and U20809 (N_20809,N_19047,N_19119);
nand U20810 (N_20810,N_19021,N_19463);
xnor U20811 (N_20811,N_19842,N_19875);
xnor U20812 (N_20812,N_19147,N_19209);
or U20813 (N_20813,N_19710,N_19350);
and U20814 (N_20814,N_19840,N_19009);
or U20815 (N_20815,N_19776,N_19470);
nor U20816 (N_20816,N_19579,N_19402);
nand U20817 (N_20817,N_19171,N_19469);
nor U20818 (N_20818,N_19945,N_19450);
nand U20819 (N_20819,N_19184,N_19913);
and U20820 (N_20820,N_19302,N_19362);
and U20821 (N_20821,N_19593,N_19147);
xnor U20822 (N_20822,N_19766,N_19959);
and U20823 (N_20823,N_19707,N_19437);
or U20824 (N_20824,N_19455,N_19270);
xnor U20825 (N_20825,N_19079,N_19238);
nand U20826 (N_20826,N_19145,N_19965);
and U20827 (N_20827,N_19187,N_19903);
nor U20828 (N_20828,N_19055,N_19484);
xor U20829 (N_20829,N_19275,N_19786);
nand U20830 (N_20830,N_19534,N_19469);
and U20831 (N_20831,N_19028,N_19872);
xor U20832 (N_20832,N_19862,N_19237);
nand U20833 (N_20833,N_19940,N_19851);
or U20834 (N_20834,N_19762,N_19907);
nor U20835 (N_20835,N_19729,N_19663);
nor U20836 (N_20836,N_19420,N_19579);
and U20837 (N_20837,N_19244,N_19254);
nand U20838 (N_20838,N_19548,N_19734);
or U20839 (N_20839,N_19395,N_19752);
or U20840 (N_20840,N_19018,N_19017);
or U20841 (N_20841,N_19734,N_19449);
xor U20842 (N_20842,N_19331,N_19218);
and U20843 (N_20843,N_19391,N_19611);
and U20844 (N_20844,N_19675,N_19302);
and U20845 (N_20845,N_19781,N_19835);
xor U20846 (N_20846,N_19623,N_19325);
or U20847 (N_20847,N_19605,N_19116);
and U20848 (N_20848,N_19693,N_19179);
nor U20849 (N_20849,N_19838,N_19988);
xor U20850 (N_20850,N_19745,N_19904);
xnor U20851 (N_20851,N_19410,N_19414);
nor U20852 (N_20852,N_19383,N_19110);
xnor U20853 (N_20853,N_19904,N_19332);
nand U20854 (N_20854,N_19749,N_19453);
and U20855 (N_20855,N_19919,N_19977);
nand U20856 (N_20856,N_19215,N_19244);
or U20857 (N_20857,N_19131,N_19495);
xnor U20858 (N_20858,N_19681,N_19590);
xnor U20859 (N_20859,N_19144,N_19058);
nor U20860 (N_20860,N_19450,N_19558);
nand U20861 (N_20861,N_19785,N_19999);
xnor U20862 (N_20862,N_19773,N_19787);
nor U20863 (N_20863,N_19989,N_19631);
and U20864 (N_20864,N_19708,N_19246);
nor U20865 (N_20865,N_19137,N_19778);
nor U20866 (N_20866,N_19333,N_19398);
nand U20867 (N_20867,N_19045,N_19777);
nor U20868 (N_20868,N_19360,N_19785);
or U20869 (N_20869,N_19169,N_19591);
and U20870 (N_20870,N_19578,N_19023);
nand U20871 (N_20871,N_19684,N_19864);
nand U20872 (N_20872,N_19400,N_19909);
or U20873 (N_20873,N_19838,N_19972);
or U20874 (N_20874,N_19390,N_19031);
or U20875 (N_20875,N_19166,N_19959);
nor U20876 (N_20876,N_19898,N_19930);
xor U20877 (N_20877,N_19534,N_19423);
and U20878 (N_20878,N_19177,N_19835);
and U20879 (N_20879,N_19826,N_19233);
nor U20880 (N_20880,N_19168,N_19197);
and U20881 (N_20881,N_19979,N_19059);
nand U20882 (N_20882,N_19079,N_19734);
nand U20883 (N_20883,N_19415,N_19793);
nor U20884 (N_20884,N_19452,N_19112);
nand U20885 (N_20885,N_19834,N_19521);
nand U20886 (N_20886,N_19588,N_19956);
and U20887 (N_20887,N_19529,N_19080);
nor U20888 (N_20888,N_19060,N_19699);
or U20889 (N_20889,N_19344,N_19540);
nor U20890 (N_20890,N_19964,N_19920);
nand U20891 (N_20891,N_19286,N_19133);
and U20892 (N_20892,N_19678,N_19046);
nand U20893 (N_20893,N_19027,N_19532);
and U20894 (N_20894,N_19753,N_19311);
and U20895 (N_20895,N_19211,N_19227);
nand U20896 (N_20896,N_19622,N_19672);
nand U20897 (N_20897,N_19030,N_19282);
nor U20898 (N_20898,N_19223,N_19231);
nor U20899 (N_20899,N_19524,N_19783);
nor U20900 (N_20900,N_19437,N_19963);
or U20901 (N_20901,N_19541,N_19720);
nand U20902 (N_20902,N_19403,N_19799);
and U20903 (N_20903,N_19951,N_19172);
or U20904 (N_20904,N_19052,N_19249);
and U20905 (N_20905,N_19103,N_19992);
nand U20906 (N_20906,N_19227,N_19558);
nand U20907 (N_20907,N_19481,N_19868);
and U20908 (N_20908,N_19127,N_19244);
nand U20909 (N_20909,N_19546,N_19940);
or U20910 (N_20910,N_19475,N_19298);
nand U20911 (N_20911,N_19628,N_19504);
and U20912 (N_20912,N_19831,N_19702);
and U20913 (N_20913,N_19864,N_19825);
xor U20914 (N_20914,N_19340,N_19488);
nand U20915 (N_20915,N_19815,N_19616);
xor U20916 (N_20916,N_19722,N_19272);
and U20917 (N_20917,N_19585,N_19132);
xnor U20918 (N_20918,N_19356,N_19361);
or U20919 (N_20919,N_19710,N_19545);
nor U20920 (N_20920,N_19481,N_19726);
nor U20921 (N_20921,N_19834,N_19401);
and U20922 (N_20922,N_19733,N_19062);
nand U20923 (N_20923,N_19642,N_19555);
nand U20924 (N_20924,N_19723,N_19060);
or U20925 (N_20925,N_19250,N_19834);
nand U20926 (N_20926,N_19835,N_19874);
nand U20927 (N_20927,N_19524,N_19188);
nor U20928 (N_20928,N_19410,N_19112);
nor U20929 (N_20929,N_19475,N_19057);
xnor U20930 (N_20930,N_19261,N_19595);
xnor U20931 (N_20931,N_19204,N_19759);
nand U20932 (N_20932,N_19288,N_19094);
and U20933 (N_20933,N_19181,N_19912);
nand U20934 (N_20934,N_19821,N_19161);
nor U20935 (N_20935,N_19110,N_19975);
or U20936 (N_20936,N_19168,N_19755);
nor U20937 (N_20937,N_19120,N_19558);
nor U20938 (N_20938,N_19237,N_19745);
or U20939 (N_20939,N_19688,N_19375);
and U20940 (N_20940,N_19855,N_19701);
xor U20941 (N_20941,N_19700,N_19529);
nand U20942 (N_20942,N_19811,N_19582);
nand U20943 (N_20943,N_19841,N_19294);
xnor U20944 (N_20944,N_19126,N_19598);
nand U20945 (N_20945,N_19270,N_19742);
nand U20946 (N_20946,N_19332,N_19029);
nand U20947 (N_20947,N_19221,N_19163);
nor U20948 (N_20948,N_19917,N_19669);
or U20949 (N_20949,N_19084,N_19458);
nand U20950 (N_20950,N_19666,N_19841);
xor U20951 (N_20951,N_19307,N_19071);
or U20952 (N_20952,N_19496,N_19958);
or U20953 (N_20953,N_19552,N_19720);
xnor U20954 (N_20954,N_19088,N_19430);
nand U20955 (N_20955,N_19430,N_19804);
nor U20956 (N_20956,N_19105,N_19403);
and U20957 (N_20957,N_19967,N_19087);
or U20958 (N_20958,N_19554,N_19419);
nor U20959 (N_20959,N_19940,N_19518);
xor U20960 (N_20960,N_19414,N_19757);
and U20961 (N_20961,N_19342,N_19226);
nand U20962 (N_20962,N_19880,N_19033);
xor U20963 (N_20963,N_19544,N_19634);
or U20964 (N_20964,N_19347,N_19516);
nand U20965 (N_20965,N_19316,N_19624);
or U20966 (N_20966,N_19698,N_19651);
nor U20967 (N_20967,N_19409,N_19810);
or U20968 (N_20968,N_19860,N_19563);
nand U20969 (N_20969,N_19152,N_19359);
xnor U20970 (N_20970,N_19865,N_19814);
xor U20971 (N_20971,N_19116,N_19487);
nor U20972 (N_20972,N_19503,N_19530);
nand U20973 (N_20973,N_19061,N_19752);
xnor U20974 (N_20974,N_19627,N_19979);
and U20975 (N_20975,N_19776,N_19396);
or U20976 (N_20976,N_19281,N_19311);
nand U20977 (N_20977,N_19927,N_19120);
xor U20978 (N_20978,N_19759,N_19199);
nand U20979 (N_20979,N_19959,N_19194);
xor U20980 (N_20980,N_19149,N_19459);
nor U20981 (N_20981,N_19729,N_19687);
nor U20982 (N_20982,N_19376,N_19597);
xnor U20983 (N_20983,N_19871,N_19880);
nor U20984 (N_20984,N_19212,N_19506);
and U20985 (N_20985,N_19283,N_19252);
nor U20986 (N_20986,N_19566,N_19907);
nor U20987 (N_20987,N_19455,N_19346);
xnor U20988 (N_20988,N_19177,N_19697);
nor U20989 (N_20989,N_19063,N_19949);
or U20990 (N_20990,N_19674,N_19240);
and U20991 (N_20991,N_19178,N_19796);
nand U20992 (N_20992,N_19136,N_19950);
nor U20993 (N_20993,N_19801,N_19380);
nand U20994 (N_20994,N_19576,N_19328);
or U20995 (N_20995,N_19877,N_19493);
and U20996 (N_20996,N_19324,N_19724);
and U20997 (N_20997,N_19638,N_19682);
and U20998 (N_20998,N_19241,N_19565);
or U20999 (N_20999,N_19416,N_19270);
and U21000 (N_21000,N_20003,N_20181);
nor U21001 (N_21001,N_20916,N_20002);
nor U21002 (N_21002,N_20231,N_20566);
nor U21003 (N_21003,N_20506,N_20540);
and U21004 (N_21004,N_20921,N_20194);
nor U21005 (N_21005,N_20375,N_20446);
or U21006 (N_21006,N_20534,N_20632);
xor U21007 (N_21007,N_20355,N_20979);
nor U21008 (N_21008,N_20106,N_20018);
nand U21009 (N_21009,N_20270,N_20338);
nand U21010 (N_21010,N_20521,N_20730);
nand U21011 (N_21011,N_20093,N_20639);
and U21012 (N_21012,N_20392,N_20843);
and U21013 (N_21013,N_20783,N_20411);
and U21014 (N_21014,N_20192,N_20102);
nand U21015 (N_21015,N_20604,N_20831);
nand U21016 (N_21016,N_20076,N_20140);
or U21017 (N_21017,N_20627,N_20918);
nor U21018 (N_21018,N_20956,N_20704);
or U21019 (N_21019,N_20924,N_20735);
and U21020 (N_21020,N_20939,N_20793);
xnor U21021 (N_21021,N_20335,N_20594);
and U21022 (N_21022,N_20298,N_20527);
xor U21023 (N_21023,N_20232,N_20949);
xor U21024 (N_21024,N_20719,N_20145);
xor U21025 (N_21025,N_20354,N_20650);
or U21026 (N_21026,N_20491,N_20655);
nand U21027 (N_21027,N_20235,N_20529);
nand U21028 (N_21028,N_20709,N_20789);
or U21029 (N_21029,N_20350,N_20778);
xor U21030 (N_21030,N_20153,N_20611);
nor U21031 (N_21031,N_20362,N_20132);
nor U21032 (N_21032,N_20160,N_20409);
nand U21033 (N_21033,N_20754,N_20171);
nor U21034 (N_21034,N_20058,N_20260);
xnor U21035 (N_21035,N_20955,N_20081);
and U21036 (N_21036,N_20937,N_20009);
nor U21037 (N_21037,N_20040,N_20244);
xnor U21038 (N_21038,N_20134,N_20114);
xnor U21039 (N_21039,N_20867,N_20385);
and U21040 (N_21040,N_20887,N_20438);
nor U21041 (N_21041,N_20431,N_20300);
or U21042 (N_21042,N_20433,N_20609);
nand U21043 (N_21043,N_20900,N_20041);
nor U21044 (N_21044,N_20673,N_20035);
nand U21045 (N_21045,N_20615,N_20349);
nor U21046 (N_21046,N_20546,N_20064);
nand U21047 (N_21047,N_20762,N_20656);
or U21048 (N_21048,N_20928,N_20873);
xnor U21049 (N_21049,N_20512,N_20562);
and U21050 (N_21050,N_20602,N_20698);
xnor U21051 (N_21051,N_20327,N_20542);
or U21052 (N_21052,N_20090,N_20832);
or U21053 (N_21053,N_20700,N_20261);
xor U21054 (N_21054,N_20773,N_20163);
or U21055 (N_21055,N_20675,N_20812);
or U21056 (N_21056,N_20858,N_20583);
xor U21057 (N_21057,N_20552,N_20470);
nand U21058 (N_21058,N_20020,N_20946);
nor U21059 (N_21059,N_20427,N_20440);
nor U21060 (N_21060,N_20404,N_20531);
or U21061 (N_21061,N_20179,N_20945);
or U21062 (N_21062,N_20087,N_20299);
nand U21063 (N_21063,N_20740,N_20084);
nor U21064 (N_21064,N_20971,N_20502);
nand U21065 (N_21065,N_20088,N_20214);
nor U21066 (N_21066,N_20897,N_20714);
nand U21067 (N_21067,N_20726,N_20795);
or U21068 (N_21068,N_20722,N_20173);
nand U21069 (N_21069,N_20280,N_20576);
nor U21070 (N_21070,N_20339,N_20008);
xnor U21071 (N_21071,N_20857,N_20712);
xor U21072 (N_21072,N_20646,N_20922);
and U21073 (N_21073,N_20803,N_20976);
nand U21074 (N_21074,N_20634,N_20985);
xnor U21075 (N_21075,N_20480,N_20652);
xor U21076 (N_21076,N_20975,N_20495);
or U21077 (N_21077,N_20026,N_20535);
and U21078 (N_21078,N_20190,N_20062);
xor U21079 (N_21079,N_20006,N_20797);
or U21080 (N_21080,N_20341,N_20238);
xor U21081 (N_21081,N_20129,N_20990);
nor U21082 (N_21082,N_20154,N_20899);
or U21083 (N_21083,N_20935,N_20051);
nand U21084 (N_21084,N_20259,N_20254);
xnor U21085 (N_21085,N_20266,N_20516);
or U21086 (N_21086,N_20091,N_20824);
and U21087 (N_21087,N_20201,N_20929);
xor U21088 (N_21088,N_20894,N_20966);
nor U21089 (N_21089,N_20965,N_20485);
xnor U21090 (N_21090,N_20997,N_20960);
nand U21091 (N_21091,N_20291,N_20188);
xor U21092 (N_21092,N_20989,N_20444);
nor U21093 (N_21093,N_20379,N_20290);
xnor U21094 (N_21094,N_20558,N_20042);
xor U21095 (N_21095,N_20511,N_20528);
nand U21096 (N_21096,N_20208,N_20834);
and U21097 (N_21097,N_20586,N_20904);
and U21098 (N_21098,N_20660,N_20988);
or U21099 (N_21099,N_20473,N_20033);
nand U21100 (N_21100,N_20418,N_20877);
nor U21101 (N_21101,N_20050,N_20209);
nor U21102 (N_21102,N_20367,N_20403);
nand U21103 (N_21103,N_20767,N_20168);
and U21104 (N_21104,N_20070,N_20371);
xor U21105 (N_21105,N_20285,N_20248);
xor U21106 (N_21106,N_20243,N_20310);
nand U21107 (N_21107,N_20913,N_20175);
and U21108 (N_21108,N_20345,N_20829);
nor U21109 (N_21109,N_20806,N_20461);
or U21110 (N_21110,N_20063,N_20449);
and U21111 (N_21111,N_20022,N_20061);
nor U21112 (N_21112,N_20896,N_20802);
nor U21113 (N_21113,N_20690,N_20768);
nor U21114 (N_21114,N_20775,N_20401);
or U21115 (N_21115,N_20980,N_20746);
and U21116 (N_21116,N_20218,N_20662);
and U21117 (N_21117,N_20610,N_20142);
or U21118 (N_21118,N_20424,N_20848);
nor U21119 (N_21119,N_20165,N_20827);
nor U21120 (N_21120,N_20413,N_20805);
and U21121 (N_21121,N_20447,N_20329);
or U21122 (N_21122,N_20891,N_20342);
or U21123 (N_21123,N_20278,N_20624);
or U21124 (N_21124,N_20237,N_20787);
nor U21125 (N_21125,N_20407,N_20784);
or U21126 (N_21126,N_20895,N_20907);
nand U21127 (N_21127,N_20023,N_20489);
nand U21128 (N_21128,N_20148,N_20236);
and U21129 (N_21129,N_20794,N_20240);
nand U21130 (N_21130,N_20464,N_20751);
xnor U21131 (N_21131,N_20230,N_20914);
nand U21132 (N_21132,N_20286,N_20068);
nand U21133 (N_21133,N_20498,N_20603);
and U21134 (N_21134,N_20573,N_20412);
and U21135 (N_21135,N_20421,N_20679);
nor U21136 (N_21136,N_20265,N_20308);
nor U21137 (N_21137,N_20920,N_20780);
xor U21138 (N_21138,N_20717,N_20469);
or U21139 (N_21139,N_20347,N_20178);
nor U21140 (N_21140,N_20809,N_20580);
and U21141 (N_21141,N_20962,N_20810);
nand U21142 (N_21142,N_20756,N_20000);
or U21143 (N_21143,N_20383,N_20432);
nor U21144 (N_21144,N_20120,N_20317);
xor U21145 (N_21145,N_20059,N_20721);
and U21146 (N_21146,N_20112,N_20731);
nor U21147 (N_21147,N_20410,N_20086);
nand U21148 (N_21148,N_20482,N_20439);
xor U21149 (N_21149,N_20055,N_20024);
nor U21150 (N_21150,N_20850,N_20222);
and U21151 (N_21151,N_20476,N_20644);
or U21152 (N_21152,N_20923,N_20680);
xnor U21153 (N_21153,N_20986,N_20964);
xnor U21154 (N_21154,N_20799,N_20189);
and U21155 (N_21155,N_20716,N_20518);
nor U21156 (N_21156,N_20402,N_20683);
or U21157 (N_21157,N_20830,N_20500);
and U21158 (N_21158,N_20283,N_20205);
nand U21159 (N_21159,N_20884,N_20919);
or U21160 (N_21160,N_20835,N_20526);
or U21161 (N_21161,N_20107,N_20908);
nand U21162 (N_21162,N_20664,N_20199);
nor U21163 (N_21163,N_20845,N_20045);
and U21164 (N_21164,N_20944,N_20926);
xnor U21165 (N_21165,N_20092,N_20519);
xor U21166 (N_21166,N_20365,N_20161);
xnor U21167 (N_21167,N_20147,N_20085);
or U21168 (N_21168,N_20555,N_20893);
nand U21169 (N_21169,N_20422,N_20868);
xor U21170 (N_21170,N_20718,N_20774);
or U21171 (N_21171,N_20781,N_20808);
xor U21172 (N_21172,N_20525,N_20110);
xnor U21173 (N_21173,N_20950,N_20465);
or U21174 (N_21174,N_20031,N_20246);
nor U21175 (N_21175,N_20130,N_20111);
and U21176 (N_21176,N_20351,N_20561);
xnor U21177 (N_21177,N_20176,N_20069);
and U21178 (N_21178,N_20874,N_20156);
nand U21179 (N_21179,N_20635,N_20359);
nor U21180 (N_21180,N_20942,N_20072);
nor U21181 (N_21181,N_20927,N_20399);
nand U21182 (N_21182,N_20826,N_20471);
nor U21183 (N_21183,N_20725,N_20816);
xnor U21184 (N_21184,N_20263,N_20890);
or U21185 (N_21185,N_20538,N_20947);
xor U21186 (N_21186,N_20258,N_20198);
and U21187 (N_21187,N_20289,N_20478);
or U21188 (N_21188,N_20141,N_20763);
or U21189 (N_21189,N_20881,N_20934);
or U21190 (N_21190,N_20079,N_20104);
xor U21191 (N_21191,N_20906,N_20545);
or U21192 (N_21192,N_20334,N_20861);
xor U21193 (N_21193,N_20551,N_20581);
or U21194 (N_21194,N_20849,N_20978);
and U21195 (N_21195,N_20115,N_20689);
or U21196 (N_21196,N_20479,N_20224);
nor U21197 (N_21197,N_20249,N_20220);
xnor U21198 (N_21198,N_20099,N_20264);
nand U21199 (N_21199,N_20430,N_20544);
nand U21200 (N_21200,N_20771,N_20174);
and U21201 (N_21201,N_20328,N_20853);
nor U21202 (N_21202,N_20435,N_20067);
and U21203 (N_21203,N_20815,N_20217);
or U21204 (N_21204,N_20322,N_20177);
nand U21205 (N_21205,N_20697,N_20702);
or U21206 (N_21206,N_20127,N_20015);
nand U21207 (N_21207,N_20150,N_20777);
and U21208 (N_21208,N_20252,N_20865);
xor U21209 (N_21209,N_20684,N_20653);
and U21210 (N_21210,N_20333,N_20614);
nor U21211 (N_21211,N_20358,N_20172);
nor U21212 (N_21212,N_20382,N_20004);
nor U21213 (N_21213,N_20723,N_20631);
xnor U21214 (N_21214,N_20094,N_20554);
nand U21215 (N_21215,N_20164,N_20348);
nand U21216 (N_21216,N_20553,N_20284);
xor U21217 (N_21217,N_20364,N_20032);
xor U21218 (N_21218,N_20738,N_20724);
nand U21219 (N_21219,N_20036,N_20822);
nand U21220 (N_21220,N_20936,N_20429);
or U21221 (N_21221,N_20082,N_20494);
and U21222 (N_21222,N_20216,N_20454);
or U21223 (N_21223,N_20619,N_20820);
xor U21224 (N_21224,N_20661,N_20159);
and U21225 (N_21225,N_20851,N_20901);
nand U21226 (N_21226,N_20488,N_20309);
nor U21227 (N_21227,N_20103,N_20612);
xnor U21228 (N_21228,N_20687,N_20608);
nor U21229 (N_21229,N_20708,N_20170);
xnor U21230 (N_21230,N_20257,N_20239);
or U21231 (N_21231,N_20373,N_20116);
nor U21232 (N_21232,N_20620,N_20269);
xor U21233 (N_21233,N_20800,N_20769);
nand U21234 (N_21234,N_20872,N_20909);
or U21235 (N_21235,N_20749,N_20353);
and U21236 (N_21236,N_20049,N_20211);
nand U21237 (N_21237,N_20999,N_20745);
xnor U21238 (N_21238,N_20665,N_20597);
or U21239 (N_21239,N_20968,N_20886);
nand U21240 (N_21240,N_20242,N_20294);
or U21241 (N_21241,N_20753,N_20352);
xnor U21242 (N_21242,N_20271,N_20303);
nor U21243 (N_21243,N_20954,N_20892);
or U21244 (N_21244,N_20911,N_20323);
nor U21245 (N_21245,N_20374,N_20011);
nor U21246 (N_21246,N_20682,N_20396);
nor U21247 (N_21247,N_20360,N_20203);
and U21248 (N_21248,N_20596,N_20706);
and U21249 (N_21249,N_20649,N_20443);
nand U21250 (N_21250,N_20757,N_20591);
xnor U21251 (N_21251,N_20996,N_20453);
and U21252 (N_21252,N_20138,N_20223);
xnor U21253 (N_21253,N_20250,N_20982);
nand U21254 (N_21254,N_20549,N_20131);
and U21255 (N_21255,N_20195,N_20507);
xor U21256 (N_21256,N_20293,N_20616);
and U21257 (N_21257,N_20860,N_20251);
nand U21258 (N_21258,N_20654,N_20785);
xnor U21259 (N_21259,N_20994,N_20095);
nand U21260 (N_21260,N_20158,N_20128);
nand U21261 (N_21261,N_20869,N_20575);
nor U21262 (N_21262,N_20623,N_20486);
and U21263 (N_21263,N_20144,N_20149);
or U21264 (N_21264,N_20277,N_20493);
nand U21265 (N_21265,N_20933,N_20543);
xor U21266 (N_21266,N_20387,N_20492);
and U21267 (N_21267,N_20613,N_20560);
and U21268 (N_21268,N_20038,N_20701);
xnor U21269 (N_21269,N_20882,N_20958);
xor U21270 (N_21270,N_20559,N_20425);
xnor U21271 (N_21271,N_20474,N_20207);
nor U21272 (N_21272,N_20484,N_20436);
and U21273 (N_21273,N_20792,N_20974);
or U21274 (N_21274,N_20537,N_20692);
or U21275 (N_21275,N_20577,N_20628);
and U21276 (N_21276,N_20056,N_20786);
nor U21277 (N_21277,N_20136,N_20047);
and U21278 (N_21278,N_20733,N_20426);
nor U21279 (N_21279,N_20197,N_20027);
and U21280 (N_21280,N_20262,N_20605);
xor U21281 (N_21281,N_20987,N_20637);
nor U21282 (N_21282,N_20667,N_20821);
and U21283 (N_21283,N_20073,N_20010);
or U21284 (N_21284,N_20316,N_20758);
and U21285 (N_21285,N_20618,N_20275);
nor U21286 (N_21286,N_20556,N_20636);
or U21287 (N_21287,N_20766,N_20255);
nand U21288 (N_21288,N_20193,N_20184);
xnor U21289 (N_21289,N_20118,N_20200);
and U21290 (N_21290,N_20951,N_20005);
nor U21291 (N_21291,N_20645,N_20080);
xnor U21292 (N_21292,N_20096,N_20245);
nand U21293 (N_21293,N_20037,N_20879);
and U21294 (N_21294,N_20539,N_20747);
xor U21295 (N_21295,N_20940,N_20057);
or U21296 (N_21296,N_20311,N_20991);
nor U21297 (N_21297,N_20221,N_20670);
xnor U21298 (N_21298,N_20267,N_20814);
xnor U21299 (N_21299,N_20463,N_20048);
and U21300 (N_21300,N_20434,N_20450);
and U21301 (N_21301,N_20441,N_20569);
and U21302 (N_21302,N_20513,N_20836);
nor U21303 (N_21303,N_20428,N_20321);
nand U21304 (N_21304,N_20305,N_20743);
nand U21305 (N_21305,N_20370,N_20419);
xnor U21306 (N_21306,N_20187,N_20589);
nor U21307 (N_21307,N_20917,N_20448);
or U21308 (N_21308,N_20640,N_20871);
or U21309 (N_21309,N_20191,N_20993);
nand U21310 (N_21310,N_20182,N_20397);
nand U21311 (N_21311,N_20852,N_20859);
and U21312 (N_21312,N_20109,N_20567);
nand U21313 (N_21313,N_20340,N_20876);
and U21314 (N_21314,N_20703,N_20372);
xor U21315 (N_21315,N_20782,N_20414);
nor U21316 (N_21316,N_20014,N_20139);
or U21317 (N_21317,N_20686,N_20776);
nor U21318 (N_21318,N_20811,N_20210);
and U21319 (N_21319,N_20643,N_20101);
xnor U21320 (N_21320,N_20393,N_20889);
or U21321 (N_21321,N_20225,N_20162);
nand U21322 (N_21322,N_20759,N_20273);
xnor U21323 (N_21323,N_20304,N_20196);
and U21324 (N_21324,N_20398,N_20970);
nand U21325 (N_21325,N_20765,N_20588);
or U21326 (N_21326,N_20274,N_20728);
nor U21327 (N_21327,N_20054,N_20016);
and U21328 (N_21328,N_20330,N_20574);
and U21329 (N_21329,N_20705,N_20394);
or U21330 (N_21330,N_20657,N_20952);
and U21331 (N_21331,N_20313,N_20408);
or U21332 (N_21332,N_20253,N_20641);
nor U21333 (N_21333,N_20856,N_20287);
or U21334 (N_21334,N_20089,N_20213);
xor U21335 (N_21335,N_20840,N_20995);
and U21336 (N_21336,N_20638,N_20417);
and U21337 (N_21337,N_20377,N_20226);
nand U21338 (N_21338,N_20622,N_20167);
xor U21339 (N_21339,N_20568,N_20406);
nor U21340 (N_21340,N_20318,N_20490);
nand U21341 (N_21341,N_20959,N_20841);
xor U21342 (N_21342,N_20301,N_20297);
nor U21343 (N_21343,N_20957,N_20572);
and U21344 (N_21344,N_20053,N_20676);
nor U21345 (N_21345,N_20981,N_20368);
xor U21346 (N_21346,N_20903,N_20466);
or U21347 (N_21347,N_20938,N_20369);
xor U21348 (N_21348,N_20750,N_20228);
nor U21349 (N_21349,N_20732,N_20455);
nor U21350 (N_21350,N_20282,N_20699);
or U21351 (N_21351,N_20630,N_20395);
xnor U21352 (N_21352,N_20391,N_20992);
and U21353 (N_21353,N_20888,N_20825);
xnor U21354 (N_21354,N_20312,N_20315);
and U21355 (N_21355,N_20442,N_20564);
or U21356 (N_21356,N_20151,N_20863);
nor U21357 (N_21357,N_20672,N_20319);
nand U21358 (N_21358,N_20752,N_20423);
nand U21359 (N_21359,N_20967,N_20791);
or U21360 (N_21360,N_20742,N_20864);
xor U21361 (N_21361,N_20515,N_20910);
xor U21362 (N_21362,N_20961,N_20666);
or U21363 (N_21363,N_20212,N_20870);
and U21364 (N_21364,N_20017,N_20452);
nand U21365 (N_21365,N_20324,N_20804);
and U21366 (N_21366,N_20314,N_20727);
and U21367 (N_21367,N_20075,N_20878);
and U21368 (N_21368,N_20113,N_20855);
xnor U21369 (N_21369,N_20117,N_20233);
and U21370 (N_21370,N_20875,N_20307);
xnor U21371 (N_21371,N_20256,N_20854);
nand U21372 (N_21372,N_20366,N_20361);
xnor U21373 (N_21373,N_20451,N_20647);
or U21374 (N_21374,N_20696,N_20941);
nor U21375 (N_21375,N_20972,N_20276);
xnor U21376 (N_21376,N_20021,N_20530);
nor U21377 (N_21377,N_20133,N_20691);
xnor U21378 (N_21378,N_20651,N_20629);
and U21379 (N_21379,N_20595,N_20905);
nand U21380 (N_21380,N_20509,N_20288);
xnor U21381 (N_21381,N_20711,N_20124);
xor U21382 (N_21382,N_20838,N_20344);
xnor U21383 (N_21383,N_20817,N_20204);
and U21384 (N_21384,N_20736,N_20592);
xnor U21385 (N_21385,N_20510,N_20607);
and U21386 (N_21386,N_20445,N_20074);
or U21387 (N_21387,N_20169,N_20590);
and U21388 (N_21388,N_20306,N_20533);
or U21389 (N_21389,N_20125,N_20514);
xnor U21390 (N_21390,N_20497,N_20621);
xnor U21391 (N_21391,N_20420,N_20157);
or U21392 (N_21392,N_20098,N_20481);
nor U21393 (N_21393,N_20547,N_20606);
nand U21394 (N_21394,N_20570,N_20504);
nand U21395 (N_21395,N_20866,N_20416);
nand U21396 (N_21396,N_20760,N_20028);
or U21397 (N_21397,N_20346,N_20524);
xor U21398 (N_21398,N_20658,N_20405);
nor U21399 (N_21399,N_20400,N_20818);
nand U21400 (N_21400,N_20185,N_20100);
or U21401 (N_21401,N_20741,N_20052);
and U21402 (N_21402,N_20522,N_20030);
and U21403 (N_21403,N_20467,N_20833);
or U21404 (N_21404,N_20790,N_20681);
and U21405 (N_21405,N_20227,N_20001);
nand U21406 (N_21406,N_20517,N_20617);
xnor U21407 (N_21407,N_20459,N_20823);
xnor U21408 (N_21408,N_20796,N_20565);
and U21409 (N_21409,N_20707,N_20121);
xnor U21410 (N_21410,N_20550,N_20685);
nor U21411 (N_21411,N_20229,N_20272);
xnor U21412 (N_21412,N_20462,N_20122);
nand U21413 (N_21413,N_20215,N_20477);
and U21414 (N_21414,N_20963,N_20029);
and U21415 (N_21415,N_20770,N_20343);
xor U21416 (N_21416,N_20801,N_20234);
nand U21417 (N_21417,N_20837,N_20532);
or U21418 (N_21418,N_20357,N_20505);
or U21419 (N_21419,N_20108,N_20520);
and U21420 (N_21420,N_20336,N_20585);
nand U21421 (N_21421,N_20499,N_20798);
nor U21422 (N_21422,N_20668,N_20071);
nand U21423 (N_21423,N_20807,N_20599);
nand U21424 (N_21424,N_20501,N_20969);
and U21425 (N_21425,N_20186,N_20813);
and U21426 (N_21426,N_20772,N_20693);
or U21427 (N_21427,N_20847,N_20548);
or U21428 (N_21428,N_20748,N_20378);
and U21429 (N_21429,N_20943,N_20626);
and U21430 (N_21430,N_20337,N_20828);
nor U21431 (N_21431,N_20483,N_20296);
nor U21432 (N_21432,N_20677,N_20043);
and U21433 (N_21433,N_20678,N_20376);
xnor U21434 (N_21434,N_20659,N_20268);
and U21435 (N_21435,N_20019,N_20457);
xnor U21436 (N_21436,N_20206,N_20219);
nand U21437 (N_21437,N_20842,N_20713);
nor U21438 (N_21438,N_20044,N_20925);
nand U21439 (N_21439,N_20363,N_20460);
and U21440 (N_21440,N_20885,N_20281);
or U21441 (N_21441,N_20295,N_20119);
or U21442 (N_21442,N_20983,N_20764);
or U21443 (N_21443,N_20761,N_20578);
or U21444 (N_21444,N_20739,N_20146);
nand U21445 (N_21445,N_20143,N_20503);
or U21446 (N_21446,N_20066,N_20931);
and U21447 (N_21447,N_20126,N_20839);
xor U21448 (N_21448,N_20737,N_20912);
nor U21449 (N_21449,N_20013,N_20734);
xnor U21450 (N_21450,N_20648,N_20180);
or U21451 (N_21451,N_20598,N_20105);
and U21452 (N_21452,N_20663,N_20202);
nor U21453 (N_21453,N_20152,N_20953);
and U21454 (N_21454,N_20137,N_20880);
nand U21455 (N_21455,N_20633,N_20984);
nor U21456 (N_21456,N_20292,N_20468);
or U21457 (N_21457,N_20720,N_20034);
and U21458 (N_21458,N_20669,N_20247);
and U21459 (N_21459,N_20846,N_20135);
and U21460 (N_21460,N_20077,N_20472);
nand U21461 (N_21461,N_20915,N_20241);
nand U21462 (N_21462,N_20593,N_20097);
nand U21463 (N_21463,N_20998,N_20541);
and U21464 (N_21464,N_20601,N_20356);
nand U21465 (N_21465,N_20563,N_20039);
and U21466 (N_21466,N_20475,N_20078);
xnor U21467 (N_21467,N_20012,N_20326);
or U21468 (N_21468,N_20536,N_20948);
or U21469 (N_21469,N_20862,N_20744);
and U21470 (N_21470,N_20065,N_20381);
nor U21471 (N_21471,N_20883,N_20932);
xnor U21472 (N_21472,N_20508,N_20844);
nand U21473 (N_21473,N_20977,N_20320);
xor U21474 (N_21474,N_20579,N_20694);
and U21475 (N_21475,N_20437,N_20331);
nand U21476 (N_21476,N_20688,N_20755);
nor U21477 (N_21477,N_20695,N_20487);
xor U21478 (N_21478,N_20390,N_20380);
and U21479 (N_21479,N_20386,N_20183);
xnor U21480 (N_21480,N_20788,N_20930);
nand U21481 (N_21481,N_20729,N_20496);
nor U21482 (N_21482,N_20557,N_20279);
nor U21483 (N_21483,N_20123,N_20674);
or U21484 (N_21484,N_20898,N_20819);
nand U21485 (N_21485,N_20046,N_20025);
xor U21486 (N_21486,N_20325,N_20166);
xor U21487 (N_21487,N_20389,N_20571);
or U21488 (N_21488,N_20388,N_20458);
xnor U21489 (N_21489,N_20582,N_20083);
nand U21490 (N_21490,N_20060,N_20671);
nand U21491 (N_21491,N_20523,N_20456);
and U21492 (N_21492,N_20007,N_20584);
and U21493 (N_21493,N_20973,N_20625);
xnor U21494 (N_21494,N_20715,N_20155);
nand U21495 (N_21495,N_20332,N_20642);
nor U21496 (N_21496,N_20302,N_20902);
xnor U21497 (N_21497,N_20587,N_20779);
nor U21498 (N_21498,N_20415,N_20384);
nor U21499 (N_21499,N_20710,N_20600);
xor U21500 (N_21500,N_20518,N_20438);
xor U21501 (N_21501,N_20688,N_20946);
xnor U21502 (N_21502,N_20455,N_20313);
nand U21503 (N_21503,N_20002,N_20474);
nand U21504 (N_21504,N_20705,N_20049);
nor U21505 (N_21505,N_20939,N_20033);
xor U21506 (N_21506,N_20124,N_20692);
or U21507 (N_21507,N_20345,N_20594);
nor U21508 (N_21508,N_20111,N_20389);
or U21509 (N_21509,N_20322,N_20853);
and U21510 (N_21510,N_20188,N_20154);
nor U21511 (N_21511,N_20739,N_20041);
nand U21512 (N_21512,N_20823,N_20016);
nand U21513 (N_21513,N_20216,N_20868);
and U21514 (N_21514,N_20581,N_20608);
nand U21515 (N_21515,N_20530,N_20867);
nor U21516 (N_21516,N_20174,N_20442);
nor U21517 (N_21517,N_20539,N_20496);
nor U21518 (N_21518,N_20224,N_20306);
or U21519 (N_21519,N_20642,N_20211);
or U21520 (N_21520,N_20828,N_20159);
and U21521 (N_21521,N_20056,N_20826);
or U21522 (N_21522,N_20419,N_20104);
or U21523 (N_21523,N_20111,N_20004);
xnor U21524 (N_21524,N_20931,N_20415);
or U21525 (N_21525,N_20896,N_20916);
nand U21526 (N_21526,N_20844,N_20644);
nor U21527 (N_21527,N_20546,N_20979);
nand U21528 (N_21528,N_20363,N_20958);
and U21529 (N_21529,N_20600,N_20156);
or U21530 (N_21530,N_20523,N_20119);
nand U21531 (N_21531,N_20275,N_20383);
nor U21532 (N_21532,N_20373,N_20104);
nand U21533 (N_21533,N_20799,N_20598);
nand U21534 (N_21534,N_20283,N_20683);
xor U21535 (N_21535,N_20261,N_20206);
nor U21536 (N_21536,N_20452,N_20586);
nand U21537 (N_21537,N_20223,N_20318);
nand U21538 (N_21538,N_20193,N_20811);
or U21539 (N_21539,N_20629,N_20122);
or U21540 (N_21540,N_20819,N_20198);
or U21541 (N_21541,N_20905,N_20830);
nor U21542 (N_21542,N_20460,N_20206);
xnor U21543 (N_21543,N_20895,N_20032);
xnor U21544 (N_21544,N_20410,N_20978);
or U21545 (N_21545,N_20561,N_20118);
and U21546 (N_21546,N_20554,N_20839);
xor U21547 (N_21547,N_20785,N_20953);
xor U21548 (N_21548,N_20054,N_20631);
xor U21549 (N_21549,N_20418,N_20426);
and U21550 (N_21550,N_20060,N_20594);
nand U21551 (N_21551,N_20179,N_20368);
xor U21552 (N_21552,N_20553,N_20660);
and U21553 (N_21553,N_20326,N_20226);
xnor U21554 (N_21554,N_20905,N_20062);
xor U21555 (N_21555,N_20342,N_20350);
or U21556 (N_21556,N_20668,N_20309);
nor U21557 (N_21557,N_20540,N_20154);
and U21558 (N_21558,N_20484,N_20415);
or U21559 (N_21559,N_20588,N_20484);
nand U21560 (N_21560,N_20672,N_20211);
and U21561 (N_21561,N_20104,N_20575);
or U21562 (N_21562,N_20522,N_20474);
nand U21563 (N_21563,N_20818,N_20676);
or U21564 (N_21564,N_20973,N_20049);
and U21565 (N_21565,N_20761,N_20163);
nand U21566 (N_21566,N_20184,N_20907);
or U21567 (N_21567,N_20559,N_20163);
or U21568 (N_21568,N_20568,N_20083);
xor U21569 (N_21569,N_20577,N_20655);
nand U21570 (N_21570,N_20668,N_20161);
nand U21571 (N_21571,N_20631,N_20168);
xor U21572 (N_21572,N_20047,N_20680);
or U21573 (N_21573,N_20781,N_20520);
and U21574 (N_21574,N_20319,N_20501);
or U21575 (N_21575,N_20550,N_20832);
and U21576 (N_21576,N_20575,N_20756);
nor U21577 (N_21577,N_20728,N_20405);
nand U21578 (N_21578,N_20575,N_20498);
nand U21579 (N_21579,N_20896,N_20092);
nand U21580 (N_21580,N_20644,N_20868);
or U21581 (N_21581,N_20971,N_20995);
nand U21582 (N_21582,N_20229,N_20212);
nor U21583 (N_21583,N_20494,N_20665);
or U21584 (N_21584,N_20832,N_20075);
or U21585 (N_21585,N_20338,N_20312);
and U21586 (N_21586,N_20673,N_20158);
or U21587 (N_21587,N_20225,N_20371);
or U21588 (N_21588,N_20089,N_20214);
xnor U21589 (N_21589,N_20321,N_20795);
nand U21590 (N_21590,N_20729,N_20875);
nor U21591 (N_21591,N_20580,N_20604);
or U21592 (N_21592,N_20679,N_20211);
nand U21593 (N_21593,N_20599,N_20555);
nand U21594 (N_21594,N_20557,N_20599);
nor U21595 (N_21595,N_20963,N_20646);
nor U21596 (N_21596,N_20190,N_20523);
or U21597 (N_21597,N_20813,N_20598);
nand U21598 (N_21598,N_20155,N_20006);
xnor U21599 (N_21599,N_20189,N_20622);
or U21600 (N_21600,N_20649,N_20910);
nor U21601 (N_21601,N_20132,N_20955);
xnor U21602 (N_21602,N_20635,N_20074);
nand U21603 (N_21603,N_20347,N_20234);
nor U21604 (N_21604,N_20952,N_20462);
xnor U21605 (N_21605,N_20978,N_20325);
nand U21606 (N_21606,N_20391,N_20621);
nor U21607 (N_21607,N_20770,N_20311);
or U21608 (N_21608,N_20645,N_20786);
xor U21609 (N_21609,N_20317,N_20445);
xnor U21610 (N_21610,N_20190,N_20051);
xnor U21611 (N_21611,N_20849,N_20517);
and U21612 (N_21612,N_20226,N_20459);
xor U21613 (N_21613,N_20303,N_20557);
nor U21614 (N_21614,N_20326,N_20891);
nand U21615 (N_21615,N_20272,N_20445);
or U21616 (N_21616,N_20088,N_20891);
nand U21617 (N_21617,N_20097,N_20681);
or U21618 (N_21618,N_20881,N_20001);
nor U21619 (N_21619,N_20205,N_20890);
nor U21620 (N_21620,N_20590,N_20207);
xor U21621 (N_21621,N_20258,N_20263);
nand U21622 (N_21622,N_20626,N_20829);
and U21623 (N_21623,N_20845,N_20213);
nor U21624 (N_21624,N_20110,N_20487);
xnor U21625 (N_21625,N_20647,N_20995);
and U21626 (N_21626,N_20100,N_20939);
xnor U21627 (N_21627,N_20212,N_20662);
xor U21628 (N_21628,N_20856,N_20496);
nand U21629 (N_21629,N_20162,N_20916);
xor U21630 (N_21630,N_20628,N_20382);
and U21631 (N_21631,N_20053,N_20781);
xnor U21632 (N_21632,N_20409,N_20477);
or U21633 (N_21633,N_20658,N_20894);
nand U21634 (N_21634,N_20285,N_20063);
xor U21635 (N_21635,N_20756,N_20680);
or U21636 (N_21636,N_20726,N_20498);
and U21637 (N_21637,N_20369,N_20420);
nor U21638 (N_21638,N_20109,N_20196);
nor U21639 (N_21639,N_20954,N_20949);
and U21640 (N_21640,N_20852,N_20394);
or U21641 (N_21641,N_20041,N_20754);
nor U21642 (N_21642,N_20232,N_20238);
nor U21643 (N_21643,N_20086,N_20340);
and U21644 (N_21644,N_20233,N_20656);
xnor U21645 (N_21645,N_20149,N_20615);
nand U21646 (N_21646,N_20703,N_20031);
xnor U21647 (N_21647,N_20068,N_20157);
and U21648 (N_21648,N_20686,N_20085);
or U21649 (N_21649,N_20516,N_20023);
and U21650 (N_21650,N_20459,N_20912);
and U21651 (N_21651,N_20638,N_20256);
or U21652 (N_21652,N_20108,N_20731);
or U21653 (N_21653,N_20238,N_20348);
nor U21654 (N_21654,N_20428,N_20860);
nand U21655 (N_21655,N_20543,N_20755);
and U21656 (N_21656,N_20294,N_20034);
xnor U21657 (N_21657,N_20138,N_20889);
or U21658 (N_21658,N_20343,N_20845);
xnor U21659 (N_21659,N_20511,N_20005);
xnor U21660 (N_21660,N_20840,N_20196);
nand U21661 (N_21661,N_20039,N_20304);
or U21662 (N_21662,N_20663,N_20591);
xnor U21663 (N_21663,N_20415,N_20411);
xor U21664 (N_21664,N_20571,N_20243);
nor U21665 (N_21665,N_20336,N_20869);
nor U21666 (N_21666,N_20825,N_20624);
xnor U21667 (N_21667,N_20934,N_20267);
nand U21668 (N_21668,N_20067,N_20809);
nand U21669 (N_21669,N_20044,N_20129);
and U21670 (N_21670,N_20306,N_20860);
nand U21671 (N_21671,N_20395,N_20273);
nor U21672 (N_21672,N_20729,N_20166);
xor U21673 (N_21673,N_20744,N_20312);
or U21674 (N_21674,N_20537,N_20818);
or U21675 (N_21675,N_20345,N_20792);
and U21676 (N_21676,N_20786,N_20964);
xnor U21677 (N_21677,N_20334,N_20342);
or U21678 (N_21678,N_20675,N_20903);
xor U21679 (N_21679,N_20737,N_20533);
nor U21680 (N_21680,N_20079,N_20648);
and U21681 (N_21681,N_20670,N_20493);
nand U21682 (N_21682,N_20152,N_20786);
xnor U21683 (N_21683,N_20843,N_20533);
xnor U21684 (N_21684,N_20884,N_20518);
nand U21685 (N_21685,N_20947,N_20846);
xnor U21686 (N_21686,N_20993,N_20118);
nand U21687 (N_21687,N_20297,N_20791);
xnor U21688 (N_21688,N_20489,N_20589);
and U21689 (N_21689,N_20813,N_20165);
or U21690 (N_21690,N_20950,N_20408);
and U21691 (N_21691,N_20466,N_20212);
xor U21692 (N_21692,N_20778,N_20587);
or U21693 (N_21693,N_20291,N_20286);
nand U21694 (N_21694,N_20832,N_20994);
nor U21695 (N_21695,N_20317,N_20525);
nor U21696 (N_21696,N_20558,N_20922);
and U21697 (N_21697,N_20576,N_20265);
nand U21698 (N_21698,N_20781,N_20004);
or U21699 (N_21699,N_20531,N_20565);
nor U21700 (N_21700,N_20738,N_20472);
nor U21701 (N_21701,N_20206,N_20825);
or U21702 (N_21702,N_20612,N_20008);
nand U21703 (N_21703,N_20759,N_20819);
nand U21704 (N_21704,N_20845,N_20699);
nand U21705 (N_21705,N_20741,N_20593);
and U21706 (N_21706,N_20597,N_20970);
or U21707 (N_21707,N_20788,N_20429);
nand U21708 (N_21708,N_20640,N_20527);
or U21709 (N_21709,N_20249,N_20284);
nor U21710 (N_21710,N_20395,N_20281);
or U21711 (N_21711,N_20836,N_20923);
xor U21712 (N_21712,N_20173,N_20343);
and U21713 (N_21713,N_20874,N_20721);
xor U21714 (N_21714,N_20058,N_20247);
or U21715 (N_21715,N_20821,N_20767);
nor U21716 (N_21716,N_20804,N_20636);
nor U21717 (N_21717,N_20384,N_20437);
or U21718 (N_21718,N_20856,N_20630);
nand U21719 (N_21719,N_20188,N_20994);
nand U21720 (N_21720,N_20100,N_20532);
or U21721 (N_21721,N_20185,N_20419);
or U21722 (N_21722,N_20844,N_20366);
xor U21723 (N_21723,N_20631,N_20556);
and U21724 (N_21724,N_20931,N_20782);
xnor U21725 (N_21725,N_20147,N_20826);
and U21726 (N_21726,N_20224,N_20132);
nor U21727 (N_21727,N_20125,N_20399);
and U21728 (N_21728,N_20925,N_20149);
xnor U21729 (N_21729,N_20437,N_20340);
nor U21730 (N_21730,N_20208,N_20407);
nor U21731 (N_21731,N_20171,N_20851);
xnor U21732 (N_21732,N_20087,N_20509);
nor U21733 (N_21733,N_20709,N_20361);
nor U21734 (N_21734,N_20923,N_20441);
or U21735 (N_21735,N_20578,N_20941);
and U21736 (N_21736,N_20771,N_20272);
nor U21737 (N_21737,N_20356,N_20434);
and U21738 (N_21738,N_20373,N_20597);
xnor U21739 (N_21739,N_20940,N_20221);
xnor U21740 (N_21740,N_20704,N_20249);
nand U21741 (N_21741,N_20294,N_20561);
nand U21742 (N_21742,N_20314,N_20955);
xnor U21743 (N_21743,N_20833,N_20915);
nor U21744 (N_21744,N_20438,N_20001);
and U21745 (N_21745,N_20261,N_20287);
or U21746 (N_21746,N_20105,N_20425);
or U21747 (N_21747,N_20863,N_20564);
or U21748 (N_21748,N_20069,N_20797);
nand U21749 (N_21749,N_20441,N_20345);
and U21750 (N_21750,N_20676,N_20936);
and U21751 (N_21751,N_20711,N_20309);
or U21752 (N_21752,N_20601,N_20544);
nor U21753 (N_21753,N_20946,N_20232);
nand U21754 (N_21754,N_20517,N_20754);
and U21755 (N_21755,N_20712,N_20228);
and U21756 (N_21756,N_20744,N_20673);
or U21757 (N_21757,N_20188,N_20886);
and U21758 (N_21758,N_20966,N_20778);
xnor U21759 (N_21759,N_20250,N_20840);
nand U21760 (N_21760,N_20143,N_20697);
and U21761 (N_21761,N_20278,N_20695);
nand U21762 (N_21762,N_20937,N_20471);
nor U21763 (N_21763,N_20416,N_20969);
xor U21764 (N_21764,N_20986,N_20838);
or U21765 (N_21765,N_20452,N_20712);
or U21766 (N_21766,N_20690,N_20395);
nor U21767 (N_21767,N_20178,N_20075);
nand U21768 (N_21768,N_20929,N_20320);
and U21769 (N_21769,N_20874,N_20524);
xnor U21770 (N_21770,N_20067,N_20173);
xor U21771 (N_21771,N_20733,N_20450);
nand U21772 (N_21772,N_20671,N_20435);
nor U21773 (N_21773,N_20258,N_20813);
nor U21774 (N_21774,N_20496,N_20056);
or U21775 (N_21775,N_20935,N_20288);
nor U21776 (N_21776,N_20543,N_20768);
xnor U21777 (N_21777,N_20706,N_20065);
nor U21778 (N_21778,N_20906,N_20728);
xor U21779 (N_21779,N_20874,N_20232);
or U21780 (N_21780,N_20280,N_20033);
xor U21781 (N_21781,N_20410,N_20742);
nor U21782 (N_21782,N_20450,N_20331);
xor U21783 (N_21783,N_20675,N_20017);
nand U21784 (N_21784,N_20109,N_20893);
nor U21785 (N_21785,N_20292,N_20240);
and U21786 (N_21786,N_20970,N_20786);
xnor U21787 (N_21787,N_20887,N_20443);
xnor U21788 (N_21788,N_20583,N_20280);
and U21789 (N_21789,N_20521,N_20756);
and U21790 (N_21790,N_20492,N_20182);
nor U21791 (N_21791,N_20737,N_20290);
and U21792 (N_21792,N_20711,N_20622);
nor U21793 (N_21793,N_20365,N_20207);
xor U21794 (N_21794,N_20595,N_20460);
nor U21795 (N_21795,N_20440,N_20757);
or U21796 (N_21796,N_20653,N_20303);
and U21797 (N_21797,N_20117,N_20265);
nor U21798 (N_21798,N_20800,N_20655);
xnor U21799 (N_21799,N_20201,N_20276);
nor U21800 (N_21800,N_20897,N_20359);
nor U21801 (N_21801,N_20633,N_20412);
and U21802 (N_21802,N_20708,N_20996);
or U21803 (N_21803,N_20519,N_20142);
or U21804 (N_21804,N_20969,N_20044);
and U21805 (N_21805,N_20271,N_20045);
nand U21806 (N_21806,N_20984,N_20502);
or U21807 (N_21807,N_20514,N_20900);
or U21808 (N_21808,N_20619,N_20346);
nor U21809 (N_21809,N_20314,N_20799);
nor U21810 (N_21810,N_20890,N_20790);
nor U21811 (N_21811,N_20465,N_20014);
xor U21812 (N_21812,N_20545,N_20026);
nand U21813 (N_21813,N_20917,N_20237);
nand U21814 (N_21814,N_20864,N_20744);
and U21815 (N_21815,N_20629,N_20754);
nand U21816 (N_21816,N_20742,N_20383);
and U21817 (N_21817,N_20848,N_20478);
nand U21818 (N_21818,N_20302,N_20388);
xnor U21819 (N_21819,N_20971,N_20734);
or U21820 (N_21820,N_20914,N_20467);
nand U21821 (N_21821,N_20750,N_20203);
nand U21822 (N_21822,N_20934,N_20036);
nor U21823 (N_21823,N_20133,N_20110);
nand U21824 (N_21824,N_20729,N_20608);
nor U21825 (N_21825,N_20349,N_20334);
nor U21826 (N_21826,N_20269,N_20487);
and U21827 (N_21827,N_20791,N_20650);
xor U21828 (N_21828,N_20225,N_20646);
nand U21829 (N_21829,N_20004,N_20118);
or U21830 (N_21830,N_20971,N_20146);
and U21831 (N_21831,N_20872,N_20899);
or U21832 (N_21832,N_20520,N_20032);
nand U21833 (N_21833,N_20959,N_20895);
nand U21834 (N_21834,N_20394,N_20346);
nor U21835 (N_21835,N_20061,N_20072);
nand U21836 (N_21836,N_20244,N_20296);
xor U21837 (N_21837,N_20659,N_20059);
or U21838 (N_21838,N_20764,N_20767);
or U21839 (N_21839,N_20840,N_20479);
or U21840 (N_21840,N_20876,N_20391);
nor U21841 (N_21841,N_20508,N_20312);
nand U21842 (N_21842,N_20238,N_20210);
nand U21843 (N_21843,N_20128,N_20830);
nor U21844 (N_21844,N_20949,N_20153);
nor U21845 (N_21845,N_20856,N_20214);
or U21846 (N_21846,N_20269,N_20672);
or U21847 (N_21847,N_20099,N_20903);
nor U21848 (N_21848,N_20755,N_20082);
nand U21849 (N_21849,N_20626,N_20397);
xnor U21850 (N_21850,N_20352,N_20985);
and U21851 (N_21851,N_20839,N_20248);
xor U21852 (N_21852,N_20900,N_20797);
nand U21853 (N_21853,N_20947,N_20331);
nand U21854 (N_21854,N_20368,N_20933);
xor U21855 (N_21855,N_20240,N_20132);
nand U21856 (N_21856,N_20417,N_20137);
xnor U21857 (N_21857,N_20762,N_20567);
nand U21858 (N_21858,N_20614,N_20843);
xnor U21859 (N_21859,N_20796,N_20224);
xnor U21860 (N_21860,N_20510,N_20203);
nor U21861 (N_21861,N_20377,N_20846);
or U21862 (N_21862,N_20270,N_20048);
nor U21863 (N_21863,N_20334,N_20929);
nor U21864 (N_21864,N_20449,N_20040);
xnor U21865 (N_21865,N_20032,N_20085);
nor U21866 (N_21866,N_20033,N_20758);
xnor U21867 (N_21867,N_20135,N_20874);
and U21868 (N_21868,N_20499,N_20146);
and U21869 (N_21869,N_20339,N_20785);
nor U21870 (N_21870,N_20888,N_20677);
and U21871 (N_21871,N_20063,N_20964);
nand U21872 (N_21872,N_20562,N_20713);
or U21873 (N_21873,N_20179,N_20969);
nor U21874 (N_21874,N_20854,N_20146);
xnor U21875 (N_21875,N_20659,N_20726);
xor U21876 (N_21876,N_20851,N_20163);
and U21877 (N_21877,N_20020,N_20679);
xnor U21878 (N_21878,N_20066,N_20356);
nor U21879 (N_21879,N_20839,N_20546);
nand U21880 (N_21880,N_20894,N_20215);
xnor U21881 (N_21881,N_20996,N_20901);
or U21882 (N_21882,N_20403,N_20730);
or U21883 (N_21883,N_20180,N_20809);
nand U21884 (N_21884,N_20650,N_20901);
nor U21885 (N_21885,N_20562,N_20422);
nor U21886 (N_21886,N_20531,N_20803);
xor U21887 (N_21887,N_20562,N_20274);
and U21888 (N_21888,N_20238,N_20707);
and U21889 (N_21889,N_20145,N_20993);
xnor U21890 (N_21890,N_20645,N_20305);
and U21891 (N_21891,N_20091,N_20012);
nand U21892 (N_21892,N_20060,N_20124);
nand U21893 (N_21893,N_20959,N_20353);
nand U21894 (N_21894,N_20571,N_20026);
or U21895 (N_21895,N_20812,N_20736);
nor U21896 (N_21896,N_20069,N_20047);
nor U21897 (N_21897,N_20644,N_20324);
and U21898 (N_21898,N_20052,N_20429);
nand U21899 (N_21899,N_20082,N_20371);
and U21900 (N_21900,N_20704,N_20631);
nand U21901 (N_21901,N_20923,N_20856);
nor U21902 (N_21902,N_20270,N_20440);
and U21903 (N_21903,N_20623,N_20339);
nand U21904 (N_21904,N_20592,N_20828);
xor U21905 (N_21905,N_20283,N_20874);
xnor U21906 (N_21906,N_20591,N_20430);
or U21907 (N_21907,N_20548,N_20505);
nor U21908 (N_21908,N_20617,N_20737);
and U21909 (N_21909,N_20526,N_20555);
or U21910 (N_21910,N_20264,N_20061);
or U21911 (N_21911,N_20458,N_20754);
xor U21912 (N_21912,N_20414,N_20064);
nand U21913 (N_21913,N_20504,N_20983);
nor U21914 (N_21914,N_20141,N_20664);
nand U21915 (N_21915,N_20955,N_20234);
xor U21916 (N_21916,N_20831,N_20145);
xnor U21917 (N_21917,N_20348,N_20925);
or U21918 (N_21918,N_20770,N_20518);
nand U21919 (N_21919,N_20589,N_20672);
or U21920 (N_21920,N_20869,N_20515);
nand U21921 (N_21921,N_20495,N_20831);
or U21922 (N_21922,N_20052,N_20694);
xor U21923 (N_21923,N_20093,N_20775);
nand U21924 (N_21924,N_20004,N_20503);
or U21925 (N_21925,N_20222,N_20391);
nor U21926 (N_21926,N_20207,N_20469);
xor U21927 (N_21927,N_20296,N_20722);
xnor U21928 (N_21928,N_20201,N_20638);
or U21929 (N_21929,N_20450,N_20108);
nand U21930 (N_21930,N_20934,N_20509);
and U21931 (N_21931,N_20890,N_20283);
xnor U21932 (N_21932,N_20248,N_20877);
xnor U21933 (N_21933,N_20458,N_20608);
nand U21934 (N_21934,N_20239,N_20234);
xor U21935 (N_21935,N_20121,N_20667);
or U21936 (N_21936,N_20889,N_20074);
nand U21937 (N_21937,N_20453,N_20608);
nand U21938 (N_21938,N_20429,N_20256);
nor U21939 (N_21939,N_20679,N_20296);
and U21940 (N_21940,N_20956,N_20463);
nand U21941 (N_21941,N_20215,N_20229);
xor U21942 (N_21942,N_20662,N_20786);
nand U21943 (N_21943,N_20892,N_20282);
and U21944 (N_21944,N_20974,N_20774);
and U21945 (N_21945,N_20829,N_20708);
nand U21946 (N_21946,N_20065,N_20991);
and U21947 (N_21947,N_20601,N_20347);
xnor U21948 (N_21948,N_20752,N_20879);
nand U21949 (N_21949,N_20528,N_20021);
and U21950 (N_21950,N_20363,N_20757);
and U21951 (N_21951,N_20452,N_20425);
xnor U21952 (N_21952,N_20989,N_20398);
nor U21953 (N_21953,N_20854,N_20232);
or U21954 (N_21954,N_20614,N_20168);
xor U21955 (N_21955,N_20849,N_20005);
or U21956 (N_21956,N_20401,N_20413);
or U21957 (N_21957,N_20632,N_20420);
nand U21958 (N_21958,N_20188,N_20433);
nor U21959 (N_21959,N_20070,N_20352);
or U21960 (N_21960,N_20522,N_20421);
and U21961 (N_21961,N_20514,N_20695);
xor U21962 (N_21962,N_20184,N_20298);
xnor U21963 (N_21963,N_20308,N_20856);
and U21964 (N_21964,N_20545,N_20729);
xnor U21965 (N_21965,N_20284,N_20147);
nor U21966 (N_21966,N_20709,N_20528);
xnor U21967 (N_21967,N_20286,N_20786);
or U21968 (N_21968,N_20966,N_20312);
nand U21969 (N_21969,N_20853,N_20269);
xor U21970 (N_21970,N_20788,N_20623);
xnor U21971 (N_21971,N_20450,N_20756);
xnor U21972 (N_21972,N_20827,N_20658);
xnor U21973 (N_21973,N_20110,N_20715);
nand U21974 (N_21974,N_20792,N_20534);
nand U21975 (N_21975,N_20499,N_20747);
xnor U21976 (N_21976,N_20841,N_20327);
xor U21977 (N_21977,N_20911,N_20788);
xor U21978 (N_21978,N_20543,N_20852);
xor U21979 (N_21979,N_20423,N_20509);
or U21980 (N_21980,N_20975,N_20138);
or U21981 (N_21981,N_20901,N_20728);
and U21982 (N_21982,N_20284,N_20218);
xor U21983 (N_21983,N_20951,N_20110);
nor U21984 (N_21984,N_20005,N_20123);
or U21985 (N_21985,N_20973,N_20352);
nand U21986 (N_21986,N_20516,N_20168);
nand U21987 (N_21987,N_20213,N_20114);
and U21988 (N_21988,N_20165,N_20608);
xor U21989 (N_21989,N_20169,N_20978);
or U21990 (N_21990,N_20667,N_20887);
xnor U21991 (N_21991,N_20960,N_20529);
or U21992 (N_21992,N_20805,N_20819);
nand U21993 (N_21993,N_20177,N_20304);
nand U21994 (N_21994,N_20258,N_20957);
xnor U21995 (N_21995,N_20364,N_20854);
xor U21996 (N_21996,N_20145,N_20614);
nor U21997 (N_21997,N_20138,N_20715);
nand U21998 (N_21998,N_20417,N_20688);
nand U21999 (N_21999,N_20748,N_20565);
or U22000 (N_22000,N_21661,N_21716);
nor U22001 (N_22001,N_21428,N_21441);
and U22002 (N_22002,N_21787,N_21700);
and U22003 (N_22003,N_21597,N_21745);
nor U22004 (N_22004,N_21276,N_21409);
nor U22005 (N_22005,N_21968,N_21375);
or U22006 (N_22006,N_21182,N_21359);
xnor U22007 (N_22007,N_21269,N_21030);
and U22008 (N_22008,N_21041,N_21087);
xor U22009 (N_22009,N_21010,N_21645);
xor U22010 (N_22010,N_21226,N_21086);
and U22011 (N_22011,N_21176,N_21130);
xor U22012 (N_22012,N_21563,N_21635);
nor U22013 (N_22013,N_21647,N_21803);
nand U22014 (N_22014,N_21321,N_21111);
nor U22015 (N_22015,N_21728,N_21495);
nand U22016 (N_22016,N_21806,N_21225);
and U22017 (N_22017,N_21117,N_21627);
nor U22018 (N_22018,N_21501,N_21574);
nor U22019 (N_22019,N_21699,N_21653);
nand U22020 (N_22020,N_21222,N_21953);
nand U22021 (N_22021,N_21917,N_21392);
or U22022 (N_22022,N_21984,N_21673);
nand U22023 (N_22023,N_21457,N_21108);
and U22024 (N_22024,N_21474,N_21139);
xor U22025 (N_22025,N_21196,N_21521);
and U22026 (N_22026,N_21398,N_21383);
nor U22027 (N_22027,N_21259,N_21790);
nor U22028 (N_22028,N_21303,N_21748);
xor U22029 (N_22029,N_21994,N_21159);
xor U22030 (N_22030,N_21479,N_21028);
nor U22031 (N_22031,N_21289,N_21496);
xnor U22032 (N_22032,N_21761,N_21184);
nand U22033 (N_22033,N_21911,N_21942);
or U22034 (N_22034,N_21508,N_21333);
and U22035 (N_22035,N_21444,N_21672);
nand U22036 (N_22036,N_21788,N_21809);
nand U22037 (N_22037,N_21224,N_21245);
nor U22038 (N_22038,N_21915,N_21737);
xor U22039 (N_22039,N_21529,N_21843);
and U22040 (N_22040,N_21988,N_21304);
and U22041 (N_22041,N_21499,N_21912);
xor U22042 (N_22042,N_21533,N_21577);
and U22043 (N_22043,N_21698,N_21373);
xor U22044 (N_22044,N_21660,N_21893);
nand U22045 (N_22045,N_21171,N_21920);
or U22046 (N_22046,N_21881,N_21278);
and U22047 (N_22047,N_21177,N_21578);
and U22048 (N_22048,N_21435,N_21561);
and U22049 (N_22049,N_21784,N_21418);
nor U22050 (N_22050,N_21361,N_21121);
nor U22051 (N_22051,N_21683,N_21460);
and U22052 (N_22052,N_21058,N_21534);
nor U22053 (N_22053,N_21451,N_21467);
xor U22054 (N_22054,N_21465,N_21341);
nor U22055 (N_22055,N_21610,N_21674);
nand U22056 (N_22056,N_21762,N_21816);
xor U22057 (N_22057,N_21141,N_21078);
nand U22058 (N_22058,N_21899,N_21879);
and U22059 (N_22059,N_21584,N_21972);
nor U22060 (N_22060,N_21997,N_21875);
xor U22061 (N_22061,N_21016,N_21414);
or U22062 (N_22062,N_21264,N_21270);
xor U22063 (N_22063,N_21487,N_21831);
or U22064 (N_22064,N_21828,N_21400);
and U22065 (N_22065,N_21516,N_21604);
xnor U22066 (N_22066,N_21100,N_21046);
and U22067 (N_22067,N_21931,N_21832);
or U22068 (N_22068,N_21725,N_21892);
and U22069 (N_22069,N_21151,N_21093);
nor U22070 (N_22070,N_21743,N_21147);
and U22071 (N_22071,N_21782,N_21128);
nor U22072 (N_22072,N_21913,N_21318);
and U22073 (N_22073,N_21693,N_21646);
and U22074 (N_22074,N_21985,N_21199);
nand U22075 (N_22075,N_21957,N_21658);
or U22076 (N_22076,N_21909,N_21345);
nand U22077 (N_22077,N_21613,N_21551);
nor U22078 (N_22078,N_21977,N_21554);
and U22079 (N_22079,N_21891,N_21694);
or U22080 (N_22080,N_21379,N_21498);
and U22081 (N_22081,N_21186,N_21095);
and U22082 (N_22082,N_21163,N_21466);
and U22083 (N_22083,N_21071,N_21509);
nor U22084 (N_22084,N_21288,N_21083);
nand U22085 (N_22085,N_21181,N_21003);
xor U22086 (N_22086,N_21277,N_21773);
nor U22087 (N_22087,N_21290,N_21742);
nand U22088 (N_22088,N_21475,N_21324);
xnor U22089 (N_22089,N_21120,N_21943);
or U22090 (N_22090,N_21469,N_21449);
or U22091 (N_22091,N_21328,N_21008);
xnor U22092 (N_22092,N_21011,N_21564);
nand U22093 (N_22093,N_21314,N_21999);
and U22094 (N_22094,N_21544,N_21013);
and U22095 (N_22095,N_21295,N_21824);
and U22096 (N_22096,N_21654,N_21160);
xor U22097 (N_22097,N_21037,N_21230);
nor U22098 (N_22098,N_21072,N_21812);
or U22099 (N_22099,N_21402,N_21884);
and U22100 (N_22100,N_21679,N_21097);
and U22101 (N_22101,N_21692,N_21726);
nor U22102 (N_22102,N_21265,N_21778);
nor U22103 (N_22103,N_21998,N_21014);
or U22104 (N_22104,N_21123,N_21894);
or U22105 (N_22105,N_21753,N_21520);
or U22106 (N_22106,N_21719,N_21606);
or U22107 (N_22107,N_21134,N_21174);
and U22108 (N_22108,N_21536,N_21631);
nor U22109 (N_22109,N_21591,N_21944);
nor U22110 (N_22110,N_21150,N_21585);
nand U22111 (N_22111,N_21396,N_21306);
and U22112 (N_22112,N_21919,N_21482);
xor U22113 (N_22113,N_21191,N_21914);
or U22114 (N_22114,N_21811,N_21838);
or U22115 (N_22115,N_21344,N_21488);
and U22116 (N_22116,N_21842,N_21101);
and U22117 (N_22117,N_21539,N_21161);
nor U22118 (N_22118,N_21808,N_21625);
xnor U22119 (N_22119,N_21605,N_21316);
nor U22120 (N_22120,N_21137,N_21733);
xor U22121 (N_22121,N_21330,N_21589);
xnor U22122 (N_22122,N_21395,N_21556);
xnor U22123 (N_22123,N_21109,N_21628);
nand U22124 (N_22124,N_21413,N_21966);
xor U22125 (N_22125,N_21031,N_21805);
nor U22126 (N_22126,N_21840,N_21979);
xor U22127 (N_22127,N_21619,N_21922);
nor U22128 (N_22128,N_21900,N_21401);
xor U22129 (N_22129,N_21601,N_21708);
xnor U22130 (N_22130,N_21547,N_21165);
or U22131 (N_22131,N_21193,N_21908);
and U22132 (N_22132,N_21019,N_21065);
nor U22133 (N_22133,N_21649,N_21676);
and U22134 (N_22134,N_21443,N_21995);
xor U22135 (N_22135,N_21667,N_21081);
nand U22136 (N_22136,N_21027,N_21825);
nor U22137 (N_22137,N_21924,N_21354);
nand U22138 (N_22138,N_21764,N_21731);
nor U22139 (N_22139,N_21242,N_21523);
nor U22140 (N_22140,N_21573,N_21009);
or U22141 (N_22141,N_21846,N_21369);
and U22142 (N_22142,N_21424,N_21727);
or U22143 (N_22143,N_21596,N_21455);
nand U22144 (N_22144,N_21056,N_21593);
nand U22145 (N_22145,N_21207,N_21655);
or U22146 (N_22146,N_21657,N_21696);
nor U22147 (N_22147,N_21091,N_21221);
xor U22148 (N_22148,N_21861,N_21143);
or U22149 (N_22149,N_21273,N_21140);
and U22150 (N_22150,N_21867,N_21734);
xnor U22151 (N_22151,N_21052,N_21180);
nor U22152 (N_22152,N_21490,N_21088);
xor U22153 (N_22153,N_21127,N_21680);
or U22154 (N_22154,N_21862,N_21412);
or U22155 (N_22155,N_21036,N_21153);
or U22156 (N_22156,N_21149,N_21434);
nor U22157 (N_22157,N_21371,N_21298);
xor U22158 (N_22158,N_21865,N_21335);
nand U22159 (N_22159,N_21067,N_21665);
nand U22160 (N_22160,N_21946,N_21374);
xnor U22161 (N_22161,N_21408,N_21952);
nand U22162 (N_22162,N_21659,N_21910);
and U22163 (N_22163,N_21332,N_21874);
or U22164 (N_22164,N_21257,N_21889);
nand U22165 (N_22165,N_21319,N_21292);
nand U22166 (N_22166,N_21210,N_21810);
xnor U22167 (N_22167,N_21393,N_21955);
or U22168 (N_22168,N_21029,N_21633);
xnor U22169 (N_22169,N_21850,N_21772);
nor U22170 (N_22170,N_21497,N_21993);
or U22171 (N_22171,N_21187,N_21250);
nor U22172 (N_22172,N_21632,N_21981);
or U22173 (N_22173,N_21722,N_21484);
and U22174 (N_22174,N_21602,N_21493);
xor U22175 (N_22175,N_21367,N_21172);
and U22176 (N_22176,N_21735,N_21525);
nor U22177 (N_22177,N_21550,N_21543);
nor U22178 (N_22178,N_21334,N_21962);
or U22179 (N_22179,N_21705,N_21930);
nor U22180 (N_22180,N_21815,N_21426);
and U22181 (N_22181,N_21399,N_21548);
or U22182 (N_22182,N_21611,N_21403);
nor U22183 (N_22183,N_21526,N_21820);
nand U22184 (N_22184,N_21220,N_21656);
and U22185 (N_22185,N_21779,N_21059);
xnor U22186 (N_22186,N_21144,N_21205);
xor U22187 (N_22187,N_21935,N_21253);
or U22188 (N_22188,N_21229,N_21795);
xnor U22189 (N_22189,N_21947,N_21362);
or U22190 (N_22190,N_21666,N_21410);
and U22191 (N_22191,N_21405,N_21928);
and U22192 (N_22192,N_21430,N_21559);
nand U22193 (N_22193,N_21387,N_21157);
nand U22194 (N_22194,N_21821,N_21975);
nor U22195 (N_22195,N_21723,N_21939);
nor U22196 (N_22196,N_21307,N_21063);
nor U22197 (N_22197,N_21118,N_21586);
nor U22198 (N_22198,N_21852,N_21471);
nand U22199 (N_22199,N_21427,N_21044);
and U22200 (N_22200,N_21227,N_21603);
xnor U22201 (N_22201,N_21446,N_21256);
or U22202 (N_22202,N_21886,N_21217);
nor U22203 (N_22203,N_21098,N_21974);
nor U22204 (N_22204,N_21807,N_21351);
xnor U22205 (N_22205,N_21888,N_21568);
or U22206 (N_22206,N_21080,N_21105);
xnor U22207 (N_22207,N_21670,N_21178);
and U22208 (N_22208,N_21195,N_21476);
and U22209 (N_22209,N_21348,N_21099);
nand U22210 (N_22210,N_21237,N_21706);
nand U22211 (N_22211,N_21480,N_21201);
and U22212 (N_22212,N_21185,N_21407);
nand U22213 (N_22213,N_21864,N_21051);
nor U22214 (N_22214,N_21263,N_21781);
and U22215 (N_22215,N_21916,N_21043);
xor U22216 (N_22216,N_21794,N_21204);
nand U22217 (N_22217,N_21189,N_21074);
or U22218 (N_22218,N_21459,N_21336);
nor U22219 (N_22219,N_21595,N_21829);
or U22220 (N_22220,N_21462,N_21156);
nor U22221 (N_22221,N_21464,N_21765);
and U22222 (N_22222,N_21858,N_21620);
nand U22223 (N_22223,N_21859,N_21502);
and U22224 (N_22224,N_21802,N_21154);
or U22225 (N_22225,N_21372,N_21384);
and U22226 (N_22226,N_21990,N_21394);
xor U22227 (N_22227,N_21510,N_21382);
nand U22228 (N_22228,N_21774,N_21724);
or U22229 (N_22229,N_21796,N_21949);
and U22230 (N_22230,N_21110,N_21869);
nor U22231 (N_22231,N_21114,N_21075);
nand U22232 (N_22232,N_21651,N_21976);
xnor U22233 (N_22233,N_21200,N_21769);
nand U22234 (N_22234,N_21125,N_21183);
or U22235 (N_22235,N_21209,N_21937);
xnor U22236 (N_22236,N_21094,N_21827);
or U22237 (N_22237,N_21575,N_21609);
xor U22238 (N_22238,N_21863,N_21729);
and U22239 (N_22239,N_21798,N_21518);
nor U22240 (N_22240,N_21311,N_21905);
and U22241 (N_22241,N_21126,N_21206);
nand U22242 (N_22242,N_21066,N_21793);
nor U22243 (N_22243,N_21901,N_21280);
nand U22244 (N_22244,N_21898,N_21702);
nor U22245 (N_22245,N_21662,N_21425);
and U22246 (N_22246,N_21356,N_21562);
or U22247 (N_22247,N_21388,N_21907);
nand U22248 (N_22248,N_21420,N_21238);
nor U22249 (N_22249,N_21638,N_21135);
xnor U22250 (N_22250,N_21983,N_21873);
nor U22251 (N_22251,N_21218,N_21216);
nor U22252 (N_22252,N_21818,N_21054);
or U22253 (N_22253,N_21274,N_21112);
nor U22254 (N_22254,N_21749,N_21040);
nor U22255 (N_22255,N_21223,N_21833);
xor U22256 (N_22256,N_21524,N_21145);
nand U22257 (N_22257,N_21079,N_21313);
nand U22258 (N_22258,N_21572,N_21535);
or U22259 (N_22259,N_21327,N_21755);
nor U22260 (N_22260,N_21717,N_21730);
and U22261 (N_22261,N_21844,N_21570);
xor U22262 (N_22262,N_21770,N_21678);
xnor U22263 (N_22263,N_21489,N_21323);
xnor U22264 (N_22264,N_21262,N_21823);
or U22265 (N_22265,N_21581,N_21275);
nor U22266 (N_22266,N_21004,N_21866);
nor U22267 (N_22267,N_21279,N_21255);
xnor U22268 (N_22268,N_21642,N_21712);
xnor U22269 (N_22269,N_21243,N_21050);
xor U22270 (N_22270,N_21532,N_21675);
nand U22271 (N_22271,N_21558,N_21624);
xnor U22272 (N_22272,N_21355,N_21945);
and U22273 (N_22273,N_21215,N_21309);
or U22274 (N_22274,N_21598,N_21709);
and U22275 (N_22275,N_21732,N_21337);
or U22276 (N_22276,N_21630,N_21073);
and U22277 (N_22277,N_21017,N_21799);
xor U22278 (N_22278,N_21517,N_21416);
nand U22279 (N_22279,N_21048,N_21148);
nor U22280 (N_22280,N_21569,N_21190);
nor U22281 (N_22281,N_21146,N_21880);
nand U22282 (N_22282,N_21677,N_21107);
or U22283 (N_22283,N_21018,N_21695);
or U22284 (N_22284,N_21877,N_21092);
xor U22285 (N_22285,N_21038,N_21233);
and U22286 (N_22286,N_21938,N_21251);
nor U22287 (N_22287,N_21515,N_21890);
or U22288 (N_22288,N_21545,N_21346);
nand U22289 (N_22289,N_21883,N_21214);
nand U22290 (N_22290,N_21167,N_21188);
nor U22291 (N_22291,N_21759,N_21711);
or U22292 (N_22292,N_21932,N_21576);
xnor U22293 (N_22293,N_21261,N_21357);
or U22294 (N_22294,N_21133,N_21791);
nor U22295 (N_22295,N_21514,N_21973);
nor U22296 (N_22296,N_21310,N_21049);
nand U22297 (N_22297,N_21197,N_21830);
xnor U22298 (N_22298,N_21746,N_21365);
nor U22299 (N_22299,N_21738,N_21583);
nor U22300 (N_22300,N_21115,N_21461);
and U22301 (N_22301,N_21084,N_21870);
nor U22302 (N_22302,N_21851,N_21228);
nand U22303 (N_22303,N_21352,N_21315);
xor U22304 (N_22304,N_21885,N_21347);
nand U22305 (N_22305,N_21353,N_21442);
nand U22306 (N_22306,N_21959,N_21904);
and U22307 (N_22307,N_21391,N_21964);
and U22308 (N_22308,N_21053,N_21194);
nor U22309 (N_22309,N_21540,N_21021);
xnor U22310 (N_22310,N_21485,N_21363);
nand U22311 (N_22311,N_21297,N_21232);
or U22312 (N_22312,N_21565,N_21042);
and U22313 (N_22313,N_21608,N_21234);
and U22314 (N_22314,N_21432,N_21338);
or U22315 (N_22315,N_21240,N_21339);
nor U22316 (N_22316,N_21438,N_21370);
nor U22317 (N_22317,N_21721,N_21247);
and U22318 (N_22318,N_21839,N_21211);
nor U22319 (N_22319,N_21744,N_21618);
xor U22320 (N_22320,N_21582,N_21213);
nand U22321 (N_22321,N_21389,N_21989);
or U22322 (N_22322,N_21329,N_21168);
xor U22323 (N_22323,N_21639,N_21640);
xnor U22324 (N_22324,N_21326,N_21766);
or U22325 (N_22325,N_21868,N_21445);
or U22326 (N_22326,N_21085,N_21106);
and U22327 (N_22327,N_21896,N_21077);
nand U22328 (N_22328,N_21854,N_21463);
nand U22329 (N_22329,N_21715,N_21267);
or U22330 (N_22330,N_21560,N_21248);
xor U22331 (N_22331,N_21650,N_21006);
nor U22332 (N_22332,N_21090,N_21697);
and U22333 (N_22333,N_21045,N_21923);
and U22334 (N_22334,N_21637,N_21477);
nor U22335 (N_22335,N_21797,N_21473);
nand U22336 (N_22336,N_21927,N_21948);
nor U22337 (N_22337,N_21668,N_21033);
or U22338 (N_22338,N_21713,N_21614);
nand U22339 (N_22339,N_21629,N_21486);
or U22340 (N_22340,N_21856,N_21012);
nor U22341 (N_22341,N_21785,N_21961);
nor U22342 (N_22342,N_21754,N_21024);
xor U22343 (N_22343,N_21644,N_21305);
xnor U22344 (N_22344,N_21836,N_21241);
and U22345 (N_22345,N_21138,N_21763);
or U22346 (N_22346,N_21512,N_21173);
or U22347 (N_22347,N_21537,N_21513);
xnor U22348 (N_22348,N_21057,N_21266);
nor U22349 (N_22349,N_21001,N_21505);
nand U22350 (N_22350,N_21268,N_21271);
xor U22351 (N_22351,N_21343,N_21690);
nor U22352 (N_22352,N_21192,N_21522);
or U22353 (N_22353,N_21129,N_21448);
nand U22354 (N_22354,N_21933,N_21982);
nor U22355 (N_22355,N_21720,N_21980);
or U22356 (N_22356,N_21136,N_21284);
nand U22357 (N_22357,N_21978,N_21320);
or U22358 (N_22358,N_21652,N_21047);
nor U22359 (N_22359,N_21579,N_21340);
and U22360 (N_22360,N_21062,N_21454);
nor U22361 (N_22361,N_21158,N_21992);
xor U22362 (N_22362,N_21623,N_21358);
nand U22363 (N_22363,N_21739,N_21089);
and U22364 (N_22364,N_21122,N_21934);
xor U22365 (N_22365,N_21847,N_21478);
nand U22366 (N_22366,N_21272,N_21260);
nand U22367 (N_22367,N_21022,N_21686);
xnor U22368 (N_22368,N_21710,N_21612);
or U22369 (N_22369,N_21929,N_21360);
xnor U22370 (N_22370,N_21826,N_21951);
or U22371 (N_22371,N_21542,N_21780);
nor U22372 (N_22372,N_21906,N_21950);
xor U22373 (N_22373,N_21747,N_21511);
and U22374 (N_22374,N_21860,N_21385);
or U22375 (N_22375,N_21472,N_21528);
xor U22376 (N_22376,N_21453,N_21350);
nand U22377 (N_22377,N_21895,N_21566);
nor U22378 (N_22378,N_21786,N_21504);
xnor U22379 (N_22379,N_21068,N_21538);
nand U22380 (N_22380,N_21817,N_21131);
xnor U22381 (N_22381,N_21855,N_21903);
or U22382 (N_22382,N_21622,N_21142);
or U22383 (N_22383,N_21155,N_21553);
and U22384 (N_22384,N_21882,N_21918);
or U22385 (N_22385,N_21804,N_21322);
and U22386 (N_22386,N_21835,N_21837);
and U22387 (N_22387,N_21671,N_21124);
nand U22388 (N_22388,N_21967,N_21617);
xor U22389 (N_22389,N_21249,N_21231);
xor U22390 (N_22390,N_21380,N_21299);
or U22391 (N_22391,N_21000,N_21703);
or U22392 (N_22392,N_21419,N_21246);
xor U22393 (N_22393,N_21740,N_21607);
nor U22394 (N_22394,N_21555,N_21281);
and U22395 (N_22395,N_21023,N_21116);
xor U22396 (N_22396,N_21636,N_21468);
nor U22397 (N_22397,N_21580,N_21039);
nand U22398 (N_22398,N_21494,N_21317);
xnor U22399 (N_22399,N_21119,N_21082);
nand U22400 (N_22400,N_21458,N_21404);
and U22401 (N_22401,N_21750,N_21055);
nand U22402 (N_22402,N_21258,N_21691);
and U22403 (N_22403,N_21175,N_21682);
xor U22404 (N_22404,N_21406,N_21594);
nand U22405 (N_22405,N_21431,N_21878);
and U22406 (N_22406,N_21969,N_21287);
xnor U22407 (N_22407,N_21368,N_21685);
nand U22408 (N_22408,N_21244,N_21102);
nor U22409 (N_22409,N_21312,N_21571);
nand U22410 (N_22410,N_21546,N_21198);
xor U22411 (N_22411,N_21848,N_21235);
nor U22412 (N_22412,N_21308,N_21436);
xnor U22413 (N_22413,N_21252,N_21113);
or U22414 (N_22414,N_21007,N_21549);
or U22415 (N_22415,N_21756,N_21301);
xnor U22416 (N_22416,N_21801,N_21887);
xnor U22417 (N_22417,N_21203,N_21970);
and U22418 (N_22418,N_21152,N_21587);
nor U22419 (N_22419,N_21688,N_21567);
and U22420 (N_22420,N_21871,N_21681);
or U22421 (N_22421,N_21777,N_21936);
xnor U22422 (N_22422,N_21364,N_21440);
or U22423 (N_22423,N_21751,N_21456);
and U22424 (N_22424,N_21776,N_21965);
xnor U22425 (N_22425,N_21902,N_21987);
or U22426 (N_22426,N_21069,N_21491);
or U22427 (N_22427,N_21437,N_21503);
nor U22428 (N_22428,N_21971,N_21684);
nand U22429 (N_22429,N_21789,N_21689);
xnor U22430 (N_22430,N_21701,N_21849);
xnor U22431 (N_22431,N_21822,N_21166);
nand U22432 (N_22432,N_21296,N_21954);
or U22433 (N_22433,N_21634,N_21897);
nor U22434 (N_22434,N_21219,N_21506);
nor U22435 (N_22435,N_21026,N_21282);
and U22436 (N_22436,N_21376,N_21669);
xor U22437 (N_22437,N_21519,N_21718);
xnor U22438 (N_22438,N_21300,N_21588);
nand U22439 (N_22439,N_21325,N_21590);
nor U22440 (N_22440,N_21792,N_21767);
or U22441 (N_22441,N_21857,N_21164);
or U22442 (N_22442,N_21283,N_21349);
nor U22443 (N_22443,N_21599,N_21294);
xnor U22444 (N_22444,N_21342,N_21845);
nor U22445 (N_22445,N_21104,N_21958);
or U22446 (N_22446,N_21500,N_21061);
or U22447 (N_22447,N_21530,N_21429);
nor U22448 (N_22448,N_21991,N_21507);
nand U22449 (N_22449,N_21390,N_21415);
nand U22450 (N_22450,N_21291,N_21926);
nor U22451 (N_22451,N_21212,N_21592);
xor U22452 (N_22452,N_21956,N_21447);
xor U22453 (N_22453,N_21819,N_21963);
and U22454 (N_22454,N_21236,N_21423);
xor U22455 (N_22455,N_21925,N_21421);
and U22456 (N_22456,N_21378,N_21616);
or U22457 (N_22457,N_21921,N_21664);
nand U22458 (N_22458,N_21621,N_21433);
or U22459 (N_22459,N_21381,N_21020);
nand U22460 (N_22460,N_21557,N_21814);
nand U22461 (N_22461,N_21752,N_21736);
and U22462 (N_22462,N_21872,N_21331);
or U22463 (N_22463,N_21417,N_21834);
nand U22464 (N_22464,N_21239,N_21202);
nand U22465 (N_22465,N_21876,N_21015);
nor U22466 (N_22466,N_21483,N_21103);
nand U22467 (N_22467,N_21768,N_21552);
nor U22468 (N_22468,N_21940,N_21254);
nand U22469 (N_22469,N_21470,N_21386);
xnor U22470 (N_22470,N_21450,N_21760);
nand U22471 (N_22471,N_21002,N_21452);
xnor U22472 (N_22472,N_21775,N_21841);
and U22473 (N_22473,N_21741,N_21064);
nor U22474 (N_22474,N_21169,N_21025);
xnor U22475 (N_22475,N_21531,N_21162);
xnor U22476 (N_22476,N_21663,N_21366);
xor U22477 (N_22477,N_21704,N_21757);
nor U22478 (N_22478,N_21179,N_21035);
nor U22479 (N_22479,N_21411,N_21286);
xor U22480 (N_22480,N_21377,N_21208);
and U22481 (N_22481,N_21714,N_21132);
or U22482 (N_22482,N_21783,N_21397);
nor U22483 (N_22483,N_21615,N_21481);
nor U22484 (N_22484,N_21302,N_21070);
xnor U22485 (N_22485,N_21960,N_21285);
nor U22486 (N_22486,N_21032,N_21813);
nor U22487 (N_22487,N_21492,N_21626);
or U22488 (N_22488,N_21527,N_21941);
and U22489 (N_22489,N_21600,N_21293);
nor U22490 (N_22490,N_21758,N_21060);
or U22491 (N_22491,N_21439,N_21771);
xor U22492 (N_22492,N_21853,N_21005);
nor U22493 (N_22493,N_21076,N_21648);
xnor U22494 (N_22494,N_21643,N_21707);
nor U22495 (N_22495,N_21641,N_21422);
nor U22496 (N_22496,N_21687,N_21986);
or U22497 (N_22497,N_21800,N_21996);
and U22498 (N_22498,N_21034,N_21096);
or U22499 (N_22499,N_21541,N_21170);
nand U22500 (N_22500,N_21184,N_21216);
xor U22501 (N_22501,N_21886,N_21352);
or U22502 (N_22502,N_21973,N_21264);
nand U22503 (N_22503,N_21377,N_21141);
and U22504 (N_22504,N_21302,N_21993);
xor U22505 (N_22505,N_21980,N_21046);
xor U22506 (N_22506,N_21095,N_21655);
xor U22507 (N_22507,N_21157,N_21167);
nand U22508 (N_22508,N_21291,N_21898);
nand U22509 (N_22509,N_21061,N_21668);
xor U22510 (N_22510,N_21399,N_21255);
nand U22511 (N_22511,N_21220,N_21364);
nor U22512 (N_22512,N_21400,N_21532);
nand U22513 (N_22513,N_21013,N_21437);
and U22514 (N_22514,N_21589,N_21730);
or U22515 (N_22515,N_21807,N_21344);
and U22516 (N_22516,N_21256,N_21291);
xnor U22517 (N_22517,N_21922,N_21701);
nand U22518 (N_22518,N_21106,N_21395);
or U22519 (N_22519,N_21895,N_21819);
xor U22520 (N_22520,N_21681,N_21962);
or U22521 (N_22521,N_21682,N_21311);
xor U22522 (N_22522,N_21993,N_21477);
nand U22523 (N_22523,N_21307,N_21557);
nand U22524 (N_22524,N_21060,N_21216);
or U22525 (N_22525,N_21972,N_21830);
xnor U22526 (N_22526,N_21469,N_21535);
and U22527 (N_22527,N_21413,N_21081);
nor U22528 (N_22528,N_21475,N_21886);
nand U22529 (N_22529,N_21753,N_21746);
and U22530 (N_22530,N_21903,N_21579);
nand U22531 (N_22531,N_21610,N_21716);
or U22532 (N_22532,N_21981,N_21778);
nand U22533 (N_22533,N_21458,N_21204);
or U22534 (N_22534,N_21239,N_21499);
nor U22535 (N_22535,N_21787,N_21422);
and U22536 (N_22536,N_21294,N_21760);
and U22537 (N_22537,N_21404,N_21751);
or U22538 (N_22538,N_21076,N_21072);
or U22539 (N_22539,N_21137,N_21623);
xnor U22540 (N_22540,N_21671,N_21370);
nand U22541 (N_22541,N_21093,N_21092);
or U22542 (N_22542,N_21634,N_21955);
nor U22543 (N_22543,N_21194,N_21866);
xnor U22544 (N_22544,N_21318,N_21575);
and U22545 (N_22545,N_21809,N_21939);
and U22546 (N_22546,N_21445,N_21938);
xor U22547 (N_22547,N_21246,N_21237);
or U22548 (N_22548,N_21547,N_21509);
xnor U22549 (N_22549,N_21577,N_21414);
and U22550 (N_22550,N_21485,N_21424);
or U22551 (N_22551,N_21649,N_21954);
nor U22552 (N_22552,N_21884,N_21621);
nor U22553 (N_22553,N_21368,N_21789);
nand U22554 (N_22554,N_21425,N_21401);
xor U22555 (N_22555,N_21961,N_21365);
and U22556 (N_22556,N_21805,N_21311);
nor U22557 (N_22557,N_21670,N_21645);
xor U22558 (N_22558,N_21276,N_21466);
nor U22559 (N_22559,N_21290,N_21488);
nor U22560 (N_22560,N_21520,N_21149);
nor U22561 (N_22561,N_21810,N_21671);
xnor U22562 (N_22562,N_21406,N_21217);
nand U22563 (N_22563,N_21374,N_21098);
or U22564 (N_22564,N_21958,N_21164);
or U22565 (N_22565,N_21318,N_21538);
or U22566 (N_22566,N_21393,N_21363);
nor U22567 (N_22567,N_21305,N_21672);
nor U22568 (N_22568,N_21157,N_21392);
nor U22569 (N_22569,N_21673,N_21772);
nand U22570 (N_22570,N_21331,N_21488);
xor U22571 (N_22571,N_21018,N_21951);
or U22572 (N_22572,N_21054,N_21111);
and U22573 (N_22573,N_21890,N_21417);
nor U22574 (N_22574,N_21259,N_21027);
nor U22575 (N_22575,N_21321,N_21468);
nand U22576 (N_22576,N_21541,N_21034);
or U22577 (N_22577,N_21734,N_21300);
nor U22578 (N_22578,N_21494,N_21160);
nand U22579 (N_22579,N_21683,N_21400);
and U22580 (N_22580,N_21169,N_21167);
and U22581 (N_22581,N_21521,N_21146);
nand U22582 (N_22582,N_21959,N_21471);
nand U22583 (N_22583,N_21158,N_21568);
nand U22584 (N_22584,N_21850,N_21028);
nor U22585 (N_22585,N_21425,N_21253);
and U22586 (N_22586,N_21235,N_21909);
xnor U22587 (N_22587,N_21845,N_21048);
or U22588 (N_22588,N_21235,N_21777);
nor U22589 (N_22589,N_21031,N_21184);
xnor U22590 (N_22590,N_21344,N_21725);
and U22591 (N_22591,N_21221,N_21878);
and U22592 (N_22592,N_21252,N_21937);
nor U22593 (N_22593,N_21928,N_21089);
or U22594 (N_22594,N_21616,N_21626);
nor U22595 (N_22595,N_21543,N_21049);
xnor U22596 (N_22596,N_21936,N_21401);
nor U22597 (N_22597,N_21044,N_21535);
or U22598 (N_22598,N_21298,N_21402);
nand U22599 (N_22599,N_21183,N_21936);
nor U22600 (N_22600,N_21529,N_21917);
or U22601 (N_22601,N_21504,N_21738);
nand U22602 (N_22602,N_21321,N_21571);
or U22603 (N_22603,N_21164,N_21636);
and U22604 (N_22604,N_21887,N_21102);
and U22605 (N_22605,N_21098,N_21113);
nor U22606 (N_22606,N_21723,N_21993);
xnor U22607 (N_22607,N_21019,N_21853);
xnor U22608 (N_22608,N_21024,N_21545);
and U22609 (N_22609,N_21831,N_21858);
and U22610 (N_22610,N_21709,N_21592);
or U22611 (N_22611,N_21841,N_21139);
or U22612 (N_22612,N_21530,N_21404);
xor U22613 (N_22613,N_21039,N_21584);
nor U22614 (N_22614,N_21818,N_21540);
nor U22615 (N_22615,N_21711,N_21176);
and U22616 (N_22616,N_21546,N_21932);
nand U22617 (N_22617,N_21285,N_21624);
nand U22618 (N_22618,N_21135,N_21916);
or U22619 (N_22619,N_21494,N_21203);
and U22620 (N_22620,N_21349,N_21816);
and U22621 (N_22621,N_21324,N_21310);
and U22622 (N_22622,N_21031,N_21924);
nand U22623 (N_22623,N_21257,N_21232);
xnor U22624 (N_22624,N_21800,N_21357);
and U22625 (N_22625,N_21578,N_21306);
nor U22626 (N_22626,N_21248,N_21355);
or U22627 (N_22627,N_21844,N_21342);
xnor U22628 (N_22628,N_21572,N_21781);
and U22629 (N_22629,N_21048,N_21627);
xnor U22630 (N_22630,N_21027,N_21662);
nor U22631 (N_22631,N_21487,N_21136);
nor U22632 (N_22632,N_21623,N_21740);
xnor U22633 (N_22633,N_21080,N_21468);
xor U22634 (N_22634,N_21003,N_21510);
nor U22635 (N_22635,N_21672,N_21599);
nor U22636 (N_22636,N_21043,N_21789);
xor U22637 (N_22637,N_21332,N_21477);
nand U22638 (N_22638,N_21015,N_21509);
nor U22639 (N_22639,N_21314,N_21316);
and U22640 (N_22640,N_21361,N_21729);
or U22641 (N_22641,N_21230,N_21079);
and U22642 (N_22642,N_21147,N_21924);
and U22643 (N_22643,N_21155,N_21060);
or U22644 (N_22644,N_21442,N_21011);
and U22645 (N_22645,N_21520,N_21033);
nand U22646 (N_22646,N_21037,N_21920);
or U22647 (N_22647,N_21344,N_21838);
or U22648 (N_22648,N_21969,N_21020);
or U22649 (N_22649,N_21143,N_21630);
nand U22650 (N_22650,N_21794,N_21265);
nor U22651 (N_22651,N_21174,N_21374);
xnor U22652 (N_22652,N_21473,N_21810);
nand U22653 (N_22653,N_21178,N_21562);
or U22654 (N_22654,N_21444,N_21061);
and U22655 (N_22655,N_21578,N_21041);
and U22656 (N_22656,N_21731,N_21169);
xnor U22657 (N_22657,N_21995,N_21718);
xor U22658 (N_22658,N_21198,N_21130);
nor U22659 (N_22659,N_21325,N_21132);
and U22660 (N_22660,N_21202,N_21017);
and U22661 (N_22661,N_21823,N_21389);
xor U22662 (N_22662,N_21298,N_21112);
or U22663 (N_22663,N_21672,N_21762);
nor U22664 (N_22664,N_21591,N_21786);
nand U22665 (N_22665,N_21394,N_21005);
and U22666 (N_22666,N_21433,N_21503);
nand U22667 (N_22667,N_21623,N_21559);
and U22668 (N_22668,N_21870,N_21823);
or U22669 (N_22669,N_21605,N_21132);
nand U22670 (N_22670,N_21592,N_21837);
nor U22671 (N_22671,N_21512,N_21222);
or U22672 (N_22672,N_21700,N_21524);
and U22673 (N_22673,N_21696,N_21114);
xnor U22674 (N_22674,N_21470,N_21703);
or U22675 (N_22675,N_21767,N_21239);
nor U22676 (N_22676,N_21901,N_21644);
xor U22677 (N_22677,N_21439,N_21046);
and U22678 (N_22678,N_21388,N_21197);
xor U22679 (N_22679,N_21332,N_21986);
or U22680 (N_22680,N_21532,N_21788);
xor U22681 (N_22681,N_21905,N_21269);
or U22682 (N_22682,N_21374,N_21914);
xor U22683 (N_22683,N_21855,N_21283);
nand U22684 (N_22684,N_21403,N_21728);
nand U22685 (N_22685,N_21874,N_21999);
nand U22686 (N_22686,N_21966,N_21050);
and U22687 (N_22687,N_21854,N_21706);
xnor U22688 (N_22688,N_21256,N_21749);
xor U22689 (N_22689,N_21294,N_21669);
nor U22690 (N_22690,N_21047,N_21306);
nand U22691 (N_22691,N_21482,N_21998);
nand U22692 (N_22692,N_21745,N_21791);
and U22693 (N_22693,N_21158,N_21112);
nand U22694 (N_22694,N_21000,N_21764);
or U22695 (N_22695,N_21019,N_21252);
or U22696 (N_22696,N_21806,N_21829);
nor U22697 (N_22697,N_21730,N_21075);
and U22698 (N_22698,N_21728,N_21501);
or U22699 (N_22699,N_21941,N_21514);
and U22700 (N_22700,N_21069,N_21184);
nand U22701 (N_22701,N_21865,N_21696);
and U22702 (N_22702,N_21000,N_21133);
nand U22703 (N_22703,N_21473,N_21195);
xor U22704 (N_22704,N_21143,N_21935);
or U22705 (N_22705,N_21271,N_21330);
nand U22706 (N_22706,N_21594,N_21435);
nor U22707 (N_22707,N_21367,N_21808);
and U22708 (N_22708,N_21284,N_21963);
xnor U22709 (N_22709,N_21913,N_21857);
nand U22710 (N_22710,N_21220,N_21259);
and U22711 (N_22711,N_21036,N_21767);
xnor U22712 (N_22712,N_21002,N_21822);
and U22713 (N_22713,N_21509,N_21179);
xor U22714 (N_22714,N_21549,N_21350);
or U22715 (N_22715,N_21910,N_21998);
and U22716 (N_22716,N_21691,N_21190);
xnor U22717 (N_22717,N_21905,N_21784);
nand U22718 (N_22718,N_21851,N_21560);
nor U22719 (N_22719,N_21400,N_21719);
xnor U22720 (N_22720,N_21865,N_21882);
or U22721 (N_22721,N_21489,N_21979);
nand U22722 (N_22722,N_21688,N_21275);
nand U22723 (N_22723,N_21666,N_21084);
xnor U22724 (N_22724,N_21803,N_21101);
and U22725 (N_22725,N_21272,N_21987);
nor U22726 (N_22726,N_21793,N_21185);
xnor U22727 (N_22727,N_21777,N_21609);
and U22728 (N_22728,N_21156,N_21747);
or U22729 (N_22729,N_21427,N_21112);
nand U22730 (N_22730,N_21828,N_21544);
or U22731 (N_22731,N_21338,N_21890);
nor U22732 (N_22732,N_21736,N_21525);
xor U22733 (N_22733,N_21371,N_21995);
or U22734 (N_22734,N_21827,N_21931);
nor U22735 (N_22735,N_21585,N_21315);
xnor U22736 (N_22736,N_21183,N_21362);
and U22737 (N_22737,N_21805,N_21616);
and U22738 (N_22738,N_21543,N_21815);
nor U22739 (N_22739,N_21262,N_21333);
nand U22740 (N_22740,N_21644,N_21296);
nor U22741 (N_22741,N_21214,N_21029);
xnor U22742 (N_22742,N_21905,N_21880);
xor U22743 (N_22743,N_21766,N_21277);
or U22744 (N_22744,N_21428,N_21914);
nand U22745 (N_22745,N_21032,N_21055);
xnor U22746 (N_22746,N_21962,N_21083);
xnor U22747 (N_22747,N_21918,N_21144);
or U22748 (N_22748,N_21665,N_21158);
and U22749 (N_22749,N_21538,N_21549);
and U22750 (N_22750,N_21040,N_21456);
and U22751 (N_22751,N_21134,N_21589);
or U22752 (N_22752,N_21249,N_21238);
xor U22753 (N_22753,N_21627,N_21473);
nor U22754 (N_22754,N_21443,N_21858);
nor U22755 (N_22755,N_21023,N_21009);
nor U22756 (N_22756,N_21679,N_21978);
xor U22757 (N_22757,N_21590,N_21887);
or U22758 (N_22758,N_21622,N_21123);
nand U22759 (N_22759,N_21651,N_21458);
and U22760 (N_22760,N_21559,N_21507);
nand U22761 (N_22761,N_21905,N_21116);
xor U22762 (N_22762,N_21191,N_21373);
or U22763 (N_22763,N_21587,N_21421);
nor U22764 (N_22764,N_21476,N_21007);
nand U22765 (N_22765,N_21146,N_21124);
nor U22766 (N_22766,N_21006,N_21295);
xor U22767 (N_22767,N_21504,N_21374);
or U22768 (N_22768,N_21866,N_21801);
nand U22769 (N_22769,N_21418,N_21707);
and U22770 (N_22770,N_21818,N_21660);
nand U22771 (N_22771,N_21110,N_21442);
and U22772 (N_22772,N_21726,N_21460);
or U22773 (N_22773,N_21238,N_21323);
or U22774 (N_22774,N_21325,N_21966);
nor U22775 (N_22775,N_21716,N_21425);
xor U22776 (N_22776,N_21205,N_21178);
or U22777 (N_22777,N_21376,N_21086);
or U22778 (N_22778,N_21238,N_21258);
nand U22779 (N_22779,N_21637,N_21780);
xor U22780 (N_22780,N_21550,N_21315);
xnor U22781 (N_22781,N_21561,N_21317);
xnor U22782 (N_22782,N_21835,N_21202);
and U22783 (N_22783,N_21888,N_21944);
and U22784 (N_22784,N_21637,N_21524);
and U22785 (N_22785,N_21226,N_21773);
and U22786 (N_22786,N_21467,N_21808);
xnor U22787 (N_22787,N_21391,N_21324);
nand U22788 (N_22788,N_21764,N_21771);
nor U22789 (N_22789,N_21937,N_21343);
and U22790 (N_22790,N_21806,N_21925);
nand U22791 (N_22791,N_21973,N_21266);
xor U22792 (N_22792,N_21757,N_21861);
nand U22793 (N_22793,N_21483,N_21345);
xor U22794 (N_22794,N_21848,N_21020);
nand U22795 (N_22795,N_21799,N_21182);
and U22796 (N_22796,N_21159,N_21860);
nand U22797 (N_22797,N_21286,N_21238);
or U22798 (N_22798,N_21462,N_21006);
nand U22799 (N_22799,N_21074,N_21077);
nor U22800 (N_22800,N_21268,N_21854);
nor U22801 (N_22801,N_21986,N_21235);
xnor U22802 (N_22802,N_21013,N_21283);
nor U22803 (N_22803,N_21773,N_21696);
nand U22804 (N_22804,N_21244,N_21225);
nor U22805 (N_22805,N_21833,N_21172);
or U22806 (N_22806,N_21742,N_21225);
nand U22807 (N_22807,N_21019,N_21814);
nand U22808 (N_22808,N_21644,N_21870);
or U22809 (N_22809,N_21817,N_21583);
and U22810 (N_22810,N_21087,N_21855);
nand U22811 (N_22811,N_21492,N_21972);
nor U22812 (N_22812,N_21896,N_21095);
nand U22813 (N_22813,N_21419,N_21344);
nor U22814 (N_22814,N_21283,N_21615);
nor U22815 (N_22815,N_21706,N_21194);
nand U22816 (N_22816,N_21891,N_21381);
xor U22817 (N_22817,N_21256,N_21789);
nand U22818 (N_22818,N_21886,N_21175);
nand U22819 (N_22819,N_21747,N_21939);
and U22820 (N_22820,N_21980,N_21025);
and U22821 (N_22821,N_21674,N_21471);
nor U22822 (N_22822,N_21585,N_21905);
nor U22823 (N_22823,N_21915,N_21135);
or U22824 (N_22824,N_21713,N_21217);
xor U22825 (N_22825,N_21616,N_21529);
or U22826 (N_22826,N_21231,N_21174);
and U22827 (N_22827,N_21290,N_21634);
and U22828 (N_22828,N_21301,N_21036);
nand U22829 (N_22829,N_21532,N_21765);
nor U22830 (N_22830,N_21481,N_21050);
or U22831 (N_22831,N_21254,N_21721);
and U22832 (N_22832,N_21599,N_21264);
nor U22833 (N_22833,N_21461,N_21341);
and U22834 (N_22834,N_21299,N_21550);
xor U22835 (N_22835,N_21951,N_21737);
or U22836 (N_22836,N_21934,N_21600);
xor U22837 (N_22837,N_21380,N_21470);
and U22838 (N_22838,N_21194,N_21319);
or U22839 (N_22839,N_21160,N_21679);
xnor U22840 (N_22840,N_21351,N_21014);
nor U22841 (N_22841,N_21723,N_21974);
xnor U22842 (N_22842,N_21731,N_21145);
nor U22843 (N_22843,N_21866,N_21013);
nor U22844 (N_22844,N_21205,N_21075);
xor U22845 (N_22845,N_21627,N_21284);
nand U22846 (N_22846,N_21863,N_21540);
nor U22847 (N_22847,N_21522,N_21928);
and U22848 (N_22848,N_21359,N_21729);
or U22849 (N_22849,N_21531,N_21992);
and U22850 (N_22850,N_21975,N_21994);
xnor U22851 (N_22851,N_21374,N_21893);
and U22852 (N_22852,N_21801,N_21569);
nand U22853 (N_22853,N_21851,N_21297);
xnor U22854 (N_22854,N_21412,N_21984);
and U22855 (N_22855,N_21074,N_21423);
nand U22856 (N_22856,N_21112,N_21873);
and U22857 (N_22857,N_21032,N_21586);
xnor U22858 (N_22858,N_21302,N_21824);
nand U22859 (N_22859,N_21823,N_21237);
xnor U22860 (N_22860,N_21370,N_21622);
xor U22861 (N_22861,N_21571,N_21075);
nand U22862 (N_22862,N_21525,N_21415);
nand U22863 (N_22863,N_21728,N_21326);
and U22864 (N_22864,N_21199,N_21883);
nand U22865 (N_22865,N_21451,N_21554);
nor U22866 (N_22866,N_21244,N_21054);
or U22867 (N_22867,N_21651,N_21598);
xor U22868 (N_22868,N_21388,N_21974);
nand U22869 (N_22869,N_21123,N_21609);
nand U22870 (N_22870,N_21528,N_21430);
xnor U22871 (N_22871,N_21516,N_21960);
nand U22872 (N_22872,N_21014,N_21472);
xor U22873 (N_22873,N_21061,N_21091);
nand U22874 (N_22874,N_21519,N_21207);
or U22875 (N_22875,N_21806,N_21916);
nand U22876 (N_22876,N_21350,N_21243);
nand U22877 (N_22877,N_21686,N_21499);
nor U22878 (N_22878,N_21290,N_21925);
xnor U22879 (N_22879,N_21084,N_21882);
nand U22880 (N_22880,N_21916,N_21856);
or U22881 (N_22881,N_21734,N_21018);
or U22882 (N_22882,N_21565,N_21535);
nor U22883 (N_22883,N_21655,N_21249);
xor U22884 (N_22884,N_21515,N_21596);
nor U22885 (N_22885,N_21320,N_21211);
and U22886 (N_22886,N_21160,N_21746);
nand U22887 (N_22887,N_21505,N_21191);
or U22888 (N_22888,N_21526,N_21598);
nand U22889 (N_22889,N_21839,N_21447);
xnor U22890 (N_22890,N_21605,N_21299);
xor U22891 (N_22891,N_21527,N_21347);
nor U22892 (N_22892,N_21961,N_21537);
xor U22893 (N_22893,N_21062,N_21619);
or U22894 (N_22894,N_21062,N_21054);
nand U22895 (N_22895,N_21748,N_21518);
xnor U22896 (N_22896,N_21269,N_21528);
nand U22897 (N_22897,N_21849,N_21069);
or U22898 (N_22898,N_21331,N_21390);
or U22899 (N_22899,N_21348,N_21241);
or U22900 (N_22900,N_21937,N_21132);
nand U22901 (N_22901,N_21277,N_21492);
nor U22902 (N_22902,N_21883,N_21285);
xor U22903 (N_22903,N_21272,N_21704);
nand U22904 (N_22904,N_21497,N_21385);
nor U22905 (N_22905,N_21226,N_21423);
nor U22906 (N_22906,N_21586,N_21006);
or U22907 (N_22907,N_21302,N_21607);
or U22908 (N_22908,N_21991,N_21472);
or U22909 (N_22909,N_21856,N_21491);
nand U22910 (N_22910,N_21645,N_21581);
nand U22911 (N_22911,N_21420,N_21052);
nor U22912 (N_22912,N_21912,N_21701);
xnor U22913 (N_22913,N_21737,N_21608);
xor U22914 (N_22914,N_21157,N_21160);
nand U22915 (N_22915,N_21252,N_21291);
nand U22916 (N_22916,N_21073,N_21511);
or U22917 (N_22917,N_21303,N_21735);
xnor U22918 (N_22918,N_21373,N_21642);
nand U22919 (N_22919,N_21365,N_21448);
nand U22920 (N_22920,N_21640,N_21741);
nor U22921 (N_22921,N_21426,N_21888);
and U22922 (N_22922,N_21547,N_21435);
nor U22923 (N_22923,N_21180,N_21080);
nor U22924 (N_22924,N_21974,N_21628);
and U22925 (N_22925,N_21895,N_21232);
nand U22926 (N_22926,N_21301,N_21528);
nand U22927 (N_22927,N_21000,N_21740);
nor U22928 (N_22928,N_21885,N_21350);
nor U22929 (N_22929,N_21869,N_21832);
xnor U22930 (N_22930,N_21417,N_21365);
and U22931 (N_22931,N_21416,N_21689);
or U22932 (N_22932,N_21840,N_21879);
and U22933 (N_22933,N_21297,N_21353);
nor U22934 (N_22934,N_21541,N_21548);
xnor U22935 (N_22935,N_21263,N_21900);
xnor U22936 (N_22936,N_21989,N_21347);
or U22937 (N_22937,N_21287,N_21639);
or U22938 (N_22938,N_21575,N_21454);
nor U22939 (N_22939,N_21564,N_21938);
nand U22940 (N_22940,N_21883,N_21810);
and U22941 (N_22941,N_21571,N_21680);
and U22942 (N_22942,N_21685,N_21000);
xnor U22943 (N_22943,N_21377,N_21406);
nor U22944 (N_22944,N_21915,N_21298);
or U22945 (N_22945,N_21886,N_21703);
or U22946 (N_22946,N_21524,N_21352);
nand U22947 (N_22947,N_21607,N_21357);
and U22948 (N_22948,N_21535,N_21829);
nor U22949 (N_22949,N_21916,N_21286);
nand U22950 (N_22950,N_21471,N_21948);
nand U22951 (N_22951,N_21925,N_21945);
nand U22952 (N_22952,N_21242,N_21467);
nor U22953 (N_22953,N_21816,N_21284);
and U22954 (N_22954,N_21946,N_21311);
and U22955 (N_22955,N_21301,N_21186);
or U22956 (N_22956,N_21305,N_21740);
xnor U22957 (N_22957,N_21649,N_21610);
and U22958 (N_22958,N_21037,N_21096);
nand U22959 (N_22959,N_21061,N_21190);
or U22960 (N_22960,N_21296,N_21595);
or U22961 (N_22961,N_21691,N_21557);
nor U22962 (N_22962,N_21187,N_21065);
or U22963 (N_22963,N_21746,N_21132);
nand U22964 (N_22964,N_21299,N_21980);
and U22965 (N_22965,N_21198,N_21104);
xnor U22966 (N_22966,N_21343,N_21634);
and U22967 (N_22967,N_21544,N_21035);
or U22968 (N_22968,N_21009,N_21470);
nand U22969 (N_22969,N_21371,N_21416);
nor U22970 (N_22970,N_21296,N_21637);
and U22971 (N_22971,N_21403,N_21316);
nor U22972 (N_22972,N_21947,N_21729);
nor U22973 (N_22973,N_21740,N_21229);
nand U22974 (N_22974,N_21723,N_21892);
nor U22975 (N_22975,N_21635,N_21552);
and U22976 (N_22976,N_21971,N_21138);
or U22977 (N_22977,N_21034,N_21109);
nor U22978 (N_22978,N_21492,N_21591);
and U22979 (N_22979,N_21563,N_21787);
and U22980 (N_22980,N_21701,N_21306);
nor U22981 (N_22981,N_21919,N_21264);
xor U22982 (N_22982,N_21681,N_21931);
or U22983 (N_22983,N_21337,N_21663);
xor U22984 (N_22984,N_21925,N_21736);
and U22985 (N_22985,N_21866,N_21619);
nor U22986 (N_22986,N_21345,N_21297);
xor U22987 (N_22987,N_21646,N_21633);
or U22988 (N_22988,N_21301,N_21066);
nor U22989 (N_22989,N_21908,N_21236);
and U22990 (N_22990,N_21712,N_21095);
xnor U22991 (N_22991,N_21663,N_21388);
nand U22992 (N_22992,N_21473,N_21742);
nor U22993 (N_22993,N_21406,N_21856);
and U22994 (N_22994,N_21713,N_21704);
xnor U22995 (N_22995,N_21456,N_21254);
and U22996 (N_22996,N_21372,N_21916);
nor U22997 (N_22997,N_21592,N_21798);
xnor U22998 (N_22998,N_21667,N_21530);
nand U22999 (N_22999,N_21309,N_21701);
and U23000 (N_23000,N_22590,N_22246);
nor U23001 (N_23001,N_22913,N_22504);
xnor U23002 (N_23002,N_22624,N_22593);
nand U23003 (N_23003,N_22135,N_22976);
or U23004 (N_23004,N_22533,N_22148);
nor U23005 (N_23005,N_22880,N_22337);
or U23006 (N_23006,N_22000,N_22923);
nor U23007 (N_23007,N_22037,N_22437);
or U23008 (N_23008,N_22832,N_22274);
xnor U23009 (N_23009,N_22256,N_22393);
nor U23010 (N_23010,N_22189,N_22397);
nor U23011 (N_23011,N_22086,N_22546);
and U23012 (N_23012,N_22157,N_22562);
nor U23013 (N_23013,N_22782,N_22443);
nor U23014 (N_23014,N_22937,N_22664);
xor U23015 (N_23015,N_22527,N_22772);
nor U23016 (N_23016,N_22183,N_22260);
nand U23017 (N_23017,N_22795,N_22843);
nor U23018 (N_23018,N_22060,N_22431);
nand U23019 (N_23019,N_22739,N_22052);
xnor U23020 (N_23020,N_22817,N_22126);
or U23021 (N_23021,N_22534,N_22839);
or U23022 (N_23022,N_22366,N_22182);
nand U23023 (N_23023,N_22849,N_22522);
nor U23024 (N_23024,N_22545,N_22237);
nand U23025 (N_23025,N_22088,N_22804);
nor U23026 (N_23026,N_22700,N_22422);
nor U23027 (N_23027,N_22800,N_22160);
and U23028 (N_23028,N_22973,N_22446);
nor U23029 (N_23029,N_22673,N_22385);
xor U23030 (N_23030,N_22865,N_22899);
and U23031 (N_23031,N_22760,N_22144);
nand U23032 (N_23032,N_22398,N_22945);
nand U23033 (N_23033,N_22611,N_22910);
or U23034 (N_23034,N_22672,N_22621);
xor U23035 (N_23035,N_22978,N_22436);
nand U23036 (N_23036,N_22339,N_22459);
and U23037 (N_23037,N_22289,N_22348);
nand U23038 (N_23038,N_22616,N_22073);
or U23039 (N_23039,N_22582,N_22379);
or U23040 (N_23040,N_22821,N_22654);
and U23041 (N_23041,N_22044,N_22234);
or U23042 (N_23042,N_22685,N_22479);
or U23043 (N_23043,N_22131,N_22346);
or U23044 (N_23044,N_22262,N_22215);
nor U23045 (N_23045,N_22888,N_22136);
xnor U23046 (N_23046,N_22854,N_22404);
and U23047 (N_23047,N_22302,N_22474);
nand U23048 (N_23048,N_22396,N_22592);
nand U23049 (N_23049,N_22637,N_22402);
nor U23050 (N_23050,N_22021,N_22958);
and U23051 (N_23051,N_22884,N_22036);
and U23052 (N_23052,N_22569,N_22738);
or U23053 (N_23053,N_22894,N_22075);
nand U23054 (N_23054,N_22934,N_22585);
xor U23055 (N_23055,N_22373,N_22825);
and U23056 (N_23056,N_22505,N_22626);
nand U23057 (N_23057,N_22689,N_22120);
nor U23058 (N_23058,N_22241,N_22803);
or U23059 (N_23059,N_22191,N_22208);
nand U23060 (N_23060,N_22190,N_22315);
nand U23061 (N_23061,N_22407,N_22158);
or U23062 (N_23062,N_22648,N_22147);
and U23063 (N_23063,N_22567,N_22311);
nand U23064 (N_23064,N_22478,N_22283);
nor U23065 (N_23065,N_22779,N_22740);
or U23066 (N_23066,N_22362,N_22501);
or U23067 (N_23067,N_22046,N_22969);
xnor U23068 (N_23068,N_22496,N_22460);
or U23069 (N_23069,N_22439,N_22091);
or U23070 (N_23070,N_22391,N_22461);
nand U23071 (N_23071,N_22635,N_22330);
xor U23072 (N_23072,N_22902,N_22040);
nor U23073 (N_23073,N_22508,N_22276);
nor U23074 (N_23074,N_22336,N_22642);
nand U23075 (N_23075,N_22809,N_22494);
nand U23076 (N_23076,N_22956,N_22462);
xor U23077 (N_23077,N_22892,N_22758);
nand U23078 (N_23078,N_22333,N_22823);
nand U23079 (N_23079,N_22442,N_22070);
xnor U23080 (N_23080,N_22889,N_22032);
or U23081 (N_23081,N_22759,N_22149);
or U23082 (N_23082,N_22993,N_22098);
nor U23083 (N_23083,N_22565,N_22087);
or U23084 (N_23084,N_22503,N_22952);
nor U23085 (N_23085,N_22445,N_22519);
or U23086 (N_23086,N_22798,N_22658);
nand U23087 (N_23087,N_22702,N_22187);
xor U23088 (N_23088,N_22376,N_22007);
xnor U23089 (N_23089,N_22080,N_22513);
xor U23090 (N_23090,N_22690,N_22421);
nor U23091 (N_23091,N_22216,N_22159);
xor U23092 (N_23092,N_22145,N_22206);
nor U23093 (N_23093,N_22022,N_22555);
or U23094 (N_23094,N_22763,N_22155);
nor U23095 (N_23095,N_22859,N_22451);
or U23096 (N_23096,N_22946,N_22855);
xor U23097 (N_23097,N_22473,N_22925);
xor U23098 (N_23098,N_22105,N_22343);
xor U23099 (N_23099,N_22423,N_22631);
and U23100 (N_23100,N_22467,N_22778);
nor U23101 (N_23101,N_22805,N_22982);
and U23102 (N_23102,N_22417,N_22477);
xnor U23103 (N_23103,N_22570,N_22305);
and U23104 (N_23104,N_22563,N_22099);
and U23105 (N_23105,N_22320,N_22224);
nand U23106 (N_23106,N_22677,N_22649);
and U23107 (N_23107,N_22598,N_22568);
xnor U23108 (N_23108,N_22537,N_22701);
nand U23109 (N_23109,N_22202,N_22604);
or U23110 (N_23110,N_22143,N_22222);
xnor U23111 (N_23111,N_22847,N_22742);
nor U23112 (N_23112,N_22732,N_22180);
xor U23113 (N_23113,N_22788,N_22801);
xnor U23114 (N_23114,N_22656,N_22510);
and U23115 (N_23115,N_22205,N_22990);
or U23116 (N_23116,N_22811,N_22428);
or U23117 (N_23117,N_22752,N_22295);
nor U23118 (N_23118,N_22725,N_22324);
and U23119 (N_23119,N_22253,N_22622);
nor U23120 (N_23120,N_22650,N_22786);
nand U23121 (N_23121,N_22067,N_22128);
or U23122 (N_23122,N_22651,N_22048);
xor U23123 (N_23123,N_22970,N_22612);
xor U23124 (N_23124,N_22613,N_22671);
nor U23125 (N_23125,N_22981,N_22317);
xnor U23126 (N_23126,N_22850,N_22053);
or U23127 (N_23127,N_22257,N_22543);
or U23128 (N_23128,N_22652,N_22620);
and U23129 (N_23129,N_22198,N_22254);
nand U23130 (N_23130,N_22367,N_22259);
nand U23131 (N_23131,N_22245,N_22242);
or U23132 (N_23132,N_22166,N_22172);
and U23133 (N_23133,N_22574,N_22340);
nand U23134 (N_23134,N_22369,N_22481);
or U23135 (N_23135,N_22281,N_22578);
xnor U23136 (N_23136,N_22907,N_22193);
xnor U23137 (N_23137,N_22667,N_22118);
nand U23138 (N_23138,N_22090,N_22056);
xor U23139 (N_23139,N_22390,N_22223);
and U23140 (N_23140,N_22236,N_22077);
xor U23141 (N_23141,N_22863,N_22600);
and U23142 (N_23142,N_22587,N_22065);
nor U23143 (N_23143,N_22525,N_22108);
xnor U23144 (N_23144,N_22745,N_22818);
xor U23145 (N_23145,N_22916,N_22948);
or U23146 (N_23146,N_22139,N_22867);
nor U23147 (N_23147,N_22006,N_22589);
and U23148 (N_23148,N_22718,N_22845);
nor U23149 (N_23149,N_22230,N_22140);
and U23150 (N_23150,N_22532,N_22174);
and U23151 (N_23151,N_22872,N_22416);
and U23152 (N_23152,N_22908,N_22175);
or U23153 (N_23153,N_22614,N_22235);
nor U23154 (N_23154,N_22171,N_22017);
xor U23155 (N_23155,N_22928,N_22030);
or U23156 (N_23156,N_22917,N_22432);
xor U23157 (N_23157,N_22891,N_22729);
or U23158 (N_23158,N_22703,N_22829);
nor U23159 (N_23159,N_22394,N_22146);
xor U23160 (N_23160,N_22848,N_22015);
nand U23161 (N_23161,N_22680,N_22350);
nand U23162 (N_23162,N_22777,N_22749);
nor U23163 (N_23163,N_22433,N_22392);
nand U23164 (N_23164,N_22342,N_22449);
nand U23165 (N_23165,N_22231,N_22607);
and U23166 (N_23166,N_22188,N_22399);
and U23167 (N_23167,N_22325,N_22711);
nand U23168 (N_23168,N_22453,N_22411);
or U23169 (N_23169,N_22409,N_22873);
nor U23170 (N_23170,N_22676,N_22045);
nand U23171 (N_23171,N_22291,N_22802);
and U23172 (N_23172,N_22258,N_22270);
nand U23173 (N_23173,N_22529,N_22357);
or U23174 (N_23174,N_22356,N_22168);
nor U23175 (N_23175,N_22141,N_22345);
xor U23176 (N_23176,N_22016,N_22783);
and U23177 (N_23177,N_22014,N_22535);
xnor U23178 (N_23178,N_22360,N_22034);
xor U23179 (N_23179,N_22864,N_22674);
and U23180 (N_23180,N_22542,N_22999);
and U23181 (N_23181,N_22435,N_22964);
and U23182 (N_23182,N_22294,N_22985);
and U23183 (N_23183,N_22893,N_22789);
xnor U23184 (N_23184,N_22430,N_22822);
nor U23185 (N_23185,N_22881,N_22837);
nand U23186 (N_23186,N_22192,N_22492);
or U23187 (N_23187,N_22933,N_22413);
or U23188 (N_23188,N_22748,N_22009);
and U23189 (N_23189,N_22214,N_22374);
xor U23190 (N_23190,N_22002,N_22349);
nor U23191 (N_23191,N_22735,N_22704);
nor U23192 (N_23192,N_22842,N_22418);
xnor U23193 (N_23193,N_22719,N_22544);
and U23194 (N_23194,N_22662,N_22572);
or U23195 (N_23195,N_22164,N_22733);
nand U23196 (N_23196,N_22887,N_22785);
xnor U23197 (N_23197,N_22408,N_22988);
nor U23198 (N_23198,N_22344,N_22271);
or U23199 (N_23199,N_22341,N_22723);
nand U23200 (N_23200,N_22915,N_22942);
and U23201 (N_23201,N_22039,N_22526);
nor U23202 (N_23202,N_22041,N_22914);
or U23203 (N_23203,N_22469,N_22475);
xnor U23204 (N_23204,N_22440,N_22996);
nand U23205 (N_23205,N_22316,N_22512);
and U23206 (N_23206,N_22554,N_22820);
nor U23207 (N_23207,N_22249,N_22815);
or U23208 (N_23208,N_22977,N_22401);
and U23209 (N_23209,N_22196,N_22661);
or U23210 (N_23210,N_22548,N_22938);
nand U23211 (N_23211,N_22035,N_22714);
or U23212 (N_23212,N_22744,N_22781);
nor U23213 (N_23213,N_22010,N_22290);
xor U23214 (N_23214,N_22628,N_22197);
or U23215 (N_23215,N_22233,N_22211);
xnor U23216 (N_23216,N_22100,N_22944);
and U23217 (N_23217,N_22365,N_22666);
xor U23218 (N_23218,N_22903,N_22247);
and U23219 (N_23219,N_22272,N_22476);
nor U23220 (N_23220,N_22874,N_22471);
nor U23221 (N_23221,N_22954,N_22886);
nand U23222 (N_23222,N_22943,N_22991);
or U23223 (N_23223,N_22737,N_22828);
or U23224 (N_23224,N_22636,N_22498);
and U23225 (N_23225,N_22328,N_22713);
or U23226 (N_23226,N_22728,N_22116);
or U23227 (N_23227,N_22113,N_22212);
and U23228 (N_23228,N_22152,N_22688);
and U23229 (N_23229,N_22826,N_22868);
and U23230 (N_23230,N_22008,N_22107);
xor U23231 (N_23231,N_22064,N_22071);
nand U23232 (N_23232,N_22178,N_22922);
nand U23233 (N_23233,N_22441,N_22655);
nand U23234 (N_23234,N_22581,N_22617);
xor U23235 (N_23235,N_22997,N_22594);
and U23236 (N_23236,N_22285,N_22757);
or U23237 (N_23237,N_22878,N_22921);
xnor U23238 (N_23238,N_22054,N_22074);
nor U23239 (N_23239,N_22455,N_22971);
nand U23240 (N_23240,N_22500,N_22089);
and U23241 (N_23241,N_22314,N_22059);
xor U23242 (N_23242,N_22687,N_22736);
nor U23243 (N_23243,N_22521,N_22905);
nor U23244 (N_23244,N_22250,N_22154);
or U23245 (N_23245,N_22406,N_22297);
or U23246 (N_23246,N_22615,N_22994);
xnor U23247 (N_23247,N_22967,N_22630);
and U23248 (N_23248,N_22601,N_22286);
xnor U23249 (N_23249,N_22480,N_22707);
or U23250 (N_23250,N_22151,N_22683);
xor U23251 (N_23251,N_22588,N_22860);
xor U23252 (N_23252,N_22097,N_22775);
nand U23253 (N_23253,N_22995,N_22632);
xor U23254 (N_23254,N_22103,N_22605);
xor U23255 (N_23255,N_22117,N_22659);
or U23256 (N_23256,N_22919,N_22576);
nor U23257 (N_23257,N_22361,N_22304);
or U23258 (N_23258,N_22063,N_22472);
and U23259 (N_23259,N_22493,N_22807);
xnor U23260 (N_23260,N_22110,N_22866);
xnor U23261 (N_23261,N_22382,N_22061);
and U23262 (N_23262,N_22571,N_22043);
xor U23263 (N_23263,N_22452,N_22012);
nand U23264 (N_23264,N_22055,N_22833);
xnor U23265 (N_23265,N_22808,N_22011);
xnor U23266 (N_23266,N_22918,N_22643);
xnor U23267 (N_23267,N_22653,N_22420);
nand U23268 (N_23268,N_22083,N_22835);
nand U23269 (N_23269,N_22024,N_22112);
nand U23270 (N_23270,N_22722,N_22799);
and U23271 (N_23271,N_22213,N_22966);
nor U23272 (N_23272,N_22912,N_22114);
or U23273 (N_23273,N_22218,N_22531);
and U23274 (N_23274,N_22068,N_22960);
nor U23275 (N_23275,N_22608,N_22470);
nor U23276 (N_23276,N_22388,N_22627);
nor U23277 (N_23277,N_22380,N_22026);
and U23278 (N_23278,N_22221,N_22766);
or U23279 (N_23279,N_22559,N_22633);
and U23280 (N_23280,N_22927,N_22194);
and U23281 (N_23281,N_22950,N_22490);
nand U23282 (N_23282,N_22909,N_22623);
nand U23283 (N_23283,N_22920,N_22106);
nand U23284 (N_23284,N_22911,N_22025);
nor U23285 (N_23285,N_22558,N_22583);
xor U23286 (N_23286,N_22355,N_22705);
xor U23287 (N_23287,N_22227,N_22338);
nand U23288 (N_23288,N_22184,N_22057);
nor U23289 (N_23289,N_22170,N_22368);
and U23290 (N_23290,N_22104,N_22530);
or U23291 (N_23291,N_22381,N_22384);
and U23292 (N_23292,N_22323,N_22890);
nand U23293 (N_23293,N_22463,N_22185);
or U23294 (N_23294,N_22939,N_22507);
nor U23295 (N_23295,N_22038,N_22499);
or U23296 (N_23296,N_22895,N_22482);
nor U23297 (N_23297,N_22844,N_22599);
nor U23298 (N_23298,N_22634,N_22949);
or U23299 (N_23299,N_22906,N_22596);
xnor U23300 (N_23300,N_22307,N_22896);
or U23301 (N_23301,N_22840,N_22326);
xnor U23302 (N_23302,N_22209,N_22931);
or U23303 (N_23303,N_22806,N_22491);
nand U23304 (N_23304,N_22790,N_22424);
or U23305 (N_23305,N_22541,N_22142);
xnor U23306 (N_23306,N_22458,N_22303);
nand U23307 (N_23307,N_22827,N_22965);
nand U23308 (N_23308,N_22313,N_22298);
or U23309 (N_23309,N_22217,N_22553);
and U23310 (N_23310,N_22836,N_22414);
or U23311 (N_23311,N_22207,N_22426);
nand U23312 (N_23312,N_22983,N_22641);
nor U23313 (N_23313,N_22095,N_22968);
nand U23314 (N_23314,N_22084,N_22846);
and U23315 (N_23315,N_22386,N_22647);
nand U23316 (N_23316,N_22852,N_22502);
and U23317 (N_23317,N_22228,N_22727);
nand U23318 (N_23318,N_22448,N_22287);
nand U23319 (N_23319,N_22756,N_22998);
xnor U23320 (N_23320,N_22762,N_22549);
xnor U23321 (N_23321,N_22591,N_22625);
nor U23322 (N_23322,N_22962,N_22638);
and U23323 (N_23323,N_22004,N_22639);
or U23324 (N_23324,N_22792,N_22769);
xnor U23325 (N_23325,N_22177,N_22780);
nor U23326 (N_23326,N_22301,N_22699);
and U23327 (N_23327,N_22841,N_22796);
xor U23328 (N_23328,N_22686,N_22101);
nand U23329 (N_23329,N_22812,N_22838);
or U23330 (N_23330,N_22288,N_22353);
or U23331 (N_23331,N_22280,N_22708);
nor U23332 (N_23332,N_22179,N_22883);
nor U23333 (N_23333,N_22584,N_22539);
nor U23334 (N_23334,N_22322,N_22679);
xnor U23335 (N_23335,N_22951,N_22869);
and U23336 (N_23336,N_22243,N_22163);
xor U23337 (N_23337,N_22468,N_22755);
xnor U23338 (N_23338,N_22768,N_22042);
or U23339 (N_23339,N_22536,N_22875);
or U23340 (N_23340,N_22019,N_22540);
nand U23341 (N_23341,N_22447,N_22743);
and U23342 (N_23342,N_22425,N_22400);
nor U23343 (N_23343,N_22329,N_22516);
or U23344 (N_23344,N_22359,N_22419);
xor U23345 (N_23345,N_22047,N_22484);
nor U23346 (N_23346,N_22248,N_22266);
xor U23347 (N_23347,N_22932,N_22602);
and U23348 (N_23348,N_22444,N_22308);
nand U23349 (N_23349,N_22963,N_22610);
xnor U23350 (N_23350,N_22364,N_22225);
or U23351 (N_23351,N_22961,N_22682);
and U23352 (N_23352,N_22123,N_22309);
xnor U23353 (N_23353,N_22957,N_22127);
nand U23354 (N_23354,N_22566,N_22358);
xnor U23355 (N_23355,N_22831,N_22856);
and U23356 (N_23356,N_22870,N_22879);
and U23357 (N_23357,N_22684,N_22564);
or U23358 (N_23358,N_22986,N_22940);
or U23359 (N_23359,N_22791,N_22132);
xor U23360 (N_23360,N_22371,N_22595);
or U23361 (N_23361,N_22200,N_22619);
xnor U23362 (N_23362,N_22560,N_22646);
nor U23363 (N_23363,N_22776,N_22058);
and U23364 (N_23364,N_22334,N_22122);
or U23365 (N_23365,N_22268,N_22706);
and U23366 (N_23366,N_22240,N_22352);
nor U23367 (N_23367,N_22715,N_22987);
or U23368 (N_23368,N_22137,N_22877);
or U23369 (N_23369,N_22434,N_22618);
nor U23370 (N_23370,N_22851,N_22121);
and U23371 (N_23371,N_22784,N_22109);
and U23372 (N_23372,N_22318,N_22277);
and U23373 (N_23373,N_22263,N_22765);
nand U23374 (N_23374,N_22031,N_22517);
and U23375 (N_23375,N_22941,N_22485);
xor U23376 (N_23376,N_22165,N_22861);
nor U23377 (N_23377,N_22028,N_22857);
nand U23378 (N_23378,N_22427,N_22495);
xnor U23379 (N_23379,N_22751,N_22279);
nor U23380 (N_23380,N_22239,N_22538);
xor U23381 (N_23381,N_22111,N_22665);
or U23382 (N_23382,N_22753,N_22747);
or U23383 (N_23383,N_22195,N_22787);
nor U23384 (N_23384,N_22310,N_22457);
nand U23385 (N_23385,N_22900,N_22293);
nand U23386 (N_23386,N_22082,N_22694);
nor U23387 (N_23387,N_22085,N_22306);
or U23388 (N_23388,N_22984,N_22936);
xnor U23389 (N_23389,N_22347,N_22681);
nand U23390 (N_23390,N_22331,N_22229);
nor U23391 (N_23391,N_22520,N_22410);
nor U23392 (N_23392,N_22102,N_22275);
xor U23393 (N_23393,N_22813,N_22528);
xnor U23394 (N_23394,N_22746,N_22050);
and U23395 (N_23395,N_22754,N_22354);
xnor U23396 (N_23396,N_22093,N_22924);
or U23397 (N_23397,N_22678,N_22199);
nand U23398 (N_23398,N_22771,N_22001);
nand U23399 (N_23399,N_22454,N_22953);
and U23400 (N_23400,N_22173,N_22824);
or U23401 (N_23401,N_22657,N_22720);
and U23402 (N_23402,N_22974,N_22489);
nor U23403 (N_23403,N_22710,N_22018);
and U23404 (N_23404,N_22292,N_22695);
xor U23405 (N_23405,N_22712,N_22816);
and U23406 (N_23406,N_22013,N_22547);
nand U23407 (N_23407,N_22094,N_22675);
and U23408 (N_23408,N_22269,N_22403);
and U23409 (N_23409,N_22130,N_22834);
xnor U23410 (N_23410,N_22220,N_22351);
nand U23411 (N_23411,N_22129,N_22989);
nand U23412 (N_23412,N_22603,N_22669);
or U23413 (N_23413,N_22265,N_22049);
nand U23414 (N_23414,N_22935,N_22134);
xnor U23415 (N_23415,N_22640,N_22261);
and U23416 (N_23416,N_22335,N_22550);
and U23417 (N_23417,N_22405,N_22926);
nor U23418 (N_23418,N_22668,N_22979);
xor U23419 (N_23419,N_22586,N_22696);
nor U23420 (N_23420,N_22955,N_22124);
nand U23421 (N_23421,N_22814,N_22556);
nand U23422 (N_23422,N_22518,N_22959);
xor U23423 (N_23423,N_22273,N_22697);
nor U23424 (N_23424,N_22660,N_22162);
nand U23425 (N_23425,N_22876,N_22079);
and U23426 (N_23426,N_22387,N_22858);
nor U23427 (N_23427,N_22514,N_22415);
nor U23428 (N_23428,N_22332,N_22201);
nand U23429 (N_23429,N_22794,N_22370);
nand U23430 (N_23430,N_22862,N_22138);
xor U23431 (N_23431,N_22204,N_22515);
xor U23432 (N_23432,N_22552,N_22020);
xnor U23433 (N_23433,N_22487,N_22300);
or U23434 (N_23434,N_22509,N_22488);
or U23435 (N_23435,N_22580,N_22483);
and U23436 (N_23436,N_22465,N_22264);
nand U23437 (N_23437,N_22267,N_22372);
nand U23438 (N_23438,N_22629,N_22663);
nor U23439 (N_23439,N_22076,N_22389);
xor U23440 (N_23440,N_22561,N_22312);
nor U23441 (N_23441,N_22027,N_22299);
and U23442 (N_23442,N_22078,N_22450);
nand U23443 (N_23443,N_22670,N_22810);
and U23444 (N_23444,N_22551,N_22161);
and U23445 (N_23445,N_22296,N_22597);
nand U23446 (N_23446,N_22726,N_22003);
or U23447 (N_23447,N_22575,N_22606);
nand U23448 (N_23448,N_22609,N_22523);
nor U23449 (N_23449,N_22731,N_22897);
and U23450 (N_23450,N_22115,N_22252);
and U23451 (N_23451,N_22975,N_22023);
xor U23452 (N_23452,N_22203,N_22062);
xor U23453 (N_23453,N_22029,N_22383);
nand U23454 (N_23454,N_22377,N_22167);
xor U23455 (N_23455,N_22069,N_22721);
and U23456 (N_23456,N_22992,N_22819);
and U23457 (N_23457,N_22226,N_22119);
xnor U23458 (N_23458,N_22282,N_22464);
nand U23459 (N_23459,N_22573,N_22750);
or U23460 (N_23460,N_22767,N_22456);
nor U23461 (N_23461,N_22797,N_22980);
or U23462 (N_23462,N_22770,N_22692);
nor U23463 (N_23463,N_22238,N_22005);
and U23464 (N_23464,N_22724,N_22133);
nand U23465 (N_23465,N_22947,N_22255);
nor U23466 (N_23466,N_22774,N_22375);
and U23467 (N_23467,N_22176,N_22698);
or U23468 (N_23468,N_22321,N_22764);
or U23469 (N_23469,N_22885,N_22066);
xor U23470 (N_23470,N_22644,N_22901);
xnor U23471 (N_23471,N_22186,N_22579);
or U23472 (N_23472,N_22081,N_22741);
nor U23473 (N_23473,N_22251,N_22092);
xnor U23474 (N_23474,N_22898,N_22327);
xnor U23475 (N_23475,N_22363,N_22853);
xnor U23476 (N_23476,N_22466,N_22761);
nand U23477 (N_23477,N_22904,N_22730);
nor U23478 (N_23478,N_22645,N_22169);
or U23479 (N_23479,N_22232,N_22716);
xor U23480 (N_23480,N_22709,N_22524);
and U23481 (N_23481,N_22051,N_22278);
or U23482 (N_23482,N_22181,N_22972);
nand U23483 (N_23483,N_22378,N_22219);
nor U23484 (N_23484,N_22319,N_22497);
and U23485 (N_23485,N_22930,N_22693);
xor U23486 (N_23486,N_22429,N_22511);
nor U23487 (N_23487,N_22153,N_22096);
or U23488 (N_23488,N_22717,N_22557);
nor U23489 (N_23489,N_22033,N_22830);
nor U23490 (N_23490,N_22506,N_22438);
and U23491 (N_23491,N_22577,N_22773);
xnor U23492 (N_23492,N_22156,N_22150);
xor U23493 (N_23493,N_22284,N_22125);
and U23494 (N_23494,N_22734,N_22486);
or U23495 (N_23495,N_22929,N_22412);
and U23496 (N_23496,N_22072,N_22871);
or U23497 (N_23497,N_22395,N_22244);
xnor U23498 (N_23498,N_22210,N_22691);
xor U23499 (N_23499,N_22793,N_22882);
or U23500 (N_23500,N_22469,N_22458);
nand U23501 (N_23501,N_22470,N_22232);
or U23502 (N_23502,N_22559,N_22006);
nand U23503 (N_23503,N_22417,N_22093);
xnor U23504 (N_23504,N_22640,N_22795);
nand U23505 (N_23505,N_22837,N_22655);
nor U23506 (N_23506,N_22701,N_22992);
nor U23507 (N_23507,N_22940,N_22291);
and U23508 (N_23508,N_22114,N_22146);
nand U23509 (N_23509,N_22816,N_22751);
nor U23510 (N_23510,N_22649,N_22410);
and U23511 (N_23511,N_22581,N_22862);
nand U23512 (N_23512,N_22174,N_22046);
xnor U23513 (N_23513,N_22018,N_22354);
xor U23514 (N_23514,N_22794,N_22982);
or U23515 (N_23515,N_22334,N_22755);
or U23516 (N_23516,N_22442,N_22379);
and U23517 (N_23517,N_22011,N_22292);
xnor U23518 (N_23518,N_22617,N_22409);
nand U23519 (N_23519,N_22352,N_22329);
nand U23520 (N_23520,N_22421,N_22810);
xnor U23521 (N_23521,N_22409,N_22015);
or U23522 (N_23522,N_22724,N_22691);
nor U23523 (N_23523,N_22232,N_22164);
xor U23524 (N_23524,N_22252,N_22887);
and U23525 (N_23525,N_22085,N_22604);
nand U23526 (N_23526,N_22492,N_22122);
or U23527 (N_23527,N_22390,N_22177);
nand U23528 (N_23528,N_22524,N_22060);
or U23529 (N_23529,N_22440,N_22103);
and U23530 (N_23530,N_22443,N_22687);
and U23531 (N_23531,N_22798,N_22973);
nor U23532 (N_23532,N_22917,N_22339);
or U23533 (N_23533,N_22934,N_22917);
or U23534 (N_23534,N_22680,N_22407);
nand U23535 (N_23535,N_22420,N_22910);
nor U23536 (N_23536,N_22722,N_22882);
and U23537 (N_23537,N_22436,N_22643);
nor U23538 (N_23538,N_22072,N_22190);
nand U23539 (N_23539,N_22513,N_22992);
nor U23540 (N_23540,N_22536,N_22098);
nand U23541 (N_23541,N_22727,N_22275);
or U23542 (N_23542,N_22893,N_22150);
nor U23543 (N_23543,N_22363,N_22093);
nand U23544 (N_23544,N_22939,N_22872);
or U23545 (N_23545,N_22011,N_22000);
nor U23546 (N_23546,N_22370,N_22119);
and U23547 (N_23547,N_22597,N_22048);
nor U23548 (N_23548,N_22139,N_22436);
xnor U23549 (N_23549,N_22603,N_22270);
or U23550 (N_23550,N_22005,N_22675);
or U23551 (N_23551,N_22062,N_22357);
nor U23552 (N_23552,N_22292,N_22477);
or U23553 (N_23553,N_22934,N_22469);
nand U23554 (N_23554,N_22626,N_22212);
xnor U23555 (N_23555,N_22670,N_22401);
or U23556 (N_23556,N_22473,N_22819);
nor U23557 (N_23557,N_22675,N_22736);
xor U23558 (N_23558,N_22222,N_22406);
and U23559 (N_23559,N_22040,N_22407);
or U23560 (N_23560,N_22116,N_22254);
xnor U23561 (N_23561,N_22960,N_22469);
nor U23562 (N_23562,N_22036,N_22621);
nor U23563 (N_23563,N_22836,N_22094);
or U23564 (N_23564,N_22437,N_22156);
xnor U23565 (N_23565,N_22690,N_22243);
or U23566 (N_23566,N_22773,N_22126);
or U23567 (N_23567,N_22771,N_22619);
xor U23568 (N_23568,N_22097,N_22447);
xor U23569 (N_23569,N_22876,N_22935);
nand U23570 (N_23570,N_22863,N_22964);
or U23571 (N_23571,N_22688,N_22359);
or U23572 (N_23572,N_22318,N_22159);
or U23573 (N_23573,N_22156,N_22778);
nand U23574 (N_23574,N_22373,N_22067);
xor U23575 (N_23575,N_22770,N_22138);
nor U23576 (N_23576,N_22273,N_22701);
nand U23577 (N_23577,N_22724,N_22482);
and U23578 (N_23578,N_22237,N_22022);
or U23579 (N_23579,N_22188,N_22812);
xor U23580 (N_23580,N_22173,N_22181);
nand U23581 (N_23581,N_22095,N_22552);
nor U23582 (N_23582,N_22350,N_22182);
nor U23583 (N_23583,N_22055,N_22078);
nor U23584 (N_23584,N_22788,N_22338);
nand U23585 (N_23585,N_22804,N_22764);
and U23586 (N_23586,N_22235,N_22145);
and U23587 (N_23587,N_22976,N_22378);
nor U23588 (N_23588,N_22579,N_22324);
nor U23589 (N_23589,N_22997,N_22749);
and U23590 (N_23590,N_22517,N_22689);
and U23591 (N_23591,N_22808,N_22335);
xor U23592 (N_23592,N_22690,N_22772);
nor U23593 (N_23593,N_22889,N_22738);
or U23594 (N_23594,N_22219,N_22350);
nand U23595 (N_23595,N_22681,N_22132);
and U23596 (N_23596,N_22951,N_22589);
nor U23597 (N_23597,N_22868,N_22358);
nand U23598 (N_23598,N_22932,N_22747);
or U23599 (N_23599,N_22551,N_22767);
nor U23600 (N_23600,N_22789,N_22295);
nand U23601 (N_23601,N_22008,N_22132);
or U23602 (N_23602,N_22064,N_22860);
xor U23603 (N_23603,N_22940,N_22373);
nand U23604 (N_23604,N_22269,N_22259);
xnor U23605 (N_23605,N_22922,N_22581);
or U23606 (N_23606,N_22503,N_22364);
nor U23607 (N_23607,N_22031,N_22911);
xnor U23608 (N_23608,N_22449,N_22003);
or U23609 (N_23609,N_22464,N_22584);
nand U23610 (N_23610,N_22740,N_22136);
and U23611 (N_23611,N_22939,N_22736);
nand U23612 (N_23612,N_22446,N_22858);
or U23613 (N_23613,N_22140,N_22997);
or U23614 (N_23614,N_22251,N_22455);
nor U23615 (N_23615,N_22672,N_22775);
nor U23616 (N_23616,N_22653,N_22202);
xnor U23617 (N_23617,N_22267,N_22808);
nor U23618 (N_23618,N_22803,N_22548);
or U23619 (N_23619,N_22922,N_22935);
xnor U23620 (N_23620,N_22795,N_22384);
xnor U23621 (N_23621,N_22762,N_22455);
xor U23622 (N_23622,N_22581,N_22425);
nand U23623 (N_23623,N_22905,N_22662);
nand U23624 (N_23624,N_22437,N_22591);
and U23625 (N_23625,N_22699,N_22487);
xor U23626 (N_23626,N_22266,N_22509);
and U23627 (N_23627,N_22393,N_22301);
or U23628 (N_23628,N_22878,N_22065);
nor U23629 (N_23629,N_22059,N_22810);
and U23630 (N_23630,N_22447,N_22488);
or U23631 (N_23631,N_22235,N_22783);
or U23632 (N_23632,N_22217,N_22876);
or U23633 (N_23633,N_22483,N_22335);
nor U23634 (N_23634,N_22725,N_22681);
xnor U23635 (N_23635,N_22002,N_22410);
xor U23636 (N_23636,N_22369,N_22219);
nand U23637 (N_23637,N_22487,N_22667);
and U23638 (N_23638,N_22727,N_22538);
xnor U23639 (N_23639,N_22935,N_22549);
xor U23640 (N_23640,N_22539,N_22286);
nor U23641 (N_23641,N_22316,N_22078);
nor U23642 (N_23642,N_22130,N_22067);
and U23643 (N_23643,N_22779,N_22301);
xnor U23644 (N_23644,N_22739,N_22554);
and U23645 (N_23645,N_22107,N_22414);
and U23646 (N_23646,N_22536,N_22426);
nor U23647 (N_23647,N_22657,N_22143);
nand U23648 (N_23648,N_22967,N_22081);
nand U23649 (N_23649,N_22679,N_22903);
nand U23650 (N_23650,N_22019,N_22218);
or U23651 (N_23651,N_22607,N_22962);
or U23652 (N_23652,N_22782,N_22627);
or U23653 (N_23653,N_22440,N_22752);
nand U23654 (N_23654,N_22542,N_22160);
nor U23655 (N_23655,N_22113,N_22968);
xnor U23656 (N_23656,N_22161,N_22717);
and U23657 (N_23657,N_22057,N_22534);
or U23658 (N_23658,N_22845,N_22818);
or U23659 (N_23659,N_22718,N_22195);
nor U23660 (N_23660,N_22522,N_22995);
or U23661 (N_23661,N_22506,N_22659);
xor U23662 (N_23662,N_22090,N_22024);
xnor U23663 (N_23663,N_22966,N_22903);
or U23664 (N_23664,N_22594,N_22934);
or U23665 (N_23665,N_22632,N_22311);
xor U23666 (N_23666,N_22861,N_22796);
nor U23667 (N_23667,N_22546,N_22121);
and U23668 (N_23668,N_22225,N_22397);
nand U23669 (N_23669,N_22846,N_22289);
or U23670 (N_23670,N_22240,N_22005);
nor U23671 (N_23671,N_22670,N_22321);
and U23672 (N_23672,N_22700,N_22564);
or U23673 (N_23673,N_22288,N_22017);
nor U23674 (N_23674,N_22791,N_22783);
nor U23675 (N_23675,N_22326,N_22923);
or U23676 (N_23676,N_22605,N_22078);
xnor U23677 (N_23677,N_22300,N_22955);
and U23678 (N_23678,N_22243,N_22385);
or U23679 (N_23679,N_22211,N_22308);
nand U23680 (N_23680,N_22070,N_22829);
xnor U23681 (N_23681,N_22228,N_22493);
and U23682 (N_23682,N_22677,N_22279);
or U23683 (N_23683,N_22309,N_22607);
xnor U23684 (N_23684,N_22028,N_22938);
and U23685 (N_23685,N_22417,N_22528);
nand U23686 (N_23686,N_22164,N_22394);
nand U23687 (N_23687,N_22417,N_22083);
or U23688 (N_23688,N_22776,N_22604);
nor U23689 (N_23689,N_22647,N_22121);
and U23690 (N_23690,N_22719,N_22811);
xor U23691 (N_23691,N_22618,N_22890);
nand U23692 (N_23692,N_22927,N_22292);
or U23693 (N_23693,N_22176,N_22473);
nand U23694 (N_23694,N_22206,N_22394);
and U23695 (N_23695,N_22816,N_22681);
and U23696 (N_23696,N_22750,N_22715);
and U23697 (N_23697,N_22125,N_22537);
or U23698 (N_23698,N_22020,N_22983);
or U23699 (N_23699,N_22254,N_22353);
or U23700 (N_23700,N_22602,N_22451);
nor U23701 (N_23701,N_22594,N_22692);
and U23702 (N_23702,N_22923,N_22943);
nand U23703 (N_23703,N_22389,N_22667);
and U23704 (N_23704,N_22868,N_22888);
nor U23705 (N_23705,N_22033,N_22224);
xnor U23706 (N_23706,N_22945,N_22504);
xnor U23707 (N_23707,N_22701,N_22589);
nand U23708 (N_23708,N_22384,N_22270);
nand U23709 (N_23709,N_22796,N_22615);
xnor U23710 (N_23710,N_22981,N_22602);
and U23711 (N_23711,N_22572,N_22348);
nand U23712 (N_23712,N_22667,N_22871);
nor U23713 (N_23713,N_22699,N_22789);
xnor U23714 (N_23714,N_22302,N_22417);
nand U23715 (N_23715,N_22686,N_22562);
and U23716 (N_23716,N_22674,N_22433);
and U23717 (N_23717,N_22996,N_22145);
xnor U23718 (N_23718,N_22026,N_22878);
xnor U23719 (N_23719,N_22176,N_22605);
nand U23720 (N_23720,N_22125,N_22446);
and U23721 (N_23721,N_22874,N_22299);
nor U23722 (N_23722,N_22082,N_22061);
or U23723 (N_23723,N_22944,N_22707);
or U23724 (N_23724,N_22871,N_22960);
xor U23725 (N_23725,N_22515,N_22047);
nor U23726 (N_23726,N_22684,N_22929);
and U23727 (N_23727,N_22354,N_22633);
nor U23728 (N_23728,N_22228,N_22674);
and U23729 (N_23729,N_22610,N_22007);
or U23730 (N_23730,N_22128,N_22446);
or U23731 (N_23731,N_22263,N_22867);
nand U23732 (N_23732,N_22575,N_22196);
xor U23733 (N_23733,N_22839,N_22641);
or U23734 (N_23734,N_22185,N_22613);
nand U23735 (N_23735,N_22735,N_22290);
xor U23736 (N_23736,N_22750,N_22082);
nor U23737 (N_23737,N_22757,N_22206);
or U23738 (N_23738,N_22608,N_22099);
nand U23739 (N_23739,N_22482,N_22036);
nor U23740 (N_23740,N_22988,N_22443);
and U23741 (N_23741,N_22392,N_22015);
and U23742 (N_23742,N_22683,N_22399);
nor U23743 (N_23743,N_22101,N_22790);
and U23744 (N_23744,N_22287,N_22414);
or U23745 (N_23745,N_22293,N_22930);
xnor U23746 (N_23746,N_22211,N_22331);
and U23747 (N_23747,N_22328,N_22820);
xnor U23748 (N_23748,N_22057,N_22956);
xnor U23749 (N_23749,N_22580,N_22359);
nor U23750 (N_23750,N_22392,N_22522);
and U23751 (N_23751,N_22923,N_22563);
and U23752 (N_23752,N_22577,N_22014);
nor U23753 (N_23753,N_22971,N_22478);
xor U23754 (N_23754,N_22796,N_22179);
and U23755 (N_23755,N_22308,N_22663);
or U23756 (N_23756,N_22531,N_22010);
and U23757 (N_23757,N_22481,N_22286);
or U23758 (N_23758,N_22579,N_22735);
xnor U23759 (N_23759,N_22954,N_22138);
nor U23760 (N_23760,N_22503,N_22832);
nand U23761 (N_23761,N_22456,N_22865);
xnor U23762 (N_23762,N_22391,N_22699);
xor U23763 (N_23763,N_22501,N_22985);
and U23764 (N_23764,N_22745,N_22022);
nand U23765 (N_23765,N_22549,N_22905);
or U23766 (N_23766,N_22759,N_22996);
or U23767 (N_23767,N_22320,N_22469);
nor U23768 (N_23768,N_22319,N_22323);
nand U23769 (N_23769,N_22438,N_22329);
nand U23770 (N_23770,N_22417,N_22543);
xor U23771 (N_23771,N_22080,N_22725);
or U23772 (N_23772,N_22070,N_22459);
nor U23773 (N_23773,N_22861,N_22944);
nor U23774 (N_23774,N_22984,N_22851);
nor U23775 (N_23775,N_22135,N_22296);
or U23776 (N_23776,N_22019,N_22497);
nand U23777 (N_23777,N_22325,N_22841);
nor U23778 (N_23778,N_22284,N_22788);
nand U23779 (N_23779,N_22483,N_22122);
nor U23780 (N_23780,N_22273,N_22943);
nand U23781 (N_23781,N_22047,N_22066);
or U23782 (N_23782,N_22718,N_22875);
nor U23783 (N_23783,N_22572,N_22945);
and U23784 (N_23784,N_22532,N_22419);
nand U23785 (N_23785,N_22575,N_22601);
and U23786 (N_23786,N_22043,N_22853);
nor U23787 (N_23787,N_22648,N_22333);
nand U23788 (N_23788,N_22315,N_22913);
or U23789 (N_23789,N_22030,N_22910);
xor U23790 (N_23790,N_22338,N_22085);
nor U23791 (N_23791,N_22067,N_22673);
and U23792 (N_23792,N_22388,N_22418);
or U23793 (N_23793,N_22819,N_22585);
nand U23794 (N_23794,N_22450,N_22896);
nor U23795 (N_23795,N_22730,N_22358);
or U23796 (N_23796,N_22698,N_22320);
xnor U23797 (N_23797,N_22860,N_22398);
nor U23798 (N_23798,N_22255,N_22137);
or U23799 (N_23799,N_22650,N_22641);
nand U23800 (N_23800,N_22431,N_22403);
nor U23801 (N_23801,N_22635,N_22093);
nand U23802 (N_23802,N_22744,N_22199);
or U23803 (N_23803,N_22344,N_22238);
xnor U23804 (N_23804,N_22018,N_22058);
nand U23805 (N_23805,N_22311,N_22991);
and U23806 (N_23806,N_22326,N_22480);
xor U23807 (N_23807,N_22482,N_22618);
and U23808 (N_23808,N_22852,N_22627);
nor U23809 (N_23809,N_22448,N_22809);
xnor U23810 (N_23810,N_22607,N_22192);
or U23811 (N_23811,N_22102,N_22663);
or U23812 (N_23812,N_22601,N_22712);
or U23813 (N_23813,N_22519,N_22955);
and U23814 (N_23814,N_22830,N_22402);
nor U23815 (N_23815,N_22689,N_22003);
nand U23816 (N_23816,N_22616,N_22336);
xor U23817 (N_23817,N_22141,N_22209);
nor U23818 (N_23818,N_22420,N_22732);
or U23819 (N_23819,N_22541,N_22307);
xnor U23820 (N_23820,N_22898,N_22350);
and U23821 (N_23821,N_22066,N_22343);
nand U23822 (N_23822,N_22081,N_22998);
and U23823 (N_23823,N_22721,N_22958);
xnor U23824 (N_23824,N_22917,N_22222);
and U23825 (N_23825,N_22127,N_22766);
nand U23826 (N_23826,N_22096,N_22772);
and U23827 (N_23827,N_22621,N_22384);
xor U23828 (N_23828,N_22662,N_22309);
xor U23829 (N_23829,N_22845,N_22344);
nor U23830 (N_23830,N_22808,N_22775);
xor U23831 (N_23831,N_22927,N_22796);
or U23832 (N_23832,N_22067,N_22452);
and U23833 (N_23833,N_22656,N_22364);
xor U23834 (N_23834,N_22065,N_22327);
and U23835 (N_23835,N_22608,N_22694);
xor U23836 (N_23836,N_22216,N_22274);
or U23837 (N_23837,N_22137,N_22011);
nor U23838 (N_23838,N_22140,N_22424);
and U23839 (N_23839,N_22303,N_22514);
xnor U23840 (N_23840,N_22487,N_22521);
xnor U23841 (N_23841,N_22525,N_22493);
nand U23842 (N_23842,N_22493,N_22899);
xnor U23843 (N_23843,N_22495,N_22888);
xor U23844 (N_23844,N_22028,N_22117);
nand U23845 (N_23845,N_22242,N_22590);
or U23846 (N_23846,N_22792,N_22580);
nor U23847 (N_23847,N_22695,N_22087);
or U23848 (N_23848,N_22209,N_22122);
nand U23849 (N_23849,N_22938,N_22048);
nand U23850 (N_23850,N_22912,N_22263);
or U23851 (N_23851,N_22139,N_22737);
nand U23852 (N_23852,N_22283,N_22324);
and U23853 (N_23853,N_22752,N_22101);
nor U23854 (N_23854,N_22822,N_22436);
and U23855 (N_23855,N_22315,N_22535);
nor U23856 (N_23856,N_22864,N_22587);
nor U23857 (N_23857,N_22771,N_22583);
nand U23858 (N_23858,N_22675,N_22886);
and U23859 (N_23859,N_22443,N_22818);
and U23860 (N_23860,N_22409,N_22075);
xnor U23861 (N_23861,N_22390,N_22418);
or U23862 (N_23862,N_22489,N_22999);
nor U23863 (N_23863,N_22942,N_22211);
nor U23864 (N_23864,N_22549,N_22159);
or U23865 (N_23865,N_22425,N_22202);
nor U23866 (N_23866,N_22364,N_22836);
and U23867 (N_23867,N_22489,N_22615);
nand U23868 (N_23868,N_22040,N_22655);
or U23869 (N_23869,N_22460,N_22555);
nor U23870 (N_23870,N_22090,N_22495);
xnor U23871 (N_23871,N_22216,N_22097);
xnor U23872 (N_23872,N_22312,N_22904);
xnor U23873 (N_23873,N_22226,N_22326);
nand U23874 (N_23874,N_22796,N_22030);
xor U23875 (N_23875,N_22017,N_22426);
nand U23876 (N_23876,N_22466,N_22435);
nand U23877 (N_23877,N_22683,N_22776);
nand U23878 (N_23878,N_22880,N_22775);
nor U23879 (N_23879,N_22205,N_22831);
and U23880 (N_23880,N_22838,N_22792);
and U23881 (N_23881,N_22154,N_22712);
and U23882 (N_23882,N_22832,N_22626);
nand U23883 (N_23883,N_22508,N_22039);
nor U23884 (N_23884,N_22658,N_22463);
or U23885 (N_23885,N_22327,N_22090);
nand U23886 (N_23886,N_22285,N_22235);
nand U23887 (N_23887,N_22047,N_22372);
nand U23888 (N_23888,N_22200,N_22839);
and U23889 (N_23889,N_22758,N_22746);
nor U23890 (N_23890,N_22704,N_22011);
and U23891 (N_23891,N_22233,N_22886);
and U23892 (N_23892,N_22613,N_22994);
nor U23893 (N_23893,N_22249,N_22812);
nor U23894 (N_23894,N_22066,N_22320);
nand U23895 (N_23895,N_22933,N_22017);
xor U23896 (N_23896,N_22408,N_22513);
xor U23897 (N_23897,N_22327,N_22542);
nor U23898 (N_23898,N_22710,N_22061);
nand U23899 (N_23899,N_22947,N_22040);
nor U23900 (N_23900,N_22848,N_22929);
nand U23901 (N_23901,N_22950,N_22862);
and U23902 (N_23902,N_22179,N_22152);
and U23903 (N_23903,N_22625,N_22372);
nor U23904 (N_23904,N_22205,N_22077);
and U23905 (N_23905,N_22805,N_22708);
and U23906 (N_23906,N_22835,N_22055);
nand U23907 (N_23907,N_22153,N_22241);
nor U23908 (N_23908,N_22790,N_22604);
nor U23909 (N_23909,N_22153,N_22615);
and U23910 (N_23910,N_22817,N_22160);
xnor U23911 (N_23911,N_22835,N_22794);
xor U23912 (N_23912,N_22891,N_22532);
nor U23913 (N_23913,N_22796,N_22147);
or U23914 (N_23914,N_22521,N_22959);
xor U23915 (N_23915,N_22635,N_22782);
nand U23916 (N_23916,N_22834,N_22228);
or U23917 (N_23917,N_22097,N_22348);
nand U23918 (N_23918,N_22450,N_22845);
nand U23919 (N_23919,N_22505,N_22533);
and U23920 (N_23920,N_22934,N_22750);
or U23921 (N_23921,N_22884,N_22151);
xnor U23922 (N_23922,N_22725,N_22110);
xor U23923 (N_23923,N_22825,N_22361);
xor U23924 (N_23924,N_22132,N_22067);
nand U23925 (N_23925,N_22974,N_22693);
or U23926 (N_23926,N_22487,N_22181);
xnor U23927 (N_23927,N_22786,N_22706);
nor U23928 (N_23928,N_22598,N_22501);
nand U23929 (N_23929,N_22522,N_22045);
nand U23930 (N_23930,N_22631,N_22786);
or U23931 (N_23931,N_22534,N_22296);
or U23932 (N_23932,N_22335,N_22466);
nand U23933 (N_23933,N_22356,N_22073);
xor U23934 (N_23934,N_22257,N_22482);
xor U23935 (N_23935,N_22472,N_22777);
xnor U23936 (N_23936,N_22559,N_22492);
nor U23937 (N_23937,N_22536,N_22213);
xor U23938 (N_23938,N_22439,N_22692);
and U23939 (N_23939,N_22305,N_22437);
nor U23940 (N_23940,N_22413,N_22397);
or U23941 (N_23941,N_22556,N_22085);
nor U23942 (N_23942,N_22448,N_22481);
and U23943 (N_23943,N_22961,N_22733);
or U23944 (N_23944,N_22136,N_22757);
and U23945 (N_23945,N_22229,N_22828);
and U23946 (N_23946,N_22404,N_22447);
nor U23947 (N_23947,N_22016,N_22376);
nor U23948 (N_23948,N_22951,N_22324);
nand U23949 (N_23949,N_22910,N_22722);
nor U23950 (N_23950,N_22589,N_22542);
nor U23951 (N_23951,N_22200,N_22409);
xor U23952 (N_23952,N_22997,N_22878);
xor U23953 (N_23953,N_22651,N_22732);
and U23954 (N_23954,N_22984,N_22877);
nand U23955 (N_23955,N_22598,N_22879);
xnor U23956 (N_23956,N_22428,N_22441);
nor U23957 (N_23957,N_22518,N_22094);
nor U23958 (N_23958,N_22866,N_22697);
and U23959 (N_23959,N_22511,N_22396);
nor U23960 (N_23960,N_22612,N_22922);
nand U23961 (N_23961,N_22747,N_22005);
nand U23962 (N_23962,N_22688,N_22329);
nor U23963 (N_23963,N_22748,N_22450);
or U23964 (N_23964,N_22638,N_22281);
and U23965 (N_23965,N_22637,N_22046);
or U23966 (N_23966,N_22094,N_22469);
or U23967 (N_23967,N_22487,N_22555);
nand U23968 (N_23968,N_22226,N_22138);
xor U23969 (N_23969,N_22898,N_22481);
or U23970 (N_23970,N_22618,N_22616);
and U23971 (N_23971,N_22817,N_22411);
nand U23972 (N_23972,N_22899,N_22817);
and U23973 (N_23973,N_22106,N_22976);
or U23974 (N_23974,N_22481,N_22270);
or U23975 (N_23975,N_22001,N_22039);
or U23976 (N_23976,N_22156,N_22120);
or U23977 (N_23977,N_22430,N_22721);
and U23978 (N_23978,N_22514,N_22053);
and U23979 (N_23979,N_22145,N_22867);
xnor U23980 (N_23980,N_22362,N_22107);
nor U23981 (N_23981,N_22171,N_22596);
and U23982 (N_23982,N_22121,N_22070);
xor U23983 (N_23983,N_22237,N_22835);
and U23984 (N_23984,N_22169,N_22122);
nor U23985 (N_23985,N_22589,N_22643);
and U23986 (N_23986,N_22970,N_22348);
or U23987 (N_23987,N_22604,N_22748);
and U23988 (N_23988,N_22412,N_22716);
and U23989 (N_23989,N_22607,N_22097);
nand U23990 (N_23990,N_22090,N_22724);
xnor U23991 (N_23991,N_22003,N_22163);
and U23992 (N_23992,N_22521,N_22107);
and U23993 (N_23993,N_22822,N_22574);
xor U23994 (N_23994,N_22093,N_22570);
nor U23995 (N_23995,N_22925,N_22221);
and U23996 (N_23996,N_22064,N_22049);
xor U23997 (N_23997,N_22643,N_22395);
nand U23998 (N_23998,N_22565,N_22391);
nand U23999 (N_23999,N_22528,N_22699);
or U24000 (N_24000,N_23836,N_23290);
nand U24001 (N_24001,N_23779,N_23778);
and U24002 (N_24002,N_23175,N_23336);
nor U24003 (N_24003,N_23994,N_23472);
nand U24004 (N_24004,N_23435,N_23546);
nand U24005 (N_24005,N_23252,N_23268);
nor U24006 (N_24006,N_23124,N_23273);
nor U24007 (N_24007,N_23674,N_23938);
and U24008 (N_24008,N_23131,N_23105);
and U24009 (N_24009,N_23693,N_23507);
and U24010 (N_24010,N_23888,N_23889);
and U24011 (N_24011,N_23917,N_23303);
or U24012 (N_24012,N_23455,N_23071);
and U24013 (N_24013,N_23618,N_23732);
xor U24014 (N_24014,N_23275,N_23081);
or U24015 (N_24015,N_23774,N_23093);
or U24016 (N_24016,N_23670,N_23390);
xnor U24017 (N_24017,N_23863,N_23680);
xor U24018 (N_24018,N_23285,N_23387);
xnor U24019 (N_24019,N_23091,N_23024);
or U24020 (N_24020,N_23983,N_23521);
xor U24021 (N_24021,N_23001,N_23531);
and U24022 (N_24022,N_23029,N_23254);
and U24023 (N_24023,N_23735,N_23748);
nand U24024 (N_24024,N_23504,N_23788);
nand U24025 (N_24025,N_23960,N_23567);
or U24026 (N_24026,N_23031,N_23980);
or U24027 (N_24027,N_23964,N_23659);
nor U24028 (N_24028,N_23734,N_23032);
nand U24029 (N_24029,N_23054,N_23266);
and U24030 (N_24030,N_23699,N_23761);
xor U24031 (N_24031,N_23347,N_23536);
xnor U24032 (N_24032,N_23775,N_23798);
nor U24033 (N_24033,N_23743,N_23510);
or U24034 (N_24034,N_23467,N_23762);
nor U24035 (N_24035,N_23215,N_23292);
and U24036 (N_24036,N_23700,N_23556);
and U24037 (N_24037,N_23601,N_23664);
nor U24038 (N_24038,N_23607,N_23453);
and U24039 (N_24039,N_23084,N_23030);
and U24040 (N_24040,N_23428,N_23009);
nor U24041 (N_24041,N_23978,N_23391);
and U24042 (N_24042,N_23548,N_23053);
nand U24043 (N_24043,N_23138,N_23544);
and U24044 (N_24044,N_23006,N_23906);
and U24045 (N_24045,N_23865,N_23361);
xnor U24046 (N_24046,N_23140,N_23595);
xor U24047 (N_24047,N_23499,N_23324);
nor U24048 (N_24048,N_23924,N_23702);
nand U24049 (N_24049,N_23620,N_23224);
or U24050 (N_24050,N_23585,N_23394);
nor U24051 (N_24051,N_23474,N_23117);
xnor U24052 (N_24052,N_23401,N_23231);
nor U24053 (N_24053,N_23015,N_23627);
nand U24054 (N_24054,N_23156,N_23405);
and U24055 (N_24055,N_23457,N_23259);
nor U24056 (N_24056,N_23027,N_23979);
nand U24057 (N_24057,N_23223,N_23957);
nor U24058 (N_24058,N_23195,N_23461);
nor U24059 (N_24059,N_23118,N_23250);
or U24060 (N_24060,N_23639,N_23654);
nand U24061 (N_24061,N_23820,N_23602);
nor U24062 (N_24062,N_23817,N_23803);
and U24063 (N_24063,N_23725,N_23039);
nand U24064 (N_24064,N_23711,N_23642);
nor U24065 (N_24065,N_23513,N_23615);
nand U24066 (N_24066,N_23524,N_23534);
nand U24067 (N_24067,N_23814,N_23241);
nor U24068 (N_24068,N_23777,N_23299);
and U24069 (N_24069,N_23959,N_23885);
xnor U24070 (N_24070,N_23806,N_23897);
or U24071 (N_24071,N_23393,N_23306);
and U24072 (N_24072,N_23500,N_23826);
or U24073 (N_24073,N_23272,N_23184);
xor U24074 (N_24074,N_23289,N_23102);
xnor U24075 (N_24075,N_23929,N_23776);
nand U24076 (N_24076,N_23133,N_23831);
nor U24077 (N_24077,N_23695,N_23229);
or U24078 (N_24078,N_23203,N_23416);
xnor U24079 (N_24079,N_23116,N_23878);
nand U24080 (N_24080,N_23846,N_23996);
xor U24081 (N_24081,N_23907,N_23334);
xnor U24082 (N_24082,N_23770,N_23549);
xor U24083 (N_24083,N_23904,N_23284);
nand U24084 (N_24084,N_23017,N_23271);
and U24085 (N_24085,N_23781,N_23600);
nand U24086 (N_24086,N_23819,N_23611);
nand U24087 (N_24087,N_23570,N_23025);
or U24088 (N_24088,N_23976,N_23191);
xnor U24089 (N_24089,N_23095,N_23921);
nor U24090 (N_24090,N_23824,N_23446);
or U24091 (N_24091,N_23818,N_23301);
nand U24092 (N_24092,N_23380,N_23676);
nor U24093 (N_24093,N_23608,N_23562);
xor U24094 (N_24094,N_23715,N_23218);
and U24095 (N_24095,N_23059,N_23640);
xnor U24096 (N_24096,N_23941,N_23211);
nand U24097 (N_24097,N_23645,N_23099);
nor U24098 (N_24098,N_23028,N_23288);
nor U24099 (N_24099,N_23076,N_23316);
nand U24100 (N_24100,N_23760,N_23772);
and U24101 (N_24101,N_23129,N_23167);
nand U24102 (N_24102,N_23657,N_23975);
nor U24103 (N_24103,N_23687,N_23898);
or U24104 (N_24104,N_23731,N_23082);
or U24105 (N_24105,N_23182,N_23368);
nand U24106 (N_24106,N_23243,N_23033);
nand U24107 (N_24107,N_23555,N_23479);
nand U24108 (N_24108,N_23582,N_23858);
xor U24109 (N_24109,N_23940,N_23578);
nand U24110 (N_24110,N_23431,N_23796);
or U24111 (N_24111,N_23718,N_23552);
and U24112 (N_24112,N_23744,N_23988);
nor U24113 (N_24113,N_23945,N_23753);
and U24114 (N_24114,N_23111,N_23438);
nand U24115 (N_24115,N_23739,N_23062);
xor U24116 (N_24116,N_23236,N_23847);
nor U24117 (N_24117,N_23974,N_23330);
xor U24118 (N_24118,N_23297,N_23125);
and U24119 (N_24119,N_23351,N_23142);
nor U24120 (N_24120,N_23650,N_23782);
and U24121 (N_24121,N_23573,N_23327);
or U24122 (N_24122,N_23230,N_23190);
and U24123 (N_24123,N_23557,N_23369);
nand U24124 (N_24124,N_23597,N_23061);
and U24125 (N_24125,N_23646,N_23527);
xor U24126 (N_24126,N_23020,N_23989);
nor U24127 (N_24127,N_23890,N_23870);
and U24128 (N_24128,N_23622,N_23848);
or U24129 (N_24129,N_23247,N_23412);
nor U24130 (N_24130,N_23204,N_23415);
xnor U24131 (N_24131,N_23923,N_23305);
nor U24132 (N_24132,N_23074,N_23644);
nand U24133 (N_24133,N_23649,N_23388);
nand U24134 (N_24134,N_23568,N_23799);
xnor U24135 (N_24135,N_23874,N_23651);
xnor U24136 (N_24136,N_23932,N_23837);
nand U24137 (N_24137,N_23669,N_23379);
and U24138 (N_24138,N_23371,N_23962);
xnor U24139 (N_24139,N_23942,N_23855);
nor U24140 (N_24140,N_23469,N_23356);
xor U24141 (N_24141,N_23026,N_23698);
nand U24142 (N_24142,N_23011,N_23736);
xor U24143 (N_24143,N_23193,N_23311);
or U24144 (N_24144,N_23248,N_23234);
nand U24145 (N_24145,N_23543,N_23764);
nand U24146 (N_24146,N_23496,N_23352);
xnor U24147 (N_24147,N_23358,N_23969);
nand U24148 (N_24148,N_23648,N_23815);
or U24149 (N_24149,N_23127,N_23377);
nor U24150 (N_24150,N_23171,N_23068);
xor U24151 (N_24151,N_23750,N_23309);
nor U24152 (N_24152,N_23905,N_23954);
nand U24153 (N_24153,N_23257,N_23302);
or U24154 (N_24154,N_23842,N_23660);
xor U24155 (N_24155,N_23321,N_23485);
and U24156 (N_24156,N_23196,N_23692);
xor U24157 (N_24157,N_23563,N_23077);
nor U24158 (N_24158,N_23579,N_23008);
xnor U24159 (N_24159,N_23495,N_23227);
or U24160 (N_24160,N_23592,N_23375);
nand U24161 (N_24161,N_23064,N_23366);
and U24162 (N_24162,N_23591,N_23364);
xnor U24163 (N_24163,N_23765,N_23867);
or U24164 (N_24164,N_23294,N_23786);
nand U24165 (N_24165,N_23261,N_23714);
xnor U24166 (N_24166,N_23007,N_23882);
and U24167 (N_24167,N_23681,N_23466);
and U24168 (N_24168,N_23443,N_23862);
or U24169 (N_24169,N_23464,N_23314);
xnor U24170 (N_24170,N_23922,N_23217);
or U24171 (N_24171,N_23427,N_23633);
or U24172 (N_24172,N_23916,N_23569);
nand U24173 (N_24173,N_23547,N_23018);
nand U24174 (N_24174,N_23048,N_23946);
xnor U24175 (N_24175,N_23386,N_23866);
and U24176 (N_24176,N_23235,N_23201);
nand U24177 (N_24177,N_23183,N_23849);
and U24178 (N_24178,N_23448,N_23286);
nor U24179 (N_24179,N_23487,N_23802);
nor U24180 (N_24180,N_23147,N_23838);
xor U24181 (N_24181,N_23130,N_23807);
nor U24182 (N_24182,N_23995,N_23049);
nand U24183 (N_24183,N_23220,N_23345);
nor U24184 (N_24184,N_23139,N_23636);
nor U24185 (N_24185,N_23797,N_23189);
nor U24186 (N_24186,N_23484,N_23035);
nand U24187 (N_24187,N_23566,N_23320);
or U24188 (N_24188,N_23354,N_23086);
nand U24189 (N_24189,N_23409,N_23722);
nand U24190 (N_24190,N_23948,N_23476);
xor U24191 (N_24191,N_23545,N_23926);
and U24192 (N_24192,N_23318,N_23065);
and U24193 (N_24193,N_23766,N_23841);
nand U24194 (N_24194,N_23784,N_23523);
or U24195 (N_24195,N_23165,N_23755);
nor U24196 (N_24196,N_23370,N_23492);
nand U24197 (N_24197,N_23704,N_23073);
nor U24198 (N_24198,N_23844,N_23903);
nand U24199 (N_24199,N_23551,N_23135);
nor U24200 (N_24200,N_23335,N_23637);
or U24201 (N_24201,N_23861,N_23016);
xnor U24202 (N_24202,N_23575,N_23440);
xnor U24203 (N_24203,N_23098,N_23720);
or U24204 (N_24204,N_23791,N_23100);
nor U24205 (N_24205,N_23389,N_23434);
and U24206 (N_24206,N_23221,N_23561);
and U24207 (N_24207,N_23088,N_23756);
or U24208 (N_24208,N_23880,N_23853);
and U24209 (N_24209,N_23280,N_23310);
or U24210 (N_24210,N_23643,N_23696);
nand U24211 (N_24211,N_23613,N_23925);
nand U24212 (N_24212,N_23883,N_23690);
or U24213 (N_24213,N_23331,N_23668);
and U24214 (N_24214,N_23442,N_23589);
xor U24215 (N_24215,N_23933,N_23216);
xor U24216 (N_24216,N_23688,N_23308);
and U24217 (N_24217,N_23603,N_23629);
xor U24218 (N_24218,N_23353,N_23399);
nor U24219 (N_24219,N_23423,N_23329);
or U24220 (N_24220,N_23860,N_23202);
or U24221 (N_24221,N_23955,N_23367);
xor U24222 (N_24222,N_23382,N_23063);
nor U24223 (N_24223,N_23475,N_23768);
xnor U24224 (N_24224,N_23200,N_23460);
nor U24225 (N_24225,N_23708,N_23517);
and U24226 (N_24226,N_23985,N_23881);
xor U24227 (N_24227,N_23827,N_23058);
or U24228 (N_24228,N_23333,N_23868);
nand U24229 (N_24229,N_23101,N_23805);
nand U24230 (N_24230,N_23604,N_23751);
nand U24231 (N_24231,N_23804,N_23228);
nor U24232 (N_24232,N_23478,N_23287);
nor U24233 (N_24233,N_23180,N_23830);
nand U24234 (N_24234,N_23877,N_23021);
nor U24235 (N_24235,N_23928,N_23754);
nor U24236 (N_24236,N_23360,N_23176);
and U24237 (N_24237,N_23539,N_23206);
xnor U24238 (N_24238,N_23205,N_23537);
nand U24239 (N_24239,N_23468,N_23406);
xor U24240 (N_24240,N_23430,N_23214);
nand U24241 (N_24241,N_23576,N_23145);
nand U24242 (N_24242,N_23956,N_23307);
nand U24243 (N_24243,N_23993,N_23584);
and U24244 (N_24244,N_23624,N_23459);
xnor U24245 (N_24245,N_23132,N_23554);
nand U24246 (N_24246,N_23991,N_23533);
nand U24247 (N_24247,N_23936,N_23747);
xor U24248 (N_24248,N_23502,N_23493);
nor U24249 (N_24249,N_23328,N_23322);
and U24250 (N_24250,N_23671,N_23719);
xnor U24251 (N_24251,N_23445,N_23914);
or U24252 (N_24252,N_23835,N_23372);
nor U24253 (N_24253,N_23686,N_23843);
nor U24254 (N_24254,N_23628,N_23871);
nor U24255 (N_24255,N_23652,N_23465);
xor U24256 (N_24256,N_23385,N_23583);
and U24257 (N_24257,N_23408,N_23003);
or U24258 (N_24258,N_23970,N_23298);
nor U24259 (N_24259,N_23509,N_23808);
xor U24260 (N_24260,N_23022,N_23886);
or U24261 (N_24261,N_23490,N_23737);
nand U24262 (N_24262,N_23729,N_23850);
nor U24263 (N_24263,N_23143,N_23717);
nor U24264 (N_24264,N_23733,N_23514);
and U24265 (N_24265,N_23488,N_23365);
and U24266 (N_24266,N_23625,N_23452);
and U24267 (N_24267,N_23056,N_23721);
nor U24268 (N_24268,N_23411,N_23078);
nand U24269 (N_24269,N_23864,N_23152);
or U24270 (N_24270,N_23966,N_23471);
xnor U24271 (N_24271,N_23647,N_23896);
or U24272 (N_24272,N_23398,N_23113);
xnor U24273 (N_24273,N_23034,N_23279);
and U24274 (N_24274,N_23242,N_23179);
nor U24275 (N_24275,N_23051,N_23421);
nor U24276 (N_24276,N_23161,N_23730);
or U24277 (N_24277,N_23363,N_23300);
nor U24278 (N_24278,N_23458,N_23973);
nand U24279 (N_24279,N_23337,N_23256);
or U24280 (N_24280,N_23771,N_23304);
xnor U24281 (N_24281,N_23376,N_23454);
and U24282 (N_24282,N_23107,N_23450);
nor U24283 (N_24283,N_23580,N_23420);
nor U24284 (N_24284,N_23893,N_23128);
xnor U24285 (N_24285,N_23678,N_23278);
and U24286 (N_24286,N_23342,N_23822);
and U24287 (N_24287,N_23588,N_23894);
xor U24288 (N_24288,N_23169,N_23374);
nand U24289 (N_24289,N_23134,N_23968);
nand U24290 (N_24290,N_23505,N_23002);
nor U24291 (N_24291,N_23141,N_23491);
xor U24292 (N_24292,N_23436,N_23901);
nand U24293 (N_24293,N_23809,N_23115);
nor U24294 (N_24294,N_23158,N_23952);
nor U24295 (N_24295,N_23194,N_23323);
xnor U24296 (N_24296,N_23173,N_23689);
nand U24297 (N_24297,N_23931,N_23269);
and U24298 (N_24298,N_23178,N_23172);
nand U24299 (N_24299,N_23825,N_23746);
xor U24300 (N_24300,N_23258,N_23512);
nand U24301 (N_24301,N_23079,N_23682);
and U24302 (N_24302,N_23998,N_23096);
xor U24303 (N_24303,N_23697,N_23168);
nand U24304 (N_24304,N_23723,N_23939);
or U24305 (N_24305,N_23449,N_23947);
nand U24306 (N_24306,N_23293,N_23037);
nor U24307 (N_24307,N_23684,N_23019);
or U24308 (N_24308,N_23759,N_23155);
and U24309 (N_24309,N_23402,N_23137);
xor U24310 (N_24310,N_23012,N_23800);
nand U24311 (N_24311,N_23617,N_23630);
nand U24312 (N_24312,N_23789,N_23341);
nand U24313 (N_24313,N_23456,N_23769);
or U24314 (N_24314,N_23041,N_23535);
nor U24315 (N_24315,N_23444,N_23949);
or U24316 (N_24316,N_23085,N_23550);
nand U24317 (N_24317,N_23587,N_23057);
nor U24318 (N_24318,N_23529,N_23667);
nand U24319 (N_24319,N_23793,N_23373);
xor U24320 (N_24320,N_23508,N_23610);
nand U24321 (N_24321,N_23727,N_23977);
xnor U24322 (N_24322,N_23596,N_23075);
and U24323 (N_24323,N_23277,N_23869);
nand U24324 (N_24324,N_23656,N_23501);
nand U24325 (N_24325,N_23912,N_23199);
and U24326 (N_24326,N_23482,N_23123);
or U24327 (N_24327,N_23150,N_23050);
nor U24328 (N_24328,N_23785,N_23662);
and U24329 (N_24329,N_23823,N_23122);
nand U24330 (N_24330,N_23344,N_23251);
and U24331 (N_24331,N_23516,N_23511);
xnor U24332 (N_24332,N_23419,N_23833);
and U24333 (N_24333,N_23590,N_23665);
and U24334 (N_24334,N_23477,N_23892);
or U24335 (N_24335,N_23349,N_23992);
nand U24336 (N_24336,N_23902,N_23422);
nand U24337 (N_24337,N_23951,N_23738);
or U24338 (N_24338,N_23210,N_23260);
and U24339 (N_24339,N_23972,N_23441);
nand U24340 (N_24340,N_23934,N_23110);
xnor U24341 (N_24341,N_23821,N_23950);
or U24342 (N_24342,N_23767,N_23635);
or U24343 (N_24343,N_23780,N_23362);
or U24344 (N_24344,N_23357,N_23166);
xor U24345 (N_24345,N_23414,N_23560);
nor U24346 (N_24346,N_23963,N_23151);
nand U24347 (N_24347,N_23429,N_23013);
xor U24348 (N_24348,N_23055,N_23565);
xnor U24349 (N_24349,N_23481,N_23913);
or U24350 (N_24350,N_23763,N_23532);
nand U24351 (N_24351,N_23087,N_23873);
nand U24352 (N_24352,N_23162,N_23944);
xnor U24353 (N_24353,N_23232,N_23999);
xnor U24354 (N_24354,N_23103,N_23213);
nor U24355 (N_24355,N_23875,N_23515);
or U24356 (N_24356,N_23599,N_23891);
nand U24357 (N_24357,N_23170,N_23348);
xnor U24358 (N_24358,N_23810,N_23192);
or U24359 (N_24359,N_23813,N_23572);
nor U24360 (N_24360,N_23417,N_23094);
and U24361 (N_24361,N_23919,N_23177);
and U24362 (N_24362,N_23726,N_23834);
or U24363 (N_24363,N_23915,N_23222);
nand U24364 (N_24364,N_23483,N_23619);
and U24365 (N_24365,N_23879,N_23282);
and U24366 (N_24366,N_23840,N_23745);
xor U24367 (N_24367,N_23574,N_23967);
and U24368 (N_24368,N_23558,N_23181);
nand U24369 (N_24369,N_23473,N_23270);
or U24370 (N_24370,N_23710,N_23742);
xnor U24371 (N_24371,N_23355,N_23790);
and U24372 (N_24372,N_23707,N_23070);
xor U24373 (N_24373,N_23519,N_23119);
or U24374 (N_24374,N_23641,N_23854);
nand U24375 (N_24375,N_23226,N_23990);
xnor U24376 (N_24376,N_23326,N_23792);
xnor U24377 (N_24377,N_23672,N_23313);
nand U24378 (N_24378,N_23069,N_23047);
and U24379 (N_24379,N_23981,N_23148);
nand U24380 (N_24380,N_23638,N_23961);
nor U24381 (N_24381,N_23295,N_23185);
nor U24382 (N_24382,N_23586,N_23447);
nand U24383 (N_24383,N_23245,N_23494);
nand U24384 (N_24384,N_23935,N_23887);
or U24385 (N_24385,N_23497,N_23413);
xor U24386 (N_24386,N_23984,N_23403);
nand U24387 (N_24387,N_23439,N_23705);
xor U24388 (N_24388,N_23605,N_23614);
xnor U24389 (N_24389,N_23598,N_23264);
xor U24390 (N_24390,N_23462,N_23042);
and U24391 (N_24391,N_23149,N_23694);
and U24392 (N_24392,N_23564,N_23381);
nor U24393 (N_24393,N_23685,N_23040);
nand U24394 (N_24394,N_23503,N_23263);
xor U24395 (N_24395,N_23498,N_23239);
xor U24396 (N_24396,N_23856,N_23080);
and U24397 (N_24397,N_23899,N_23325);
nor U24398 (N_24398,N_23432,N_23383);
nand U24399 (N_24399,N_23872,N_23724);
or U24400 (N_24400,N_23249,N_23233);
or U24401 (N_24401,N_23090,N_23010);
nor U24402 (N_24402,N_23186,N_23982);
or U24403 (N_24403,N_23312,N_23225);
nand U24404 (N_24404,N_23706,N_23159);
and U24405 (N_24405,N_23400,N_23593);
and U24406 (N_24406,N_23758,N_23174);
and U24407 (N_24407,N_23136,N_23092);
and U24408 (N_24408,N_23197,N_23291);
nor U24409 (N_24409,N_23240,N_23188);
xor U24410 (N_24410,N_23839,N_23000);
xor U24411 (N_24411,N_23106,N_23038);
nand U24412 (N_24412,N_23395,N_23631);
nand U24413 (N_24413,N_23773,N_23317);
nor U24414 (N_24414,N_23319,N_23046);
and U24415 (N_24415,N_23014,N_23609);
nor U24416 (N_24416,N_23208,N_23052);
and U24417 (N_24417,N_23424,N_23023);
and U24418 (N_24418,N_23281,N_23274);
and U24419 (N_24419,N_23626,N_23522);
and U24420 (N_24420,N_23953,N_23392);
nand U24421 (N_24421,N_23691,N_23623);
xnor U24422 (N_24422,N_23121,N_23219);
nor U24423 (N_24423,N_23426,N_23060);
nand U24424 (N_24424,N_23701,N_23920);
or U24425 (N_24425,N_23036,N_23616);
and U24426 (N_24426,N_23378,N_23187);
or U24427 (N_24427,N_23404,N_23816);
and U24428 (N_24428,N_23757,N_23163);
xor U24429 (N_24429,N_23908,N_23930);
and U24430 (N_24430,N_23852,N_23741);
nand U24431 (N_24431,N_23716,N_23713);
and U24432 (N_24432,N_23658,N_23900);
xnor U24433 (N_24433,N_23965,N_23884);
nor U24434 (N_24434,N_23634,N_23709);
and U24435 (N_24435,N_23811,N_23540);
nand U24436 (N_24436,N_23340,N_23787);
nand U24437 (N_24437,N_23104,N_23845);
nor U24438 (N_24438,N_23783,N_23997);
or U24439 (N_24439,N_23752,N_23518);
xnor U24440 (N_24440,N_23359,N_23506);
and U24441 (N_24441,N_23740,N_23910);
and U24442 (N_24442,N_23114,N_23253);
xor U24443 (N_24443,N_23433,N_23343);
and U24444 (N_24444,N_23857,N_23661);
xor U24445 (N_24445,N_23525,N_23801);
or U24446 (N_24446,N_23655,N_23212);
xnor U24447 (N_24447,N_23244,N_23987);
nand U24448 (N_24448,N_23728,N_23004);
or U24449 (N_24449,N_23986,N_23126);
nor U24450 (N_24450,N_23120,N_23238);
nand U24451 (N_24451,N_23683,N_23198);
and U24452 (N_24452,N_23237,N_23267);
or U24453 (N_24453,N_23296,N_23520);
xnor U24454 (N_24454,N_23338,N_23918);
or U24455 (N_24455,N_23209,N_23246);
nor U24456 (N_24456,N_23144,N_23276);
nor U24457 (N_24457,N_23350,N_23146);
and U24458 (N_24458,N_23943,N_23528);
xnor U24459 (N_24459,N_23911,N_23526);
or U24460 (N_24460,N_23971,N_23937);
nand U24461 (N_24461,N_23153,N_23612);
nand U24462 (N_24462,N_23470,N_23425);
or U24463 (N_24463,N_23463,N_23397);
and U24464 (N_24464,N_23089,N_23489);
or U24465 (N_24465,N_23712,N_23437);
xnor U24466 (N_24466,N_23653,N_23571);
nand U24467 (N_24467,N_23679,N_23666);
or U24468 (N_24468,N_23480,N_23541);
nor U24469 (N_24469,N_23339,N_23396);
nor U24470 (N_24470,N_23410,N_23530);
and U24471 (N_24471,N_23581,N_23559);
xor U24472 (N_24472,N_23829,N_23703);
and U24473 (N_24473,N_23109,N_23164);
xnor U24474 (N_24474,N_23486,N_23332);
or U24475 (N_24475,N_23851,N_23832);
and U24476 (N_24476,N_23112,N_23108);
xor U24477 (N_24477,N_23262,N_23384);
or U24478 (N_24478,N_23154,N_23909);
nor U24479 (N_24479,N_23538,N_23160);
nand U24480 (N_24480,N_23828,N_23958);
xor U24481 (N_24481,N_23045,N_23157);
or U24482 (N_24482,N_23553,N_23265);
and U24483 (N_24483,N_23632,N_23749);
nor U24484 (N_24484,N_23005,N_23066);
and U24485 (N_24485,N_23255,N_23044);
and U24486 (N_24486,N_23283,N_23812);
and U24487 (N_24487,N_23663,N_23083);
or U24488 (N_24488,N_23067,N_23097);
or U24489 (N_24489,N_23594,N_23673);
nand U24490 (N_24490,N_23315,N_23606);
xnor U24491 (N_24491,N_23542,N_23072);
nand U24492 (N_24492,N_23407,N_23895);
nor U24493 (N_24493,N_23207,N_23927);
nand U24494 (N_24494,N_23346,N_23677);
xnor U24495 (N_24495,N_23418,N_23621);
nand U24496 (N_24496,N_23043,N_23577);
and U24497 (N_24497,N_23795,N_23876);
nand U24498 (N_24498,N_23794,N_23859);
and U24499 (N_24499,N_23451,N_23675);
xor U24500 (N_24500,N_23323,N_23177);
and U24501 (N_24501,N_23384,N_23430);
and U24502 (N_24502,N_23006,N_23522);
nand U24503 (N_24503,N_23873,N_23161);
nor U24504 (N_24504,N_23302,N_23568);
nand U24505 (N_24505,N_23600,N_23475);
or U24506 (N_24506,N_23541,N_23180);
nor U24507 (N_24507,N_23201,N_23665);
or U24508 (N_24508,N_23535,N_23829);
and U24509 (N_24509,N_23615,N_23034);
and U24510 (N_24510,N_23186,N_23752);
nand U24511 (N_24511,N_23405,N_23476);
xor U24512 (N_24512,N_23958,N_23497);
and U24513 (N_24513,N_23962,N_23780);
or U24514 (N_24514,N_23628,N_23074);
and U24515 (N_24515,N_23410,N_23003);
or U24516 (N_24516,N_23141,N_23929);
xnor U24517 (N_24517,N_23063,N_23779);
or U24518 (N_24518,N_23040,N_23852);
or U24519 (N_24519,N_23872,N_23589);
and U24520 (N_24520,N_23607,N_23109);
xor U24521 (N_24521,N_23608,N_23762);
nand U24522 (N_24522,N_23948,N_23051);
xor U24523 (N_24523,N_23100,N_23321);
nand U24524 (N_24524,N_23069,N_23922);
or U24525 (N_24525,N_23910,N_23241);
xnor U24526 (N_24526,N_23303,N_23189);
xor U24527 (N_24527,N_23348,N_23370);
nor U24528 (N_24528,N_23765,N_23317);
nand U24529 (N_24529,N_23459,N_23217);
xnor U24530 (N_24530,N_23189,N_23322);
xor U24531 (N_24531,N_23666,N_23010);
nor U24532 (N_24532,N_23800,N_23772);
nand U24533 (N_24533,N_23670,N_23728);
and U24534 (N_24534,N_23461,N_23515);
xor U24535 (N_24535,N_23802,N_23449);
and U24536 (N_24536,N_23592,N_23983);
nand U24537 (N_24537,N_23013,N_23488);
and U24538 (N_24538,N_23113,N_23925);
or U24539 (N_24539,N_23689,N_23322);
nor U24540 (N_24540,N_23593,N_23696);
xnor U24541 (N_24541,N_23750,N_23675);
or U24542 (N_24542,N_23945,N_23619);
nand U24543 (N_24543,N_23787,N_23128);
or U24544 (N_24544,N_23337,N_23829);
or U24545 (N_24545,N_23499,N_23129);
xor U24546 (N_24546,N_23897,N_23422);
xnor U24547 (N_24547,N_23930,N_23383);
xor U24548 (N_24548,N_23644,N_23251);
xnor U24549 (N_24549,N_23510,N_23040);
nand U24550 (N_24550,N_23538,N_23355);
and U24551 (N_24551,N_23281,N_23723);
and U24552 (N_24552,N_23687,N_23933);
nor U24553 (N_24553,N_23309,N_23648);
nor U24554 (N_24554,N_23862,N_23340);
and U24555 (N_24555,N_23684,N_23340);
or U24556 (N_24556,N_23979,N_23919);
or U24557 (N_24557,N_23417,N_23543);
or U24558 (N_24558,N_23372,N_23767);
or U24559 (N_24559,N_23997,N_23019);
xor U24560 (N_24560,N_23819,N_23582);
nor U24561 (N_24561,N_23612,N_23578);
and U24562 (N_24562,N_23002,N_23560);
and U24563 (N_24563,N_23173,N_23095);
xor U24564 (N_24564,N_23755,N_23356);
nand U24565 (N_24565,N_23351,N_23772);
and U24566 (N_24566,N_23590,N_23034);
and U24567 (N_24567,N_23304,N_23031);
and U24568 (N_24568,N_23672,N_23323);
nand U24569 (N_24569,N_23252,N_23151);
xor U24570 (N_24570,N_23222,N_23391);
and U24571 (N_24571,N_23200,N_23953);
nor U24572 (N_24572,N_23091,N_23098);
xnor U24573 (N_24573,N_23218,N_23885);
nor U24574 (N_24574,N_23298,N_23040);
or U24575 (N_24575,N_23298,N_23699);
nand U24576 (N_24576,N_23803,N_23182);
and U24577 (N_24577,N_23903,N_23754);
nand U24578 (N_24578,N_23656,N_23578);
nor U24579 (N_24579,N_23311,N_23701);
nor U24580 (N_24580,N_23406,N_23539);
or U24581 (N_24581,N_23827,N_23385);
and U24582 (N_24582,N_23911,N_23261);
nor U24583 (N_24583,N_23970,N_23171);
xnor U24584 (N_24584,N_23176,N_23926);
nand U24585 (N_24585,N_23659,N_23025);
or U24586 (N_24586,N_23061,N_23178);
or U24587 (N_24587,N_23917,N_23937);
nand U24588 (N_24588,N_23094,N_23587);
or U24589 (N_24589,N_23607,N_23269);
nand U24590 (N_24590,N_23000,N_23209);
nand U24591 (N_24591,N_23011,N_23439);
xnor U24592 (N_24592,N_23287,N_23008);
nand U24593 (N_24593,N_23520,N_23961);
nor U24594 (N_24594,N_23338,N_23011);
and U24595 (N_24595,N_23494,N_23830);
nand U24596 (N_24596,N_23400,N_23362);
nand U24597 (N_24597,N_23207,N_23849);
and U24598 (N_24598,N_23414,N_23687);
or U24599 (N_24599,N_23926,N_23398);
or U24600 (N_24600,N_23260,N_23540);
nor U24601 (N_24601,N_23493,N_23016);
and U24602 (N_24602,N_23505,N_23888);
nor U24603 (N_24603,N_23284,N_23180);
nand U24604 (N_24604,N_23735,N_23076);
nor U24605 (N_24605,N_23167,N_23044);
and U24606 (N_24606,N_23926,N_23834);
nand U24607 (N_24607,N_23898,N_23103);
nand U24608 (N_24608,N_23463,N_23262);
xor U24609 (N_24609,N_23993,N_23110);
or U24610 (N_24610,N_23136,N_23567);
nor U24611 (N_24611,N_23394,N_23207);
nand U24612 (N_24612,N_23069,N_23889);
nand U24613 (N_24613,N_23461,N_23171);
and U24614 (N_24614,N_23173,N_23545);
xnor U24615 (N_24615,N_23666,N_23572);
or U24616 (N_24616,N_23992,N_23215);
and U24617 (N_24617,N_23927,N_23974);
nor U24618 (N_24618,N_23553,N_23611);
xnor U24619 (N_24619,N_23314,N_23473);
xor U24620 (N_24620,N_23574,N_23760);
xor U24621 (N_24621,N_23850,N_23730);
and U24622 (N_24622,N_23154,N_23705);
and U24623 (N_24623,N_23896,N_23438);
and U24624 (N_24624,N_23267,N_23056);
and U24625 (N_24625,N_23557,N_23640);
nand U24626 (N_24626,N_23032,N_23688);
nand U24627 (N_24627,N_23134,N_23053);
and U24628 (N_24628,N_23388,N_23286);
nand U24629 (N_24629,N_23354,N_23751);
xnor U24630 (N_24630,N_23077,N_23833);
nand U24631 (N_24631,N_23429,N_23040);
and U24632 (N_24632,N_23628,N_23120);
nor U24633 (N_24633,N_23326,N_23726);
nor U24634 (N_24634,N_23922,N_23323);
or U24635 (N_24635,N_23280,N_23268);
nand U24636 (N_24636,N_23789,N_23430);
and U24637 (N_24637,N_23479,N_23888);
nor U24638 (N_24638,N_23835,N_23819);
nor U24639 (N_24639,N_23044,N_23843);
nand U24640 (N_24640,N_23420,N_23291);
nand U24641 (N_24641,N_23332,N_23431);
nor U24642 (N_24642,N_23288,N_23812);
or U24643 (N_24643,N_23983,N_23331);
or U24644 (N_24644,N_23838,N_23029);
nor U24645 (N_24645,N_23831,N_23360);
nand U24646 (N_24646,N_23205,N_23587);
nor U24647 (N_24647,N_23276,N_23566);
nand U24648 (N_24648,N_23401,N_23321);
nand U24649 (N_24649,N_23261,N_23029);
nor U24650 (N_24650,N_23802,N_23153);
xor U24651 (N_24651,N_23329,N_23891);
nor U24652 (N_24652,N_23256,N_23321);
xor U24653 (N_24653,N_23239,N_23510);
xor U24654 (N_24654,N_23542,N_23242);
nor U24655 (N_24655,N_23683,N_23385);
nor U24656 (N_24656,N_23668,N_23739);
nand U24657 (N_24657,N_23241,N_23966);
and U24658 (N_24658,N_23976,N_23971);
and U24659 (N_24659,N_23009,N_23416);
nor U24660 (N_24660,N_23288,N_23811);
and U24661 (N_24661,N_23050,N_23573);
xor U24662 (N_24662,N_23363,N_23081);
and U24663 (N_24663,N_23165,N_23462);
and U24664 (N_24664,N_23901,N_23738);
or U24665 (N_24665,N_23782,N_23930);
or U24666 (N_24666,N_23658,N_23521);
or U24667 (N_24667,N_23899,N_23977);
nand U24668 (N_24668,N_23671,N_23292);
xnor U24669 (N_24669,N_23968,N_23403);
or U24670 (N_24670,N_23960,N_23335);
xor U24671 (N_24671,N_23472,N_23773);
and U24672 (N_24672,N_23653,N_23263);
nand U24673 (N_24673,N_23202,N_23728);
xor U24674 (N_24674,N_23161,N_23743);
xor U24675 (N_24675,N_23631,N_23083);
and U24676 (N_24676,N_23705,N_23287);
nand U24677 (N_24677,N_23339,N_23591);
and U24678 (N_24678,N_23001,N_23887);
nand U24679 (N_24679,N_23421,N_23251);
or U24680 (N_24680,N_23573,N_23717);
or U24681 (N_24681,N_23262,N_23568);
and U24682 (N_24682,N_23771,N_23983);
nand U24683 (N_24683,N_23384,N_23468);
and U24684 (N_24684,N_23858,N_23823);
nor U24685 (N_24685,N_23602,N_23693);
and U24686 (N_24686,N_23572,N_23281);
xor U24687 (N_24687,N_23767,N_23845);
nand U24688 (N_24688,N_23470,N_23133);
or U24689 (N_24689,N_23908,N_23401);
nand U24690 (N_24690,N_23119,N_23889);
xnor U24691 (N_24691,N_23348,N_23994);
or U24692 (N_24692,N_23968,N_23915);
and U24693 (N_24693,N_23436,N_23374);
and U24694 (N_24694,N_23345,N_23136);
nor U24695 (N_24695,N_23276,N_23699);
xnor U24696 (N_24696,N_23293,N_23471);
or U24697 (N_24697,N_23976,N_23168);
nor U24698 (N_24698,N_23284,N_23679);
nand U24699 (N_24699,N_23816,N_23542);
nand U24700 (N_24700,N_23061,N_23746);
nand U24701 (N_24701,N_23095,N_23346);
nor U24702 (N_24702,N_23828,N_23141);
nor U24703 (N_24703,N_23528,N_23602);
nor U24704 (N_24704,N_23056,N_23793);
xnor U24705 (N_24705,N_23171,N_23992);
or U24706 (N_24706,N_23961,N_23199);
xnor U24707 (N_24707,N_23808,N_23083);
nor U24708 (N_24708,N_23588,N_23787);
xnor U24709 (N_24709,N_23438,N_23152);
nand U24710 (N_24710,N_23547,N_23408);
nand U24711 (N_24711,N_23477,N_23494);
nor U24712 (N_24712,N_23770,N_23539);
xnor U24713 (N_24713,N_23755,N_23256);
and U24714 (N_24714,N_23500,N_23433);
nand U24715 (N_24715,N_23208,N_23463);
nor U24716 (N_24716,N_23163,N_23389);
or U24717 (N_24717,N_23731,N_23798);
nor U24718 (N_24718,N_23399,N_23760);
nand U24719 (N_24719,N_23136,N_23369);
or U24720 (N_24720,N_23715,N_23068);
xnor U24721 (N_24721,N_23336,N_23886);
nor U24722 (N_24722,N_23616,N_23921);
and U24723 (N_24723,N_23006,N_23914);
nand U24724 (N_24724,N_23937,N_23593);
nor U24725 (N_24725,N_23376,N_23658);
nor U24726 (N_24726,N_23174,N_23514);
nand U24727 (N_24727,N_23335,N_23344);
nor U24728 (N_24728,N_23880,N_23283);
nand U24729 (N_24729,N_23674,N_23129);
or U24730 (N_24730,N_23683,N_23772);
nor U24731 (N_24731,N_23787,N_23339);
xnor U24732 (N_24732,N_23073,N_23571);
xnor U24733 (N_24733,N_23146,N_23181);
xor U24734 (N_24734,N_23023,N_23711);
and U24735 (N_24735,N_23427,N_23554);
xnor U24736 (N_24736,N_23307,N_23168);
or U24737 (N_24737,N_23643,N_23906);
and U24738 (N_24738,N_23507,N_23481);
and U24739 (N_24739,N_23275,N_23141);
or U24740 (N_24740,N_23320,N_23970);
nor U24741 (N_24741,N_23312,N_23003);
nor U24742 (N_24742,N_23172,N_23769);
or U24743 (N_24743,N_23666,N_23798);
and U24744 (N_24744,N_23551,N_23085);
nand U24745 (N_24745,N_23034,N_23448);
nand U24746 (N_24746,N_23943,N_23748);
or U24747 (N_24747,N_23824,N_23393);
xnor U24748 (N_24748,N_23972,N_23625);
or U24749 (N_24749,N_23439,N_23177);
or U24750 (N_24750,N_23230,N_23889);
nor U24751 (N_24751,N_23132,N_23486);
and U24752 (N_24752,N_23601,N_23683);
and U24753 (N_24753,N_23592,N_23935);
and U24754 (N_24754,N_23734,N_23145);
nor U24755 (N_24755,N_23734,N_23266);
and U24756 (N_24756,N_23549,N_23086);
nor U24757 (N_24757,N_23980,N_23666);
nor U24758 (N_24758,N_23486,N_23617);
nand U24759 (N_24759,N_23022,N_23247);
nand U24760 (N_24760,N_23982,N_23064);
nand U24761 (N_24761,N_23286,N_23330);
and U24762 (N_24762,N_23357,N_23897);
nand U24763 (N_24763,N_23187,N_23314);
or U24764 (N_24764,N_23306,N_23340);
nand U24765 (N_24765,N_23979,N_23321);
nand U24766 (N_24766,N_23440,N_23817);
nand U24767 (N_24767,N_23159,N_23890);
nand U24768 (N_24768,N_23605,N_23720);
nor U24769 (N_24769,N_23902,N_23612);
and U24770 (N_24770,N_23273,N_23839);
or U24771 (N_24771,N_23100,N_23477);
xnor U24772 (N_24772,N_23707,N_23037);
nand U24773 (N_24773,N_23358,N_23001);
xnor U24774 (N_24774,N_23576,N_23516);
or U24775 (N_24775,N_23448,N_23738);
and U24776 (N_24776,N_23745,N_23088);
xnor U24777 (N_24777,N_23207,N_23720);
or U24778 (N_24778,N_23613,N_23174);
nand U24779 (N_24779,N_23693,N_23585);
and U24780 (N_24780,N_23061,N_23834);
nor U24781 (N_24781,N_23605,N_23531);
nand U24782 (N_24782,N_23647,N_23178);
xor U24783 (N_24783,N_23066,N_23169);
xnor U24784 (N_24784,N_23518,N_23873);
nand U24785 (N_24785,N_23483,N_23075);
or U24786 (N_24786,N_23926,N_23871);
and U24787 (N_24787,N_23361,N_23540);
xnor U24788 (N_24788,N_23144,N_23612);
nand U24789 (N_24789,N_23611,N_23823);
or U24790 (N_24790,N_23911,N_23662);
nand U24791 (N_24791,N_23311,N_23734);
and U24792 (N_24792,N_23663,N_23978);
or U24793 (N_24793,N_23104,N_23087);
nand U24794 (N_24794,N_23606,N_23881);
xor U24795 (N_24795,N_23242,N_23540);
nor U24796 (N_24796,N_23125,N_23427);
xor U24797 (N_24797,N_23613,N_23205);
and U24798 (N_24798,N_23941,N_23901);
nor U24799 (N_24799,N_23673,N_23284);
nand U24800 (N_24800,N_23129,N_23433);
nor U24801 (N_24801,N_23623,N_23019);
and U24802 (N_24802,N_23230,N_23253);
nand U24803 (N_24803,N_23829,N_23669);
or U24804 (N_24804,N_23281,N_23824);
xor U24805 (N_24805,N_23931,N_23534);
nor U24806 (N_24806,N_23973,N_23276);
or U24807 (N_24807,N_23164,N_23414);
nor U24808 (N_24808,N_23846,N_23308);
or U24809 (N_24809,N_23934,N_23200);
nand U24810 (N_24810,N_23932,N_23020);
nand U24811 (N_24811,N_23515,N_23702);
and U24812 (N_24812,N_23311,N_23983);
nor U24813 (N_24813,N_23567,N_23253);
nor U24814 (N_24814,N_23329,N_23771);
xnor U24815 (N_24815,N_23070,N_23040);
and U24816 (N_24816,N_23062,N_23386);
or U24817 (N_24817,N_23067,N_23407);
xnor U24818 (N_24818,N_23929,N_23314);
nor U24819 (N_24819,N_23947,N_23685);
and U24820 (N_24820,N_23734,N_23639);
or U24821 (N_24821,N_23877,N_23225);
and U24822 (N_24822,N_23439,N_23457);
nor U24823 (N_24823,N_23506,N_23715);
nand U24824 (N_24824,N_23827,N_23888);
nor U24825 (N_24825,N_23052,N_23262);
xor U24826 (N_24826,N_23540,N_23681);
nand U24827 (N_24827,N_23865,N_23180);
or U24828 (N_24828,N_23871,N_23642);
xor U24829 (N_24829,N_23357,N_23632);
xnor U24830 (N_24830,N_23213,N_23542);
and U24831 (N_24831,N_23760,N_23911);
nand U24832 (N_24832,N_23508,N_23693);
nor U24833 (N_24833,N_23872,N_23982);
or U24834 (N_24834,N_23223,N_23390);
nor U24835 (N_24835,N_23708,N_23377);
or U24836 (N_24836,N_23563,N_23027);
xnor U24837 (N_24837,N_23804,N_23511);
or U24838 (N_24838,N_23144,N_23223);
nand U24839 (N_24839,N_23570,N_23527);
or U24840 (N_24840,N_23796,N_23157);
nor U24841 (N_24841,N_23517,N_23655);
nor U24842 (N_24842,N_23346,N_23941);
nand U24843 (N_24843,N_23665,N_23280);
xor U24844 (N_24844,N_23039,N_23853);
and U24845 (N_24845,N_23057,N_23256);
nand U24846 (N_24846,N_23896,N_23146);
or U24847 (N_24847,N_23258,N_23124);
xor U24848 (N_24848,N_23441,N_23487);
xnor U24849 (N_24849,N_23504,N_23866);
nor U24850 (N_24850,N_23409,N_23664);
nor U24851 (N_24851,N_23855,N_23444);
and U24852 (N_24852,N_23967,N_23299);
nand U24853 (N_24853,N_23770,N_23598);
xnor U24854 (N_24854,N_23495,N_23237);
or U24855 (N_24855,N_23271,N_23029);
nand U24856 (N_24856,N_23509,N_23258);
or U24857 (N_24857,N_23969,N_23885);
xnor U24858 (N_24858,N_23090,N_23508);
and U24859 (N_24859,N_23947,N_23857);
and U24860 (N_24860,N_23424,N_23384);
and U24861 (N_24861,N_23698,N_23386);
nand U24862 (N_24862,N_23192,N_23763);
and U24863 (N_24863,N_23818,N_23362);
xnor U24864 (N_24864,N_23458,N_23746);
and U24865 (N_24865,N_23749,N_23013);
nand U24866 (N_24866,N_23916,N_23797);
xnor U24867 (N_24867,N_23332,N_23730);
or U24868 (N_24868,N_23251,N_23701);
nand U24869 (N_24869,N_23516,N_23662);
or U24870 (N_24870,N_23358,N_23929);
nand U24871 (N_24871,N_23645,N_23953);
nand U24872 (N_24872,N_23505,N_23869);
xnor U24873 (N_24873,N_23611,N_23562);
xor U24874 (N_24874,N_23827,N_23474);
or U24875 (N_24875,N_23665,N_23176);
or U24876 (N_24876,N_23848,N_23970);
nor U24877 (N_24877,N_23566,N_23078);
and U24878 (N_24878,N_23823,N_23691);
and U24879 (N_24879,N_23938,N_23254);
or U24880 (N_24880,N_23791,N_23702);
nor U24881 (N_24881,N_23144,N_23950);
and U24882 (N_24882,N_23197,N_23569);
nand U24883 (N_24883,N_23070,N_23569);
nand U24884 (N_24884,N_23383,N_23754);
or U24885 (N_24885,N_23701,N_23537);
nor U24886 (N_24886,N_23263,N_23153);
or U24887 (N_24887,N_23415,N_23695);
nand U24888 (N_24888,N_23706,N_23055);
xor U24889 (N_24889,N_23939,N_23674);
xor U24890 (N_24890,N_23807,N_23141);
or U24891 (N_24891,N_23287,N_23388);
or U24892 (N_24892,N_23584,N_23348);
xor U24893 (N_24893,N_23924,N_23067);
nand U24894 (N_24894,N_23130,N_23822);
or U24895 (N_24895,N_23108,N_23259);
nor U24896 (N_24896,N_23496,N_23668);
nand U24897 (N_24897,N_23581,N_23599);
or U24898 (N_24898,N_23080,N_23905);
nor U24899 (N_24899,N_23691,N_23779);
or U24900 (N_24900,N_23653,N_23659);
and U24901 (N_24901,N_23809,N_23389);
and U24902 (N_24902,N_23865,N_23505);
nor U24903 (N_24903,N_23984,N_23918);
and U24904 (N_24904,N_23004,N_23085);
nor U24905 (N_24905,N_23344,N_23818);
or U24906 (N_24906,N_23151,N_23004);
nand U24907 (N_24907,N_23850,N_23557);
and U24908 (N_24908,N_23386,N_23927);
and U24909 (N_24909,N_23757,N_23794);
nor U24910 (N_24910,N_23880,N_23642);
and U24911 (N_24911,N_23400,N_23801);
nor U24912 (N_24912,N_23610,N_23746);
nand U24913 (N_24913,N_23794,N_23484);
nand U24914 (N_24914,N_23703,N_23040);
and U24915 (N_24915,N_23257,N_23277);
xnor U24916 (N_24916,N_23538,N_23356);
and U24917 (N_24917,N_23072,N_23441);
or U24918 (N_24918,N_23695,N_23987);
and U24919 (N_24919,N_23334,N_23314);
or U24920 (N_24920,N_23804,N_23748);
xnor U24921 (N_24921,N_23538,N_23125);
nor U24922 (N_24922,N_23857,N_23030);
xor U24923 (N_24923,N_23779,N_23436);
and U24924 (N_24924,N_23777,N_23560);
or U24925 (N_24925,N_23280,N_23201);
xnor U24926 (N_24926,N_23426,N_23311);
nor U24927 (N_24927,N_23082,N_23018);
xor U24928 (N_24928,N_23339,N_23004);
xnor U24929 (N_24929,N_23935,N_23403);
or U24930 (N_24930,N_23192,N_23491);
or U24931 (N_24931,N_23522,N_23365);
nor U24932 (N_24932,N_23724,N_23044);
nand U24933 (N_24933,N_23292,N_23218);
xnor U24934 (N_24934,N_23374,N_23398);
or U24935 (N_24935,N_23250,N_23819);
nor U24936 (N_24936,N_23736,N_23709);
nor U24937 (N_24937,N_23482,N_23048);
nand U24938 (N_24938,N_23166,N_23486);
nor U24939 (N_24939,N_23186,N_23872);
xnor U24940 (N_24940,N_23717,N_23790);
or U24941 (N_24941,N_23110,N_23570);
xnor U24942 (N_24942,N_23264,N_23329);
nor U24943 (N_24943,N_23348,N_23342);
xor U24944 (N_24944,N_23504,N_23378);
or U24945 (N_24945,N_23261,N_23188);
or U24946 (N_24946,N_23166,N_23103);
or U24947 (N_24947,N_23876,N_23513);
or U24948 (N_24948,N_23271,N_23583);
nor U24949 (N_24949,N_23498,N_23214);
xnor U24950 (N_24950,N_23944,N_23758);
nor U24951 (N_24951,N_23573,N_23397);
or U24952 (N_24952,N_23924,N_23330);
nor U24953 (N_24953,N_23864,N_23551);
nand U24954 (N_24954,N_23470,N_23516);
xor U24955 (N_24955,N_23918,N_23996);
nand U24956 (N_24956,N_23140,N_23364);
xnor U24957 (N_24957,N_23704,N_23366);
or U24958 (N_24958,N_23331,N_23449);
xnor U24959 (N_24959,N_23838,N_23231);
xor U24960 (N_24960,N_23731,N_23900);
or U24961 (N_24961,N_23406,N_23722);
xnor U24962 (N_24962,N_23266,N_23505);
nand U24963 (N_24963,N_23527,N_23892);
xnor U24964 (N_24964,N_23133,N_23997);
nor U24965 (N_24965,N_23702,N_23546);
xnor U24966 (N_24966,N_23925,N_23856);
and U24967 (N_24967,N_23988,N_23365);
xnor U24968 (N_24968,N_23919,N_23867);
nor U24969 (N_24969,N_23554,N_23499);
or U24970 (N_24970,N_23888,N_23053);
xor U24971 (N_24971,N_23169,N_23392);
and U24972 (N_24972,N_23427,N_23380);
xnor U24973 (N_24973,N_23210,N_23424);
nor U24974 (N_24974,N_23016,N_23620);
nor U24975 (N_24975,N_23361,N_23135);
nand U24976 (N_24976,N_23634,N_23232);
or U24977 (N_24977,N_23772,N_23457);
xnor U24978 (N_24978,N_23912,N_23432);
xnor U24979 (N_24979,N_23470,N_23662);
nor U24980 (N_24980,N_23541,N_23441);
and U24981 (N_24981,N_23863,N_23288);
nor U24982 (N_24982,N_23161,N_23883);
nand U24983 (N_24983,N_23933,N_23295);
nand U24984 (N_24984,N_23378,N_23229);
nor U24985 (N_24985,N_23034,N_23416);
xor U24986 (N_24986,N_23654,N_23102);
nand U24987 (N_24987,N_23463,N_23148);
or U24988 (N_24988,N_23323,N_23252);
xnor U24989 (N_24989,N_23852,N_23678);
nand U24990 (N_24990,N_23497,N_23226);
nor U24991 (N_24991,N_23511,N_23226);
or U24992 (N_24992,N_23439,N_23876);
and U24993 (N_24993,N_23270,N_23596);
nand U24994 (N_24994,N_23556,N_23057);
and U24995 (N_24995,N_23626,N_23101);
xnor U24996 (N_24996,N_23666,N_23268);
xnor U24997 (N_24997,N_23142,N_23710);
and U24998 (N_24998,N_23964,N_23918);
and U24999 (N_24999,N_23532,N_23046);
xnor U25000 (N_25000,N_24067,N_24623);
nor U25001 (N_25001,N_24754,N_24040);
nand U25002 (N_25002,N_24625,N_24440);
xor U25003 (N_25003,N_24948,N_24113);
and U25004 (N_25004,N_24962,N_24845);
or U25005 (N_25005,N_24798,N_24468);
nand U25006 (N_25006,N_24816,N_24888);
nand U25007 (N_25007,N_24227,N_24146);
or U25008 (N_25008,N_24240,N_24528);
xor U25009 (N_25009,N_24525,N_24839);
nor U25010 (N_25010,N_24865,N_24426);
nand U25011 (N_25011,N_24870,N_24460);
or U25012 (N_25012,N_24725,N_24813);
nor U25013 (N_25013,N_24297,N_24098);
and U25014 (N_25014,N_24666,N_24614);
xnor U25015 (N_25015,N_24309,N_24521);
xor U25016 (N_25016,N_24230,N_24781);
or U25017 (N_25017,N_24351,N_24716);
nor U25018 (N_25018,N_24689,N_24663);
and U25019 (N_25019,N_24021,N_24852);
or U25020 (N_25020,N_24171,N_24041);
and U25021 (N_25021,N_24779,N_24758);
nand U25022 (N_25022,N_24403,N_24670);
nand U25023 (N_25023,N_24883,N_24286);
nor U25024 (N_25024,N_24767,N_24189);
nor U25025 (N_25025,N_24029,N_24952);
or U25026 (N_25026,N_24488,N_24137);
or U25027 (N_25027,N_24047,N_24081);
nor U25028 (N_25028,N_24773,N_24596);
and U25029 (N_25029,N_24511,N_24943);
nand U25030 (N_25030,N_24919,N_24937);
nand U25031 (N_25031,N_24165,N_24875);
or U25032 (N_25032,N_24369,N_24025);
nand U25033 (N_25033,N_24475,N_24750);
or U25034 (N_25034,N_24885,N_24386);
or U25035 (N_25035,N_24533,N_24751);
or U25036 (N_25036,N_24517,N_24244);
nand U25037 (N_25037,N_24495,N_24008);
nor U25038 (N_25038,N_24539,N_24688);
and U25039 (N_25039,N_24134,N_24616);
nor U25040 (N_25040,N_24748,N_24258);
nor U25041 (N_25041,N_24201,N_24215);
xor U25042 (N_25042,N_24929,N_24967);
or U25043 (N_25043,N_24178,N_24209);
nor U25044 (N_25044,N_24484,N_24994);
nor U25045 (N_25045,N_24062,N_24699);
nand U25046 (N_25046,N_24785,N_24589);
nand U25047 (N_25047,N_24945,N_24043);
or U25048 (N_25048,N_24465,N_24375);
or U25049 (N_25049,N_24551,N_24974);
nor U25050 (N_25050,N_24678,N_24114);
or U25051 (N_25051,N_24195,N_24064);
nand U25052 (N_25052,N_24391,N_24438);
xor U25053 (N_25053,N_24661,N_24708);
and U25054 (N_25054,N_24541,N_24478);
or U25055 (N_25055,N_24420,N_24355);
and U25056 (N_25056,N_24574,N_24556);
nor U25057 (N_25057,N_24103,N_24977);
xor U25058 (N_25058,N_24404,N_24272);
nand U25059 (N_25059,N_24602,N_24190);
nor U25060 (N_25060,N_24612,N_24322);
nor U25061 (N_25061,N_24480,N_24807);
nand U25062 (N_25062,N_24848,N_24712);
xor U25063 (N_25063,N_24173,N_24153);
nand U25064 (N_25064,N_24519,N_24471);
nor U25065 (N_25065,N_24953,N_24808);
nor U25066 (N_25066,N_24193,N_24925);
nand U25067 (N_25067,N_24504,N_24439);
xor U25068 (N_25068,N_24594,N_24859);
xor U25069 (N_25069,N_24547,N_24010);
xor U25070 (N_25070,N_24128,N_24806);
and U25071 (N_25071,N_24166,N_24985);
or U25072 (N_25072,N_24874,N_24986);
and U25073 (N_25073,N_24609,N_24995);
xor U25074 (N_25074,N_24646,N_24879);
or U25075 (N_25075,N_24829,N_24815);
nor U25076 (N_25076,N_24123,N_24847);
nor U25077 (N_25077,N_24109,N_24045);
or U25078 (N_25078,N_24867,N_24301);
nand U25079 (N_25079,N_24409,N_24151);
nand U25080 (N_25080,N_24464,N_24503);
nand U25081 (N_25081,N_24655,N_24685);
xor U25082 (N_25082,N_24431,N_24674);
or U25083 (N_25083,N_24940,N_24778);
or U25084 (N_25084,N_24347,N_24901);
or U25085 (N_25085,N_24833,N_24760);
or U25086 (N_25086,N_24357,N_24882);
nor U25087 (N_25087,N_24631,N_24342);
or U25088 (N_25088,N_24991,N_24690);
nor U25089 (N_25089,N_24555,N_24553);
nand U25090 (N_25090,N_24296,N_24881);
nand U25091 (N_25091,N_24110,N_24142);
or U25092 (N_25092,N_24711,N_24163);
or U25093 (N_25093,N_24115,N_24837);
nand U25094 (N_25094,N_24639,N_24120);
and U25095 (N_25095,N_24963,N_24158);
nor U25096 (N_25096,N_24030,N_24950);
and U25097 (N_25097,N_24263,N_24376);
and U25098 (N_25098,N_24841,N_24621);
xor U25099 (N_25099,N_24695,N_24709);
nor U25100 (N_25100,N_24014,N_24513);
and U25101 (N_25101,N_24105,N_24789);
and U25102 (N_25102,N_24292,N_24753);
nand U25103 (N_25103,N_24942,N_24673);
nand U25104 (N_25104,N_24472,N_24584);
nor U25105 (N_25105,N_24486,N_24518);
nand U25106 (N_25106,N_24020,N_24252);
or U25107 (N_25107,N_24324,N_24824);
and U25108 (N_25108,N_24918,N_24400);
and U25109 (N_25109,N_24065,N_24433);
nor U25110 (N_25110,N_24900,N_24500);
xnor U25111 (N_25111,N_24122,N_24392);
nand U25112 (N_25112,N_24473,N_24580);
or U25113 (N_25113,N_24540,N_24809);
xor U25114 (N_25114,N_24745,N_24117);
nand U25115 (N_25115,N_24566,N_24361);
or U25116 (N_25116,N_24229,N_24761);
or U25117 (N_25117,N_24191,N_24922);
xnor U25118 (N_25118,N_24213,N_24780);
nor U25119 (N_25119,N_24615,N_24279);
and U25120 (N_25120,N_24455,N_24176);
and U25121 (N_25121,N_24184,N_24320);
or U25122 (N_25122,N_24707,N_24493);
xor U25123 (N_25123,N_24838,N_24331);
nand U25124 (N_25124,N_24291,N_24397);
nand U25125 (N_25125,N_24415,N_24659);
nand U25126 (N_25126,N_24572,N_24742);
or U25127 (N_25127,N_24933,N_24759);
or U25128 (N_25128,N_24786,N_24703);
and U25129 (N_25129,N_24335,N_24267);
nor U25130 (N_25130,N_24914,N_24526);
nor U25131 (N_25131,N_24198,N_24763);
and U25132 (N_25132,N_24164,N_24152);
nor U25133 (N_25133,N_24696,N_24731);
and U25134 (N_25134,N_24450,N_24958);
nor U25135 (N_25135,N_24034,N_24293);
or U25136 (N_25136,N_24340,N_24319);
nor U25137 (N_25137,N_24980,N_24474);
and U25138 (N_25138,N_24370,N_24441);
nor U25139 (N_25139,N_24443,N_24532);
and U25140 (N_25140,N_24905,N_24204);
nand U25141 (N_25141,N_24805,N_24633);
nand U25142 (N_25142,N_24315,N_24212);
nand U25143 (N_25143,N_24728,N_24428);
nand U25144 (N_25144,N_24740,N_24636);
and U25145 (N_25145,N_24095,N_24871);
and U25146 (N_25146,N_24048,N_24333);
nand U25147 (N_25147,N_24321,N_24565);
or U25148 (N_25148,N_24920,N_24238);
xor U25149 (N_25149,N_24931,N_24714);
and U25150 (N_25150,N_24070,N_24219);
and U25151 (N_25151,N_24592,N_24573);
and U25152 (N_25152,N_24013,N_24973);
nor U25153 (N_25153,N_24821,N_24372);
xor U25154 (N_25154,N_24393,N_24262);
or U25155 (N_25155,N_24650,N_24956);
or U25156 (N_25156,N_24097,N_24481);
xnor U25157 (N_25157,N_24307,N_24436);
xnor U25158 (N_25158,N_24652,N_24329);
nor U25159 (N_25159,N_24687,N_24924);
nor U25160 (N_25160,N_24700,N_24864);
or U25161 (N_25161,N_24003,N_24583);
nand U25162 (N_25162,N_24358,N_24456);
nand U25163 (N_25163,N_24903,N_24494);
and U25164 (N_25164,N_24089,N_24832);
or U25165 (N_25165,N_24599,N_24776);
xor U25166 (N_25166,N_24162,N_24237);
and U25167 (N_25167,N_24782,N_24463);
nor U25168 (N_25168,N_24039,N_24733);
and U25169 (N_25169,N_24851,N_24457);
or U25170 (N_25170,N_24271,N_24537);
nand U25171 (N_25171,N_24476,N_24298);
or U25172 (N_25172,N_24990,N_24242);
nor U25173 (N_25173,N_24111,N_24591);
and U25174 (N_25174,N_24487,N_24080);
xnor U25175 (N_25175,N_24445,N_24765);
and U25176 (N_25176,N_24529,N_24796);
or U25177 (N_25177,N_24857,N_24660);
nand U25178 (N_25178,N_24314,N_24846);
and U25179 (N_25179,N_24068,N_24453);
or U25180 (N_25180,N_24112,N_24434);
nand U25181 (N_25181,N_24417,N_24414);
or U25182 (N_25182,N_24278,N_24218);
or U25183 (N_25183,N_24777,N_24299);
nor U25184 (N_25184,N_24693,N_24011);
nor U25185 (N_25185,N_24275,N_24647);
nor U25186 (N_25186,N_24266,N_24124);
and U25187 (N_25187,N_24645,N_24288);
and U25188 (N_25188,N_24969,N_24175);
and U25189 (N_25189,N_24934,N_24031);
xor U25190 (N_25190,N_24015,N_24345);
xnor U25191 (N_25191,N_24601,N_24738);
nand U25192 (N_25192,N_24233,N_24531);
and U25193 (N_25193,N_24643,N_24515);
xor U25194 (N_25194,N_24385,N_24603);
xor U25195 (N_25195,N_24447,N_24578);
nand U25196 (N_25196,N_24641,N_24667);
or U25197 (N_25197,N_24160,N_24721);
xor U25198 (N_25198,N_24524,N_24954);
and U25199 (N_25199,N_24087,N_24133);
xnor U25200 (N_25200,N_24657,N_24843);
xor U25201 (N_25201,N_24033,N_24383);
nor U25202 (N_25202,N_24066,N_24886);
nand U25203 (N_25203,N_24125,N_24167);
nand U25204 (N_25204,N_24715,N_24605);
xor U25205 (N_25205,N_24268,N_24828);
and U25206 (N_25206,N_24961,N_24944);
and U25207 (N_25207,N_24069,N_24568);
and U25208 (N_25208,N_24844,N_24390);
nand U25209 (N_25209,N_24817,N_24059);
and U25210 (N_25210,N_24577,N_24235);
xor U25211 (N_25211,N_24516,N_24662);
nand U25212 (N_25212,N_24294,N_24410);
and U25213 (N_25213,N_24698,N_24970);
nand U25214 (N_25214,N_24570,N_24091);
xnor U25215 (N_25215,N_24073,N_24211);
nor U25216 (N_25216,N_24895,N_24979);
nor U25217 (N_25217,N_24527,N_24788);
nor U25218 (N_25218,N_24827,N_24968);
nand U25219 (N_25219,N_24251,N_24199);
and U25220 (N_25220,N_24648,N_24581);
or U25221 (N_25221,N_24339,N_24972);
nor U25222 (N_25222,N_24446,N_24630);
nor U25223 (N_25223,N_24597,N_24156);
xnor U25224 (N_25224,N_24261,N_24717);
xnor U25225 (N_25225,N_24629,N_24022);
nand U25226 (N_25226,N_24228,N_24971);
or U25227 (N_25227,N_24873,N_24334);
xor U25228 (N_25228,N_24395,N_24150);
and U25229 (N_25229,N_24856,N_24260);
nand U25230 (N_25230,N_24326,N_24810);
or U25231 (N_25231,N_24653,N_24889);
nor U25232 (N_25232,N_24665,N_24401);
or U25233 (N_25233,N_24206,N_24382);
xnor U25234 (N_25234,N_24203,N_24935);
or U25235 (N_25235,N_24019,N_24564);
nor U25236 (N_25236,N_24850,N_24510);
and U25237 (N_25237,N_24672,N_24181);
nor U25238 (N_25238,N_24567,N_24202);
nand U25239 (N_25239,N_24530,N_24437);
or U25240 (N_25240,N_24604,N_24380);
xor U25241 (N_25241,N_24042,N_24887);
and U25242 (N_25242,N_24576,N_24939);
or U25243 (N_25243,N_24811,N_24477);
or U25244 (N_25244,N_24100,N_24902);
or U25245 (N_25245,N_24651,N_24136);
or U25246 (N_25246,N_24793,N_24394);
nand U25247 (N_25247,N_24571,N_24543);
and U25248 (N_25248,N_24496,N_24139);
or U25249 (N_25249,N_24752,N_24732);
or U25250 (N_25250,N_24200,N_24622);
xor U25251 (N_25251,N_24444,N_24536);
or U25252 (N_25252,N_24050,N_24960);
xor U25253 (N_25253,N_24017,N_24452);
nor U25254 (N_25254,N_24823,N_24305);
and U25255 (N_25255,N_24966,N_24826);
and U25256 (N_25256,N_24911,N_24989);
nand U25257 (N_25257,N_24220,N_24412);
nand U25258 (N_25258,N_24285,N_24317);
nand U25259 (N_25259,N_24787,N_24144);
and U25260 (N_25260,N_24544,N_24454);
nand U25261 (N_25261,N_24791,N_24469);
xor U25262 (N_25262,N_24627,N_24757);
nor U25263 (N_25263,N_24327,N_24365);
and U25264 (N_25264,N_24044,N_24897);
nand U25265 (N_25265,N_24046,N_24884);
nand U25266 (N_25266,N_24007,N_24722);
and U25267 (N_25267,N_24619,N_24161);
or U25268 (N_25268,N_24637,N_24634);
xnor U25269 (N_25269,N_24702,N_24949);
nand U25270 (N_25270,N_24264,N_24035);
or U25271 (N_25271,N_24729,N_24978);
nand U25272 (N_25272,N_24534,N_24490);
and U25273 (N_25273,N_24726,N_24099);
nand U25274 (N_25274,N_24684,N_24669);
or U25275 (N_25275,N_24277,N_24255);
nand U25276 (N_25276,N_24951,N_24032);
nor U25277 (N_25277,N_24096,N_24304);
xnor U25278 (N_25278,N_24746,N_24877);
and U25279 (N_25279,N_24273,N_24535);
and U25280 (N_25280,N_24483,N_24701);
nor U25281 (N_25281,N_24135,N_24054);
nor U25282 (N_25282,N_24632,N_24938);
nand U25283 (N_25283,N_24074,N_24587);
nor U25284 (N_25284,N_24381,N_24668);
xnor U25285 (N_25285,N_24104,N_24774);
or U25286 (N_25286,N_24155,N_24179);
or U25287 (N_25287,N_24399,N_24502);
nor U25288 (N_25288,N_24367,N_24281);
xor U25289 (N_25289,N_24620,N_24679);
nor U25290 (N_25290,N_24232,N_24613);
or U25291 (N_25291,N_24343,N_24427);
nand U25292 (N_25292,N_24975,N_24253);
and U25293 (N_25293,N_24101,N_24312);
nand U25294 (N_25294,N_24349,N_24554);
xnor U25295 (N_25295,N_24835,N_24718);
nand U25296 (N_25296,N_24308,N_24311);
or U25297 (N_25297,N_24697,N_24461);
nand U25298 (N_25298,N_24545,N_24893);
nand U25299 (N_25299,N_24058,N_24177);
nand U25300 (N_25300,N_24056,N_24224);
nor U25301 (N_25301,N_24507,N_24223);
and U25302 (N_25302,N_24368,N_24790);
nand U25303 (N_25303,N_24143,N_24470);
and U25304 (N_25304,N_24234,N_24004);
or U25305 (N_25305,N_24586,N_24849);
nor U25306 (N_25306,N_24770,N_24585);
nand U25307 (N_25307,N_24520,N_24449);
or U25308 (N_25308,N_24353,N_24231);
xor U25309 (N_25309,N_24820,N_24598);
and U25310 (N_25310,N_24834,N_24140);
nor U25311 (N_25311,N_24055,N_24006);
or U25312 (N_25312,N_24088,N_24141);
and U25313 (N_25313,N_24421,N_24344);
xor U25314 (N_25314,N_24964,N_24860);
xor U25315 (N_25315,N_24996,N_24563);
or U25316 (N_25316,N_24287,N_24723);
or U25317 (N_25317,N_24898,N_24241);
and U25318 (N_25318,N_24378,N_24741);
and U25319 (N_25319,N_24492,N_24027);
xnor U25320 (N_25320,N_24772,N_24280);
and U25321 (N_25321,N_24057,N_24649);
nor U25322 (N_25322,N_24549,N_24270);
xnor U25323 (N_25323,N_24656,N_24318);
nand U25324 (N_25324,N_24559,N_24965);
nand U25325 (N_25325,N_24664,N_24910);
or U25326 (N_25326,N_24710,N_24071);
nor U25327 (N_25327,N_24082,N_24356);
and U25328 (N_25328,N_24051,N_24799);
and U25329 (N_25329,N_24462,N_24691);
or U25330 (N_25330,N_24747,N_24254);
nand U25331 (N_25331,N_24677,N_24768);
or U25332 (N_25332,N_24127,N_24290);
nor U25333 (N_25333,N_24611,N_24131);
and U25334 (N_25334,N_24694,N_24595);
and U25335 (N_25335,N_24466,N_24222);
xor U25336 (N_25336,N_24499,N_24138);
nor U25337 (N_25337,N_24265,N_24947);
xor U25338 (N_25338,N_24498,N_24187);
or U25339 (N_25339,N_24987,N_24946);
xnor U25340 (N_25340,N_24988,N_24430);
nand U25341 (N_25341,N_24398,N_24388);
and U25342 (N_25342,N_24562,N_24245);
or U25343 (N_25343,N_24932,N_24330);
nor U25344 (N_25344,N_24210,N_24997);
and U25345 (N_25345,N_24090,N_24276);
xor U25346 (N_25346,N_24590,N_24917);
and U25347 (N_25347,N_24862,N_24075);
xnor U25348 (N_25348,N_24724,N_24078);
nor U25349 (N_25349,N_24310,N_24217);
and U25350 (N_25350,N_24825,N_24891);
and U25351 (N_25351,N_24274,N_24323);
nor U25352 (N_25352,N_24077,N_24283);
nand U25353 (N_25353,N_24814,N_24797);
nor U25354 (N_25354,N_24755,N_24418);
xnor U25355 (N_25355,N_24121,N_24624);
nand U25356 (N_25356,N_24289,N_24366);
xnor U25357 (N_25357,N_24744,N_24792);
nor U25358 (N_25358,N_24295,N_24955);
nor U25359 (N_25359,N_24675,N_24192);
nand U25360 (N_25360,N_24130,N_24106);
or U25361 (N_25361,N_24569,N_24916);
nor U25362 (N_25362,N_24626,N_24243);
nor U25363 (N_25363,N_24734,N_24681);
xor U25364 (N_25364,N_24159,N_24352);
nand U25365 (N_25365,N_24053,N_24802);
nor U25366 (N_25366,N_24593,N_24557);
nand U25367 (N_25367,N_24442,N_24148);
nor U25368 (N_25368,N_24610,N_24226);
nor U25369 (N_25369,N_24350,N_24561);
and U25370 (N_25370,N_24076,N_24915);
xnor U25371 (N_25371,N_24912,N_24804);
nor U25372 (N_25372,N_24981,N_24558);
nor U25373 (N_25373,N_24923,N_24256);
xor U25374 (N_25374,N_24683,N_24313);
and U25375 (N_25375,N_24467,N_24771);
nand U25376 (N_25376,N_24941,N_24126);
nor U25377 (N_25377,N_24063,N_24482);
xor U25378 (N_25378,N_24154,N_24416);
xnor U25379 (N_25379,N_24435,N_24913);
and U25380 (N_25380,N_24706,N_24384);
nor U25381 (N_25381,N_24107,N_24061);
nor U25382 (N_25382,N_24617,N_24908);
or U25383 (N_25383,N_24016,N_24379);
nand U25384 (N_25384,N_24998,N_24840);
nand U25385 (N_25385,N_24743,N_24546);
nand U25386 (N_25386,N_24085,N_24575);
and U25387 (N_25387,N_24855,N_24406);
nand U25388 (N_25388,N_24364,N_24522);
nand U25389 (N_25389,N_24906,N_24818);
xnor U25390 (N_25390,N_24899,N_24374);
or U25391 (N_25391,N_24506,N_24928);
xnor U25392 (N_25392,N_24079,N_24337);
nor U25393 (N_25393,N_24419,N_24992);
nor U25394 (N_25394,N_24086,N_24197);
nor U25395 (N_25395,N_24719,N_24214);
nor U25396 (N_25396,N_24775,N_24682);
xor U25397 (N_25397,N_24360,N_24982);
nand U25398 (N_25398,N_24373,N_24582);
or U25399 (N_25399,N_24005,N_24239);
nor U25400 (N_25400,N_24028,N_24896);
nor U25401 (N_25401,N_24514,N_24936);
xor U25402 (N_25402,N_24387,N_24560);
nor U25403 (N_25403,N_24550,N_24676);
nor U25404 (N_25404,N_24249,N_24921);
nand U25405 (N_25405,N_24654,N_24842);
xnor U25406 (N_25406,N_24102,N_24092);
and U25407 (N_25407,N_24225,N_24692);
xnor U25408 (N_25408,N_24284,N_24411);
xor U25409 (N_25409,N_24036,N_24306);
or U25410 (N_25410,N_24432,N_24730);
and U25411 (N_25411,N_24812,N_24783);
nor U25412 (N_25412,N_24930,N_24423);
or U25413 (N_25413,N_24926,N_24269);
nand U25414 (N_25414,N_24038,N_24523);
nand U25415 (N_25415,N_24168,N_24145);
xor U25416 (N_25416,N_24188,N_24858);
nor U25417 (N_25417,N_24705,N_24854);
nor U25418 (N_25418,N_24316,N_24861);
xor U25419 (N_25419,N_24282,N_24425);
and U25420 (N_25420,N_24907,N_24332);
or U25421 (N_25421,N_24377,N_24037);
xor U25422 (N_25422,N_24491,N_24853);
nand U25423 (N_25423,N_24894,N_24300);
nor U25424 (N_25424,N_24194,N_24756);
and U25425 (N_25425,N_24408,N_24868);
and U25426 (N_25426,N_24083,N_24250);
nand U25427 (N_25427,N_24246,N_24094);
nand U25428 (N_25428,N_24644,N_24248);
and U25429 (N_25429,N_24405,N_24303);
nor U25430 (N_25430,N_24422,N_24221);
xnor U25431 (N_25431,N_24800,N_24459);
and U25432 (N_25432,N_24640,N_24764);
xnor U25433 (N_25433,N_24671,N_24402);
xor U25434 (N_25434,N_24129,N_24512);
or U25435 (N_25435,N_24362,N_24749);
nand U25436 (N_25436,N_24739,N_24371);
nand U25437 (N_25437,N_24658,N_24170);
xnor U25438 (N_25438,N_24052,N_24588);
xnor U25439 (N_25439,N_24119,N_24993);
or U25440 (N_25440,N_24205,N_24208);
nor U25441 (N_25441,N_24999,N_24132);
xnor U25442 (N_25442,N_24257,N_24359);
and U25443 (N_25443,N_24023,N_24009);
nor U25444 (N_25444,N_24769,N_24822);
xor U25445 (N_25445,N_24424,N_24720);
nand U25446 (N_25446,N_24762,N_24346);
and U25447 (N_25447,N_24766,N_24169);
or U25448 (N_25448,N_24451,N_24325);
or U25449 (N_25449,N_24892,N_24983);
nor U25450 (N_25450,N_24348,N_24863);
xor U25451 (N_25451,N_24976,N_24338);
and U25452 (N_25452,N_24084,N_24328);
or U25453 (N_25453,N_24784,N_24407);
or U25454 (N_25454,N_24413,N_24819);
or U25455 (N_25455,N_24341,N_24497);
or U25456 (N_25456,N_24904,N_24542);
nand U25457 (N_25457,N_24302,N_24429);
xor U25458 (N_25458,N_24116,N_24927);
nand U25459 (N_25459,N_24485,N_24890);
or U25460 (N_25460,N_24149,N_24183);
or U25461 (N_25461,N_24600,N_24866);
or U25462 (N_25462,N_24354,N_24869);
nor U25463 (N_25463,N_24207,N_24458);
nand U25464 (N_25464,N_24185,N_24489);
and U25465 (N_25465,N_24735,N_24638);
nand U25466 (N_25466,N_24247,N_24736);
and U25467 (N_25467,N_24336,N_24093);
nor U25468 (N_25468,N_24060,N_24108);
xor U25469 (N_25469,N_24727,N_24795);
and U25470 (N_25470,N_24216,N_24831);
nand U25471 (N_25471,N_24180,N_24579);
xnor U25472 (N_25472,N_24552,N_24801);
or U25473 (N_25473,N_24172,N_24878);
and U25474 (N_25474,N_24836,N_24396);
nor U25475 (N_25475,N_24024,N_24049);
and U25476 (N_25476,N_24002,N_24236);
nand U25477 (N_25477,N_24876,N_24196);
nor U25478 (N_25478,N_24872,N_24001);
nand U25479 (N_25479,N_24501,N_24880);
nor U25480 (N_25480,N_24147,N_24538);
or U25481 (N_25481,N_24363,N_24389);
or U25482 (N_25482,N_24157,N_24909);
nand U25483 (N_25483,N_24635,N_24704);
and U25484 (N_25484,N_24713,N_24072);
nand U25485 (N_25485,N_24182,N_24642);
nor U25486 (N_25486,N_24606,N_24505);
nand U25487 (N_25487,N_24686,N_24259);
xnor U25488 (N_25488,N_24957,N_24508);
or U25489 (N_25489,N_24479,N_24509);
nor U25490 (N_25490,N_24680,N_24628);
and U25491 (N_25491,N_24012,N_24026);
nor U25492 (N_25492,N_24018,N_24174);
or U25493 (N_25493,N_24803,N_24794);
or U25494 (N_25494,N_24607,N_24118);
nand U25495 (N_25495,N_24737,N_24618);
nand U25496 (N_25496,N_24186,N_24608);
nand U25497 (N_25497,N_24959,N_24984);
or U25498 (N_25498,N_24830,N_24548);
or U25499 (N_25499,N_24000,N_24448);
xor U25500 (N_25500,N_24696,N_24643);
and U25501 (N_25501,N_24280,N_24766);
nand U25502 (N_25502,N_24305,N_24005);
and U25503 (N_25503,N_24795,N_24462);
xnor U25504 (N_25504,N_24905,N_24449);
and U25505 (N_25505,N_24854,N_24072);
or U25506 (N_25506,N_24866,N_24468);
nor U25507 (N_25507,N_24426,N_24789);
nor U25508 (N_25508,N_24384,N_24174);
nand U25509 (N_25509,N_24054,N_24612);
or U25510 (N_25510,N_24814,N_24971);
and U25511 (N_25511,N_24619,N_24071);
xor U25512 (N_25512,N_24184,N_24609);
and U25513 (N_25513,N_24363,N_24269);
and U25514 (N_25514,N_24427,N_24797);
xnor U25515 (N_25515,N_24191,N_24193);
xor U25516 (N_25516,N_24993,N_24928);
or U25517 (N_25517,N_24118,N_24724);
nand U25518 (N_25518,N_24058,N_24879);
xor U25519 (N_25519,N_24042,N_24028);
or U25520 (N_25520,N_24112,N_24448);
or U25521 (N_25521,N_24249,N_24382);
nor U25522 (N_25522,N_24215,N_24803);
or U25523 (N_25523,N_24326,N_24627);
xnor U25524 (N_25524,N_24746,N_24039);
nor U25525 (N_25525,N_24761,N_24094);
nand U25526 (N_25526,N_24110,N_24317);
xor U25527 (N_25527,N_24405,N_24703);
nand U25528 (N_25528,N_24102,N_24363);
xor U25529 (N_25529,N_24810,N_24207);
xor U25530 (N_25530,N_24811,N_24197);
or U25531 (N_25531,N_24121,N_24001);
or U25532 (N_25532,N_24968,N_24522);
or U25533 (N_25533,N_24883,N_24981);
and U25534 (N_25534,N_24264,N_24839);
or U25535 (N_25535,N_24329,N_24544);
or U25536 (N_25536,N_24231,N_24934);
or U25537 (N_25537,N_24927,N_24659);
nor U25538 (N_25538,N_24102,N_24636);
nand U25539 (N_25539,N_24837,N_24998);
nor U25540 (N_25540,N_24236,N_24388);
nor U25541 (N_25541,N_24499,N_24747);
xnor U25542 (N_25542,N_24258,N_24350);
xor U25543 (N_25543,N_24274,N_24220);
nor U25544 (N_25544,N_24703,N_24991);
xor U25545 (N_25545,N_24183,N_24077);
nor U25546 (N_25546,N_24102,N_24156);
nand U25547 (N_25547,N_24033,N_24643);
nand U25548 (N_25548,N_24454,N_24697);
or U25549 (N_25549,N_24899,N_24754);
and U25550 (N_25550,N_24467,N_24505);
and U25551 (N_25551,N_24022,N_24628);
or U25552 (N_25552,N_24993,N_24516);
xor U25553 (N_25553,N_24454,N_24260);
nand U25554 (N_25554,N_24692,N_24189);
xnor U25555 (N_25555,N_24229,N_24732);
or U25556 (N_25556,N_24788,N_24347);
and U25557 (N_25557,N_24877,N_24465);
nor U25558 (N_25558,N_24878,N_24543);
and U25559 (N_25559,N_24186,N_24142);
xor U25560 (N_25560,N_24613,N_24803);
nor U25561 (N_25561,N_24129,N_24985);
xnor U25562 (N_25562,N_24512,N_24151);
and U25563 (N_25563,N_24821,N_24922);
nand U25564 (N_25564,N_24049,N_24818);
nor U25565 (N_25565,N_24901,N_24458);
xor U25566 (N_25566,N_24164,N_24922);
or U25567 (N_25567,N_24506,N_24881);
and U25568 (N_25568,N_24820,N_24222);
and U25569 (N_25569,N_24584,N_24947);
nand U25570 (N_25570,N_24527,N_24045);
nand U25571 (N_25571,N_24487,N_24258);
nor U25572 (N_25572,N_24089,N_24324);
nand U25573 (N_25573,N_24822,N_24653);
nand U25574 (N_25574,N_24426,N_24991);
nand U25575 (N_25575,N_24395,N_24047);
nand U25576 (N_25576,N_24925,N_24982);
nand U25577 (N_25577,N_24156,N_24357);
xnor U25578 (N_25578,N_24551,N_24645);
xnor U25579 (N_25579,N_24422,N_24180);
and U25580 (N_25580,N_24695,N_24217);
nor U25581 (N_25581,N_24266,N_24618);
and U25582 (N_25582,N_24776,N_24192);
nor U25583 (N_25583,N_24631,N_24480);
and U25584 (N_25584,N_24827,N_24457);
or U25585 (N_25585,N_24656,N_24268);
or U25586 (N_25586,N_24298,N_24067);
or U25587 (N_25587,N_24326,N_24069);
nand U25588 (N_25588,N_24598,N_24587);
nand U25589 (N_25589,N_24715,N_24978);
and U25590 (N_25590,N_24998,N_24926);
nand U25591 (N_25591,N_24477,N_24340);
nand U25592 (N_25592,N_24425,N_24442);
xnor U25593 (N_25593,N_24867,N_24126);
nand U25594 (N_25594,N_24661,N_24433);
nor U25595 (N_25595,N_24488,N_24084);
xnor U25596 (N_25596,N_24751,N_24635);
nand U25597 (N_25597,N_24624,N_24857);
or U25598 (N_25598,N_24419,N_24380);
and U25599 (N_25599,N_24732,N_24337);
nand U25600 (N_25600,N_24725,N_24587);
or U25601 (N_25601,N_24928,N_24018);
nor U25602 (N_25602,N_24822,N_24764);
or U25603 (N_25603,N_24875,N_24271);
or U25604 (N_25604,N_24138,N_24974);
xor U25605 (N_25605,N_24467,N_24914);
or U25606 (N_25606,N_24221,N_24643);
xor U25607 (N_25607,N_24391,N_24877);
or U25608 (N_25608,N_24756,N_24774);
or U25609 (N_25609,N_24169,N_24082);
xnor U25610 (N_25610,N_24712,N_24998);
nor U25611 (N_25611,N_24981,N_24596);
nor U25612 (N_25612,N_24264,N_24871);
and U25613 (N_25613,N_24911,N_24721);
xor U25614 (N_25614,N_24177,N_24523);
and U25615 (N_25615,N_24227,N_24772);
or U25616 (N_25616,N_24556,N_24396);
xnor U25617 (N_25617,N_24521,N_24842);
nor U25618 (N_25618,N_24485,N_24878);
xor U25619 (N_25619,N_24889,N_24212);
or U25620 (N_25620,N_24447,N_24939);
nand U25621 (N_25621,N_24741,N_24757);
nand U25622 (N_25622,N_24616,N_24186);
nor U25623 (N_25623,N_24757,N_24206);
or U25624 (N_25624,N_24895,N_24806);
nor U25625 (N_25625,N_24820,N_24149);
xnor U25626 (N_25626,N_24948,N_24480);
and U25627 (N_25627,N_24097,N_24792);
and U25628 (N_25628,N_24251,N_24678);
nor U25629 (N_25629,N_24361,N_24835);
xor U25630 (N_25630,N_24729,N_24615);
or U25631 (N_25631,N_24002,N_24756);
nor U25632 (N_25632,N_24299,N_24915);
xnor U25633 (N_25633,N_24733,N_24318);
nor U25634 (N_25634,N_24262,N_24211);
xor U25635 (N_25635,N_24537,N_24472);
nor U25636 (N_25636,N_24033,N_24950);
and U25637 (N_25637,N_24879,N_24545);
nand U25638 (N_25638,N_24210,N_24694);
or U25639 (N_25639,N_24799,N_24330);
nor U25640 (N_25640,N_24352,N_24645);
xor U25641 (N_25641,N_24362,N_24969);
nand U25642 (N_25642,N_24332,N_24289);
xnor U25643 (N_25643,N_24369,N_24641);
or U25644 (N_25644,N_24317,N_24899);
and U25645 (N_25645,N_24258,N_24791);
xor U25646 (N_25646,N_24806,N_24045);
or U25647 (N_25647,N_24838,N_24224);
nand U25648 (N_25648,N_24218,N_24870);
nor U25649 (N_25649,N_24403,N_24107);
xor U25650 (N_25650,N_24101,N_24376);
nor U25651 (N_25651,N_24730,N_24820);
and U25652 (N_25652,N_24485,N_24161);
or U25653 (N_25653,N_24648,N_24043);
nand U25654 (N_25654,N_24312,N_24546);
nand U25655 (N_25655,N_24868,N_24829);
nor U25656 (N_25656,N_24864,N_24129);
nor U25657 (N_25657,N_24889,N_24114);
nor U25658 (N_25658,N_24251,N_24856);
and U25659 (N_25659,N_24481,N_24290);
and U25660 (N_25660,N_24330,N_24779);
xnor U25661 (N_25661,N_24773,N_24614);
and U25662 (N_25662,N_24252,N_24491);
nand U25663 (N_25663,N_24025,N_24907);
or U25664 (N_25664,N_24946,N_24879);
nor U25665 (N_25665,N_24952,N_24056);
xor U25666 (N_25666,N_24602,N_24026);
nand U25667 (N_25667,N_24440,N_24093);
or U25668 (N_25668,N_24840,N_24412);
or U25669 (N_25669,N_24061,N_24159);
nor U25670 (N_25670,N_24407,N_24940);
or U25671 (N_25671,N_24990,N_24430);
xor U25672 (N_25672,N_24841,N_24819);
nor U25673 (N_25673,N_24098,N_24241);
and U25674 (N_25674,N_24853,N_24298);
or U25675 (N_25675,N_24018,N_24726);
nand U25676 (N_25676,N_24131,N_24046);
or U25677 (N_25677,N_24151,N_24742);
and U25678 (N_25678,N_24540,N_24876);
or U25679 (N_25679,N_24096,N_24539);
and U25680 (N_25680,N_24668,N_24179);
and U25681 (N_25681,N_24904,N_24117);
nor U25682 (N_25682,N_24765,N_24629);
or U25683 (N_25683,N_24310,N_24247);
xnor U25684 (N_25684,N_24709,N_24718);
or U25685 (N_25685,N_24659,N_24441);
and U25686 (N_25686,N_24803,N_24462);
xor U25687 (N_25687,N_24580,N_24998);
nand U25688 (N_25688,N_24150,N_24017);
and U25689 (N_25689,N_24692,N_24150);
xor U25690 (N_25690,N_24610,N_24836);
nand U25691 (N_25691,N_24934,N_24801);
nand U25692 (N_25692,N_24774,N_24424);
and U25693 (N_25693,N_24292,N_24328);
or U25694 (N_25694,N_24758,N_24449);
nor U25695 (N_25695,N_24814,N_24458);
and U25696 (N_25696,N_24642,N_24087);
xnor U25697 (N_25697,N_24658,N_24069);
and U25698 (N_25698,N_24091,N_24126);
xor U25699 (N_25699,N_24179,N_24216);
or U25700 (N_25700,N_24050,N_24396);
xor U25701 (N_25701,N_24422,N_24155);
xor U25702 (N_25702,N_24722,N_24030);
or U25703 (N_25703,N_24262,N_24927);
and U25704 (N_25704,N_24422,N_24017);
and U25705 (N_25705,N_24375,N_24126);
and U25706 (N_25706,N_24917,N_24950);
and U25707 (N_25707,N_24444,N_24337);
nand U25708 (N_25708,N_24631,N_24401);
nor U25709 (N_25709,N_24355,N_24635);
or U25710 (N_25710,N_24176,N_24621);
nand U25711 (N_25711,N_24196,N_24729);
or U25712 (N_25712,N_24784,N_24218);
nand U25713 (N_25713,N_24145,N_24932);
xnor U25714 (N_25714,N_24613,N_24320);
or U25715 (N_25715,N_24994,N_24614);
or U25716 (N_25716,N_24105,N_24943);
xor U25717 (N_25717,N_24917,N_24075);
xor U25718 (N_25718,N_24514,N_24611);
nand U25719 (N_25719,N_24047,N_24848);
nor U25720 (N_25720,N_24770,N_24418);
xor U25721 (N_25721,N_24796,N_24580);
or U25722 (N_25722,N_24484,N_24239);
xnor U25723 (N_25723,N_24630,N_24295);
nor U25724 (N_25724,N_24165,N_24163);
xor U25725 (N_25725,N_24047,N_24584);
nand U25726 (N_25726,N_24411,N_24671);
and U25727 (N_25727,N_24982,N_24384);
nand U25728 (N_25728,N_24677,N_24415);
or U25729 (N_25729,N_24581,N_24964);
xor U25730 (N_25730,N_24466,N_24640);
or U25731 (N_25731,N_24213,N_24264);
xor U25732 (N_25732,N_24473,N_24579);
or U25733 (N_25733,N_24367,N_24094);
xor U25734 (N_25734,N_24117,N_24915);
nand U25735 (N_25735,N_24654,N_24551);
nor U25736 (N_25736,N_24021,N_24404);
nand U25737 (N_25737,N_24875,N_24247);
nor U25738 (N_25738,N_24579,N_24765);
nor U25739 (N_25739,N_24583,N_24566);
and U25740 (N_25740,N_24146,N_24625);
and U25741 (N_25741,N_24852,N_24627);
nor U25742 (N_25742,N_24156,N_24943);
or U25743 (N_25743,N_24428,N_24108);
nand U25744 (N_25744,N_24866,N_24195);
nor U25745 (N_25745,N_24782,N_24798);
xnor U25746 (N_25746,N_24763,N_24768);
xor U25747 (N_25747,N_24596,N_24869);
nand U25748 (N_25748,N_24306,N_24854);
and U25749 (N_25749,N_24407,N_24564);
or U25750 (N_25750,N_24874,N_24327);
xor U25751 (N_25751,N_24399,N_24347);
nor U25752 (N_25752,N_24431,N_24855);
or U25753 (N_25753,N_24494,N_24896);
nor U25754 (N_25754,N_24295,N_24862);
or U25755 (N_25755,N_24539,N_24484);
nor U25756 (N_25756,N_24041,N_24507);
nand U25757 (N_25757,N_24347,N_24786);
and U25758 (N_25758,N_24060,N_24242);
nand U25759 (N_25759,N_24317,N_24785);
or U25760 (N_25760,N_24466,N_24601);
nor U25761 (N_25761,N_24570,N_24668);
nand U25762 (N_25762,N_24814,N_24507);
or U25763 (N_25763,N_24367,N_24899);
xor U25764 (N_25764,N_24766,N_24525);
or U25765 (N_25765,N_24781,N_24098);
nand U25766 (N_25766,N_24253,N_24520);
and U25767 (N_25767,N_24858,N_24389);
and U25768 (N_25768,N_24517,N_24195);
and U25769 (N_25769,N_24708,N_24655);
nor U25770 (N_25770,N_24518,N_24541);
or U25771 (N_25771,N_24893,N_24618);
nor U25772 (N_25772,N_24921,N_24636);
nand U25773 (N_25773,N_24574,N_24315);
nor U25774 (N_25774,N_24809,N_24730);
or U25775 (N_25775,N_24188,N_24221);
nand U25776 (N_25776,N_24470,N_24894);
and U25777 (N_25777,N_24190,N_24441);
and U25778 (N_25778,N_24618,N_24674);
nand U25779 (N_25779,N_24254,N_24281);
and U25780 (N_25780,N_24217,N_24842);
nand U25781 (N_25781,N_24453,N_24586);
or U25782 (N_25782,N_24338,N_24699);
or U25783 (N_25783,N_24704,N_24254);
or U25784 (N_25784,N_24451,N_24187);
nand U25785 (N_25785,N_24000,N_24566);
and U25786 (N_25786,N_24177,N_24760);
nand U25787 (N_25787,N_24274,N_24653);
xnor U25788 (N_25788,N_24607,N_24580);
or U25789 (N_25789,N_24486,N_24223);
nor U25790 (N_25790,N_24845,N_24321);
and U25791 (N_25791,N_24800,N_24478);
xor U25792 (N_25792,N_24102,N_24572);
or U25793 (N_25793,N_24152,N_24318);
nand U25794 (N_25794,N_24486,N_24610);
xor U25795 (N_25795,N_24841,N_24812);
or U25796 (N_25796,N_24279,N_24649);
xor U25797 (N_25797,N_24270,N_24056);
nand U25798 (N_25798,N_24324,N_24392);
nor U25799 (N_25799,N_24885,N_24381);
or U25800 (N_25800,N_24706,N_24979);
or U25801 (N_25801,N_24870,N_24265);
xnor U25802 (N_25802,N_24062,N_24013);
xnor U25803 (N_25803,N_24549,N_24776);
xor U25804 (N_25804,N_24920,N_24234);
nor U25805 (N_25805,N_24451,N_24495);
xnor U25806 (N_25806,N_24213,N_24562);
and U25807 (N_25807,N_24340,N_24492);
and U25808 (N_25808,N_24784,N_24510);
nor U25809 (N_25809,N_24376,N_24756);
or U25810 (N_25810,N_24477,N_24024);
xor U25811 (N_25811,N_24120,N_24380);
and U25812 (N_25812,N_24855,N_24593);
and U25813 (N_25813,N_24865,N_24405);
nor U25814 (N_25814,N_24919,N_24143);
nor U25815 (N_25815,N_24426,N_24147);
or U25816 (N_25816,N_24149,N_24144);
and U25817 (N_25817,N_24632,N_24810);
nand U25818 (N_25818,N_24185,N_24236);
xor U25819 (N_25819,N_24491,N_24476);
or U25820 (N_25820,N_24469,N_24586);
and U25821 (N_25821,N_24204,N_24108);
xnor U25822 (N_25822,N_24110,N_24880);
xnor U25823 (N_25823,N_24031,N_24455);
xor U25824 (N_25824,N_24581,N_24069);
or U25825 (N_25825,N_24207,N_24656);
nand U25826 (N_25826,N_24141,N_24545);
xor U25827 (N_25827,N_24424,N_24559);
nor U25828 (N_25828,N_24131,N_24677);
xnor U25829 (N_25829,N_24004,N_24151);
or U25830 (N_25830,N_24079,N_24935);
nand U25831 (N_25831,N_24970,N_24354);
and U25832 (N_25832,N_24641,N_24709);
and U25833 (N_25833,N_24586,N_24148);
xor U25834 (N_25834,N_24106,N_24564);
and U25835 (N_25835,N_24167,N_24033);
nand U25836 (N_25836,N_24326,N_24454);
xor U25837 (N_25837,N_24590,N_24346);
and U25838 (N_25838,N_24214,N_24251);
xor U25839 (N_25839,N_24990,N_24850);
and U25840 (N_25840,N_24458,N_24460);
or U25841 (N_25841,N_24867,N_24830);
or U25842 (N_25842,N_24341,N_24961);
xor U25843 (N_25843,N_24033,N_24134);
nor U25844 (N_25844,N_24863,N_24779);
nand U25845 (N_25845,N_24493,N_24383);
xor U25846 (N_25846,N_24916,N_24002);
nand U25847 (N_25847,N_24125,N_24564);
nand U25848 (N_25848,N_24233,N_24080);
nor U25849 (N_25849,N_24911,N_24085);
or U25850 (N_25850,N_24687,N_24711);
or U25851 (N_25851,N_24435,N_24099);
nor U25852 (N_25852,N_24923,N_24003);
nand U25853 (N_25853,N_24244,N_24755);
or U25854 (N_25854,N_24446,N_24200);
nor U25855 (N_25855,N_24086,N_24082);
nor U25856 (N_25856,N_24990,N_24073);
or U25857 (N_25857,N_24082,N_24786);
nand U25858 (N_25858,N_24361,N_24186);
nand U25859 (N_25859,N_24012,N_24981);
nor U25860 (N_25860,N_24657,N_24126);
nor U25861 (N_25861,N_24868,N_24833);
or U25862 (N_25862,N_24534,N_24561);
nor U25863 (N_25863,N_24901,N_24871);
nor U25864 (N_25864,N_24914,N_24728);
or U25865 (N_25865,N_24519,N_24190);
nand U25866 (N_25866,N_24099,N_24485);
nand U25867 (N_25867,N_24461,N_24754);
nand U25868 (N_25868,N_24872,N_24360);
nor U25869 (N_25869,N_24896,N_24451);
xor U25870 (N_25870,N_24982,N_24459);
and U25871 (N_25871,N_24125,N_24601);
nand U25872 (N_25872,N_24153,N_24435);
and U25873 (N_25873,N_24183,N_24216);
and U25874 (N_25874,N_24375,N_24975);
nor U25875 (N_25875,N_24878,N_24737);
or U25876 (N_25876,N_24426,N_24950);
or U25877 (N_25877,N_24993,N_24393);
and U25878 (N_25878,N_24604,N_24130);
nand U25879 (N_25879,N_24116,N_24577);
nor U25880 (N_25880,N_24831,N_24360);
xnor U25881 (N_25881,N_24217,N_24481);
nor U25882 (N_25882,N_24353,N_24808);
or U25883 (N_25883,N_24141,N_24349);
nand U25884 (N_25884,N_24631,N_24825);
nand U25885 (N_25885,N_24305,N_24495);
nand U25886 (N_25886,N_24295,N_24481);
nor U25887 (N_25887,N_24067,N_24392);
or U25888 (N_25888,N_24475,N_24733);
or U25889 (N_25889,N_24581,N_24278);
nand U25890 (N_25890,N_24399,N_24005);
and U25891 (N_25891,N_24780,N_24874);
xor U25892 (N_25892,N_24231,N_24569);
or U25893 (N_25893,N_24000,N_24517);
or U25894 (N_25894,N_24815,N_24766);
nor U25895 (N_25895,N_24422,N_24402);
nor U25896 (N_25896,N_24498,N_24065);
or U25897 (N_25897,N_24263,N_24785);
xnor U25898 (N_25898,N_24716,N_24194);
or U25899 (N_25899,N_24331,N_24365);
and U25900 (N_25900,N_24391,N_24256);
nor U25901 (N_25901,N_24507,N_24459);
or U25902 (N_25902,N_24617,N_24900);
nor U25903 (N_25903,N_24734,N_24563);
or U25904 (N_25904,N_24484,N_24700);
nor U25905 (N_25905,N_24044,N_24904);
nand U25906 (N_25906,N_24076,N_24299);
or U25907 (N_25907,N_24308,N_24827);
and U25908 (N_25908,N_24966,N_24331);
nand U25909 (N_25909,N_24394,N_24090);
nand U25910 (N_25910,N_24002,N_24182);
nor U25911 (N_25911,N_24747,N_24491);
nand U25912 (N_25912,N_24610,N_24590);
nand U25913 (N_25913,N_24487,N_24588);
or U25914 (N_25914,N_24327,N_24385);
xnor U25915 (N_25915,N_24081,N_24566);
nor U25916 (N_25916,N_24929,N_24971);
xnor U25917 (N_25917,N_24038,N_24764);
xor U25918 (N_25918,N_24832,N_24556);
and U25919 (N_25919,N_24942,N_24637);
nand U25920 (N_25920,N_24760,N_24059);
nor U25921 (N_25921,N_24700,N_24908);
or U25922 (N_25922,N_24428,N_24634);
nor U25923 (N_25923,N_24560,N_24831);
xnor U25924 (N_25924,N_24916,N_24956);
xor U25925 (N_25925,N_24826,N_24034);
nor U25926 (N_25926,N_24468,N_24200);
xor U25927 (N_25927,N_24019,N_24149);
or U25928 (N_25928,N_24845,N_24867);
or U25929 (N_25929,N_24923,N_24985);
nor U25930 (N_25930,N_24844,N_24243);
or U25931 (N_25931,N_24900,N_24019);
or U25932 (N_25932,N_24254,N_24466);
xnor U25933 (N_25933,N_24532,N_24355);
or U25934 (N_25934,N_24526,N_24691);
nor U25935 (N_25935,N_24487,N_24495);
xor U25936 (N_25936,N_24206,N_24585);
and U25937 (N_25937,N_24755,N_24668);
nor U25938 (N_25938,N_24266,N_24833);
and U25939 (N_25939,N_24309,N_24000);
and U25940 (N_25940,N_24107,N_24079);
or U25941 (N_25941,N_24508,N_24629);
and U25942 (N_25942,N_24542,N_24171);
xnor U25943 (N_25943,N_24989,N_24069);
or U25944 (N_25944,N_24773,N_24851);
and U25945 (N_25945,N_24595,N_24403);
or U25946 (N_25946,N_24003,N_24109);
xnor U25947 (N_25947,N_24985,N_24260);
nand U25948 (N_25948,N_24879,N_24680);
and U25949 (N_25949,N_24796,N_24957);
nor U25950 (N_25950,N_24357,N_24238);
and U25951 (N_25951,N_24597,N_24891);
xnor U25952 (N_25952,N_24870,N_24624);
and U25953 (N_25953,N_24889,N_24506);
nand U25954 (N_25954,N_24454,N_24464);
or U25955 (N_25955,N_24827,N_24559);
nor U25956 (N_25956,N_24537,N_24181);
nand U25957 (N_25957,N_24031,N_24921);
xor U25958 (N_25958,N_24499,N_24192);
and U25959 (N_25959,N_24867,N_24699);
xor U25960 (N_25960,N_24489,N_24592);
and U25961 (N_25961,N_24649,N_24727);
and U25962 (N_25962,N_24948,N_24167);
or U25963 (N_25963,N_24699,N_24696);
and U25964 (N_25964,N_24956,N_24551);
and U25965 (N_25965,N_24806,N_24932);
nor U25966 (N_25966,N_24697,N_24188);
and U25967 (N_25967,N_24683,N_24254);
and U25968 (N_25968,N_24282,N_24448);
nand U25969 (N_25969,N_24015,N_24433);
xor U25970 (N_25970,N_24469,N_24370);
or U25971 (N_25971,N_24358,N_24224);
nor U25972 (N_25972,N_24496,N_24116);
nand U25973 (N_25973,N_24471,N_24573);
nor U25974 (N_25974,N_24978,N_24250);
xor U25975 (N_25975,N_24340,N_24919);
and U25976 (N_25976,N_24148,N_24011);
or U25977 (N_25977,N_24873,N_24505);
and U25978 (N_25978,N_24236,N_24630);
nor U25979 (N_25979,N_24135,N_24909);
or U25980 (N_25980,N_24353,N_24228);
or U25981 (N_25981,N_24910,N_24916);
xnor U25982 (N_25982,N_24435,N_24802);
nand U25983 (N_25983,N_24974,N_24124);
or U25984 (N_25984,N_24143,N_24624);
nor U25985 (N_25985,N_24651,N_24878);
nand U25986 (N_25986,N_24309,N_24180);
xor U25987 (N_25987,N_24249,N_24024);
and U25988 (N_25988,N_24962,N_24754);
and U25989 (N_25989,N_24854,N_24362);
xnor U25990 (N_25990,N_24412,N_24068);
nor U25991 (N_25991,N_24621,N_24872);
and U25992 (N_25992,N_24203,N_24223);
xor U25993 (N_25993,N_24015,N_24800);
or U25994 (N_25994,N_24990,N_24939);
xnor U25995 (N_25995,N_24076,N_24490);
xor U25996 (N_25996,N_24931,N_24812);
or U25997 (N_25997,N_24560,N_24731);
xnor U25998 (N_25998,N_24885,N_24573);
or U25999 (N_25999,N_24775,N_24136);
nand U26000 (N_26000,N_25709,N_25480);
and U26001 (N_26001,N_25939,N_25267);
and U26002 (N_26002,N_25720,N_25315);
and U26003 (N_26003,N_25955,N_25252);
nand U26004 (N_26004,N_25577,N_25590);
and U26005 (N_26005,N_25591,N_25484);
nor U26006 (N_26006,N_25877,N_25820);
and U26007 (N_26007,N_25189,N_25175);
xnor U26008 (N_26008,N_25755,N_25722);
nand U26009 (N_26009,N_25675,N_25422);
and U26010 (N_26010,N_25646,N_25676);
xor U26011 (N_26011,N_25151,N_25684);
or U26012 (N_26012,N_25573,N_25089);
xnor U26013 (N_26013,N_25423,N_25533);
nor U26014 (N_26014,N_25524,N_25688);
xnor U26015 (N_26015,N_25201,N_25313);
nor U26016 (N_26016,N_25585,N_25377);
or U26017 (N_26017,N_25016,N_25127);
nand U26018 (N_26018,N_25233,N_25110);
and U26019 (N_26019,N_25203,N_25657);
xnor U26020 (N_26020,N_25703,N_25586);
nand U26021 (N_26021,N_25804,N_25496);
and U26022 (N_26022,N_25772,N_25176);
or U26023 (N_26023,N_25965,N_25236);
and U26024 (N_26024,N_25753,N_25924);
xnor U26025 (N_26025,N_25025,N_25521);
or U26026 (N_26026,N_25083,N_25019);
and U26027 (N_26027,N_25882,N_25697);
xnor U26028 (N_26028,N_25084,N_25476);
nand U26029 (N_26029,N_25119,N_25731);
nand U26030 (N_26030,N_25013,N_25736);
xor U26031 (N_26031,N_25711,N_25562);
or U26032 (N_26032,N_25331,N_25656);
nor U26033 (N_26033,N_25557,N_25050);
nand U26034 (N_26034,N_25705,N_25730);
or U26035 (N_26035,N_25005,N_25283);
xor U26036 (N_26036,N_25715,N_25088);
xnor U26037 (N_26037,N_25260,N_25015);
nand U26038 (N_26038,N_25985,N_25274);
xnor U26039 (N_26039,N_25485,N_25692);
xnor U26040 (N_26040,N_25263,N_25404);
nand U26041 (N_26041,N_25474,N_25909);
or U26042 (N_26042,N_25850,N_25165);
and U26043 (N_26043,N_25883,N_25426);
or U26044 (N_26044,N_25744,N_25038);
nor U26045 (N_26045,N_25919,N_25589);
or U26046 (N_26046,N_25707,N_25011);
nor U26047 (N_26047,N_25397,N_25946);
xnor U26048 (N_26048,N_25219,N_25527);
or U26049 (N_26049,N_25543,N_25229);
nand U26050 (N_26050,N_25196,N_25477);
or U26051 (N_26051,N_25662,N_25704);
xor U26052 (N_26052,N_25440,N_25729);
and U26053 (N_26053,N_25205,N_25538);
nand U26054 (N_26054,N_25942,N_25362);
xnor U26055 (N_26055,N_25216,N_25545);
xor U26056 (N_26056,N_25858,N_25262);
nor U26057 (N_26057,N_25981,N_25462);
nand U26058 (N_26058,N_25978,N_25861);
xnor U26059 (N_26059,N_25246,N_25987);
and U26060 (N_26060,N_25359,N_25328);
nor U26061 (N_26061,N_25580,N_25624);
or U26062 (N_26062,N_25568,N_25375);
xor U26063 (N_26063,N_25797,N_25154);
or U26064 (N_26064,N_25152,N_25217);
and U26065 (N_26065,N_25493,N_25444);
or U26066 (N_26066,N_25596,N_25340);
or U26067 (N_26067,N_25643,N_25010);
and U26068 (N_26068,N_25598,N_25275);
xor U26069 (N_26069,N_25342,N_25391);
nor U26070 (N_26070,N_25846,N_25364);
nor U26071 (N_26071,N_25380,N_25872);
xnor U26072 (N_26072,N_25413,N_25035);
nor U26073 (N_26073,N_25650,N_25706);
or U26074 (N_26074,N_25698,N_25660);
xor U26075 (N_26075,N_25895,N_25158);
or U26076 (N_26076,N_25323,N_25728);
xor U26077 (N_26077,N_25156,N_25523);
and U26078 (N_26078,N_25139,N_25424);
nor U26079 (N_26079,N_25183,N_25501);
and U26080 (N_26080,N_25007,N_25979);
or U26081 (N_26081,N_25756,N_25266);
xor U26082 (N_26082,N_25102,N_25220);
nand U26083 (N_26083,N_25876,N_25137);
nor U26084 (N_26084,N_25320,N_25504);
nand U26085 (N_26085,N_25925,N_25750);
and U26086 (N_26086,N_25164,N_25917);
nand U26087 (N_26087,N_25746,N_25531);
nand U26088 (N_26088,N_25178,N_25180);
nor U26089 (N_26089,N_25901,N_25309);
and U26090 (N_26090,N_25109,N_25579);
or U26091 (N_26091,N_25487,N_25392);
nor U26092 (N_26092,N_25051,N_25247);
and U26093 (N_26093,N_25295,N_25903);
or U26094 (N_26094,N_25108,N_25930);
nor U26095 (N_26095,N_25992,N_25206);
nor U26096 (N_26096,N_25214,N_25161);
and U26097 (N_26097,N_25285,N_25499);
nor U26098 (N_26098,N_25608,N_25291);
or U26099 (N_26099,N_25818,N_25450);
or U26100 (N_26100,N_25814,N_25481);
xor U26101 (N_26101,N_25649,N_25542);
nor U26102 (N_26102,N_25115,N_25685);
and U26103 (N_26103,N_25078,N_25251);
and U26104 (N_26104,N_25854,N_25502);
xnor U26105 (N_26105,N_25467,N_25918);
or U26106 (N_26106,N_25963,N_25767);
nor U26107 (N_26107,N_25594,N_25672);
and U26108 (N_26108,N_25036,N_25149);
or U26109 (N_26109,N_25223,N_25922);
or U26110 (N_26110,N_25126,N_25635);
or U26111 (N_26111,N_25076,N_25099);
nand U26112 (N_26112,N_25582,N_25966);
or U26113 (N_26113,N_25620,N_25202);
or U26114 (N_26114,N_25130,N_25425);
xor U26115 (N_26115,N_25864,N_25230);
nand U26116 (N_26116,N_25337,N_25498);
or U26117 (N_26117,N_25983,N_25798);
xnor U26118 (N_26118,N_25863,N_25244);
or U26119 (N_26119,N_25836,N_25609);
nand U26120 (N_26120,N_25689,N_25757);
nand U26121 (N_26121,N_25443,N_25588);
or U26122 (N_26122,N_25610,N_25072);
nand U26123 (N_26123,N_25103,N_25254);
xnor U26124 (N_26124,N_25301,N_25973);
xnor U26125 (N_26125,N_25014,N_25454);
and U26126 (N_26126,N_25446,N_25314);
and U26127 (N_26127,N_25781,N_25002);
or U26128 (N_26128,N_25349,N_25293);
or U26129 (N_26129,N_25435,N_25827);
nor U26130 (N_26130,N_25079,N_25256);
xor U26131 (N_26131,N_25506,N_25823);
nand U26132 (N_26132,N_25682,N_25511);
or U26133 (N_26133,N_25592,N_25517);
xnor U26134 (N_26134,N_25897,N_25461);
nor U26135 (N_26135,N_25896,N_25259);
or U26136 (N_26136,N_25940,N_25522);
nand U26137 (N_26137,N_25224,N_25373);
and U26138 (N_26138,N_25638,N_25242);
or U26139 (N_26139,N_25037,N_25228);
and U26140 (N_26140,N_25075,N_25612);
xnor U26141 (N_26141,N_25875,N_25419);
or U26142 (N_26142,N_25761,N_25106);
xor U26143 (N_26143,N_25564,N_25700);
nor U26144 (N_26144,N_25209,N_25428);
and U26145 (N_26145,N_25352,N_25004);
or U26146 (N_26146,N_25032,N_25546);
and U26147 (N_26147,N_25647,N_25021);
or U26148 (N_26148,N_25621,N_25341);
or U26149 (N_26149,N_25681,N_25600);
nor U26150 (N_26150,N_25497,N_25500);
nor U26151 (N_26151,N_25411,N_25438);
or U26152 (N_26152,N_25702,N_25654);
nor U26153 (N_26153,N_25311,N_25358);
nor U26154 (N_26154,N_25353,N_25994);
nand U26155 (N_26155,N_25475,N_25408);
nand U26156 (N_26156,N_25257,N_25599);
xnor U26157 (N_26157,N_25033,N_25226);
or U26158 (N_26158,N_25794,N_25911);
or U26159 (N_26159,N_25355,N_25677);
or U26160 (N_26160,N_25733,N_25250);
or U26161 (N_26161,N_25881,N_25410);
or U26162 (N_26162,N_25748,N_25350);
nor U26163 (N_26163,N_25515,N_25095);
and U26164 (N_26164,N_25418,N_25416);
nand U26165 (N_26165,N_25017,N_25726);
nor U26166 (N_26166,N_25184,N_25210);
nor U26167 (N_26167,N_25607,N_25304);
nand U26168 (N_26168,N_25721,N_25764);
or U26169 (N_26169,N_25322,N_25473);
nand U26170 (N_26170,N_25009,N_25800);
nand U26171 (N_26171,N_25382,N_25991);
nand U26172 (N_26172,N_25128,N_25988);
or U26173 (N_26173,N_25125,N_25952);
nand U26174 (N_26174,N_25305,N_25751);
xor U26175 (N_26175,N_25330,N_25563);
nor U26176 (N_26176,N_25111,N_25817);
nand U26177 (N_26177,N_25822,N_25270);
xnor U26178 (N_26178,N_25551,N_25300);
nor U26179 (N_26179,N_25972,N_25347);
or U26180 (N_26180,N_25540,N_25695);
or U26181 (N_26181,N_25860,N_25316);
nor U26182 (N_26182,N_25121,N_25796);
xnor U26183 (N_26183,N_25276,N_25063);
or U26184 (N_26184,N_25307,N_25921);
or U26185 (N_26185,N_25041,N_25970);
nor U26186 (N_26186,N_25890,N_25948);
nand U26187 (N_26187,N_25363,N_25690);
xnor U26188 (N_26188,N_25082,N_25029);
or U26189 (N_26189,N_25891,N_25759);
nor U26190 (N_26190,N_25949,N_25777);
and U26191 (N_26191,N_25466,N_25554);
xor U26192 (N_26192,N_25699,N_25792);
nor U26193 (N_26193,N_25652,N_25775);
xnor U26194 (N_26194,N_25844,N_25616);
nand U26195 (N_26195,N_25144,N_25281);
nand U26196 (N_26196,N_25779,N_25490);
or U26197 (N_26197,N_25980,N_25287);
nand U26198 (N_26198,N_25514,N_25321);
and U26199 (N_26199,N_25866,N_25225);
and U26200 (N_26200,N_25296,N_25548);
xnor U26201 (N_26201,N_25054,N_25964);
nand U26202 (N_26202,N_25138,N_25336);
or U26203 (N_26203,N_25631,N_25566);
or U26204 (N_26204,N_25833,N_25665);
xor U26205 (N_26205,N_25837,N_25483);
nand U26206 (N_26206,N_25874,N_25625);
xor U26207 (N_26207,N_25302,N_25163);
or U26208 (N_26208,N_25951,N_25065);
nor U26209 (N_26209,N_25006,N_25085);
and U26210 (N_26210,N_25795,N_25583);
and U26211 (N_26211,N_25787,N_25603);
and U26212 (N_26212,N_25122,N_25606);
nand U26213 (N_26213,N_25478,N_25989);
or U26214 (N_26214,N_25146,N_25819);
or U26215 (N_26215,N_25414,N_25264);
or U26216 (N_26216,N_25813,N_25816);
or U26217 (N_26217,N_25329,N_25995);
nand U26218 (N_26218,N_25071,N_25031);
and U26219 (N_26219,N_25034,N_25519);
nand U26220 (N_26220,N_25464,N_25303);
and U26221 (N_26221,N_25859,N_25834);
nor U26222 (N_26222,N_25100,N_25288);
nand U26223 (N_26223,N_25143,N_25441);
xnor U26224 (N_26224,N_25830,N_25198);
nor U26225 (N_26225,N_25055,N_25962);
nand U26226 (N_26226,N_25537,N_25943);
xor U26227 (N_26227,N_25402,N_25576);
and U26228 (N_26228,N_25332,N_25788);
xnor U26229 (N_26229,N_25098,N_25213);
nor U26230 (N_26230,N_25191,N_25870);
xor U26231 (N_26231,N_25286,N_25935);
or U26232 (N_26232,N_25086,N_25388);
xnor U26233 (N_26233,N_25920,N_25857);
nor U26234 (N_26234,N_25243,N_25693);
nand U26235 (N_26235,N_25384,N_25871);
xor U26236 (N_26236,N_25740,N_25671);
nor U26237 (N_26237,N_25207,N_25162);
or U26238 (N_26238,N_25237,N_25701);
and U26239 (N_26239,N_25645,N_25070);
xnor U26240 (N_26240,N_25905,N_25471);
and U26241 (N_26241,N_25026,N_25843);
nor U26242 (N_26242,N_25640,N_25674);
nor U26243 (N_26243,N_25713,N_25190);
nand U26244 (N_26244,N_25773,N_25766);
or U26245 (N_26245,N_25595,N_25718);
nand U26246 (N_26246,N_25835,N_25512);
or U26247 (N_26247,N_25208,N_25786);
xor U26248 (N_26248,N_25299,N_25604);
nand U26249 (N_26249,N_25714,N_25436);
nor U26250 (N_26250,N_25298,N_25136);
nor U26251 (N_26251,N_25027,N_25459);
xnor U26252 (N_26252,N_25453,N_25123);
xnor U26253 (N_26253,N_25437,N_25601);
xnor U26254 (N_26254,N_25782,N_25663);
nand U26255 (N_26255,N_25494,N_25648);
xor U26256 (N_26256,N_25977,N_25280);
xnor U26257 (N_26257,N_25231,N_25087);
nand U26258 (N_26258,N_25996,N_25957);
xnor U26259 (N_26259,N_25687,N_25632);
or U26260 (N_26260,N_25308,N_25150);
nand U26261 (N_26261,N_25018,N_25101);
or U26262 (N_26262,N_25194,N_25181);
nand U26263 (N_26263,N_25926,N_25407);
xor U26264 (N_26264,N_25094,N_25294);
nor U26265 (N_26265,N_25869,N_25403);
xor U26266 (N_26266,N_25096,N_25354);
xor U26267 (N_26267,N_25971,N_25389);
xor U26268 (N_26268,N_25365,N_25113);
nor U26269 (N_26269,N_25003,N_25651);
nand U26270 (N_26270,N_25039,N_25914);
nor U26271 (N_26271,N_25140,N_25587);
nor U26272 (N_26272,N_25998,N_25628);
xnor U26273 (N_26273,N_25265,N_25449);
nor U26274 (N_26274,N_25581,N_25776);
and U26275 (N_26275,N_25838,N_25434);
nand U26276 (N_26276,N_25928,N_25145);
nor U26277 (N_26277,N_25908,N_25735);
nand U26278 (N_26278,N_25975,N_25763);
nand U26279 (N_26279,N_25240,N_25468);
or U26280 (N_26280,N_25912,N_25451);
xnor U26281 (N_26281,N_25742,N_25893);
xnor U26282 (N_26282,N_25062,N_25765);
and U26283 (N_26283,N_25052,N_25769);
nand U26284 (N_26284,N_25556,N_25778);
nor U26285 (N_26285,N_25399,N_25204);
nand U26286 (N_26286,N_25617,N_25661);
xnor U26287 (N_26287,N_25659,N_25048);
or U26288 (N_26288,N_25068,N_25001);
nor U26289 (N_26289,N_25169,N_25356);
or U26290 (N_26290,N_25547,N_25452);
and U26291 (N_26291,N_25578,N_25749);
and U26292 (N_26292,N_25944,N_25771);
nand U26293 (N_26293,N_25719,N_25218);
or U26294 (N_26294,N_25370,N_25986);
or U26295 (N_26295,N_25486,N_25241);
and U26296 (N_26296,N_25815,N_25999);
or U26297 (N_26297,N_25878,N_25310);
or U26298 (N_26298,N_25116,N_25694);
nand U26299 (N_26299,N_25560,N_25369);
nor U26300 (N_26300,N_25134,N_25915);
and U26301 (N_26301,N_25530,N_25064);
nand U26302 (N_26302,N_25770,N_25887);
and U26303 (N_26303,N_25712,N_25345);
nor U26304 (N_26304,N_25541,N_25852);
nand U26305 (N_26305,N_25458,N_25249);
or U26306 (N_26306,N_25567,N_25505);
nor U26307 (N_26307,N_25147,N_25832);
nor U26308 (N_26308,N_25465,N_25059);
nor U26309 (N_26309,N_25023,N_25529);
and U26310 (N_26310,N_25611,N_25160);
and U26311 (N_26311,N_25398,N_25385);
nand U26312 (N_26312,N_25880,N_25780);
or U26313 (N_26313,N_25862,N_25066);
and U26314 (N_26314,N_25976,N_25509);
xnor U26315 (N_26315,N_25442,N_25811);
nand U26316 (N_26316,N_25752,N_25167);
nand U26317 (N_26317,N_25679,N_25417);
or U26318 (N_26318,N_25405,N_25171);
and U26319 (N_26319,N_25723,N_25351);
nand U26320 (N_26320,N_25990,N_25653);
nand U26321 (N_26321,N_25664,N_25374);
and U26322 (N_26322,N_25326,N_25539);
nand U26323 (N_26323,N_25848,N_25574);
and U26324 (N_26324,N_25049,N_25785);
nand U26325 (N_26325,N_25069,N_25107);
xor U26326 (N_26326,N_25215,N_25636);
nand U26327 (N_26327,N_25555,N_25809);
or U26328 (N_26328,N_25325,N_25741);
and U26329 (N_26329,N_25544,N_25024);
nor U26330 (N_26330,N_25284,N_25271);
nand U26331 (N_26331,N_25383,N_25460);
nand U26332 (N_26332,N_25093,N_25269);
and U26333 (N_26333,N_25774,N_25810);
or U26334 (N_26334,N_25510,N_25124);
xnor U26335 (N_26335,N_25187,N_25894);
nor U26336 (N_26336,N_25784,N_25680);
xnor U26337 (N_26337,N_25367,N_25378);
xnor U26338 (N_26338,N_25867,N_25982);
nand U26339 (N_26339,N_25668,N_25802);
nor U26340 (N_26340,N_25916,N_25406);
nor U26341 (N_26341,N_25793,N_25950);
nand U26342 (N_26342,N_25348,N_25807);
or U26343 (N_26343,N_25170,N_25532);
nand U26344 (N_26344,N_25132,N_25826);
nor U26345 (N_26345,N_25053,N_25118);
nor U26346 (N_26346,N_25840,N_25536);
xnor U26347 (N_26347,N_25724,N_25691);
and U26348 (N_26348,N_25520,N_25327);
nor U26349 (N_26349,N_25470,N_25923);
and U26350 (N_26350,N_25457,N_25012);
xor U26351 (N_26351,N_25552,N_25945);
nand U26352 (N_26352,N_25421,N_25849);
and U26353 (N_26353,N_25993,N_25934);
xor U26354 (N_26354,N_25941,N_25339);
xnor U26355 (N_26355,N_25805,N_25630);
nand U26356 (N_26356,N_25448,N_25077);
xor U26357 (N_26357,N_25629,N_25297);
or U26358 (N_26358,N_25155,N_25045);
nand U26359 (N_26359,N_25879,N_25456);
or U26360 (N_26360,N_25758,N_25008);
and U26361 (N_26361,N_25953,N_25873);
and U26362 (N_26362,N_25197,N_25503);
nor U26363 (N_26363,N_25495,N_25239);
xnor U26364 (N_26364,N_25090,N_25614);
or U26365 (N_26365,N_25080,N_25186);
nand U26366 (N_26366,N_25227,N_25028);
nand U26367 (N_26367,N_25222,N_25431);
or U26368 (N_26368,N_25931,N_25831);
nor U26369 (N_26369,N_25984,N_25046);
and U26370 (N_26370,N_25899,N_25129);
nor U26371 (N_26371,N_25381,N_25278);
xor U26372 (N_26372,N_25710,N_25120);
or U26373 (N_26373,N_25273,N_25221);
xor U26374 (N_26374,N_25185,N_25969);
or U26375 (N_26375,N_25081,N_25235);
or U26376 (N_26376,N_25847,N_25074);
and U26377 (N_26377,N_25559,N_25754);
and U26378 (N_26378,N_25633,N_25390);
xor U26379 (N_26379,N_25334,N_25768);
and U26380 (N_26380,N_25200,N_25900);
nor U26381 (N_26381,N_25958,N_25174);
nor U26382 (N_26382,N_25371,N_25429);
nand U26383 (N_26383,N_25828,N_25067);
and U26384 (N_26384,N_25289,N_25360);
or U26385 (N_26385,N_25433,N_25439);
and U26386 (N_26386,N_25114,N_25727);
or U26387 (N_26387,N_25936,N_25892);
or U26388 (N_26388,N_25575,N_25131);
nand U26389 (N_26389,N_25199,N_25821);
nor U26390 (N_26390,N_25073,N_25042);
nor U26391 (N_26391,N_25829,N_25211);
xnor U26392 (N_26392,N_25550,N_25317);
and U26393 (N_26393,N_25622,N_25961);
nor U26394 (N_26394,N_25333,N_25841);
xor U26395 (N_26395,N_25762,N_25104);
nor U26396 (N_26396,N_25518,N_25279);
nor U26397 (N_26397,N_25386,N_25412);
and U26398 (N_26398,N_25683,N_25799);
or U26399 (N_26399,N_25553,N_25974);
and U26400 (N_26400,N_25376,N_25602);
xor U26401 (N_26401,N_25043,N_25558);
nor U26402 (N_26402,N_25669,N_25343);
nor U26403 (N_26403,N_25292,N_25627);
nand U26404 (N_26404,N_25904,N_25686);
nor U26405 (N_26405,N_25133,N_25745);
nor U26406 (N_26406,N_25569,N_25022);
xnor U26407 (N_26407,N_25868,N_25142);
or U26408 (N_26408,N_25626,N_25097);
nor U26409 (N_26409,N_25482,N_25166);
nand U26410 (N_26410,N_25179,N_25491);
and U26411 (N_26411,N_25234,N_25248);
and U26412 (N_26412,N_25489,N_25855);
nor U26413 (N_26413,N_25839,N_25565);
and U26414 (N_26414,N_25615,N_25513);
xor U26415 (N_26415,N_25357,N_25889);
and U26416 (N_26416,N_25056,N_25112);
and U26417 (N_26417,N_25312,N_25856);
nor U26418 (N_26418,N_25667,N_25888);
and U26419 (N_26419,N_25886,N_25245);
nand U26420 (N_26420,N_25658,N_25061);
and U26421 (N_26421,N_25670,N_25584);
or U26422 (N_26422,N_25516,N_25678);
nand U26423 (N_26423,N_25387,N_25060);
nand U26424 (N_26424,N_25535,N_25865);
xnor U26425 (N_26425,N_25725,N_25938);
nor U26426 (N_26426,N_25047,N_25913);
and U26427 (N_26427,N_25193,N_25335);
nand U26428 (N_26428,N_25789,N_25716);
xor U26429 (N_26429,N_25808,N_25644);
nand U26430 (N_26430,N_25572,N_25153);
xnor U26431 (N_26431,N_25395,N_25997);
nor U26432 (N_26432,N_25534,N_25157);
xnor U26433 (N_26433,N_25195,N_25409);
or U26434 (N_26434,N_25737,N_25253);
xnor U26435 (N_26435,N_25372,N_25401);
nor U26436 (N_26436,N_25238,N_25368);
or U26437 (N_26437,N_25927,N_25933);
and U26438 (N_26438,N_25277,N_25324);
nor U26439 (N_26439,N_25783,N_25760);
or U26440 (N_26440,N_25488,N_25791);
and U26441 (N_26441,N_25907,N_25623);
xnor U26442 (N_26442,N_25306,N_25057);
nor U26443 (N_26443,N_25954,N_25379);
and U26444 (N_26444,N_25427,N_25570);
or U26445 (N_26445,N_25020,N_25708);
or U26446 (N_26446,N_25177,N_25338);
and U26447 (N_26447,N_25641,N_25947);
nand U26448 (N_26448,N_25666,N_25597);
and U26449 (N_26449,N_25141,N_25092);
xnor U26450 (N_26450,N_25282,N_25853);
nor U26451 (N_26451,N_25168,N_25508);
or U26452 (N_26452,N_25430,N_25272);
and U26453 (N_26453,N_25812,N_25824);
nor U26454 (N_26454,N_25344,N_25618);
xor U26455 (N_26455,N_25319,N_25906);
or U26456 (N_26456,N_25549,N_25717);
nand U26457 (N_26457,N_25845,N_25159);
xnor U26458 (N_26458,N_25605,N_25884);
nor U26459 (N_26459,N_25959,N_25561);
nor U26460 (N_26460,N_25739,N_25040);
nand U26461 (N_26461,N_25902,N_25188);
nor U26462 (N_26462,N_25447,N_25634);
nor U26463 (N_26463,N_25696,N_25734);
nand U26464 (N_26464,N_25135,N_25885);
nand U26465 (N_26465,N_25091,N_25148);
or U26466 (N_26466,N_25268,N_25469);
and U26467 (N_26467,N_25613,N_25842);
xnor U26468 (N_26468,N_25673,N_25655);
nand U26469 (N_26469,N_25639,N_25910);
or U26470 (N_26470,N_25642,N_25117);
and U26471 (N_26471,N_25182,N_25851);
nor U26472 (N_26472,N_25507,N_25463);
or U26473 (N_26473,N_25420,N_25258);
nor U26474 (N_26474,N_25415,N_25044);
nand U26475 (N_26475,N_25479,N_25105);
and U26476 (N_26476,N_25212,N_25825);
nand U26477 (N_26477,N_25192,N_25738);
nand U26478 (N_26478,N_25801,N_25472);
and U26479 (N_26479,N_25732,N_25366);
nor U26480 (N_26480,N_25030,N_25290);
nor U26481 (N_26481,N_25593,N_25743);
nand U26482 (N_26482,N_25455,N_25261);
nor U26483 (N_26483,N_25898,N_25528);
or U26484 (N_26484,N_25526,N_25967);
and U26485 (N_26485,N_25790,N_25932);
nor U26486 (N_26486,N_25173,N_25806);
and U26487 (N_26487,N_25400,N_25492);
xnor U26488 (N_26488,N_25000,N_25747);
xnor U26489 (N_26489,N_25361,N_25571);
nor U26490 (N_26490,N_25956,N_25232);
nor U26491 (N_26491,N_25318,N_25396);
nand U26492 (N_26492,N_25929,N_25525);
xor U26493 (N_26493,N_25960,N_25445);
nand U26494 (N_26494,N_25255,N_25432);
nor U26495 (N_26495,N_25346,N_25619);
and U26496 (N_26496,N_25803,N_25172);
nand U26497 (N_26497,N_25394,N_25937);
nor U26498 (N_26498,N_25058,N_25393);
or U26499 (N_26499,N_25637,N_25968);
nand U26500 (N_26500,N_25548,N_25703);
nand U26501 (N_26501,N_25746,N_25395);
or U26502 (N_26502,N_25228,N_25515);
nor U26503 (N_26503,N_25489,N_25624);
or U26504 (N_26504,N_25008,N_25887);
or U26505 (N_26505,N_25456,N_25630);
nor U26506 (N_26506,N_25370,N_25000);
and U26507 (N_26507,N_25749,N_25857);
nand U26508 (N_26508,N_25227,N_25458);
xnor U26509 (N_26509,N_25827,N_25612);
or U26510 (N_26510,N_25819,N_25637);
xor U26511 (N_26511,N_25766,N_25919);
xor U26512 (N_26512,N_25568,N_25552);
nor U26513 (N_26513,N_25094,N_25398);
and U26514 (N_26514,N_25315,N_25681);
xor U26515 (N_26515,N_25645,N_25929);
nor U26516 (N_26516,N_25466,N_25735);
nor U26517 (N_26517,N_25503,N_25744);
and U26518 (N_26518,N_25960,N_25530);
or U26519 (N_26519,N_25335,N_25318);
xnor U26520 (N_26520,N_25048,N_25080);
or U26521 (N_26521,N_25923,N_25115);
nand U26522 (N_26522,N_25260,N_25458);
and U26523 (N_26523,N_25103,N_25256);
nand U26524 (N_26524,N_25599,N_25102);
nor U26525 (N_26525,N_25129,N_25736);
xor U26526 (N_26526,N_25939,N_25485);
nor U26527 (N_26527,N_25911,N_25896);
nand U26528 (N_26528,N_25678,N_25366);
nand U26529 (N_26529,N_25590,N_25373);
nand U26530 (N_26530,N_25455,N_25792);
nor U26531 (N_26531,N_25089,N_25549);
nor U26532 (N_26532,N_25793,N_25140);
and U26533 (N_26533,N_25314,N_25866);
or U26534 (N_26534,N_25766,N_25788);
or U26535 (N_26535,N_25946,N_25973);
and U26536 (N_26536,N_25652,N_25165);
nand U26537 (N_26537,N_25057,N_25118);
or U26538 (N_26538,N_25516,N_25259);
or U26539 (N_26539,N_25579,N_25960);
or U26540 (N_26540,N_25889,N_25121);
and U26541 (N_26541,N_25358,N_25017);
nor U26542 (N_26542,N_25249,N_25234);
or U26543 (N_26543,N_25066,N_25507);
and U26544 (N_26544,N_25233,N_25974);
and U26545 (N_26545,N_25472,N_25501);
or U26546 (N_26546,N_25805,N_25256);
nor U26547 (N_26547,N_25153,N_25994);
nor U26548 (N_26548,N_25240,N_25817);
or U26549 (N_26549,N_25833,N_25117);
or U26550 (N_26550,N_25545,N_25473);
xnor U26551 (N_26551,N_25493,N_25823);
nand U26552 (N_26552,N_25434,N_25816);
nand U26553 (N_26553,N_25282,N_25354);
and U26554 (N_26554,N_25556,N_25348);
nor U26555 (N_26555,N_25964,N_25047);
or U26556 (N_26556,N_25484,N_25830);
nor U26557 (N_26557,N_25055,N_25166);
nand U26558 (N_26558,N_25509,N_25333);
nor U26559 (N_26559,N_25616,N_25483);
or U26560 (N_26560,N_25273,N_25266);
or U26561 (N_26561,N_25568,N_25126);
nand U26562 (N_26562,N_25939,N_25442);
nor U26563 (N_26563,N_25286,N_25453);
or U26564 (N_26564,N_25888,N_25829);
nor U26565 (N_26565,N_25996,N_25824);
nor U26566 (N_26566,N_25270,N_25977);
xnor U26567 (N_26567,N_25015,N_25168);
or U26568 (N_26568,N_25343,N_25315);
nand U26569 (N_26569,N_25067,N_25302);
or U26570 (N_26570,N_25618,N_25952);
nor U26571 (N_26571,N_25513,N_25956);
nor U26572 (N_26572,N_25326,N_25726);
nor U26573 (N_26573,N_25319,N_25810);
or U26574 (N_26574,N_25511,N_25704);
or U26575 (N_26575,N_25786,N_25485);
xnor U26576 (N_26576,N_25507,N_25020);
xnor U26577 (N_26577,N_25490,N_25231);
nand U26578 (N_26578,N_25415,N_25476);
xnor U26579 (N_26579,N_25947,N_25487);
nor U26580 (N_26580,N_25324,N_25108);
or U26581 (N_26581,N_25463,N_25192);
xor U26582 (N_26582,N_25439,N_25076);
xnor U26583 (N_26583,N_25733,N_25628);
nor U26584 (N_26584,N_25846,N_25375);
xnor U26585 (N_26585,N_25511,N_25600);
nor U26586 (N_26586,N_25088,N_25051);
nor U26587 (N_26587,N_25005,N_25676);
nor U26588 (N_26588,N_25015,N_25899);
xnor U26589 (N_26589,N_25066,N_25768);
nand U26590 (N_26590,N_25993,N_25584);
nor U26591 (N_26591,N_25677,N_25684);
or U26592 (N_26592,N_25540,N_25658);
xnor U26593 (N_26593,N_25627,N_25124);
and U26594 (N_26594,N_25394,N_25172);
xnor U26595 (N_26595,N_25909,N_25015);
and U26596 (N_26596,N_25537,N_25459);
and U26597 (N_26597,N_25714,N_25142);
xor U26598 (N_26598,N_25688,N_25872);
or U26599 (N_26599,N_25419,N_25729);
and U26600 (N_26600,N_25010,N_25471);
xnor U26601 (N_26601,N_25501,N_25620);
nand U26602 (N_26602,N_25774,N_25738);
and U26603 (N_26603,N_25328,N_25112);
or U26604 (N_26604,N_25347,N_25031);
and U26605 (N_26605,N_25387,N_25831);
or U26606 (N_26606,N_25423,N_25510);
or U26607 (N_26607,N_25168,N_25182);
or U26608 (N_26608,N_25805,N_25078);
or U26609 (N_26609,N_25303,N_25630);
and U26610 (N_26610,N_25655,N_25001);
nor U26611 (N_26611,N_25143,N_25076);
nand U26612 (N_26612,N_25812,N_25350);
xnor U26613 (N_26613,N_25953,N_25222);
or U26614 (N_26614,N_25693,N_25080);
xnor U26615 (N_26615,N_25594,N_25084);
nor U26616 (N_26616,N_25142,N_25382);
and U26617 (N_26617,N_25070,N_25135);
or U26618 (N_26618,N_25217,N_25687);
nor U26619 (N_26619,N_25180,N_25523);
nand U26620 (N_26620,N_25514,N_25825);
nor U26621 (N_26621,N_25395,N_25265);
and U26622 (N_26622,N_25859,N_25755);
and U26623 (N_26623,N_25725,N_25421);
and U26624 (N_26624,N_25422,N_25528);
nor U26625 (N_26625,N_25598,N_25224);
and U26626 (N_26626,N_25758,N_25837);
nor U26627 (N_26627,N_25320,N_25274);
or U26628 (N_26628,N_25580,N_25070);
or U26629 (N_26629,N_25595,N_25412);
or U26630 (N_26630,N_25465,N_25356);
nand U26631 (N_26631,N_25424,N_25510);
or U26632 (N_26632,N_25558,N_25492);
and U26633 (N_26633,N_25481,N_25567);
xnor U26634 (N_26634,N_25732,N_25185);
and U26635 (N_26635,N_25306,N_25562);
nor U26636 (N_26636,N_25385,N_25392);
or U26637 (N_26637,N_25474,N_25522);
xnor U26638 (N_26638,N_25184,N_25690);
nand U26639 (N_26639,N_25168,N_25252);
and U26640 (N_26640,N_25122,N_25169);
nand U26641 (N_26641,N_25048,N_25198);
or U26642 (N_26642,N_25613,N_25944);
or U26643 (N_26643,N_25762,N_25863);
and U26644 (N_26644,N_25705,N_25971);
xnor U26645 (N_26645,N_25187,N_25902);
xor U26646 (N_26646,N_25245,N_25811);
nor U26647 (N_26647,N_25322,N_25679);
nor U26648 (N_26648,N_25623,N_25004);
and U26649 (N_26649,N_25013,N_25746);
nor U26650 (N_26650,N_25987,N_25502);
xnor U26651 (N_26651,N_25191,N_25691);
nor U26652 (N_26652,N_25061,N_25058);
xnor U26653 (N_26653,N_25486,N_25764);
xor U26654 (N_26654,N_25138,N_25241);
nand U26655 (N_26655,N_25687,N_25353);
nor U26656 (N_26656,N_25182,N_25548);
nor U26657 (N_26657,N_25385,N_25934);
nand U26658 (N_26658,N_25888,N_25789);
nand U26659 (N_26659,N_25506,N_25247);
and U26660 (N_26660,N_25073,N_25723);
or U26661 (N_26661,N_25900,N_25444);
or U26662 (N_26662,N_25506,N_25047);
or U26663 (N_26663,N_25189,N_25445);
or U26664 (N_26664,N_25808,N_25691);
nand U26665 (N_26665,N_25966,N_25304);
and U26666 (N_26666,N_25972,N_25138);
nand U26667 (N_26667,N_25931,N_25746);
xor U26668 (N_26668,N_25992,N_25036);
or U26669 (N_26669,N_25899,N_25649);
nand U26670 (N_26670,N_25267,N_25283);
nand U26671 (N_26671,N_25396,N_25262);
xnor U26672 (N_26672,N_25498,N_25492);
xor U26673 (N_26673,N_25305,N_25558);
nor U26674 (N_26674,N_25614,N_25743);
nand U26675 (N_26675,N_25415,N_25546);
xnor U26676 (N_26676,N_25536,N_25193);
and U26677 (N_26677,N_25407,N_25295);
nand U26678 (N_26678,N_25650,N_25293);
xor U26679 (N_26679,N_25247,N_25834);
nor U26680 (N_26680,N_25212,N_25328);
xor U26681 (N_26681,N_25026,N_25071);
nor U26682 (N_26682,N_25937,N_25026);
or U26683 (N_26683,N_25989,N_25990);
and U26684 (N_26684,N_25818,N_25043);
nand U26685 (N_26685,N_25191,N_25753);
and U26686 (N_26686,N_25536,N_25459);
xor U26687 (N_26687,N_25930,N_25735);
nand U26688 (N_26688,N_25579,N_25302);
nand U26689 (N_26689,N_25883,N_25935);
xnor U26690 (N_26690,N_25629,N_25609);
nand U26691 (N_26691,N_25441,N_25257);
and U26692 (N_26692,N_25224,N_25904);
or U26693 (N_26693,N_25143,N_25464);
nor U26694 (N_26694,N_25411,N_25151);
and U26695 (N_26695,N_25094,N_25616);
nor U26696 (N_26696,N_25859,N_25346);
or U26697 (N_26697,N_25962,N_25995);
nor U26698 (N_26698,N_25395,N_25111);
xnor U26699 (N_26699,N_25580,N_25257);
nand U26700 (N_26700,N_25336,N_25295);
xor U26701 (N_26701,N_25303,N_25394);
and U26702 (N_26702,N_25393,N_25323);
nand U26703 (N_26703,N_25880,N_25768);
nor U26704 (N_26704,N_25849,N_25454);
xnor U26705 (N_26705,N_25797,N_25538);
nand U26706 (N_26706,N_25174,N_25974);
nand U26707 (N_26707,N_25259,N_25274);
and U26708 (N_26708,N_25763,N_25670);
nor U26709 (N_26709,N_25783,N_25461);
xor U26710 (N_26710,N_25079,N_25093);
nand U26711 (N_26711,N_25788,N_25277);
and U26712 (N_26712,N_25629,N_25998);
or U26713 (N_26713,N_25162,N_25867);
nand U26714 (N_26714,N_25212,N_25758);
or U26715 (N_26715,N_25569,N_25671);
xor U26716 (N_26716,N_25333,N_25517);
and U26717 (N_26717,N_25758,N_25600);
xnor U26718 (N_26718,N_25510,N_25892);
xnor U26719 (N_26719,N_25780,N_25113);
xnor U26720 (N_26720,N_25207,N_25287);
nor U26721 (N_26721,N_25125,N_25157);
and U26722 (N_26722,N_25458,N_25902);
or U26723 (N_26723,N_25912,N_25587);
nand U26724 (N_26724,N_25876,N_25187);
or U26725 (N_26725,N_25269,N_25367);
and U26726 (N_26726,N_25884,N_25341);
or U26727 (N_26727,N_25966,N_25862);
nor U26728 (N_26728,N_25983,N_25612);
nor U26729 (N_26729,N_25765,N_25695);
nor U26730 (N_26730,N_25858,N_25516);
nor U26731 (N_26731,N_25609,N_25695);
nor U26732 (N_26732,N_25429,N_25477);
and U26733 (N_26733,N_25785,N_25448);
and U26734 (N_26734,N_25938,N_25925);
nand U26735 (N_26735,N_25336,N_25760);
or U26736 (N_26736,N_25010,N_25393);
xor U26737 (N_26737,N_25742,N_25023);
or U26738 (N_26738,N_25449,N_25444);
and U26739 (N_26739,N_25043,N_25551);
nand U26740 (N_26740,N_25376,N_25460);
nor U26741 (N_26741,N_25344,N_25713);
nand U26742 (N_26742,N_25432,N_25747);
xnor U26743 (N_26743,N_25809,N_25483);
xnor U26744 (N_26744,N_25330,N_25147);
and U26745 (N_26745,N_25087,N_25332);
xor U26746 (N_26746,N_25396,N_25791);
nand U26747 (N_26747,N_25908,N_25830);
xor U26748 (N_26748,N_25038,N_25120);
nor U26749 (N_26749,N_25639,N_25182);
xor U26750 (N_26750,N_25957,N_25003);
xnor U26751 (N_26751,N_25320,N_25802);
nor U26752 (N_26752,N_25974,N_25831);
nand U26753 (N_26753,N_25452,N_25324);
or U26754 (N_26754,N_25776,N_25701);
or U26755 (N_26755,N_25878,N_25275);
xor U26756 (N_26756,N_25928,N_25574);
nor U26757 (N_26757,N_25747,N_25727);
nor U26758 (N_26758,N_25134,N_25571);
and U26759 (N_26759,N_25371,N_25123);
or U26760 (N_26760,N_25366,N_25368);
or U26761 (N_26761,N_25166,N_25289);
and U26762 (N_26762,N_25733,N_25620);
nor U26763 (N_26763,N_25463,N_25877);
nor U26764 (N_26764,N_25238,N_25910);
xor U26765 (N_26765,N_25742,N_25136);
nor U26766 (N_26766,N_25379,N_25021);
nor U26767 (N_26767,N_25132,N_25638);
nand U26768 (N_26768,N_25548,N_25207);
nor U26769 (N_26769,N_25463,N_25024);
or U26770 (N_26770,N_25641,N_25345);
nand U26771 (N_26771,N_25039,N_25960);
and U26772 (N_26772,N_25279,N_25262);
nand U26773 (N_26773,N_25392,N_25289);
xor U26774 (N_26774,N_25585,N_25761);
xnor U26775 (N_26775,N_25133,N_25139);
xor U26776 (N_26776,N_25650,N_25814);
xor U26777 (N_26777,N_25210,N_25336);
and U26778 (N_26778,N_25038,N_25331);
or U26779 (N_26779,N_25906,N_25572);
nor U26780 (N_26780,N_25315,N_25449);
or U26781 (N_26781,N_25631,N_25211);
and U26782 (N_26782,N_25394,N_25118);
or U26783 (N_26783,N_25396,N_25371);
or U26784 (N_26784,N_25395,N_25249);
xnor U26785 (N_26785,N_25506,N_25046);
nor U26786 (N_26786,N_25914,N_25683);
nor U26787 (N_26787,N_25227,N_25886);
and U26788 (N_26788,N_25858,N_25631);
nor U26789 (N_26789,N_25297,N_25404);
or U26790 (N_26790,N_25475,N_25981);
nand U26791 (N_26791,N_25991,N_25921);
and U26792 (N_26792,N_25482,N_25311);
nand U26793 (N_26793,N_25089,N_25849);
and U26794 (N_26794,N_25619,N_25021);
nand U26795 (N_26795,N_25639,N_25911);
xor U26796 (N_26796,N_25172,N_25386);
and U26797 (N_26797,N_25468,N_25462);
xnor U26798 (N_26798,N_25227,N_25235);
and U26799 (N_26799,N_25355,N_25344);
or U26800 (N_26800,N_25370,N_25019);
xnor U26801 (N_26801,N_25080,N_25347);
nor U26802 (N_26802,N_25653,N_25994);
nor U26803 (N_26803,N_25578,N_25086);
nand U26804 (N_26804,N_25227,N_25034);
nor U26805 (N_26805,N_25375,N_25978);
and U26806 (N_26806,N_25084,N_25411);
xnor U26807 (N_26807,N_25054,N_25987);
or U26808 (N_26808,N_25191,N_25430);
nand U26809 (N_26809,N_25332,N_25934);
xnor U26810 (N_26810,N_25433,N_25799);
nand U26811 (N_26811,N_25387,N_25197);
or U26812 (N_26812,N_25881,N_25558);
nor U26813 (N_26813,N_25810,N_25052);
nor U26814 (N_26814,N_25379,N_25362);
nor U26815 (N_26815,N_25439,N_25712);
xnor U26816 (N_26816,N_25114,N_25239);
and U26817 (N_26817,N_25603,N_25161);
nand U26818 (N_26818,N_25583,N_25890);
nand U26819 (N_26819,N_25967,N_25880);
xnor U26820 (N_26820,N_25276,N_25136);
xnor U26821 (N_26821,N_25592,N_25709);
or U26822 (N_26822,N_25361,N_25139);
or U26823 (N_26823,N_25244,N_25692);
and U26824 (N_26824,N_25431,N_25690);
nor U26825 (N_26825,N_25422,N_25792);
nor U26826 (N_26826,N_25559,N_25356);
and U26827 (N_26827,N_25490,N_25560);
nor U26828 (N_26828,N_25668,N_25775);
or U26829 (N_26829,N_25070,N_25227);
xor U26830 (N_26830,N_25147,N_25671);
xnor U26831 (N_26831,N_25711,N_25287);
xnor U26832 (N_26832,N_25025,N_25226);
or U26833 (N_26833,N_25906,N_25986);
or U26834 (N_26834,N_25314,N_25482);
nand U26835 (N_26835,N_25261,N_25247);
xor U26836 (N_26836,N_25000,N_25093);
or U26837 (N_26837,N_25297,N_25391);
or U26838 (N_26838,N_25681,N_25601);
or U26839 (N_26839,N_25704,N_25210);
nand U26840 (N_26840,N_25096,N_25730);
xor U26841 (N_26841,N_25119,N_25463);
xnor U26842 (N_26842,N_25453,N_25962);
or U26843 (N_26843,N_25618,N_25740);
or U26844 (N_26844,N_25213,N_25273);
and U26845 (N_26845,N_25214,N_25851);
nand U26846 (N_26846,N_25412,N_25373);
nor U26847 (N_26847,N_25885,N_25924);
nor U26848 (N_26848,N_25674,N_25426);
or U26849 (N_26849,N_25083,N_25908);
xnor U26850 (N_26850,N_25971,N_25939);
nor U26851 (N_26851,N_25363,N_25529);
xnor U26852 (N_26852,N_25766,N_25739);
xor U26853 (N_26853,N_25033,N_25669);
nor U26854 (N_26854,N_25843,N_25518);
or U26855 (N_26855,N_25223,N_25479);
nand U26856 (N_26856,N_25140,N_25318);
xnor U26857 (N_26857,N_25668,N_25977);
nand U26858 (N_26858,N_25328,N_25416);
nor U26859 (N_26859,N_25278,N_25909);
or U26860 (N_26860,N_25991,N_25909);
and U26861 (N_26861,N_25246,N_25045);
nand U26862 (N_26862,N_25461,N_25259);
nor U26863 (N_26863,N_25699,N_25360);
xnor U26864 (N_26864,N_25094,N_25137);
or U26865 (N_26865,N_25139,N_25632);
nand U26866 (N_26866,N_25853,N_25394);
nor U26867 (N_26867,N_25479,N_25719);
xnor U26868 (N_26868,N_25825,N_25405);
nor U26869 (N_26869,N_25516,N_25419);
and U26870 (N_26870,N_25271,N_25380);
nor U26871 (N_26871,N_25575,N_25783);
or U26872 (N_26872,N_25704,N_25004);
xor U26873 (N_26873,N_25641,N_25552);
and U26874 (N_26874,N_25489,N_25731);
xor U26875 (N_26875,N_25715,N_25420);
nor U26876 (N_26876,N_25625,N_25794);
xnor U26877 (N_26877,N_25203,N_25115);
nor U26878 (N_26878,N_25553,N_25347);
nand U26879 (N_26879,N_25137,N_25085);
or U26880 (N_26880,N_25148,N_25399);
xnor U26881 (N_26881,N_25217,N_25769);
nor U26882 (N_26882,N_25877,N_25301);
xor U26883 (N_26883,N_25251,N_25408);
nor U26884 (N_26884,N_25553,N_25458);
or U26885 (N_26885,N_25906,N_25728);
xor U26886 (N_26886,N_25061,N_25518);
nor U26887 (N_26887,N_25364,N_25030);
and U26888 (N_26888,N_25361,N_25389);
xor U26889 (N_26889,N_25842,N_25835);
and U26890 (N_26890,N_25149,N_25266);
nor U26891 (N_26891,N_25614,N_25579);
nor U26892 (N_26892,N_25523,N_25366);
and U26893 (N_26893,N_25920,N_25016);
nand U26894 (N_26894,N_25473,N_25100);
nand U26895 (N_26895,N_25229,N_25006);
xor U26896 (N_26896,N_25368,N_25466);
and U26897 (N_26897,N_25467,N_25594);
and U26898 (N_26898,N_25427,N_25650);
and U26899 (N_26899,N_25330,N_25208);
and U26900 (N_26900,N_25238,N_25712);
and U26901 (N_26901,N_25818,N_25406);
nor U26902 (N_26902,N_25666,N_25895);
nor U26903 (N_26903,N_25291,N_25264);
nor U26904 (N_26904,N_25138,N_25220);
nand U26905 (N_26905,N_25337,N_25947);
nor U26906 (N_26906,N_25319,N_25337);
nand U26907 (N_26907,N_25539,N_25728);
nor U26908 (N_26908,N_25869,N_25660);
nor U26909 (N_26909,N_25891,N_25921);
nand U26910 (N_26910,N_25486,N_25462);
and U26911 (N_26911,N_25031,N_25469);
xnor U26912 (N_26912,N_25525,N_25839);
nor U26913 (N_26913,N_25426,N_25112);
nand U26914 (N_26914,N_25083,N_25631);
nand U26915 (N_26915,N_25990,N_25273);
and U26916 (N_26916,N_25531,N_25342);
xor U26917 (N_26917,N_25381,N_25952);
nand U26918 (N_26918,N_25118,N_25645);
and U26919 (N_26919,N_25093,N_25358);
nand U26920 (N_26920,N_25551,N_25819);
xnor U26921 (N_26921,N_25993,N_25193);
or U26922 (N_26922,N_25690,N_25239);
and U26923 (N_26923,N_25177,N_25580);
xnor U26924 (N_26924,N_25687,N_25450);
nand U26925 (N_26925,N_25664,N_25727);
nor U26926 (N_26926,N_25240,N_25966);
nor U26927 (N_26927,N_25684,N_25540);
or U26928 (N_26928,N_25402,N_25163);
nand U26929 (N_26929,N_25290,N_25859);
or U26930 (N_26930,N_25133,N_25312);
xor U26931 (N_26931,N_25490,N_25005);
or U26932 (N_26932,N_25511,N_25118);
xnor U26933 (N_26933,N_25058,N_25600);
nor U26934 (N_26934,N_25596,N_25707);
or U26935 (N_26935,N_25433,N_25838);
nand U26936 (N_26936,N_25187,N_25812);
nand U26937 (N_26937,N_25389,N_25080);
xnor U26938 (N_26938,N_25813,N_25737);
xor U26939 (N_26939,N_25057,N_25524);
and U26940 (N_26940,N_25904,N_25608);
nor U26941 (N_26941,N_25717,N_25510);
or U26942 (N_26942,N_25551,N_25795);
or U26943 (N_26943,N_25322,N_25781);
nor U26944 (N_26944,N_25260,N_25808);
xor U26945 (N_26945,N_25977,N_25894);
and U26946 (N_26946,N_25438,N_25398);
xnor U26947 (N_26947,N_25974,N_25985);
nand U26948 (N_26948,N_25545,N_25827);
nand U26949 (N_26949,N_25438,N_25031);
or U26950 (N_26950,N_25071,N_25787);
xnor U26951 (N_26951,N_25220,N_25775);
xnor U26952 (N_26952,N_25914,N_25186);
or U26953 (N_26953,N_25521,N_25479);
or U26954 (N_26954,N_25912,N_25702);
nand U26955 (N_26955,N_25322,N_25362);
nor U26956 (N_26956,N_25688,N_25622);
xor U26957 (N_26957,N_25497,N_25424);
xor U26958 (N_26958,N_25844,N_25116);
and U26959 (N_26959,N_25055,N_25499);
or U26960 (N_26960,N_25867,N_25308);
and U26961 (N_26961,N_25356,N_25308);
xnor U26962 (N_26962,N_25984,N_25101);
and U26963 (N_26963,N_25822,N_25815);
xnor U26964 (N_26964,N_25663,N_25856);
nand U26965 (N_26965,N_25462,N_25559);
xor U26966 (N_26966,N_25342,N_25487);
nand U26967 (N_26967,N_25570,N_25254);
xnor U26968 (N_26968,N_25272,N_25938);
xnor U26969 (N_26969,N_25532,N_25814);
nor U26970 (N_26970,N_25570,N_25207);
or U26971 (N_26971,N_25971,N_25243);
nor U26972 (N_26972,N_25683,N_25223);
xor U26973 (N_26973,N_25572,N_25735);
or U26974 (N_26974,N_25130,N_25734);
or U26975 (N_26975,N_25776,N_25166);
or U26976 (N_26976,N_25190,N_25411);
and U26977 (N_26977,N_25864,N_25700);
nor U26978 (N_26978,N_25130,N_25761);
nor U26979 (N_26979,N_25896,N_25335);
nor U26980 (N_26980,N_25696,N_25154);
nand U26981 (N_26981,N_25036,N_25776);
nand U26982 (N_26982,N_25890,N_25674);
or U26983 (N_26983,N_25532,N_25959);
nor U26984 (N_26984,N_25153,N_25749);
or U26985 (N_26985,N_25885,N_25701);
nand U26986 (N_26986,N_25518,N_25996);
nor U26987 (N_26987,N_25301,N_25936);
or U26988 (N_26988,N_25299,N_25831);
xor U26989 (N_26989,N_25191,N_25439);
and U26990 (N_26990,N_25371,N_25711);
nand U26991 (N_26991,N_25997,N_25678);
and U26992 (N_26992,N_25847,N_25161);
and U26993 (N_26993,N_25818,N_25900);
and U26994 (N_26994,N_25528,N_25005);
nand U26995 (N_26995,N_25155,N_25664);
nor U26996 (N_26996,N_25853,N_25626);
xor U26997 (N_26997,N_25803,N_25165);
xor U26998 (N_26998,N_25373,N_25727);
or U26999 (N_26999,N_25707,N_25384);
xor U27000 (N_27000,N_26648,N_26565);
xor U27001 (N_27001,N_26543,N_26049);
xnor U27002 (N_27002,N_26009,N_26256);
or U27003 (N_27003,N_26567,N_26766);
xnor U27004 (N_27004,N_26643,N_26966);
nor U27005 (N_27005,N_26157,N_26182);
nand U27006 (N_27006,N_26644,N_26642);
xor U27007 (N_27007,N_26133,N_26755);
or U27008 (N_27008,N_26340,N_26325);
and U27009 (N_27009,N_26839,N_26054);
nand U27010 (N_27010,N_26624,N_26029);
xor U27011 (N_27011,N_26367,N_26877);
nand U27012 (N_27012,N_26835,N_26019);
nand U27013 (N_27013,N_26456,N_26045);
and U27014 (N_27014,N_26844,N_26374);
or U27015 (N_27015,N_26968,N_26493);
xnor U27016 (N_27016,N_26812,N_26801);
and U27017 (N_27017,N_26486,N_26449);
xnor U27018 (N_27018,N_26739,N_26244);
nor U27019 (N_27019,N_26387,N_26473);
and U27020 (N_27020,N_26179,N_26251);
nand U27021 (N_27021,N_26089,N_26768);
and U27022 (N_27022,N_26266,N_26833);
nand U27023 (N_27023,N_26732,N_26665);
or U27024 (N_27024,N_26727,N_26756);
or U27025 (N_27025,N_26806,N_26993);
nor U27026 (N_27026,N_26587,N_26941);
or U27027 (N_27027,N_26464,N_26724);
and U27028 (N_27028,N_26892,N_26440);
and U27029 (N_27029,N_26479,N_26361);
and U27030 (N_27030,N_26615,N_26682);
and U27031 (N_27031,N_26669,N_26746);
nand U27032 (N_27032,N_26327,N_26524);
xor U27033 (N_27033,N_26073,N_26592);
nor U27034 (N_27034,N_26992,N_26792);
or U27035 (N_27035,N_26093,N_26646);
xnor U27036 (N_27036,N_26990,N_26043);
nor U27037 (N_27037,N_26581,N_26626);
nor U27038 (N_27038,N_26185,N_26301);
xor U27039 (N_27039,N_26427,N_26834);
nor U27040 (N_27040,N_26824,N_26509);
and U27041 (N_27041,N_26930,N_26653);
xnor U27042 (N_27042,N_26995,N_26339);
or U27043 (N_27043,N_26541,N_26106);
and U27044 (N_27044,N_26095,N_26282);
or U27045 (N_27045,N_26671,N_26603);
and U27046 (N_27046,N_26151,N_26061);
and U27047 (N_27047,N_26773,N_26243);
nand U27048 (N_27048,N_26060,N_26810);
nand U27049 (N_27049,N_26854,N_26178);
nand U27050 (N_27050,N_26032,N_26711);
xnor U27051 (N_27051,N_26690,N_26641);
nor U27052 (N_27052,N_26575,N_26666);
nand U27053 (N_27053,N_26776,N_26245);
and U27054 (N_27054,N_26111,N_26321);
and U27055 (N_27055,N_26942,N_26520);
nand U27056 (N_27056,N_26860,N_26602);
or U27057 (N_27057,N_26980,N_26584);
or U27058 (N_27058,N_26228,N_26884);
or U27059 (N_27059,N_26016,N_26475);
nor U27060 (N_27060,N_26580,N_26880);
nor U27061 (N_27061,N_26379,N_26426);
and U27062 (N_27062,N_26147,N_26199);
xor U27063 (N_27063,N_26416,N_26976);
and U27064 (N_27064,N_26637,N_26536);
nor U27065 (N_27065,N_26096,N_26752);
and U27066 (N_27066,N_26336,N_26720);
nor U27067 (N_27067,N_26809,N_26888);
nand U27068 (N_27068,N_26355,N_26700);
or U27069 (N_27069,N_26115,N_26161);
or U27070 (N_27070,N_26654,N_26769);
and U27071 (N_27071,N_26088,N_26289);
xnor U27072 (N_27072,N_26636,N_26323);
or U27073 (N_27073,N_26553,N_26136);
xnor U27074 (N_27074,N_26303,N_26476);
nor U27075 (N_27075,N_26918,N_26154);
or U27076 (N_27076,N_26905,N_26511);
nand U27077 (N_27077,N_26681,N_26840);
and U27078 (N_27078,N_26235,N_26633);
nor U27079 (N_27079,N_26530,N_26651);
xnor U27080 (N_27080,N_26948,N_26505);
or U27081 (N_27081,N_26099,N_26913);
nand U27082 (N_27082,N_26158,N_26070);
and U27083 (N_27083,N_26163,N_26242);
or U27084 (N_27084,N_26693,N_26173);
nor U27085 (N_27085,N_26529,N_26977);
nand U27086 (N_27086,N_26922,N_26398);
or U27087 (N_27087,N_26634,N_26863);
xnor U27088 (N_27088,N_26712,N_26063);
nor U27089 (N_27089,N_26431,N_26378);
xor U27090 (N_27090,N_26546,N_26687);
nor U27091 (N_27091,N_26503,N_26470);
nor U27092 (N_27092,N_26194,N_26858);
nand U27093 (N_27093,N_26613,N_26439);
nand U27094 (N_27094,N_26400,N_26443);
nor U27095 (N_27095,N_26605,N_26772);
xnor U27096 (N_27096,N_26808,N_26219);
xnor U27097 (N_27097,N_26931,N_26114);
nand U27098 (N_27098,N_26497,N_26571);
and U27099 (N_27099,N_26155,N_26310);
nand U27100 (N_27100,N_26925,N_26399);
or U27101 (N_27101,N_26939,N_26079);
nand U27102 (N_27102,N_26857,N_26261);
nand U27103 (N_27103,N_26196,N_26790);
xnor U27104 (N_27104,N_26798,N_26488);
xnor U27105 (N_27105,N_26477,N_26337);
nor U27106 (N_27106,N_26110,N_26973);
xnor U27107 (N_27107,N_26864,N_26504);
xor U27108 (N_27108,N_26388,N_26385);
or U27109 (N_27109,N_26077,N_26058);
and U27110 (N_27110,N_26326,N_26866);
xor U27111 (N_27111,N_26030,N_26177);
xor U27112 (N_27112,N_26607,N_26128);
xor U27113 (N_27113,N_26655,N_26652);
xnor U27114 (N_27114,N_26647,N_26932);
and U27115 (N_27115,N_26627,N_26225);
nand U27116 (N_27116,N_26786,N_26164);
nor U27117 (N_27117,N_26050,N_26342);
and U27118 (N_27118,N_26663,N_26532);
nand U27119 (N_27119,N_26425,N_26559);
and U27120 (N_27120,N_26501,N_26744);
and U27121 (N_27121,N_26015,N_26903);
nor U27122 (N_27122,N_26881,N_26871);
or U27123 (N_27123,N_26629,N_26238);
nand U27124 (N_27124,N_26902,N_26064);
nand U27125 (N_27125,N_26382,N_26041);
and U27126 (N_27126,N_26997,N_26991);
nand U27127 (N_27127,N_26429,N_26120);
or U27128 (N_27128,N_26468,N_26793);
and U27129 (N_27129,N_26375,N_26754);
and U27130 (N_27130,N_26038,N_26820);
xnor U27131 (N_27131,N_26344,N_26467);
or U27132 (N_27132,N_26861,N_26174);
nor U27133 (N_27133,N_26483,N_26075);
and U27134 (N_27134,N_26421,N_26356);
or U27135 (N_27135,N_26787,N_26350);
and U27136 (N_27136,N_26090,N_26999);
xnor U27137 (N_27137,N_26490,N_26287);
or U27138 (N_27138,N_26743,N_26121);
or U27139 (N_27139,N_26851,N_26923);
nor U27140 (N_27140,N_26510,N_26283);
xnor U27141 (N_27141,N_26713,N_26928);
or U27142 (N_27142,N_26152,N_26764);
and U27143 (N_27143,N_26859,N_26302);
xnor U27144 (N_27144,N_26583,N_26175);
xnor U27145 (N_27145,N_26001,N_26376);
or U27146 (N_27146,N_26577,N_26401);
xnor U27147 (N_27147,N_26292,N_26240);
nand U27148 (N_27148,N_26288,N_26940);
nor U27149 (N_27149,N_26211,N_26057);
nor U27150 (N_27150,N_26207,N_26296);
and U27151 (N_27151,N_26908,N_26481);
xor U27152 (N_27152,N_26482,N_26293);
nor U27153 (N_27153,N_26365,N_26778);
nand U27154 (N_27154,N_26679,N_26448);
xnor U27155 (N_27155,N_26684,N_26794);
nand U27156 (N_27156,N_26300,N_26869);
xor U27157 (N_27157,N_26662,N_26229);
xnor U27158 (N_27158,N_26212,N_26970);
xor U27159 (N_27159,N_26224,N_26492);
nor U27160 (N_27160,N_26703,N_26205);
and U27161 (N_27161,N_26371,N_26929);
and U27162 (N_27162,N_26558,N_26328);
or U27163 (N_27163,N_26188,N_26312);
nand U27164 (N_27164,N_26619,N_26384);
nor U27165 (N_27165,N_26522,N_26474);
nand U27166 (N_27166,N_26444,N_26614);
xor U27167 (N_27167,N_26017,N_26232);
nand U27168 (N_27168,N_26837,N_26442);
nor U27169 (N_27169,N_26363,N_26831);
or U27170 (N_27170,N_26461,N_26618);
nor U27171 (N_27171,N_26290,N_26517);
or U27172 (N_27172,N_26269,N_26085);
xor U27173 (N_27173,N_26496,N_26799);
xnor U27174 (N_27174,N_26039,N_26203);
nand U27175 (N_27175,N_26148,N_26829);
or U27176 (N_27176,N_26140,N_26975);
xnor U27177 (N_27177,N_26535,N_26286);
or U27178 (N_27178,N_26911,N_26499);
nor U27179 (N_27179,N_26206,N_26938);
nor U27180 (N_27180,N_26710,N_26515);
or U27181 (N_27181,N_26020,N_26707);
and U27182 (N_27182,N_26455,N_26714);
xnor U27183 (N_27183,N_26434,N_26391);
xor U27184 (N_27184,N_26753,N_26631);
nor U27185 (N_27185,N_26542,N_26838);
nand U27186 (N_27186,N_26471,N_26589);
nor U27187 (N_27187,N_26370,N_26156);
nand U27188 (N_27188,N_26137,N_26936);
xnor U27189 (N_27189,N_26873,N_26192);
nand U27190 (N_27190,N_26143,N_26359);
nor U27191 (N_27191,N_26953,N_26411);
and U27192 (N_27192,N_26612,N_26422);
nor U27193 (N_27193,N_26609,N_26130);
or U27194 (N_27194,N_26765,N_26625);
and U27195 (N_27195,N_26958,N_26572);
and U27196 (N_27196,N_26962,N_26112);
nand U27197 (N_27197,N_26722,N_26119);
or U27198 (N_27198,N_26215,N_26534);
nand U27199 (N_27199,N_26432,N_26390);
or U27200 (N_27200,N_26181,N_26495);
nor U27201 (N_27201,N_26308,N_26314);
and U27202 (N_27202,N_26879,N_26696);
or U27203 (N_27203,N_26048,N_26557);
nor U27204 (N_27204,N_26708,N_26569);
nand U27205 (N_27205,N_26149,N_26721);
and U27206 (N_27206,N_26927,N_26351);
nor U27207 (N_27207,N_26441,N_26162);
or U27208 (N_27208,N_26555,N_26819);
nor U27209 (N_27209,N_26804,N_26450);
nand U27210 (N_27210,N_26564,N_26022);
and U27211 (N_27211,N_26658,N_26952);
nand U27212 (N_27212,N_26200,N_26252);
xor U27213 (N_27213,N_26774,N_26322);
nand U27214 (N_27214,N_26132,N_26998);
nor U27215 (N_27215,N_26526,N_26067);
xnor U27216 (N_27216,N_26189,N_26725);
xor U27217 (N_27217,N_26981,N_26291);
xor U27218 (N_27218,N_26123,N_26987);
and U27219 (N_27219,N_26889,N_26210);
xor U27220 (N_27220,N_26352,N_26796);
and U27221 (N_27221,N_26544,N_26319);
nor U27222 (N_27222,N_26621,N_26248);
and U27223 (N_27223,N_26784,N_26920);
and U27224 (N_27224,N_26563,N_26271);
xor U27225 (N_27225,N_26412,N_26042);
nor U27226 (N_27226,N_26960,N_26066);
and U27227 (N_27227,N_26741,N_26409);
and U27228 (N_27228,N_26736,N_26628);
xnor U27229 (N_27229,N_26895,N_26538);
and U27230 (N_27230,N_26814,N_26904);
nand U27231 (N_27231,N_26898,N_26632);
or U27232 (N_27232,N_26678,N_26101);
and U27233 (N_27233,N_26317,N_26635);
or U27234 (N_27234,N_26417,N_26116);
nand U27235 (N_27235,N_26452,N_26082);
or U27236 (N_27236,N_26874,N_26608);
nor U27237 (N_27237,N_26539,N_26630);
nand U27238 (N_27238,N_26946,N_26969);
or U27239 (N_27239,N_26767,N_26909);
or U27240 (N_27240,N_26438,N_26389);
nand U27241 (N_27241,N_26453,N_26068);
nor U27242 (N_27242,N_26227,N_26836);
and U27243 (N_27243,N_26430,N_26545);
or U27244 (N_27244,N_26454,N_26435);
nand U27245 (N_27245,N_26570,N_26047);
nor U27246 (N_27246,N_26886,N_26974);
or U27247 (N_27247,N_26267,N_26280);
xor U27248 (N_27248,N_26491,N_26285);
nor U27249 (N_27249,N_26171,N_26008);
nand U27250 (N_27250,N_26113,N_26100);
and U27251 (N_27251,N_26761,N_26588);
nor U27252 (N_27252,N_26771,N_26780);
xnor U27253 (N_27253,N_26415,N_26051);
xnor U27254 (N_27254,N_26660,N_26423);
or U27255 (N_27255,N_26084,N_26978);
nor U27256 (N_27256,N_26424,N_26413);
and U27257 (N_27257,N_26601,N_26717);
nand U27258 (N_27258,N_26165,N_26268);
nand U27259 (N_27259,N_26081,N_26954);
and U27260 (N_27260,N_26318,N_26726);
or U27261 (N_27261,N_26817,N_26979);
and U27262 (N_27262,N_26000,N_26763);
nand U27263 (N_27263,N_26332,N_26947);
xor U27264 (N_27264,N_26885,N_26876);
nor U27265 (N_27265,N_26957,N_26330);
and U27266 (N_27266,N_26893,N_26396);
or U27267 (N_27267,N_26685,N_26005);
and U27268 (N_27268,N_26742,N_26264);
nor U27269 (N_27269,N_26528,N_26369);
and U27270 (N_27270,N_26349,N_26846);
and U27271 (N_27271,N_26316,N_26023);
nand U27272 (N_27272,N_26380,N_26596);
nand U27273 (N_27273,N_26297,N_26141);
nand U27274 (N_27274,N_26540,N_26273);
or U27275 (N_27275,N_26521,N_26353);
nand U27276 (N_27276,N_26853,N_26709);
and U27277 (N_27277,N_26234,N_26715);
or U27278 (N_27278,N_26279,N_26031);
and U27279 (N_27279,N_26166,N_26597);
and U27280 (N_27280,N_26305,N_26802);
nand U27281 (N_27281,N_26915,N_26190);
nor U27282 (N_27282,N_26683,N_26875);
xor U27283 (N_27283,N_26433,N_26402);
nand U27284 (N_27284,N_26697,N_26594);
and U27285 (N_27285,N_26664,N_26791);
xor U27286 (N_27286,N_26578,N_26728);
nor U27287 (N_27287,N_26445,N_26191);
nor U27288 (N_27288,N_26056,N_26582);
nand U27289 (N_27289,N_26972,N_26469);
or U27290 (N_27290,N_26983,N_26692);
or U27291 (N_27291,N_26329,N_26071);
nand U27292 (N_27292,N_26485,N_26500);
xnor U27293 (N_27293,N_26457,N_26872);
xnor U27294 (N_27294,N_26259,N_26783);
or U27295 (N_27295,N_26750,N_26815);
and U27296 (N_27296,N_26333,N_26912);
nand U27297 (N_27297,N_26357,N_26740);
nor U27298 (N_27298,N_26502,N_26735);
nand U27299 (N_27299,N_26150,N_26656);
nor U27300 (N_27300,N_26036,N_26506);
nor U27301 (N_27301,N_26103,N_26368);
xnor U27302 (N_27302,N_26018,N_26822);
nand U27303 (N_27303,N_26272,N_26865);
or U27304 (N_27304,N_26645,N_26551);
or U27305 (N_27305,N_26566,N_26487);
nand U27306 (N_27306,N_26894,N_26677);
xnor U27307 (N_27307,N_26988,N_26704);
xnor U27308 (N_27308,N_26026,N_26011);
nand U27309 (N_27309,N_26508,N_26222);
nor U27310 (N_27310,N_26014,N_26883);
xnor U27311 (N_27311,N_26788,N_26270);
and U27312 (N_27312,N_26105,N_26281);
nor U27313 (N_27313,N_26856,N_26354);
or U27314 (N_27314,N_26914,N_26549);
or U27315 (N_27315,N_26890,N_26298);
and U27316 (N_27316,N_26122,N_26102);
xor U27317 (N_27317,N_26760,N_26343);
or U27318 (N_27318,N_26358,N_26097);
nor U27319 (N_27319,N_26184,N_26598);
and U27320 (N_27320,N_26295,N_26394);
xnor U27321 (N_27321,N_26694,N_26777);
or U27322 (N_27322,N_26418,N_26574);
nor U27323 (N_27323,N_26306,N_26673);
xor U27324 (N_27324,N_26069,N_26260);
nor U27325 (N_27325,N_26169,N_26087);
or U27326 (N_27326,N_26706,N_26950);
xnor U27327 (N_27327,N_26518,N_26868);
nor U27328 (N_27328,N_26213,N_26964);
nor U27329 (N_27329,N_26770,N_26007);
xor U27330 (N_27330,N_26127,N_26489);
nor U27331 (N_27331,N_26933,N_26003);
and U27332 (N_27332,N_26118,N_26144);
and U27333 (N_27333,N_26170,N_26437);
nor U27334 (N_27334,N_26523,N_26335);
nand U27335 (N_27335,N_26218,N_26214);
xnor U27336 (N_27336,N_26153,N_26278);
and U27337 (N_27337,N_26985,N_26527);
or U27338 (N_27338,N_26393,N_26701);
and U27339 (N_27339,N_26552,N_26623);
nand U27340 (N_27340,N_26672,N_26949);
nand U27341 (N_27341,N_26847,N_26748);
nand U27342 (N_27342,N_26034,N_26963);
nand U27343 (N_27343,N_26718,N_26257);
xnor U27344 (N_27344,N_26562,N_26818);
nor U27345 (N_27345,N_26046,N_26986);
and U27346 (N_27346,N_26955,N_26098);
nand U27347 (N_27347,N_26989,N_26338);
nor U27348 (N_27348,N_26324,N_26782);
nand U27349 (N_27349,N_26254,N_26650);
xor U27350 (N_27350,N_26255,N_26956);
and U27351 (N_27351,N_26816,N_26160);
xor U27352 (N_27352,N_26674,N_26059);
or U27353 (N_27353,N_26965,N_26138);
and U27354 (N_27354,N_26217,N_26813);
and U27355 (N_27355,N_26657,N_26420);
nand U27356 (N_27356,N_26498,N_26187);
nor U27357 (N_27357,N_26145,N_26463);
nand U27358 (N_27358,N_26951,N_26702);
and U27359 (N_27359,N_26407,N_26315);
and U27360 (N_27360,N_26852,N_26494);
nand U27361 (N_27361,N_26943,N_26785);
nor U27362 (N_27362,N_26465,N_26307);
or U27363 (N_27363,N_26078,N_26404);
and U27364 (N_27364,N_26896,N_26576);
and U27365 (N_27365,N_26172,N_26617);
nor U27366 (N_27366,N_26897,N_26593);
or U27367 (N_27367,N_26944,N_26142);
and U27368 (N_27368,N_26186,N_26436);
or U27369 (N_27369,N_26104,N_26080);
or U27370 (N_27370,N_26231,N_26108);
and U27371 (N_27371,N_26878,N_26230);
nor U27372 (N_27372,N_26971,N_26334);
xor U27373 (N_27373,N_26345,N_26568);
xnor U27374 (N_27374,N_26447,N_26072);
or U27375 (N_27375,N_26241,N_26265);
and U27376 (N_27376,N_26221,N_26035);
nor U27377 (N_27377,N_26901,N_26406);
nor U27378 (N_27378,N_26331,N_26004);
nor U27379 (N_27379,N_26403,N_26841);
nand U27380 (N_27380,N_26640,N_26537);
xnor U27381 (N_27381,N_26781,N_26313);
and U27382 (N_27382,N_26758,N_26855);
or U27383 (N_27383,N_26346,N_26309);
xnor U27384 (N_27384,N_26691,N_26092);
or U27385 (N_27385,N_26519,N_26466);
and U27386 (N_27386,N_26606,N_26216);
nor U27387 (N_27387,N_26373,N_26253);
nand U27388 (N_27388,N_26299,N_26074);
xnor U27389 (N_27389,N_26446,N_26304);
or U27390 (N_27390,N_26091,N_26021);
xnor U27391 (N_27391,N_26843,N_26139);
or U27392 (N_27392,N_26320,N_26550);
and U27393 (N_27393,N_26638,N_26239);
nand U27394 (N_27394,N_26383,N_26737);
or U27395 (N_27395,N_26795,N_26392);
nand U27396 (N_27396,N_26193,N_26013);
and U27397 (N_27397,N_26226,N_26554);
and U27398 (N_27398,N_26805,N_26887);
nor U27399 (N_27399,N_26716,N_26052);
nand U27400 (N_27400,N_26937,N_26294);
nand U27401 (N_27401,N_26675,N_26745);
and U27402 (N_27402,N_26803,N_26006);
and U27403 (N_27403,N_26906,N_26996);
nor U27404 (N_27404,N_26807,N_26591);
and U27405 (N_27405,N_26600,N_26579);
nor U27406 (N_27406,N_26201,N_26410);
xnor U27407 (N_27407,N_26659,N_26237);
xor U27408 (N_27408,N_26823,N_26347);
or U27409 (N_27409,N_26377,N_26360);
and U27410 (N_27410,N_26668,N_26408);
nand U27411 (N_27411,N_26729,N_26250);
nand U27412 (N_27412,N_26197,N_26366);
nor U27413 (N_27413,N_26661,N_26276);
nor U27414 (N_27414,N_26062,N_26649);
nor U27415 (N_27415,N_26667,N_26202);
nand U27416 (N_27416,N_26311,N_26135);
nor U27417 (N_27417,N_26263,N_26168);
and U27418 (N_27418,N_26590,N_26223);
nor U27419 (N_27419,N_26599,N_26686);
or U27420 (N_27420,N_26094,N_26797);
xor U27421 (N_27421,N_26195,N_26900);
nand U27422 (N_27422,N_26723,N_26459);
or U27423 (N_27423,N_26738,N_26076);
nand U27424 (N_27424,N_26198,N_26622);
and U27425 (N_27425,N_26670,N_26533);
or U27426 (N_27426,N_26131,N_26825);
and U27427 (N_27427,N_26531,N_26381);
nor U27428 (N_27428,N_26053,N_26907);
xor U27429 (N_27429,N_26086,N_26247);
or U27430 (N_27430,N_26891,N_26428);
and U27431 (N_27431,N_26458,N_26984);
nand U27432 (N_27432,N_26757,N_26733);
and U27433 (N_27433,N_26117,N_26109);
nand U27434 (N_27434,N_26917,N_26341);
nand U27435 (N_27435,N_26134,N_26826);
and U27436 (N_27436,N_26994,N_26386);
xnor U27437 (N_27437,N_26348,N_26516);
nand U27438 (N_27438,N_26830,N_26525);
nor U27439 (N_27439,N_26620,N_26695);
or U27440 (N_27440,N_26862,N_26611);
nor U27441 (N_27441,N_26882,N_26055);
nor U27442 (N_27442,N_26126,N_26037);
nand U27443 (N_27443,N_26959,N_26451);
nor U27444 (N_27444,N_26934,N_26775);
or U27445 (N_27445,N_26249,N_26698);
xnor U27446 (N_27446,N_26033,N_26513);
or U27447 (N_27447,N_26870,N_26460);
and U27448 (N_27448,N_26842,N_26556);
or U27449 (N_27449,N_26419,N_26827);
xor U27450 (N_27450,N_26176,N_26800);
nand U27451 (N_27451,N_26167,N_26921);
xnor U27452 (N_27452,N_26789,N_26610);
nor U27453 (N_27453,N_26688,N_26083);
xnor U27454 (N_27454,N_26246,N_26945);
or U27455 (N_27455,N_26604,N_26107);
nor U27456 (N_27456,N_26044,N_26762);
and U27457 (N_27457,N_26586,N_26747);
or U27458 (N_27458,N_26204,N_26967);
xor U27459 (N_27459,N_26560,N_26040);
xnor U27460 (N_27460,N_26262,N_26484);
nand U27461 (N_27461,N_26012,N_26236);
xnor U27462 (N_27462,N_26462,N_26585);
nor U27463 (N_27463,N_26573,N_26924);
or U27464 (N_27464,N_26208,N_26183);
nor U27465 (N_27465,N_26233,N_26832);
nand U27466 (N_27466,N_26850,N_26364);
or U27467 (N_27467,N_26849,N_26751);
or U27468 (N_27468,N_26595,N_26478);
or U27469 (N_27469,N_26926,N_26867);
or U27470 (N_27470,N_26699,N_26561);
nand U27471 (N_27471,N_26159,N_26734);
nand U27472 (N_27472,N_26414,N_26731);
nand U27473 (N_27473,N_26899,N_26680);
nor U27474 (N_27474,N_26719,N_26180);
or U27475 (N_27475,N_26676,N_26275);
and U27476 (N_27476,N_26821,N_26935);
and U27477 (N_27477,N_26507,N_26028);
nand U27478 (N_27478,N_26919,N_26910);
nor U27479 (N_27479,N_26220,N_26828);
nand U27480 (N_27480,N_26705,N_26961);
nand U27481 (N_27481,N_26749,N_26480);
nor U27482 (N_27482,N_26274,N_26065);
and U27483 (N_27483,N_26845,N_26472);
and U27484 (N_27484,N_26395,N_26759);
xor U27485 (N_27485,N_26405,N_26010);
nand U27486 (N_27486,N_26124,N_26209);
nor U27487 (N_27487,N_26547,N_26024);
and U27488 (N_27488,N_26129,N_26548);
and U27489 (N_27489,N_26730,N_26514);
xor U27490 (N_27490,N_26284,N_26027);
nor U27491 (N_27491,N_26512,N_26982);
nor U27492 (N_27492,N_26258,N_26025);
xor U27493 (N_27493,N_26125,N_26362);
nor U27494 (N_27494,N_26811,N_26372);
xnor U27495 (N_27495,N_26639,N_26397);
nor U27496 (N_27496,N_26848,N_26277);
or U27497 (N_27497,N_26779,N_26689);
nand U27498 (N_27498,N_26146,N_26916);
nor U27499 (N_27499,N_26616,N_26002);
and U27500 (N_27500,N_26655,N_26192);
nor U27501 (N_27501,N_26411,N_26827);
and U27502 (N_27502,N_26520,N_26592);
and U27503 (N_27503,N_26672,N_26771);
nor U27504 (N_27504,N_26742,N_26784);
xor U27505 (N_27505,N_26309,N_26423);
nand U27506 (N_27506,N_26684,N_26341);
and U27507 (N_27507,N_26733,N_26046);
nor U27508 (N_27508,N_26558,N_26962);
or U27509 (N_27509,N_26084,N_26552);
xnor U27510 (N_27510,N_26408,N_26562);
nor U27511 (N_27511,N_26899,N_26202);
or U27512 (N_27512,N_26262,N_26887);
and U27513 (N_27513,N_26917,N_26709);
nand U27514 (N_27514,N_26054,N_26379);
or U27515 (N_27515,N_26677,N_26099);
xnor U27516 (N_27516,N_26348,N_26610);
xnor U27517 (N_27517,N_26398,N_26883);
or U27518 (N_27518,N_26842,N_26571);
nand U27519 (N_27519,N_26679,N_26737);
and U27520 (N_27520,N_26981,N_26778);
nor U27521 (N_27521,N_26022,N_26817);
nand U27522 (N_27522,N_26757,N_26217);
nor U27523 (N_27523,N_26863,N_26096);
nor U27524 (N_27524,N_26033,N_26933);
or U27525 (N_27525,N_26459,N_26211);
nor U27526 (N_27526,N_26560,N_26582);
and U27527 (N_27527,N_26394,N_26489);
xnor U27528 (N_27528,N_26715,N_26897);
and U27529 (N_27529,N_26989,N_26291);
or U27530 (N_27530,N_26434,N_26147);
nand U27531 (N_27531,N_26373,N_26212);
and U27532 (N_27532,N_26139,N_26408);
xnor U27533 (N_27533,N_26331,N_26977);
or U27534 (N_27534,N_26486,N_26527);
xnor U27535 (N_27535,N_26106,N_26395);
xnor U27536 (N_27536,N_26212,N_26416);
or U27537 (N_27537,N_26622,N_26802);
nor U27538 (N_27538,N_26646,N_26317);
and U27539 (N_27539,N_26889,N_26966);
nand U27540 (N_27540,N_26379,N_26383);
nand U27541 (N_27541,N_26617,N_26554);
xor U27542 (N_27542,N_26902,N_26874);
or U27543 (N_27543,N_26907,N_26670);
xnor U27544 (N_27544,N_26508,N_26645);
or U27545 (N_27545,N_26601,N_26302);
or U27546 (N_27546,N_26116,N_26089);
nor U27547 (N_27547,N_26472,N_26874);
xnor U27548 (N_27548,N_26356,N_26086);
xor U27549 (N_27549,N_26834,N_26098);
nor U27550 (N_27550,N_26211,N_26282);
nand U27551 (N_27551,N_26173,N_26236);
or U27552 (N_27552,N_26341,N_26752);
nor U27553 (N_27553,N_26486,N_26750);
xnor U27554 (N_27554,N_26573,N_26659);
nand U27555 (N_27555,N_26279,N_26029);
or U27556 (N_27556,N_26664,N_26383);
and U27557 (N_27557,N_26596,N_26349);
nor U27558 (N_27558,N_26236,N_26392);
nand U27559 (N_27559,N_26590,N_26719);
nand U27560 (N_27560,N_26051,N_26042);
xnor U27561 (N_27561,N_26415,N_26541);
nand U27562 (N_27562,N_26777,N_26322);
or U27563 (N_27563,N_26364,N_26959);
and U27564 (N_27564,N_26743,N_26445);
xor U27565 (N_27565,N_26659,N_26035);
and U27566 (N_27566,N_26406,N_26362);
nand U27567 (N_27567,N_26642,N_26717);
nand U27568 (N_27568,N_26759,N_26881);
or U27569 (N_27569,N_26879,N_26509);
or U27570 (N_27570,N_26403,N_26724);
nor U27571 (N_27571,N_26268,N_26975);
or U27572 (N_27572,N_26793,N_26092);
and U27573 (N_27573,N_26587,N_26430);
nand U27574 (N_27574,N_26895,N_26181);
or U27575 (N_27575,N_26846,N_26150);
nand U27576 (N_27576,N_26129,N_26440);
nor U27577 (N_27577,N_26612,N_26126);
or U27578 (N_27578,N_26998,N_26684);
nor U27579 (N_27579,N_26845,N_26587);
xnor U27580 (N_27580,N_26140,N_26321);
or U27581 (N_27581,N_26100,N_26609);
and U27582 (N_27582,N_26072,N_26065);
xnor U27583 (N_27583,N_26525,N_26074);
and U27584 (N_27584,N_26636,N_26689);
nand U27585 (N_27585,N_26576,N_26038);
nor U27586 (N_27586,N_26498,N_26106);
nand U27587 (N_27587,N_26945,N_26132);
or U27588 (N_27588,N_26499,N_26093);
nand U27589 (N_27589,N_26645,N_26950);
nor U27590 (N_27590,N_26463,N_26280);
or U27591 (N_27591,N_26111,N_26417);
nand U27592 (N_27592,N_26634,N_26287);
or U27593 (N_27593,N_26854,N_26901);
nand U27594 (N_27594,N_26287,N_26801);
and U27595 (N_27595,N_26376,N_26166);
nand U27596 (N_27596,N_26293,N_26002);
nor U27597 (N_27597,N_26851,N_26719);
xnor U27598 (N_27598,N_26855,N_26604);
or U27599 (N_27599,N_26356,N_26307);
nor U27600 (N_27600,N_26788,N_26975);
and U27601 (N_27601,N_26701,N_26861);
xnor U27602 (N_27602,N_26538,N_26609);
nand U27603 (N_27603,N_26413,N_26040);
and U27604 (N_27604,N_26938,N_26054);
and U27605 (N_27605,N_26797,N_26474);
or U27606 (N_27606,N_26767,N_26624);
nor U27607 (N_27607,N_26728,N_26867);
nand U27608 (N_27608,N_26385,N_26759);
and U27609 (N_27609,N_26873,N_26906);
xor U27610 (N_27610,N_26341,N_26087);
nor U27611 (N_27611,N_26555,N_26558);
and U27612 (N_27612,N_26681,N_26173);
nor U27613 (N_27613,N_26470,N_26159);
and U27614 (N_27614,N_26673,N_26143);
xnor U27615 (N_27615,N_26996,N_26528);
or U27616 (N_27616,N_26835,N_26317);
nand U27617 (N_27617,N_26226,N_26618);
nor U27618 (N_27618,N_26418,N_26608);
nor U27619 (N_27619,N_26017,N_26610);
nor U27620 (N_27620,N_26037,N_26824);
nand U27621 (N_27621,N_26724,N_26863);
xnor U27622 (N_27622,N_26847,N_26956);
nand U27623 (N_27623,N_26234,N_26059);
nand U27624 (N_27624,N_26803,N_26772);
nand U27625 (N_27625,N_26313,N_26922);
nand U27626 (N_27626,N_26748,N_26205);
nor U27627 (N_27627,N_26003,N_26843);
or U27628 (N_27628,N_26205,N_26156);
or U27629 (N_27629,N_26906,N_26578);
nor U27630 (N_27630,N_26398,N_26528);
nor U27631 (N_27631,N_26673,N_26798);
and U27632 (N_27632,N_26367,N_26285);
and U27633 (N_27633,N_26256,N_26071);
xor U27634 (N_27634,N_26438,N_26688);
or U27635 (N_27635,N_26966,N_26623);
nor U27636 (N_27636,N_26311,N_26982);
nor U27637 (N_27637,N_26489,N_26986);
and U27638 (N_27638,N_26125,N_26590);
and U27639 (N_27639,N_26970,N_26549);
nand U27640 (N_27640,N_26234,N_26372);
and U27641 (N_27641,N_26762,N_26634);
or U27642 (N_27642,N_26623,N_26523);
or U27643 (N_27643,N_26552,N_26686);
or U27644 (N_27644,N_26536,N_26838);
and U27645 (N_27645,N_26381,N_26475);
xnor U27646 (N_27646,N_26552,N_26577);
or U27647 (N_27647,N_26984,N_26095);
or U27648 (N_27648,N_26798,N_26381);
xnor U27649 (N_27649,N_26381,N_26705);
nand U27650 (N_27650,N_26921,N_26079);
and U27651 (N_27651,N_26380,N_26954);
nand U27652 (N_27652,N_26273,N_26407);
and U27653 (N_27653,N_26862,N_26790);
nand U27654 (N_27654,N_26372,N_26026);
and U27655 (N_27655,N_26761,N_26655);
and U27656 (N_27656,N_26321,N_26049);
or U27657 (N_27657,N_26915,N_26535);
and U27658 (N_27658,N_26130,N_26131);
or U27659 (N_27659,N_26237,N_26608);
xnor U27660 (N_27660,N_26262,N_26081);
or U27661 (N_27661,N_26811,N_26582);
and U27662 (N_27662,N_26281,N_26657);
and U27663 (N_27663,N_26143,N_26906);
or U27664 (N_27664,N_26378,N_26613);
and U27665 (N_27665,N_26862,N_26935);
xnor U27666 (N_27666,N_26354,N_26126);
nor U27667 (N_27667,N_26628,N_26973);
nor U27668 (N_27668,N_26348,N_26117);
nor U27669 (N_27669,N_26218,N_26946);
nor U27670 (N_27670,N_26884,N_26271);
and U27671 (N_27671,N_26125,N_26662);
or U27672 (N_27672,N_26016,N_26726);
nand U27673 (N_27673,N_26052,N_26365);
and U27674 (N_27674,N_26499,N_26256);
xnor U27675 (N_27675,N_26615,N_26593);
or U27676 (N_27676,N_26003,N_26068);
or U27677 (N_27677,N_26161,N_26091);
xor U27678 (N_27678,N_26227,N_26695);
or U27679 (N_27679,N_26146,N_26630);
nand U27680 (N_27680,N_26453,N_26099);
or U27681 (N_27681,N_26305,N_26903);
nand U27682 (N_27682,N_26550,N_26121);
and U27683 (N_27683,N_26685,N_26262);
nand U27684 (N_27684,N_26355,N_26595);
nand U27685 (N_27685,N_26143,N_26829);
nor U27686 (N_27686,N_26051,N_26432);
nor U27687 (N_27687,N_26492,N_26693);
nor U27688 (N_27688,N_26790,N_26566);
and U27689 (N_27689,N_26360,N_26902);
xnor U27690 (N_27690,N_26976,N_26089);
nor U27691 (N_27691,N_26344,N_26063);
and U27692 (N_27692,N_26539,N_26658);
and U27693 (N_27693,N_26454,N_26995);
xor U27694 (N_27694,N_26762,N_26091);
xor U27695 (N_27695,N_26160,N_26401);
nor U27696 (N_27696,N_26780,N_26247);
nand U27697 (N_27697,N_26284,N_26861);
or U27698 (N_27698,N_26343,N_26750);
and U27699 (N_27699,N_26252,N_26268);
nor U27700 (N_27700,N_26043,N_26852);
nor U27701 (N_27701,N_26804,N_26738);
and U27702 (N_27702,N_26203,N_26328);
xor U27703 (N_27703,N_26706,N_26692);
and U27704 (N_27704,N_26446,N_26408);
xor U27705 (N_27705,N_26207,N_26071);
nor U27706 (N_27706,N_26091,N_26958);
xnor U27707 (N_27707,N_26080,N_26985);
and U27708 (N_27708,N_26753,N_26026);
xor U27709 (N_27709,N_26563,N_26208);
or U27710 (N_27710,N_26317,N_26455);
and U27711 (N_27711,N_26433,N_26287);
nand U27712 (N_27712,N_26060,N_26842);
xnor U27713 (N_27713,N_26397,N_26617);
or U27714 (N_27714,N_26583,N_26843);
xnor U27715 (N_27715,N_26144,N_26436);
nor U27716 (N_27716,N_26494,N_26329);
nand U27717 (N_27717,N_26065,N_26118);
or U27718 (N_27718,N_26882,N_26906);
nor U27719 (N_27719,N_26045,N_26258);
nor U27720 (N_27720,N_26818,N_26555);
nor U27721 (N_27721,N_26023,N_26180);
nor U27722 (N_27722,N_26797,N_26361);
nor U27723 (N_27723,N_26413,N_26017);
nor U27724 (N_27724,N_26161,N_26457);
xor U27725 (N_27725,N_26220,N_26221);
or U27726 (N_27726,N_26012,N_26745);
or U27727 (N_27727,N_26680,N_26430);
or U27728 (N_27728,N_26687,N_26164);
and U27729 (N_27729,N_26289,N_26988);
xnor U27730 (N_27730,N_26293,N_26554);
nor U27731 (N_27731,N_26893,N_26750);
and U27732 (N_27732,N_26083,N_26638);
and U27733 (N_27733,N_26040,N_26479);
nand U27734 (N_27734,N_26177,N_26931);
or U27735 (N_27735,N_26287,N_26996);
or U27736 (N_27736,N_26567,N_26236);
nor U27737 (N_27737,N_26243,N_26882);
and U27738 (N_27738,N_26242,N_26672);
or U27739 (N_27739,N_26854,N_26435);
xnor U27740 (N_27740,N_26524,N_26068);
and U27741 (N_27741,N_26717,N_26826);
xnor U27742 (N_27742,N_26344,N_26450);
or U27743 (N_27743,N_26682,N_26093);
nor U27744 (N_27744,N_26946,N_26063);
xnor U27745 (N_27745,N_26139,N_26804);
xor U27746 (N_27746,N_26817,N_26214);
nor U27747 (N_27747,N_26850,N_26006);
and U27748 (N_27748,N_26224,N_26123);
xnor U27749 (N_27749,N_26479,N_26265);
nand U27750 (N_27750,N_26328,N_26478);
nand U27751 (N_27751,N_26947,N_26305);
xor U27752 (N_27752,N_26456,N_26435);
and U27753 (N_27753,N_26517,N_26958);
nor U27754 (N_27754,N_26001,N_26487);
nor U27755 (N_27755,N_26056,N_26895);
nand U27756 (N_27756,N_26095,N_26581);
or U27757 (N_27757,N_26135,N_26853);
nor U27758 (N_27758,N_26396,N_26675);
xnor U27759 (N_27759,N_26659,N_26909);
and U27760 (N_27760,N_26214,N_26169);
or U27761 (N_27761,N_26599,N_26972);
and U27762 (N_27762,N_26111,N_26393);
or U27763 (N_27763,N_26641,N_26196);
nand U27764 (N_27764,N_26202,N_26083);
nand U27765 (N_27765,N_26321,N_26293);
nand U27766 (N_27766,N_26109,N_26329);
or U27767 (N_27767,N_26889,N_26928);
nor U27768 (N_27768,N_26951,N_26731);
nor U27769 (N_27769,N_26690,N_26601);
nor U27770 (N_27770,N_26059,N_26706);
nor U27771 (N_27771,N_26003,N_26495);
xnor U27772 (N_27772,N_26842,N_26362);
or U27773 (N_27773,N_26776,N_26275);
and U27774 (N_27774,N_26861,N_26110);
and U27775 (N_27775,N_26461,N_26537);
or U27776 (N_27776,N_26350,N_26383);
or U27777 (N_27777,N_26940,N_26945);
xnor U27778 (N_27778,N_26010,N_26303);
or U27779 (N_27779,N_26836,N_26403);
and U27780 (N_27780,N_26139,N_26763);
nand U27781 (N_27781,N_26356,N_26661);
nor U27782 (N_27782,N_26355,N_26921);
xnor U27783 (N_27783,N_26546,N_26818);
xnor U27784 (N_27784,N_26503,N_26979);
or U27785 (N_27785,N_26465,N_26150);
nor U27786 (N_27786,N_26405,N_26100);
nand U27787 (N_27787,N_26574,N_26828);
or U27788 (N_27788,N_26692,N_26392);
nor U27789 (N_27789,N_26491,N_26876);
nand U27790 (N_27790,N_26442,N_26871);
and U27791 (N_27791,N_26718,N_26804);
nor U27792 (N_27792,N_26160,N_26683);
or U27793 (N_27793,N_26220,N_26048);
nor U27794 (N_27794,N_26152,N_26484);
and U27795 (N_27795,N_26901,N_26760);
xor U27796 (N_27796,N_26974,N_26133);
xnor U27797 (N_27797,N_26659,N_26712);
and U27798 (N_27798,N_26126,N_26547);
and U27799 (N_27799,N_26431,N_26158);
nor U27800 (N_27800,N_26375,N_26069);
xor U27801 (N_27801,N_26867,N_26128);
and U27802 (N_27802,N_26702,N_26404);
and U27803 (N_27803,N_26112,N_26013);
xor U27804 (N_27804,N_26042,N_26996);
and U27805 (N_27805,N_26107,N_26017);
nand U27806 (N_27806,N_26255,N_26959);
xnor U27807 (N_27807,N_26364,N_26197);
or U27808 (N_27808,N_26602,N_26090);
nand U27809 (N_27809,N_26579,N_26850);
and U27810 (N_27810,N_26625,N_26889);
or U27811 (N_27811,N_26800,N_26398);
nor U27812 (N_27812,N_26829,N_26710);
nor U27813 (N_27813,N_26754,N_26675);
or U27814 (N_27814,N_26068,N_26955);
xor U27815 (N_27815,N_26264,N_26913);
nand U27816 (N_27816,N_26314,N_26115);
and U27817 (N_27817,N_26798,N_26509);
nand U27818 (N_27818,N_26364,N_26800);
and U27819 (N_27819,N_26916,N_26591);
and U27820 (N_27820,N_26992,N_26297);
xor U27821 (N_27821,N_26395,N_26940);
or U27822 (N_27822,N_26053,N_26424);
nor U27823 (N_27823,N_26729,N_26348);
nor U27824 (N_27824,N_26621,N_26961);
or U27825 (N_27825,N_26928,N_26822);
nor U27826 (N_27826,N_26125,N_26855);
nor U27827 (N_27827,N_26188,N_26639);
nor U27828 (N_27828,N_26315,N_26062);
nand U27829 (N_27829,N_26742,N_26297);
and U27830 (N_27830,N_26565,N_26317);
nand U27831 (N_27831,N_26384,N_26351);
nand U27832 (N_27832,N_26316,N_26094);
nor U27833 (N_27833,N_26684,N_26663);
nor U27834 (N_27834,N_26880,N_26661);
and U27835 (N_27835,N_26337,N_26813);
nor U27836 (N_27836,N_26898,N_26473);
and U27837 (N_27837,N_26483,N_26636);
nor U27838 (N_27838,N_26088,N_26087);
xnor U27839 (N_27839,N_26509,N_26612);
nor U27840 (N_27840,N_26761,N_26836);
and U27841 (N_27841,N_26988,N_26477);
nand U27842 (N_27842,N_26659,N_26927);
nor U27843 (N_27843,N_26244,N_26298);
and U27844 (N_27844,N_26398,N_26230);
and U27845 (N_27845,N_26341,N_26787);
xnor U27846 (N_27846,N_26777,N_26939);
xnor U27847 (N_27847,N_26571,N_26981);
nor U27848 (N_27848,N_26496,N_26380);
or U27849 (N_27849,N_26444,N_26800);
and U27850 (N_27850,N_26359,N_26721);
and U27851 (N_27851,N_26999,N_26493);
and U27852 (N_27852,N_26746,N_26740);
nand U27853 (N_27853,N_26316,N_26471);
nor U27854 (N_27854,N_26864,N_26785);
xor U27855 (N_27855,N_26338,N_26075);
nor U27856 (N_27856,N_26519,N_26845);
nor U27857 (N_27857,N_26180,N_26313);
or U27858 (N_27858,N_26490,N_26174);
xnor U27859 (N_27859,N_26093,N_26249);
and U27860 (N_27860,N_26862,N_26268);
nor U27861 (N_27861,N_26099,N_26735);
nand U27862 (N_27862,N_26223,N_26071);
nor U27863 (N_27863,N_26774,N_26352);
and U27864 (N_27864,N_26740,N_26450);
nor U27865 (N_27865,N_26173,N_26825);
nand U27866 (N_27866,N_26831,N_26225);
and U27867 (N_27867,N_26862,N_26228);
or U27868 (N_27868,N_26929,N_26654);
and U27869 (N_27869,N_26898,N_26570);
xor U27870 (N_27870,N_26536,N_26534);
and U27871 (N_27871,N_26746,N_26967);
nor U27872 (N_27872,N_26226,N_26830);
xor U27873 (N_27873,N_26400,N_26848);
or U27874 (N_27874,N_26556,N_26252);
or U27875 (N_27875,N_26755,N_26252);
nor U27876 (N_27876,N_26452,N_26691);
xor U27877 (N_27877,N_26100,N_26975);
xnor U27878 (N_27878,N_26560,N_26462);
nand U27879 (N_27879,N_26112,N_26434);
xnor U27880 (N_27880,N_26016,N_26097);
nand U27881 (N_27881,N_26899,N_26536);
xnor U27882 (N_27882,N_26326,N_26796);
and U27883 (N_27883,N_26471,N_26434);
nand U27884 (N_27884,N_26425,N_26444);
and U27885 (N_27885,N_26041,N_26284);
nor U27886 (N_27886,N_26352,N_26589);
or U27887 (N_27887,N_26530,N_26718);
nor U27888 (N_27888,N_26258,N_26012);
or U27889 (N_27889,N_26953,N_26864);
and U27890 (N_27890,N_26715,N_26605);
nand U27891 (N_27891,N_26589,N_26432);
nor U27892 (N_27892,N_26771,N_26806);
or U27893 (N_27893,N_26109,N_26326);
nand U27894 (N_27894,N_26730,N_26336);
or U27895 (N_27895,N_26197,N_26230);
and U27896 (N_27896,N_26041,N_26063);
nor U27897 (N_27897,N_26234,N_26914);
xor U27898 (N_27898,N_26922,N_26062);
and U27899 (N_27899,N_26417,N_26738);
nor U27900 (N_27900,N_26943,N_26127);
xnor U27901 (N_27901,N_26358,N_26130);
and U27902 (N_27902,N_26148,N_26456);
or U27903 (N_27903,N_26180,N_26306);
nand U27904 (N_27904,N_26842,N_26365);
and U27905 (N_27905,N_26829,N_26168);
nor U27906 (N_27906,N_26226,N_26560);
xnor U27907 (N_27907,N_26691,N_26003);
nor U27908 (N_27908,N_26206,N_26638);
or U27909 (N_27909,N_26438,N_26936);
or U27910 (N_27910,N_26778,N_26211);
xnor U27911 (N_27911,N_26378,N_26518);
xor U27912 (N_27912,N_26956,N_26640);
nor U27913 (N_27913,N_26817,N_26566);
nand U27914 (N_27914,N_26757,N_26238);
or U27915 (N_27915,N_26033,N_26907);
nand U27916 (N_27916,N_26781,N_26504);
nor U27917 (N_27917,N_26930,N_26467);
or U27918 (N_27918,N_26841,N_26917);
nand U27919 (N_27919,N_26561,N_26417);
and U27920 (N_27920,N_26338,N_26803);
and U27921 (N_27921,N_26978,N_26208);
xor U27922 (N_27922,N_26432,N_26106);
nor U27923 (N_27923,N_26225,N_26090);
or U27924 (N_27924,N_26014,N_26629);
nor U27925 (N_27925,N_26798,N_26875);
and U27926 (N_27926,N_26973,N_26231);
nand U27927 (N_27927,N_26230,N_26412);
xor U27928 (N_27928,N_26152,N_26883);
and U27929 (N_27929,N_26889,N_26931);
and U27930 (N_27930,N_26446,N_26531);
and U27931 (N_27931,N_26545,N_26376);
nor U27932 (N_27932,N_26296,N_26098);
xnor U27933 (N_27933,N_26591,N_26776);
nor U27934 (N_27934,N_26279,N_26466);
xor U27935 (N_27935,N_26457,N_26606);
or U27936 (N_27936,N_26063,N_26385);
xnor U27937 (N_27937,N_26162,N_26800);
or U27938 (N_27938,N_26335,N_26708);
nor U27939 (N_27939,N_26425,N_26196);
and U27940 (N_27940,N_26192,N_26208);
xor U27941 (N_27941,N_26389,N_26701);
and U27942 (N_27942,N_26881,N_26616);
nor U27943 (N_27943,N_26668,N_26247);
and U27944 (N_27944,N_26542,N_26354);
and U27945 (N_27945,N_26605,N_26539);
xnor U27946 (N_27946,N_26747,N_26447);
nor U27947 (N_27947,N_26736,N_26095);
and U27948 (N_27948,N_26878,N_26863);
and U27949 (N_27949,N_26814,N_26603);
or U27950 (N_27950,N_26157,N_26248);
nor U27951 (N_27951,N_26232,N_26449);
xor U27952 (N_27952,N_26365,N_26088);
or U27953 (N_27953,N_26208,N_26935);
nand U27954 (N_27954,N_26470,N_26729);
or U27955 (N_27955,N_26302,N_26988);
and U27956 (N_27956,N_26925,N_26991);
and U27957 (N_27957,N_26600,N_26734);
or U27958 (N_27958,N_26677,N_26841);
nand U27959 (N_27959,N_26999,N_26797);
and U27960 (N_27960,N_26700,N_26775);
nor U27961 (N_27961,N_26148,N_26345);
xnor U27962 (N_27962,N_26357,N_26175);
and U27963 (N_27963,N_26430,N_26005);
or U27964 (N_27964,N_26945,N_26192);
nor U27965 (N_27965,N_26179,N_26767);
nor U27966 (N_27966,N_26730,N_26110);
nor U27967 (N_27967,N_26255,N_26136);
xor U27968 (N_27968,N_26024,N_26754);
nand U27969 (N_27969,N_26621,N_26546);
xor U27970 (N_27970,N_26783,N_26539);
and U27971 (N_27971,N_26143,N_26616);
nor U27972 (N_27972,N_26290,N_26094);
and U27973 (N_27973,N_26611,N_26050);
and U27974 (N_27974,N_26631,N_26132);
nor U27975 (N_27975,N_26509,N_26101);
and U27976 (N_27976,N_26623,N_26379);
nor U27977 (N_27977,N_26850,N_26008);
xnor U27978 (N_27978,N_26203,N_26381);
xnor U27979 (N_27979,N_26602,N_26400);
nand U27980 (N_27980,N_26444,N_26915);
nor U27981 (N_27981,N_26633,N_26958);
and U27982 (N_27982,N_26396,N_26295);
nor U27983 (N_27983,N_26302,N_26918);
xor U27984 (N_27984,N_26481,N_26740);
nor U27985 (N_27985,N_26793,N_26771);
and U27986 (N_27986,N_26085,N_26014);
nor U27987 (N_27987,N_26116,N_26986);
xor U27988 (N_27988,N_26771,N_26032);
xnor U27989 (N_27989,N_26201,N_26866);
nor U27990 (N_27990,N_26282,N_26128);
nand U27991 (N_27991,N_26919,N_26055);
nor U27992 (N_27992,N_26354,N_26411);
nor U27993 (N_27993,N_26479,N_26607);
xnor U27994 (N_27994,N_26490,N_26065);
xor U27995 (N_27995,N_26870,N_26170);
or U27996 (N_27996,N_26163,N_26568);
nor U27997 (N_27997,N_26080,N_26328);
or U27998 (N_27998,N_26356,N_26810);
nand U27999 (N_27999,N_26968,N_26877);
or U28000 (N_28000,N_27731,N_27460);
and U28001 (N_28001,N_27907,N_27424);
and U28002 (N_28002,N_27482,N_27880);
or U28003 (N_28003,N_27867,N_27374);
and U28004 (N_28004,N_27170,N_27008);
or U28005 (N_28005,N_27293,N_27646);
nor U28006 (N_28006,N_27135,N_27933);
xor U28007 (N_28007,N_27471,N_27048);
xor U28008 (N_28008,N_27288,N_27510);
nor U28009 (N_28009,N_27743,N_27352);
and U28010 (N_28010,N_27379,N_27409);
and U28011 (N_28011,N_27014,N_27676);
nand U28012 (N_28012,N_27000,N_27452);
and U28013 (N_28013,N_27323,N_27446);
and U28014 (N_28014,N_27702,N_27234);
and U28015 (N_28015,N_27984,N_27146);
nand U28016 (N_28016,N_27613,N_27378);
nor U28017 (N_28017,N_27227,N_27204);
nor U28018 (N_28018,N_27007,N_27531);
nor U28019 (N_28019,N_27728,N_27775);
nor U28020 (N_28020,N_27061,N_27607);
or U28021 (N_28021,N_27395,N_27079);
or U28022 (N_28022,N_27666,N_27372);
nand U28023 (N_28023,N_27337,N_27053);
xnor U28024 (N_28024,N_27756,N_27312);
nor U28025 (N_28025,N_27611,N_27050);
xnor U28026 (N_28026,N_27939,N_27035);
nand U28027 (N_28027,N_27125,N_27417);
nand U28028 (N_28028,N_27366,N_27650);
nor U28029 (N_28029,N_27967,N_27310);
and U28030 (N_28030,N_27259,N_27391);
xor U28031 (N_28031,N_27441,N_27322);
xnor U28032 (N_28032,N_27023,N_27275);
nand U28033 (N_28033,N_27506,N_27705);
nand U28034 (N_28034,N_27747,N_27104);
nand U28035 (N_28035,N_27548,N_27016);
or U28036 (N_28036,N_27997,N_27658);
nand U28037 (N_28037,N_27052,N_27484);
xor U28038 (N_28038,N_27988,N_27044);
or U28039 (N_28039,N_27265,N_27041);
xor U28040 (N_28040,N_27771,N_27464);
nand U28041 (N_28041,N_27882,N_27573);
and U28042 (N_28042,N_27225,N_27869);
nand U28043 (N_28043,N_27892,N_27586);
and U28044 (N_28044,N_27371,N_27431);
xnor U28045 (N_28045,N_27303,N_27526);
nand U28046 (N_28046,N_27049,N_27317);
xnor U28047 (N_28047,N_27752,N_27037);
and U28048 (N_28048,N_27365,N_27147);
or U28049 (N_28049,N_27924,N_27836);
nand U28050 (N_28050,N_27354,N_27885);
and U28051 (N_28051,N_27191,N_27628);
xor U28052 (N_28052,N_27179,N_27311);
nand U28053 (N_28053,N_27338,N_27358);
or U28054 (N_28054,N_27690,N_27392);
nand U28055 (N_28055,N_27339,N_27580);
xnor U28056 (N_28056,N_27797,N_27152);
nor U28057 (N_28057,N_27999,N_27544);
xor U28058 (N_28058,N_27952,N_27645);
xnor U28059 (N_28059,N_27261,N_27381);
and U28060 (N_28060,N_27958,N_27438);
nor U28061 (N_28061,N_27759,N_27746);
xnor U28062 (N_28062,N_27382,N_27272);
nand U28063 (N_28063,N_27683,N_27951);
nor U28064 (N_28064,N_27214,N_27551);
and U28065 (N_28065,N_27130,N_27782);
nand U28066 (N_28066,N_27964,N_27855);
nor U28067 (N_28067,N_27292,N_27886);
nand U28068 (N_28068,N_27300,N_27659);
or U28069 (N_28069,N_27238,N_27220);
nand U28070 (N_28070,N_27440,N_27593);
or U28071 (N_28071,N_27554,N_27149);
or U28072 (N_28072,N_27437,N_27983);
and U28073 (N_28073,N_27900,N_27282);
xnor U28074 (N_28074,N_27472,N_27533);
xor U28075 (N_28075,N_27183,N_27257);
xor U28076 (N_28076,N_27560,N_27973);
and U28077 (N_28077,N_27162,N_27725);
or U28078 (N_28078,N_27173,N_27156);
or U28079 (N_28079,N_27062,N_27218);
nor U28080 (N_28080,N_27652,N_27215);
and U28081 (N_28081,N_27477,N_27109);
nor U28082 (N_28082,N_27516,N_27271);
xnor U28083 (N_28083,N_27622,N_27080);
nor U28084 (N_28084,N_27093,N_27833);
xor U28085 (N_28085,N_27263,N_27071);
nand U28086 (N_28086,N_27821,N_27587);
nand U28087 (N_28087,N_27253,N_27945);
nor U28088 (N_28088,N_27793,N_27153);
and U28089 (N_28089,N_27298,N_27831);
and U28090 (N_28090,N_27995,N_27091);
or U28091 (N_28091,N_27588,N_27647);
nor U28092 (N_28092,N_27709,N_27333);
nor U28093 (N_28093,N_27235,N_27331);
xor U28094 (N_28094,N_27577,N_27851);
and U28095 (N_28095,N_27555,N_27631);
and U28096 (N_28096,N_27405,N_27013);
nand U28097 (N_28097,N_27115,N_27626);
xor U28098 (N_28098,N_27906,N_27154);
nor U28099 (N_28099,N_27783,N_27325);
nand U28100 (N_28100,N_27615,N_27329);
and U28101 (N_28101,N_27345,N_27285);
nor U28102 (N_28102,N_27874,N_27736);
nand U28103 (N_28103,N_27595,N_27565);
or U28104 (N_28104,N_27534,N_27066);
and U28105 (N_28105,N_27915,N_27419);
nor U28106 (N_28106,N_27639,N_27277);
nor U28107 (N_28107,N_27734,N_27972);
or U28108 (N_28108,N_27875,N_27081);
or U28109 (N_28109,N_27503,N_27667);
nand U28110 (N_28110,N_27584,N_27627);
and U28111 (N_28111,N_27180,N_27742);
or U28112 (N_28112,N_27753,N_27059);
nor U28113 (N_28113,N_27136,N_27027);
nand U28114 (N_28114,N_27530,N_27818);
xnor U28115 (N_28115,N_27456,N_27172);
nand U28116 (N_28116,N_27582,N_27523);
nand U28117 (N_28117,N_27287,N_27262);
nand U28118 (N_28118,N_27996,N_27454);
xor U28119 (N_28119,N_27351,N_27450);
nor U28120 (N_28120,N_27096,N_27612);
or U28121 (N_28121,N_27436,N_27026);
or U28122 (N_28122,N_27765,N_27617);
nor U28123 (N_28123,N_27110,N_27866);
xnor U28124 (N_28124,N_27657,N_27228);
and U28125 (N_28125,N_27737,N_27090);
or U28126 (N_28126,N_27224,N_27729);
nor U28127 (N_28127,N_27521,N_27971);
xor U28128 (N_28128,N_27192,N_27426);
xor U28129 (N_28129,N_27641,N_27633);
or U28130 (N_28130,N_27425,N_27127);
and U28131 (N_28131,N_27332,N_27935);
or U28132 (N_28132,N_27870,N_27025);
nor U28133 (N_28133,N_27844,N_27468);
or U28134 (N_28134,N_27655,N_27871);
nor U28135 (N_28135,N_27735,N_27733);
nand U28136 (N_28136,N_27769,N_27755);
and U28137 (N_28137,N_27632,N_27184);
or U28138 (N_28138,N_27202,N_27888);
nand U28139 (N_28139,N_27792,N_27175);
or U28140 (N_28140,N_27800,N_27065);
nor U28141 (N_28141,N_27363,N_27357);
and U28142 (N_28142,N_27549,N_27786);
and U28143 (N_28143,N_27400,N_27137);
nor U28144 (N_28144,N_27854,N_27126);
nor U28145 (N_28145,N_27106,N_27660);
or U28146 (N_28146,N_27910,N_27808);
and U28147 (N_28147,N_27877,N_27682);
xor U28148 (N_28148,N_27722,N_27112);
xnor U28149 (N_28149,N_27608,N_27201);
and U28150 (N_28150,N_27543,N_27922);
or U28151 (N_28151,N_27122,N_27411);
nor U28152 (N_28152,N_27036,N_27458);
and U28153 (N_28153,N_27406,N_27445);
and U28154 (N_28154,N_27809,N_27340);
or U28155 (N_28155,N_27205,N_27230);
xor U28156 (N_28156,N_27063,N_27822);
nor U28157 (N_28157,N_27969,N_27919);
and U28158 (N_28158,N_27505,N_27950);
xnor U28159 (N_28159,N_27449,N_27150);
xnor U28160 (N_28160,N_27114,N_27813);
and U28161 (N_28161,N_27562,N_27324);
xor U28162 (N_28162,N_27306,N_27605);
nor U28163 (N_28163,N_27868,N_27539);
and U28164 (N_28164,N_27087,N_27826);
or U28165 (N_28165,N_27475,N_27174);
nor U28166 (N_28166,N_27592,N_27416);
nor U28167 (N_28167,N_27828,N_27077);
nand U28168 (N_28168,N_27434,N_27414);
and U28169 (N_28169,N_27266,N_27883);
nor U28170 (N_28170,N_27221,N_27415);
xnor U28171 (N_28171,N_27802,N_27067);
or U28172 (N_28172,N_27545,N_27046);
or U28173 (N_28173,N_27019,N_27779);
or U28174 (N_28174,N_27444,N_27637);
xor U28175 (N_28175,N_27893,N_27700);
nor U28176 (N_28176,N_27740,N_27251);
nand U28177 (N_28177,N_27692,N_27120);
and U28178 (N_28178,N_27360,N_27865);
nand U28179 (N_28179,N_27909,N_27992);
or U28180 (N_28180,N_27344,N_27713);
nor U28181 (N_28181,N_27721,N_27474);
and U28182 (N_28182,N_27989,N_27912);
and U28183 (N_28183,N_27466,N_27965);
and U28184 (N_28184,N_27194,N_27520);
nor U28185 (N_28185,N_27798,N_27051);
or U28186 (N_28186,N_27789,N_27507);
and U28187 (N_28187,N_27572,N_27057);
nand U28188 (N_28188,N_27089,N_27649);
nand U28189 (N_28189,N_27567,N_27006);
and U28190 (N_28190,N_27853,N_27494);
nand U28191 (N_28191,N_27603,N_27167);
and U28192 (N_28192,N_27258,N_27124);
nand U28193 (N_28193,N_27304,N_27442);
nand U28194 (N_28194,N_27761,N_27862);
xor U28195 (N_28195,N_27461,N_27591);
and U28196 (N_28196,N_27599,N_27856);
or U28197 (N_28197,N_27791,N_27476);
nor U28198 (N_28198,N_27896,N_27579);
and U28199 (N_28199,N_27393,N_27540);
xnor U28200 (N_28200,N_27780,N_27574);
or U28201 (N_28201,N_27849,N_27522);
xnor U28202 (N_28202,N_27823,N_27487);
nand U28203 (N_28203,N_27404,N_27979);
and U28204 (N_28204,N_27914,N_27768);
nand U28205 (N_28205,N_27998,N_27182);
nor U28206 (N_28206,N_27447,N_27047);
or U28207 (N_28207,N_27547,N_27981);
and U28208 (N_28208,N_27671,N_27794);
or U28209 (N_28209,N_27313,N_27402);
and U28210 (N_28210,N_27237,N_27648);
nor U28211 (N_28211,N_27529,N_27994);
nor U28212 (N_28212,N_27872,N_27837);
xnor U28213 (N_28213,N_27255,N_27084);
or U28214 (N_28214,N_27320,N_27668);
xor U28215 (N_28215,N_27852,N_27538);
and U28216 (N_28216,N_27207,N_27576);
and U28217 (N_28217,N_27103,N_27443);
nand U28218 (N_28218,N_27166,N_27643);
xnor U28219 (N_28219,N_27168,N_27569);
nand U28220 (N_28220,N_27955,N_27042);
or U28221 (N_28221,N_27401,N_27219);
nand U28222 (N_28222,N_27428,N_27993);
xnor U28223 (N_28223,N_27663,N_27086);
xnor U28224 (N_28224,N_27478,N_27832);
nor U28225 (N_28225,N_27075,N_27398);
nor U28226 (N_28226,N_27140,N_27911);
or U28227 (N_28227,N_27467,N_27073);
and U28228 (N_28228,N_27710,N_27718);
or U28229 (N_28229,N_27850,N_27314);
nor U28230 (N_28230,N_27350,N_27032);
and U28231 (N_28231,N_27028,N_27519);
nand U28232 (N_28232,N_27376,N_27701);
or U28233 (N_28233,N_27473,N_27578);
nand U28234 (N_28234,N_27624,N_27502);
nand U28235 (N_28235,N_27824,N_27291);
and U28236 (N_28236,N_27098,N_27845);
nor U28237 (N_28237,N_27095,N_27925);
or U28238 (N_28238,N_27031,N_27515);
xor U28239 (N_28239,N_27790,N_27847);
or U28240 (N_28240,N_27327,N_27196);
and U28241 (N_28241,N_27216,N_27097);
nand U28242 (N_28242,N_27748,N_27581);
xnor U28243 (N_28243,N_27812,N_27841);
and U28244 (N_28244,N_27018,N_27767);
nor U28245 (N_28245,N_27630,N_27963);
or U28246 (N_28246,N_27898,N_27241);
nand U28247 (N_28247,N_27606,N_27088);
or U28248 (N_28248,N_27335,N_27346);
and U28249 (N_28249,N_27222,N_27664);
or U28250 (N_28250,N_27677,N_27661);
nand U28251 (N_28251,N_27913,N_27078);
and U28252 (N_28252,N_27223,N_27268);
xnor U28253 (N_28253,N_27076,N_27210);
xor U28254 (N_28254,N_27679,N_27842);
or U28255 (N_28255,N_27762,N_27693);
and U28256 (N_28256,N_27723,N_27585);
nand U28257 (N_28257,N_27039,N_27439);
nand U28258 (N_28258,N_27903,N_27699);
and U28259 (N_28259,N_27102,N_27714);
nor U28260 (N_28260,N_27662,N_27361);
xor U28261 (N_28261,N_27488,N_27695);
xor U28262 (N_28262,N_27375,N_27129);
or U28263 (N_28263,N_27399,N_27651);
nand U28264 (N_28264,N_27961,N_27189);
nor U28265 (N_28265,N_27370,N_27159);
or U28266 (N_28266,N_27155,N_27083);
or U28267 (N_28267,N_27185,N_27108);
and U28268 (N_28268,N_27396,N_27432);
nand U28269 (N_28269,N_27887,N_27448);
or U28270 (N_28270,N_27099,N_27176);
and U28271 (N_28271,N_27717,N_27111);
or U28272 (N_28272,N_27512,N_27364);
and U28273 (N_28273,N_27760,N_27489);
xor U28274 (N_28274,N_27362,N_27015);
or U28275 (N_28275,N_27094,N_27937);
xnor U28276 (N_28276,N_27956,N_27463);
nor U28277 (N_28277,N_27388,N_27318);
xor U28278 (N_28278,N_27920,N_27987);
and U28279 (N_28279,N_27348,N_27929);
xor U28280 (N_28280,N_27604,N_27541);
xnor U28281 (N_28281,N_27423,N_27139);
and U28282 (N_28282,N_27316,N_27575);
xnor U28283 (N_28283,N_27879,N_27819);
or U28284 (N_28284,N_27524,N_27601);
nand U28285 (N_28285,N_27926,N_27509);
nand U28286 (N_28286,N_27669,N_27247);
or U28287 (N_28287,N_27589,N_27349);
or U28288 (N_28288,N_27953,N_27500);
nor U28289 (N_28289,N_27686,N_27665);
nor U28290 (N_28290,N_27960,N_27236);
xor U28291 (N_28291,N_27355,N_27427);
nor U28292 (N_28292,N_27918,N_27289);
nor U28293 (N_28293,N_27315,N_27121);
nand U28294 (N_28294,N_27068,N_27429);
or U28295 (N_28295,N_27240,N_27899);
nor U28296 (N_28296,N_27001,N_27290);
nand U28297 (N_28297,N_27390,N_27299);
nand U28298 (N_28298,N_27141,N_27629);
and U28299 (N_28299,N_27817,N_27727);
nor U28300 (N_28300,N_27570,N_27260);
nand U28301 (N_28301,N_27085,N_27499);
nor U28302 (N_28302,N_27273,N_27281);
and U28303 (N_28303,N_27038,N_27732);
nand U28304 (N_28304,N_27490,N_27905);
nor U28305 (N_28305,N_27517,N_27212);
nand U28306 (N_28306,N_27597,N_27985);
and U28307 (N_28307,N_27394,N_27117);
xnor U28308 (N_28308,N_27169,N_27003);
xor U28309 (N_28309,N_27930,N_27777);
and U28310 (N_28310,N_27239,N_27481);
nand U28311 (N_28311,N_27623,N_27092);
and U28312 (N_28312,N_27766,N_27758);
nand U28313 (N_28313,N_27590,N_27511);
nor U28314 (N_28314,N_27148,N_27943);
nand U28315 (N_28315,N_27787,N_27977);
or U28316 (N_28316,N_27165,N_27757);
or U28317 (N_28317,N_27635,N_27982);
nor U28318 (N_28318,N_27895,N_27072);
nor U28319 (N_28319,N_27796,N_27616);
or U28320 (N_28320,N_27594,N_27535);
nor U28321 (N_28321,N_27485,N_27403);
nand U28322 (N_28322,N_27678,N_27462);
or U28323 (N_28323,N_27525,N_27561);
or U28324 (N_28324,N_27280,N_27835);
or U28325 (N_28325,N_27745,N_27707);
and U28326 (N_28326,N_27373,N_27640);
nand U28327 (N_28327,N_27527,N_27706);
or U28328 (N_28328,N_27422,N_27942);
xor U28329 (N_28329,N_27209,N_27583);
nor U28330 (N_28330,N_27034,N_27785);
nor U28331 (N_28331,N_27902,N_27389);
and U28332 (N_28332,N_27465,N_27248);
and U28333 (N_28333,N_27749,N_27407);
nand U28334 (N_28334,N_27772,N_27421);
nand U28335 (N_28335,N_27948,N_27142);
xnor U28336 (N_28336,N_27386,N_27101);
and U28337 (N_28337,N_27741,N_27211);
and U28338 (N_28338,N_27060,N_27321);
or U28339 (N_28339,N_27208,N_27229);
xor U28340 (N_28340,N_27070,N_27968);
nand U28341 (N_28341,N_27145,N_27550);
or U28342 (N_28342,N_27917,N_27254);
xor U28343 (N_28343,N_27932,N_27553);
xnor U28344 (N_28344,N_27687,N_27644);
nor U28345 (N_28345,N_27341,N_27784);
and U28346 (N_28346,N_27957,N_27181);
xnor U28347 (N_28347,N_27685,N_27493);
and U28348 (N_28348,N_27839,N_27128);
and U28349 (N_28349,N_27383,N_27980);
nand U28350 (N_28350,N_27483,N_27161);
nor U28351 (N_28351,N_27040,N_27413);
xnor U28352 (N_28352,N_27568,N_27256);
xor U28353 (N_28353,N_27778,N_27319);
xor U28354 (N_28354,N_27116,N_27788);
or U28355 (N_28355,N_27618,N_27217);
nand U28356 (N_28356,N_27163,N_27675);
nor U28357 (N_28357,N_27566,N_27203);
or U28358 (N_28358,N_27621,N_27359);
nand U28359 (N_28359,N_27508,N_27131);
nor U28360 (N_28360,N_27295,N_27420);
and U28361 (N_28361,N_27542,N_27469);
nand U28362 (N_28362,N_27283,N_27410);
or U28363 (N_28363,N_27171,N_27514);
nand U28364 (N_28364,N_27878,N_27901);
xnor U28365 (N_28365,N_27619,N_27064);
and U28366 (N_28366,N_27367,N_27764);
and U28367 (N_28367,N_27267,N_27654);
and U28368 (N_28368,N_27698,N_27495);
or U28369 (N_28369,N_27056,N_27730);
or U28370 (N_28370,N_27928,N_27033);
and U28371 (N_28371,N_27804,N_27636);
nand U28372 (N_28372,N_27861,N_27453);
xnor U28373 (N_28373,N_27353,N_27571);
or U28374 (N_28374,N_27133,N_27810);
xor U28375 (N_28375,N_27672,N_27751);
and U28376 (N_28376,N_27232,N_27716);
and U28377 (N_28377,N_27107,N_27055);
and U28378 (N_28378,N_27944,N_27904);
nor U28379 (N_28379,N_27164,N_27653);
nor U28380 (N_28380,N_27814,N_27342);
nand U28381 (N_28381,N_27811,N_27773);
xnor U28382 (N_28382,N_27536,N_27750);
nand U28383 (N_28383,N_27816,N_27876);
nand U28384 (N_28384,N_27936,N_27602);
or U28385 (N_28385,N_27949,N_27719);
xnor U28386 (N_28386,N_27451,N_27105);
and U28387 (N_28387,N_27532,N_27864);
and U28388 (N_28388,N_27546,N_27694);
xor U28389 (N_28389,N_27715,N_27190);
or U28390 (N_28390,N_27486,N_27848);
and U28391 (N_28391,N_27609,N_27151);
nand U28392 (N_28392,N_27610,N_27931);
xnor U28393 (N_28393,N_27563,N_27496);
nand U28394 (N_28394,N_27250,N_27673);
nor U28395 (N_28395,N_27830,N_27347);
nand U28396 (N_28396,N_27249,N_27005);
or U28397 (N_28397,N_27829,N_27962);
xor U28398 (N_28398,N_27946,N_27860);
nand U28399 (N_28399,N_27278,N_27681);
and U28400 (N_28400,N_27620,N_27480);
nor U28401 (N_28401,N_27518,N_27947);
and U28402 (N_28402,N_27160,N_27387);
nor U28403 (N_28403,N_27596,N_27975);
nand U28404 (N_28404,N_27923,N_27118);
xor U28405 (N_28405,N_27455,N_27976);
nand U28406 (N_28406,N_27328,N_27843);
xnor U28407 (N_28407,N_27246,N_27863);
xnor U28408 (N_28408,N_27552,N_27881);
nor U28409 (N_28409,N_27825,N_27157);
and U28410 (N_28410,N_27938,N_27763);
and U28411 (N_28411,N_27308,N_27143);
nor U28412 (N_28412,N_27625,N_27978);
xnor U28413 (N_28413,N_27187,N_27284);
nand U28414 (N_28414,N_27326,N_27199);
nor U28415 (N_28415,N_27859,N_27457);
nand U28416 (N_28416,N_27873,N_27356);
or U28417 (N_28417,N_27252,N_27670);
or U28418 (N_28418,N_27754,N_27691);
or U28419 (N_28419,N_27801,N_27638);
xnor U28420 (N_28420,N_27195,N_27724);
xnor U28421 (N_28421,N_27634,N_27017);
nor U28422 (N_28422,N_27642,N_27846);
or U28423 (N_28423,N_27513,N_27030);
and U28424 (N_28424,N_27274,N_27827);
nor U28425 (N_28425,N_27770,N_27795);
xor U28426 (N_28426,N_27021,N_27138);
and U28427 (N_28427,N_27336,N_27704);
or U28428 (N_28428,N_27433,N_27739);
xnor U28429 (N_28429,N_27177,N_27744);
or U28430 (N_28430,N_27774,N_27144);
and U28431 (N_28431,N_27213,N_27697);
xnor U28432 (N_28432,N_27069,N_27954);
nor U28433 (N_28433,N_27680,N_27408);
and U28434 (N_28434,N_27123,N_27297);
or U28435 (N_28435,N_27002,N_27082);
xnor U28436 (N_28436,N_27974,N_27307);
nand U28437 (N_28437,N_27799,N_27397);
and U28438 (N_28438,N_27004,N_27276);
and U28439 (N_28439,N_27264,N_27045);
xor U28440 (N_28440,N_27269,N_27776);
or U28441 (N_28441,N_27302,N_27435);
xnor U28442 (N_28442,N_27891,N_27054);
and U28443 (N_28443,N_27838,N_27296);
or U28444 (N_28444,N_27688,N_27134);
nor U28445 (N_28445,N_27206,N_27242);
or U28446 (N_28446,N_27806,N_27100);
and U28447 (N_28447,N_27074,N_27294);
nor U28448 (N_28448,N_27857,N_27934);
or U28449 (N_28449,N_27884,N_27119);
and U28450 (N_28450,N_27738,N_27479);
and U28451 (N_28451,N_27491,N_27726);
nor U28452 (N_28452,N_27815,N_27897);
and U28453 (N_28453,N_27711,N_27889);
nand U28454 (N_28454,N_27186,N_27537);
nor U28455 (N_28455,N_27970,N_27198);
and U28456 (N_28456,N_27684,N_27504);
nor U28457 (N_28457,N_27286,N_27301);
nand U28458 (N_28458,N_27674,N_27270);
or U28459 (N_28459,N_27368,N_27385);
or U28460 (N_28460,N_27894,N_27243);
nand U28461 (N_28461,N_27501,N_27708);
nand U28462 (N_28462,N_27890,N_27921);
and U28463 (N_28463,N_27600,N_27197);
nor U28464 (N_28464,N_27043,N_27022);
and U28465 (N_28465,N_27614,N_27598);
or U28466 (N_28466,N_27556,N_27990);
xnor U28467 (N_28467,N_27343,N_27696);
nand U28468 (N_28468,N_27858,N_27559);
or U28469 (N_28469,N_27245,N_27178);
nand U28470 (N_28470,N_27820,N_27158);
or U28471 (N_28471,N_27470,N_27200);
or U28472 (N_28472,N_27966,N_27803);
xor U28473 (N_28473,N_27369,N_27233);
or U28474 (N_28474,N_27492,N_27058);
or U28475 (N_28475,N_27986,N_27330);
and U28476 (N_28476,N_27279,N_27557);
nor U28477 (N_28477,N_27009,N_27834);
nor U28478 (N_28478,N_27334,N_27412);
or U28479 (N_28479,N_27805,N_27558);
or U28480 (N_28480,N_27959,N_27908);
and U28481 (N_28481,N_27528,N_27132);
or U28482 (N_28482,N_27377,N_27712);
or U28483 (N_28483,N_27927,N_27231);
xnor U28484 (N_28484,N_27024,N_27498);
or U28485 (N_28485,N_27012,N_27720);
nand U28486 (N_28486,N_27656,N_27193);
nand U28487 (N_28487,N_27497,N_27020);
xor U28488 (N_28488,N_27991,N_27305);
nor U28489 (N_28489,N_27689,N_27188);
xnor U28490 (N_28490,N_27916,N_27380);
xnor U28491 (N_28491,N_27703,N_27840);
nor U28492 (N_28492,N_27807,N_27384);
nand U28493 (N_28493,N_27430,N_27309);
nand U28494 (N_28494,N_27564,N_27940);
nor U28495 (N_28495,N_27941,N_27029);
xor U28496 (N_28496,N_27226,N_27244);
nand U28497 (N_28497,N_27781,N_27010);
nand U28498 (N_28498,N_27011,N_27418);
nand U28499 (N_28499,N_27459,N_27113);
or U28500 (N_28500,N_27426,N_27336);
and U28501 (N_28501,N_27645,N_27630);
nand U28502 (N_28502,N_27729,N_27460);
nor U28503 (N_28503,N_27947,N_27261);
and U28504 (N_28504,N_27161,N_27592);
nor U28505 (N_28505,N_27533,N_27806);
nand U28506 (N_28506,N_27610,N_27384);
nand U28507 (N_28507,N_27678,N_27115);
nand U28508 (N_28508,N_27039,N_27978);
and U28509 (N_28509,N_27216,N_27674);
and U28510 (N_28510,N_27298,N_27664);
or U28511 (N_28511,N_27814,N_27942);
nand U28512 (N_28512,N_27706,N_27180);
nand U28513 (N_28513,N_27704,N_27272);
or U28514 (N_28514,N_27179,N_27350);
and U28515 (N_28515,N_27674,N_27231);
nor U28516 (N_28516,N_27880,N_27332);
and U28517 (N_28517,N_27212,N_27795);
nor U28518 (N_28518,N_27358,N_27011);
and U28519 (N_28519,N_27760,N_27811);
nor U28520 (N_28520,N_27875,N_27119);
and U28521 (N_28521,N_27878,N_27407);
nor U28522 (N_28522,N_27610,N_27018);
nand U28523 (N_28523,N_27848,N_27905);
xnor U28524 (N_28524,N_27542,N_27585);
or U28525 (N_28525,N_27205,N_27429);
nor U28526 (N_28526,N_27874,N_27956);
nand U28527 (N_28527,N_27449,N_27452);
nand U28528 (N_28528,N_27420,N_27185);
nand U28529 (N_28529,N_27712,N_27708);
or U28530 (N_28530,N_27262,N_27867);
or U28531 (N_28531,N_27750,N_27051);
and U28532 (N_28532,N_27718,N_27620);
nand U28533 (N_28533,N_27518,N_27055);
and U28534 (N_28534,N_27919,N_27846);
or U28535 (N_28535,N_27548,N_27546);
nand U28536 (N_28536,N_27207,N_27862);
and U28537 (N_28537,N_27725,N_27424);
and U28538 (N_28538,N_27941,N_27490);
xnor U28539 (N_28539,N_27476,N_27864);
xnor U28540 (N_28540,N_27660,N_27129);
or U28541 (N_28541,N_27332,N_27261);
nor U28542 (N_28542,N_27868,N_27042);
and U28543 (N_28543,N_27676,N_27647);
nor U28544 (N_28544,N_27937,N_27293);
xor U28545 (N_28545,N_27931,N_27140);
xor U28546 (N_28546,N_27525,N_27007);
or U28547 (N_28547,N_27065,N_27949);
xnor U28548 (N_28548,N_27768,N_27443);
and U28549 (N_28549,N_27021,N_27347);
or U28550 (N_28550,N_27954,N_27284);
nor U28551 (N_28551,N_27284,N_27390);
nand U28552 (N_28552,N_27176,N_27355);
or U28553 (N_28553,N_27597,N_27460);
or U28554 (N_28554,N_27880,N_27624);
and U28555 (N_28555,N_27073,N_27486);
nand U28556 (N_28556,N_27442,N_27608);
or U28557 (N_28557,N_27379,N_27684);
nand U28558 (N_28558,N_27642,N_27727);
xor U28559 (N_28559,N_27613,N_27138);
nand U28560 (N_28560,N_27530,N_27319);
or U28561 (N_28561,N_27272,N_27859);
or U28562 (N_28562,N_27950,N_27348);
nand U28563 (N_28563,N_27337,N_27297);
nor U28564 (N_28564,N_27564,N_27878);
and U28565 (N_28565,N_27591,N_27381);
and U28566 (N_28566,N_27676,N_27490);
nor U28567 (N_28567,N_27370,N_27067);
or U28568 (N_28568,N_27372,N_27616);
nor U28569 (N_28569,N_27699,N_27484);
and U28570 (N_28570,N_27377,N_27571);
xnor U28571 (N_28571,N_27804,N_27718);
xnor U28572 (N_28572,N_27408,N_27146);
xor U28573 (N_28573,N_27793,N_27417);
xor U28574 (N_28574,N_27250,N_27210);
and U28575 (N_28575,N_27867,N_27807);
nand U28576 (N_28576,N_27862,N_27374);
and U28577 (N_28577,N_27964,N_27507);
and U28578 (N_28578,N_27904,N_27890);
and U28579 (N_28579,N_27882,N_27842);
nor U28580 (N_28580,N_27195,N_27973);
and U28581 (N_28581,N_27979,N_27727);
nor U28582 (N_28582,N_27359,N_27423);
nand U28583 (N_28583,N_27878,N_27589);
or U28584 (N_28584,N_27208,N_27147);
nand U28585 (N_28585,N_27312,N_27401);
and U28586 (N_28586,N_27326,N_27567);
nor U28587 (N_28587,N_27630,N_27962);
and U28588 (N_28588,N_27464,N_27893);
and U28589 (N_28589,N_27316,N_27636);
nand U28590 (N_28590,N_27299,N_27147);
nand U28591 (N_28591,N_27258,N_27520);
and U28592 (N_28592,N_27852,N_27527);
or U28593 (N_28593,N_27415,N_27033);
nand U28594 (N_28594,N_27023,N_27514);
xor U28595 (N_28595,N_27993,N_27965);
nand U28596 (N_28596,N_27654,N_27824);
xor U28597 (N_28597,N_27592,N_27375);
or U28598 (N_28598,N_27724,N_27106);
xor U28599 (N_28599,N_27100,N_27275);
xor U28600 (N_28600,N_27485,N_27261);
or U28601 (N_28601,N_27817,N_27982);
xnor U28602 (N_28602,N_27031,N_27209);
nor U28603 (N_28603,N_27765,N_27598);
or U28604 (N_28604,N_27508,N_27534);
nor U28605 (N_28605,N_27842,N_27265);
nand U28606 (N_28606,N_27229,N_27935);
xnor U28607 (N_28607,N_27474,N_27953);
nor U28608 (N_28608,N_27472,N_27807);
or U28609 (N_28609,N_27828,N_27649);
or U28610 (N_28610,N_27122,N_27530);
nor U28611 (N_28611,N_27170,N_27785);
nand U28612 (N_28612,N_27651,N_27944);
nand U28613 (N_28613,N_27180,N_27682);
xor U28614 (N_28614,N_27650,N_27286);
nand U28615 (N_28615,N_27380,N_27757);
nand U28616 (N_28616,N_27364,N_27580);
nor U28617 (N_28617,N_27486,N_27725);
xor U28618 (N_28618,N_27806,N_27197);
and U28619 (N_28619,N_27692,N_27277);
nand U28620 (N_28620,N_27882,N_27988);
or U28621 (N_28621,N_27143,N_27262);
or U28622 (N_28622,N_27976,N_27468);
and U28623 (N_28623,N_27644,N_27237);
nand U28624 (N_28624,N_27463,N_27373);
nor U28625 (N_28625,N_27470,N_27097);
xnor U28626 (N_28626,N_27415,N_27381);
and U28627 (N_28627,N_27375,N_27569);
xnor U28628 (N_28628,N_27834,N_27884);
and U28629 (N_28629,N_27787,N_27337);
and U28630 (N_28630,N_27616,N_27946);
or U28631 (N_28631,N_27833,N_27240);
nand U28632 (N_28632,N_27345,N_27900);
and U28633 (N_28633,N_27341,N_27750);
and U28634 (N_28634,N_27793,N_27512);
or U28635 (N_28635,N_27979,N_27250);
xnor U28636 (N_28636,N_27298,N_27064);
and U28637 (N_28637,N_27955,N_27046);
or U28638 (N_28638,N_27219,N_27602);
and U28639 (N_28639,N_27133,N_27299);
and U28640 (N_28640,N_27100,N_27308);
xor U28641 (N_28641,N_27740,N_27235);
nor U28642 (N_28642,N_27347,N_27273);
nand U28643 (N_28643,N_27714,N_27258);
or U28644 (N_28644,N_27845,N_27710);
and U28645 (N_28645,N_27049,N_27013);
nand U28646 (N_28646,N_27537,N_27076);
nor U28647 (N_28647,N_27022,N_27216);
nor U28648 (N_28648,N_27160,N_27357);
or U28649 (N_28649,N_27346,N_27244);
or U28650 (N_28650,N_27322,N_27796);
or U28651 (N_28651,N_27627,N_27072);
nand U28652 (N_28652,N_27000,N_27231);
nor U28653 (N_28653,N_27352,N_27716);
xor U28654 (N_28654,N_27798,N_27514);
or U28655 (N_28655,N_27288,N_27981);
nor U28656 (N_28656,N_27809,N_27069);
nor U28657 (N_28657,N_27058,N_27175);
xnor U28658 (N_28658,N_27214,N_27935);
and U28659 (N_28659,N_27608,N_27675);
or U28660 (N_28660,N_27651,N_27200);
nand U28661 (N_28661,N_27066,N_27720);
xnor U28662 (N_28662,N_27938,N_27538);
and U28663 (N_28663,N_27195,N_27786);
and U28664 (N_28664,N_27871,N_27130);
xor U28665 (N_28665,N_27049,N_27194);
nor U28666 (N_28666,N_27308,N_27665);
and U28667 (N_28667,N_27200,N_27003);
and U28668 (N_28668,N_27895,N_27737);
and U28669 (N_28669,N_27416,N_27482);
xor U28670 (N_28670,N_27312,N_27209);
or U28671 (N_28671,N_27638,N_27477);
or U28672 (N_28672,N_27793,N_27525);
nor U28673 (N_28673,N_27496,N_27982);
xnor U28674 (N_28674,N_27683,N_27825);
nand U28675 (N_28675,N_27818,N_27572);
or U28676 (N_28676,N_27173,N_27384);
or U28677 (N_28677,N_27461,N_27041);
nor U28678 (N_28678,N_27553,N_27667);
nor U28679 (N_28679,N_27854,N_27186);
and U28680 (N_28680,N_27670,N_27595);
nand U28681 (N_28681,N_27025,N_27516);
or U28682 (N_28682,N_27090,N_27704);
nand U28683 (N_28683,N_27848,N_27488);
nand U28684 (N_28684,N_27426,N_27509);
and U28685 (N_28685,N_27385,N_27006);
and U28686 (N_28686,N_27630,N_27783);
and U28687 (N_28687,N_27830,N_27249);
nand U28688 (N_28688,N_27258,N_27540);
and U28689 (N_28689,N_27448,N_27362);
nand U28690 (N_28690,N_27143,N_27459);
xor U28691 (N_28691,N_27908,N_27726);
nand U28692 (N_28692,N_27090,N_27686);
or U28693 (N_28693,N_27508,N_27794);
xor U28694 (N_28694,N_27935,N_27050);
and U28695 (N_28695,N_27760,N_27561);
nand U28696 (N_28696,N_27583,N_27012);
or U28697 (N_28697,N_27115,N_27556);
or U28698 (N_28698,N_27291,N_27372);
or U28699 (N_28699,N_27330,N_27023);
nand U28700 (N_28700,N_27609,N_27398);
nor U28701 (N_28701,N_27015,N_27174);
and U28702 (N_28702,N_27612,N_27496);
xor U28703 (N_28703,N_27136,N_27953);
nor U28704 (N_28704,N_27440,N_27357);
nand U28705 (N_28705,N_27428,N_27124);
nor U28706 (N_28706,N_27404,N_27189);
nand U28707 (N_28707,N_27623,N_27223);
xnor U28708 (N_28708,N_27406,N_27901);
nor U28709 (N_28709,N_27854,N_27902);
nand U28710 (N_28710,N_27822,N_27542);
and U28711 (N_28711,N_27117,N_27491);
nand U28712 (N_28712,N_27759,N_27699);
and U28713 (N_28713,N_27851,N_27056);
nor U28714 (N_28714,N_27130,N_27847);
xor U28715 (N_28715,N_27159,N_27309);
or U28716 (N_28716,N_27504,N_27393);
nor U28717 (N_28717,N_27222,N_27093);
and U28718 (N_28718,N_27864,N_27565);
nor U28719 (N_28719,N_27251,N_27984);
xor U28720 (N_28720,N_27310,N_27124);
nor U28721 (N_28721,N_27541,N_27580);
or U28722 (N_28722,N_27967,N_27208);
and U28723 (N_28723,N_27697,N_27202);
and U28724 (N_28724,N_27090,N_27177);
or U28725 (N_28725,N_27688,N_27090);
xor U28726 (N_28726,N_27217,N_27728);
and U28727 (N_28727,N_27947,N_27262);
nor U28728 (N_28728,N_27138,N_27795);
nor U28729 (N_28729,N_27801,N_27118);
nor U28730 (N_28730,N_27859,N_27414);
xor U28731 (N_28731,N_27660,N_27789);
or U28732 (N_28732,N_27553,N_27257);
or U28733 (N_28733,N_27359,N_27666);
or U28734 (N_28734,N_27562,N_27643);
xor U28735 (N_28735,N_27790,N_27300);
xor U28736 (N_28736,N_27639,N_27188);
nand U28737 (N_28737,N_27638,N_27233);
and U28738 (N_28738,N_27819,N_27133);
nand U28739 (N_28739,N_27157,N_27259);
nand U28740 (N_28740,N_27722,N_27622);
and U28741 (N_28741,N_27986,N_27525);
nand U28742 (N_28742,N_27400,N_27376);
and U28743 (N_28743,N_27057,N_27427);
nor U28744 (N_28744,N_27859,N_27989);
nor U28745 (N_28745,N_27408,N_27573);
xnor U28746 (N_28746,N_27855,N_27625);
or U28747 (N_28747,N_27670,N_27063);
or U28748 (N_28748,N_27673,N_27899);
nor U28749 (N_28749,N_27140,N_27582);
or U28750 (N_28750,N_27591,N_27367);
nor U28751 (N_28751,N_27277,N_27683);
and U28752 (N_28752,N_27139,N_27678);
and U28753 (N_28753,N_27192,N_27341);
or U28754 (N_28754,N_27773,N_27411);
and U28755 (N_28755,N_27493,N_27712);
nand U28756 (N_28756,N_27818,N_27653);
xnor U28757 (N_28757,N_27626,N_27556);
and U28758 (N_28758,N_27743,N_27436);
nand U28759 (N_28759,N_27758,N_27781);
nor U28760 (N_28760,N_27303,N_27612);
nor U28761 (N_28761,N_27760,N_27703);
nand U28762 (N_28762,N_27652,N_27720);
xor U28763 (N_28763,N_27380,N_27872);
or U28764 (N_28764,N_27671,N_27330);
and U28765 (N_28765,N_27621,N_27456);
and U28766 (N_28766,N_27615,N_27029);
xnor U28767 (N_28767,N_27792,N_27257);
and U28768 (N_28768,N_27916,N_27902);
nand U28769 (N_28769,N_27022,N_27795);
xor U28770 (N_28770,N_27003,N_27304);
or U28771 (N_28771,N_27213,N_27434);
xor U28772 (N_28772,N_27783,N_27938);
nor U28773 (N_28773,N_27331,N_27141);
nor U28774 (N_28774,N_27190,N_27918);
nand U28775 (N_28775,N_27445,N_27751);
and U28776 (N_28776,N_27939,N_27854);
nand U28777 (N_28777,N_27657,N_27215);
xnor U28778 (N_28778,N_27615,N_27204);
xor U28779 (N_28779,N_27442,N_27871);
xnor U28780 (N_28780,N_27696,N_27180);
nand U28781 (N_28781,N_27100,N_27905);
nor U28782 (N_28782,N_27161,N_27244);
xor U28783 (N_28783,N_27470,N_27652);
and U28784 (N_28784,N_27544,N_27017);
nand U28785 (N_28785,N_27200,N_27380);
nand U28786 (N_28786,N_27426,N_27626);
or U28787 (N_28787,N_27078,N_27186);
or U28788 (N_28788,N_27996,N_27250);
xnor U28789 (N_28789,N_27205,N_27723);
nand U28790 (N_28790,N_27837,N_27951);
and U28791 (N_28791,N_27813,N_27632);
xnor U28792 (N_28792,N_27619,N_27583);
nor U28793 (N_28793,N_27291,N_27858);
and U28794 (N_28794,N_27248,N_27437);
and U28795 (N_28795,N_27866,N_27120);
and U28796 (N_28796,N_27943,N_27302);
and U28797 (N_28797,N_27214,N_27800);
or U28798 (N_28798,N_27017,N_27429);
xor U28799 (N_28799,N_27169,N_27860);
xor U28800 (N_28800,N_27737,N_27502);
and U28801 (N_28801,N_27565,N_27706);
nand U28802 (N_28802,N_27271,N_27351);
or U28803 (N_28803,N_27401,N_27971);
and U28804 (N_28804,N_27133,N_27491);
or U28805 (N_28805,N_27892,N_27557);
xnor U28806 (N_28806,N_27343,N_27941);
nor U28807 (N_28807,N_27226,N_27850);
nand U28808 (N_28808,N_27417,N_27654);
or U28809 (N_28809,N_27892,N_27110);
and U28810 (N_28810,N_27647,N_27681);
xnor U28811 (N_28811,N_27735,N_27962);
nor U28812 (N_28812,N_27607,N_27847);
xnor U28813 (N_28813,N_27536,N_27225);
and U28814 (N_28814,N_27490,N_27039);
xor U28815 (N_28815,N_27635,N_27176);
nand U28816 (N_28816,N_27336,N_27709);
xor U28817 (N_28817,N_27456,N_27440);
or U28818 (N_28818,N_27561,N_27558);
or U28819 (N_28819,N_27429,N_27211);
nand U28820 (N_28820,N_27031,N_27131);
xor U28821 (N_28821,N_27715,N_27368);
nor U28822 (N_28822,N_27410,N_27419);
and U28823 (N_28823,N_27159,N_27009);
and U28824 (N_28824,N_27003,N_27027);
or U28825 (N_28825,N_27723,N_27807);
nand U28826 (N_28826,N_27187,N_27248);
nor U28827 (N_28827,N_27006,N_27889);
or U28828 (N_28828,N_27990,N_27769);
or U28829 (N_28829,N_27827,N_27936);
xor U28830 (N_28830,N_27308,N_27114);
nand U28831 (N_28831,N_27214,N_27023);
nor U28832 (N_28832,N_27673,N_27236);
xor U28833 (N_28833,N_27374,N_27028);
nor U28834 (N_28834,N_27245,N_27964);
or U28835 (N_28835,N_27610,N_27114);
or U28836 (N_28836,N_27124,N_27302);
xnor U28837 (N_28837,N_27599,N_27003);
or U28838 (N_28838,N_27020,N_27191);
nor U28839 (N_28839,N_27865,N_27818);
xor U28840 (N_28840,N_27437,N_27338);
and U28841 (N_28841,N_27213,N_27820);
or U28842 (N_28842,N_27820,N_27390);
nor U28843 (N_28843,N_27005,N_27806);
nand U28844 (N_28844,N_27964,N_27853);
nand U28845 (N_28845,N_27948,N_27512);
or U28846 (N_28846,N_27917,N_27668);
or U28847 (N_28847,N_27954,N_27465);
nor U28848 (N_28848,N_27521,N_27004);
xnor U28849 (N_28849,N_27803,N_27410);
xnor U28850 (N_28850,N_27367,N_27518);
nand U28851 (N_28851,N_27067,N_27642);
xor U28852 (N_28852,N_27700,N_27008);
nor U28853 (N_28853,N_27690,N_27949);
nand U28854 (N_28854,N_27228,N_27001);
and U28855 (N_28855,N_27378,N_27593);
nor U28856 (N_28856,N_27054,N_27602);
nand U28857 (N_28857,N_27464,N_27533);
or U28858 (N_28858,N_27726,N_27240);
and U28859 (N_28859,N_27321,N_27464);
and U28860 (N_28860,N_27783,N_27765);
or U28861 (N_28861,N_27660,N_27156);
and U28862 (N_28862,N_27541,N_27953);
nand U28863 (N_28863,N_27729,N_27893);
xor U28864 (N_28864,N_27101,N_27135);
and U28865 (N_28865,N_27556,N_27155);
xor U28866 (N_28866,N_27463,N_27798);
and U28867 (N_28867,N_27899,N_27282);
nand U28868 (N_28868,N_27199,N_27325);
xnor U28869 (N_28869,N_27656,N_27893);
nand U28870 (N_28870,N_27811,N_27222);
nor U28871 (N_28871,N_27506,N_27215);
and U28872 (N_28872,N_27547,N_27460);
nand U28873 (N_28873,N_27915,N_27289);
nor U28874 (N_28874,N_27126,N_27515);
nor U28875 (N_28875,N_27759,N_27072);
nor U28876 (N_28876,N_27776,N_27307);
or U28877 (N_28877,N_27813,N_27248);
nand U28878 (N_28878,N_27154,N_27979);
nand U28879 (N_28879,N_27245,N_27126);
or U28880 (N_28880,N_27269,N_27419);
or U28881 (N_28881,N_27016,N_27004);
or U28882 (N_28882,N_27015,N_27250);
or U28883 (N_28883,N_27386,N_27732);
and U28884 (N_28884,N_27863,N_27113);
or U28885 (N_28885,N_27291,N_27946);
nor U28886 (N_28886,N_27693,N_27818);
nand U28887 (N_28887,N_27989,N_27651);
nand U28888 (N_28888,N_27409,N_27894);
nor U28889 (N_28889,N_27674,N_27241);
and U28890 (N_28890,N_27347,N_27652);
nand U28891 (N_28891,N_27071,N_27118);
nor U28892 (N_28892,N_27479,N_27618);
or U28893 (N_28893,N_27158,N_27540);
xor U28894 (N_28894,N_27285,N_27332);
and U28895 (N_28895,N_27647,N_27082);
and U28896 (N_28896,N_27422,N_27792);
and U28897 (N_28897,N_27580,N_27384);
or U28898 (N_28898,N_27840,N_27807);
nand U28899 (N_28899,N_27070,N_27484);
or U28900 (N_28900,N_27822,N_27547);
nand U28901 (N_28901,N_27762,N_27737);
and U28902 (N_28902,N_27200,N_27166);
xor U28903 (N_28903,N_27503,N_27016);
and U28904 (N_28904,N_27184,N_27936);
xor U28905 (N_28905,N_27995,N_27808);
or U28906 (N_28906,N_27704,N_27990);
or U28907 (N_28907,N_27557,N_27227);
and U28908 (N_28908,N_27932,N_27595);
nor U28909 (N_28909,N_27398,N_27399);
or U28910 (N_28910,N_27163,N_27894);
nand U28911 (N_28911,N_27035,N_27658);
xnor U28912 (N_28912,N_27041,N_27443);
xor U28913 (N_28913,N_27802,N_27287);
xnor U28914 (N_28914,N_27866,N_27300);
xor U28915 (N_28915,N_27837,N_27407);
and U28916 (N_28916,N_27553,N_27535);
nand U28917 (N_28917,N_27915,N_27004);
nor U28918 (N_28918,N_27426,N_27969);
and U28919 (N_28919,N_27260,N_27022);
or U28920 (N_28920,N_27530,N_27131);
or U28921 (N_28921,N_27100,N_27958);
or U28922 (N_28922,N_27400,N_27345);
nor U28923 (N_28923,N_27763,N_27922);
xnor U28924 (N_28924,N_27886,N_27460);
nand U28925 (N_28925,N_27480,N_27856);
or U28926 (N_28926,N_27177,N_27345);
nor U28927 (N_28927,N_27767,N_27673);
and U28928 (N_28928,N_27114,N_27608);
nor U28929 (N_28929,N_27974,N_27888);
nor U28930 (N_28930,N_27463,N_27628);
nor U28931 (N_28931,N_27028,N_27551);
nor U28932 (N_28932,N_27449,N_27489);
or U28933 (N_28933,N_27155,N_27600);
and U28934 (N_28934,N_27576,N_27546);
nor U28935 (N_28935,N_27018,N_27890);
or U28936 (N_28936,N_27245,N_27488);
or U28937 (N_28937,N_27495,N_27433);
and U28938 (N_28938,N_27301,N_27094);
or U28939 (N_28939,N_27489,N_27158);
or U28940 (N_28940,N_27784,N_27727);
nor U28941 (N_28941,N_27906,N_27745);
xor U28942 (N_28942,N_27591,N_27608);
nand U28943 (N_28943,N_27879,N_27494);
nor U28944 (N_28944,N_27265,N_27920);
and U28945 (N_28945,N_27300,N_27052);
and U28946 (N_28946,N_27789,N_27122);
nor U28947 (N_28947,N_27282,N_27677);
nand U28948 (N_28948,N_27709,N_27164);
nor U28949 (N_28949,N_27288,N_27792);
nand U28950 (N_28950,N_27545,N_27633);
nand U28951 (N_28951,N_27306,N_27931);
nand U28952 (N_28952,N_27721,N_27307);
nand U28953 (N_28953,N_27130,N_27990);
and U28954 (N_28954,N_27229,N_27984);
and U28955 (N_28955,N_27401,N_27380);
xor U28956 (N_28956,N_27083,N_27184);
nand U28957 (N_28957,N_27272,N_27479);
nand U28958 (N_28958,N_27973,N_27987);
xor U28959 (N_28959,N_27536,N_27569);
xnor U28960 (N_28960,N_27229,N_27853);
or U28961 (N_28961,N_27611,N_27919);
xnor U28962 (N_28962,N_27359,N_27699);
nor U28963 (N_28963,N_27692,N_27746);
nor U28964 (N_28964,N_27237,N_27453);
nand U28965 (N_28965,N_27978,N_27499);
or U28966 (N_28966,N_27262,N_27896);
nand U28967 (N_28967,N_27979,N_27908);
xor U28968 (N_28968,N_27287,N_27613);
and U28969 (N_28969,N_27654,N_27784);
nand U28970 (N_28970,N_27511,N_27740);
xnor U28971 (N_28971,N_27420,N_27392);
nor U28972 (N_28972,N_27862,N_27272);
xor U28973 (N_28973,N_27663,N_27740);
nor U28974 (N_28974,N_27016,N_27664);
and U28975 (N_28975,N_27501,N_27605);
and U28976 (N_28976,N_27684,N_27925);
or U28977 (N_28977,N_27371,N_27868);
nor U28978 (N_28978,N_27913,N_27278);
or U28979 (N_28979,N_27996,N_27283);
nor U28980 (N_28980,N_27161,N_27189);
or U28981 (N_28981,N_27923,N_27563);
xor U28982 (N_28982,N_27907,N_27678);
nand U28983 (N_28983,N_27601,N_27400);
nor U28984 (N_28984,N_27880,N_27596);
xor U28985 (N_28985,N_27301,N_27388);
nand U28986 (N_28986,N_27334,N_27861);
xor U28987 (N_28987,N_27538,N_27974);
nor U28988 (N_28988,N_27726,N_27696);
nor U28989 (N_28989,N_27146,N_27841);
or U28990 (N_28990,N_27703,N_27812);
or U28991 (N_28991,N_27424,N_27059);
nor U28992 (N_28992,N_27063,N_27136);
xnor U28993 (N_28993,N_27840,N_27408);
nand U28994 (N_28994,N_27056,N_27214);
nor U28995 (N_28995,N_27762,N_27485);
nor U28996 (N_28996,N_27312,N_27801);
or U28997 (N_28997,N_27579,N_27683);
or U28998 (N_28998,N_27188,N_27587);
or U28999 (N_28999,N_27709,N_27569);
and U29000 (N_29000,N_28426,N_28268);
or U29001 (N_29001,N_28778,N_28471);
nand U29002 (N_29002,N_28877,N_28170);
xnor U29003 (N_29003,N_28896,N_28468);
nand U29004 (N_29004,N_28797,N_28027);
xor U29005 (N_29005,N_28430,N_28502);
xnor U29006 (N_29006,N_28393,N_28727);
nand U29007 (N_29007,N_28205,N_28044);
and U29008 (N_29008,N_28061,N_28334);
and U29009 (N_29009,N_28763,N_28910);
nor U29010 (N_29010,N_28386,N_28233);
or U29011 (N_29011,N_28480,N_28368);
nor U29012 (N_29012,N_28781,N_28932);
xor U29013 (N_29013,N_28382,N_28294);
xor U29014 (N_29014,N_28574,N_28737);
nor U29015 (N_29015,N_28648,N_28521);
and U29016 (N_29016,N_28167,N_28542);
xnor U29017 (N_29017,N_28094,N_28337);
nor U29018 (N_29018,N_28551,N_28228);
xnor U29019 (N_29019,N_28365,N_28056);
nand U29020 (N_29020,N_28377,N_28580);
nand U29021 (N_29021,N_28159,N_28853);
xor U29022 (N_29022,N_28138,N_28768);
or U29023 (N_29023,N_28086,N_28608);
or U29024 (N_29024,N_28692,N_28584);
and U29025 (N_29025,N_28341,N_28688);
and U29026 (N_29026,N_28078,N_28193);
nand U29027 (N_29027,N_28767,N_28133);
or U29028 (N_29028,N_28612,N_28655);
and U29029 (N_29029,N_28746,N_28090);
and U29030 (N_29030,N_28242,N_28567);
xor U29031 (N_29031,N_28474,N_28921);
nor U29032 (N_29032,N_28892,N_28192);
nand U29033 (N_29033,N_28296,N_28728);
or U29034 (N_29034,N_28554,N_28220);
xnor U29035 (N_29035,N_28911,N_28069);
or U29036 (N_29036,N_28741,N_28565);
nor U29037 (N_29037,N_28929,N_28615);
and U29038 (N_29038,N_28195,N_28861);
nor U29039 (N_29039,N_28062,N_28923);
nand U29040 (N_29040,N_28351,N_28376);
xor U29041 (N_29041,N_28844,N_28756);
nand U29042 (N_29042,N_28963,N_28941);
nand U29043 (N_29043,N_28211,N_28018);
nand U29044 (N_29044,N_28662,N_28645);
xor U29045 (N_29045,N_28774,N_28428);
and U29046 (N_29046,N_28845,N_28516);
nand U29047 (N_29047,N_28846,N_28217);
or U29048 (N_29048,N_28623,N_28080);
or U29049 (N_29049,N_28272,N_28405);
or U29050 (N_29050,N_28618,N_28966);
or U29051 (N_29051,N_28886,N_28264);
xnor U29052 (N_29052,N_28742,N_28681);
nand U29053 (N_29053,N_28253,N_28293);
or U29054 (N_29054,N_28239,N_28038);
nand U29055 (N_29055,N_28687,N_28976);
nor U29056 (N_29056,N_28917,N_28524);
nor U29057 (N_29057,N_28026,N_28012);
or U29058 (N_29058,N_28475,N_28409);
or U29059 (N_29059,N_28510,N_28826);
nand U29060 (N_29060,N_28723,N_28811);
nand U29061 (N_29061,N_28606,N_28443);
xnor U29062 (N_29062,N_28964,N_28806);
nand U29063 (N_29063,N_28665,N_28909);
or U29064 (N_29064,N_28011,N_28423);
and U29065 (N_29065,N_28406,N_28734);
nor U29066 (N_29066,N_28482,N_28593);
nand U29067 (N_29067,N_28631,N_28472);
and U29068 (N_29068,N_28749,N_28320);
nor U29069 (N_29069,N_28637,N_28936);
nand U29070 (N_29070,N_28943,N_28375);
and U29071 (N_29071,N_28558,N_28492);
nand U29072 (N_29072,N_28420,N_28547);
nor U29073 (N_29073,N_28456,N_28161);
nand U29074 (N_29074,N_28315,N_28720);
or U29075 (N_29075,N_28125,N_28200);
and U29076 (N_29076,N_28660,N_28980);
and U29077 (N_29077,N_28361,N_28557);
and U29078 (N_29078,N_28503,N_28171);
nand U29079 (N_29079,N_28156,N_28732);
nand U29080 (N_29080,N_28676,N_28336);
nor U29081 (N_29081,N_28355,N_28063);
xor U29082 (N_29082,N_28536,N_28031);
nor U29083 (N_29083,N_28479,N_28476);
xor U29084 (N_29084,N_28863,N_28089);
nor U29085 (N_29085,N_28888,N_28747);
nor U29086 (N_29086,N_28345,N_28110);
xnor U29087 (N_29087,N_28550,N_28979);
xnor U29088 (N_29088,N_28130,N_28632);
or U29089 (N_29089,N_28743,N_28578);
nand U29090 (N_29090,N_28814,N_28883);
nand U29091 (N_29091,N_28023,N_28967);
and U29092 (N_29092,N_28777,N_28391);
nand U29093 (N_29093,N_28396,N_28539);
or U29094 (N_29094,N_28649,N_28187);
and U29095 (N_29095,N_28572,N_28390);
xnor U29096 (N_29096,N_28152,N_28231);
and U29097 (N_29097,N_28962,N_28875);
xnor U29098 (N_29098,N_28893,N_28575);
xor U29099 (N_29099,N_28782,N_28956);
nand U29100 (N_29100,N_28635,N_28280);
or U29101 (N_29101,N_28642,N_28257);
xnor U29102 (N_29102,N_28988,N_28384);
xor U29103 (N_29103,N_28939,N_28537);
and U29104 (N_29104,N_28983,N_28106);
or U29105 (N_29105,N_28633,N_28843);
nor U29106 (N_29106,N_28385,N_28677);
or U29107 (N_29107,N_28650,N_28616);
xnor U29108 (N_29108,N_28670,N_28571);
nand U29109 (N_29109,N_28794,N_28041);
nand U29110 (N_29110,N_28022,N_28407);
xor U29111 (N_29111,N_28099,N_28311);
and U29112 (N_29112,N_28514,N_28952);
xor U29113 (N_29113,N_28064,N_28577);
and U29114 (N_29114,N_28721,N_28899);
nand U29115 (N_29115,N_28849,N_28255);
xnor U29116 (N_29116,N_28169,N_28147);
nand U29117 (N_29117,N_28212,N_28301);
xnor U29118 (N_29118,N_28850,N_28189);
xnor U29119 (N_29119,N_28975,N_28684);
nor U29120 (N_29120,N_28807,N_28006);
xnor U29121 (N_29121,N_28775,N_28058);
nor U29122 (N_29122,N_28517,N_28124);
or U29123 (N_29123,N_28552,N_28329);
nand U29124 (N_29124,N_28977,N_28271);
nor U29125 (N_29125,N_28267,N_28188);
or U29126 (N_29126,N_28674,N_28071);
and U29127 (N_29127,N_28981,N_28190);
or U29128 (N_29128,N_28528,N_28306);
nand U29129 (N_29129,N_28927,N_28869);
nor U29130 (N_29130,N_28278,N_28465);
nand U29131 (N_29131,N_28045,N_28215);
nor U29132 (N_29132,N_28788,N_28994);
nand U29133 (N_29133,N_28088,N_28413);
nand U29134 (N_29134,N_28113,N_28328);
nand U29135 (N_29135,N_28651,N_28411);
nand U29136 (N_29136,N_28232,N_28748);
or U29137 (N_29137,N_28180,N_28431);
xor U29138 (N_29138,N_28596,N_28715);
nor U29139 (N_29139,N_28034,N_28796);
xnor U29140 (N_29140,N_28046,N_28313);
nor U29141 (N_29141,N_28834,N_28226);
and U29142 (N_29142,N_28793,N_28809);
nand U29143 (N_29143,N_28751,N_28609);
nand U29144 (N_29144,N_28444,N_28437);
nor U29145 (N_29145,N_28096,N_28297);
nor U29146 (N_29146,N_28379,N_28639);
xnor U29147 (N_29147,N_28214,N_28820);
nand U29148 (N_29148,N_28644,N_28652);
nand U29149 (N_29149,N_28511,N_28378);
xor U29150 (N_29150,N_28252,N_28135);
nand U29151 (N_29151,N_28559,N_28039);
and U29152 (N_29152,N_28116,N_28776);
or U29153 (N_29153,N_28241,N_28965);
and U29154 (N_29154,N_28523,N_28706);
nor U29155 (N_29155,N_28166,N_28488);
and U29156 (N_29156,N_28245,N_28682);
or U29157 (N_29157,N_28837,N_28750);
nand U29158 (N_29158,N_28813,N_28592);
nand U29159 (N_29159,N_28417,N_28504);
or U29160 (N_29160,N_28455,N_28388);
nand U29161 (N_29161,N_28338,N_28050);
nand U29162 (N_29162,N_28817,N_28326);
nand U29163 (N_29163,N_28305,N_28761);
nor U29164 (N_29164,N_28082,N_28083);
and U29165 (N_29165,N_28590,N_28640);
and U29166 (N_29166,N_28999,N_28601);
nand U29167 (N_29167,N_28425,N_28604);
or U29168 (N_29168,N_28054,N_28803);
xnor U29169 (N_29169,N_28295,N_28851);
nor U29170 (N_29170,N_28597,N_28447);
xnor U29171 (N_29171,N_28889,N_28438);
xor U29172 (N_29172,N_28460,N_28546);
nand U29173 (N_29173,N_28276,N_28122);
and U29174 (N_29174,N_28238,N_28594);
nor U29175 (N_29175,N_28105,N_28172);
or U29176 (N_29176,N_28564,N_28505);
nand U29177 (N_29177,N_28364,N_28545);
and U29178 (N_29178,N_28458,N_28669);
and U29179 (N_29179,N_28408,N_28619);
or U29180 (N_29180,N_28906,N_28209);
or U29181 (N_29181,N_28340,N_28261);
or U29182 (N_29182,N_28701,N_28020);
nand U29183 (N_29183,N_28137,N_28699);
nand U29184 (N_29184,N_28289,N_28555);
or U29185 (N_29185,N_28237,N_28532);
nand U29186 (N_29186,N_28785,N_28136);
nand U29187 (N_29187,N_28191,N_28800);
or U29188 (N_29188,N_28698,N_28638);
xnor U29189 (N_29189,N_28362,N_28760);
and U29190 (N_29190,N_28733,N_28179);
or U29191 (N_29191,N_28653,N_28657);
and U29192 (N_29192,N_28014,N_28128);
nand U29193 (N_29193,N_28766,N_28403);
nand U29194 (N_29194,N_28114,N_28184);
and U29195 (N_29195,N_28835,N_28829);
xnor U29196 (N_29196,N_28867,N_28452);
xor U29197 (N_29197,N_28937,N_28828);
xnor U29198 (N_29198,N_28440,N_28079);
nand U29199 (N_29199,N_28015,N_28881);
xnor U29200 (N_29200,N_28959,N_28779);
xor U29201 (N_29201,N_28387,N_28145);
nor U29202 (N_29202,N_28515,N_28076);
or U29203 (N_29203,N_28954,N_28548);
nand U29204 (N_29204,N_28040,N_28908);
nand U29205 (N_29205,N_28696,N_28489);
xor U29206 (N_29206,N_28412,N_28634);
xor U29207 (N_29207,N_28714,N_28808);
nand U29208 (N_29208,N_28925,N_28483);
nor U29209 (N_29209,N_28501,N_28984);
xor U29210 (N_29210,N_28028,N_28769);
and U29211 (N_29211,N_28628,N_28229);
xnor U29212 (N_29212,N_28816,N_28757);
and U29213 (N_29213,N_28392,N_28182);
and U29214 (N_29214,N_28525,N_28507);
nor U29215 (N_29215,N_28562,N_28993);
and U29216 (N_29216,N_28887,N_28201);
nand U29217 (N_29217,N_28146,N_28457);
nand U29218 (N_29218,N_28541,N_28155);
nor U29219 (N_29219,N_28754,N_28284);
nand U29220 (N_29220,N_28726,N_28093);
nor U29221 (N_29221,N_28569,N_28092);
nand U29222 (N_29222,N_28019,N_28944);
xnor U29223 (N_29223,N_28694,N_28491);
and U29224 (N_29224,N_28581,N_28758);
nand U29225 (N_29225,N_28225,N_28544);
nor U29226 (N_29226,N_28174,N_28711);
or U29227 (N_29227,N_28357,N_28931);
nor U29228 (N_29228,N_28065,N_28010);
or U29229 (N_29229,N_28433,N_28918);
xnor U29230 (N_29230,N_28540,N_28494);
or U29231 (N_29231,N_28697,N_28473);
and U29232 (N_29232,N_28335,N_28947);
and U29233 (N_29233,N_28224,N_28860);
and U29234 (N_29234,N_28266,N_28924);
nor U29235 (N_29235,N_28583,N_28478);
or U29236 (N_29236,N_28589,N_28247);
or U29237 (N_29237,N_28825,N_28804);
xor U29238 (N_29238,N_28907,N_28827);
or U29239 (N_29239,N_28024,N_28210);
xor U29240 (N_29240,N_28163,N_28611);
or U29241 (N_29241,N_28177,N_28422);
and U29242 (N_29242,N_28576,N_28989);
xnor U29243 (N_29243,N_28531,N_28535);
or U29244 (N_29244,N_28709,N_28745);
or U29245 (N_29245,N_28416,N_28350);
xor U29246 (N_29246,N_28765,N_28216);
nor U29247 (N_29247,N_28852,N_28933);
and U29248 (N_29248,N_28500,N_28771);
and U29249 (N_29249,N_28198,N_28705);
xor U29250 (N_29250,N_28968,N_28081);
nand U29251 (N_29251,N_28702,N_28185);
nand U29252 (N_29252,N_28922,N_28996);
or U29253 (N_29253,N_28770,N_28270);
nor U29254 (N_29254,N_28248,N_28970);
nor U29255 (N_29255,N_28493,N_28363);
nor U29256 (N_29256,N_28399,N_28389);
xor U29257 (N_29257,N_28913,N_28207);
and U29258 (N_29258,N_28052,N_28316);
nand U29259 (N_29259,N_28029,N_28928);
nor U29260 (N_29260,N_28486,N_28667);
and U29261 (N_29261,N_28900,N_28453);
and U29262 (N_29262,N_28129,N_28509);
or U29263 (N_29263,N_28288,N_28414);
xnor U29264 (N_29264,N_28789,N_28464);
nor U29265 (N_29265,N_28141,N_28822);
or U29266 (N_29266,N_28495,N_28673);
and U29267 (N_29267,N_28030,N_28077);
and U29268 (N_29268,N_28862,N_28042);
xnor U29269 (N_29269,N_28561,N_28882);
and U29270 (N_29270,N_28343,N_28878);
or U29271 (N_29271,N_28049,N_28281);
and U29272 (N_29272,N_28181,N_28360);
and U29273 (N_29273,N_28973,N_28534);
xor U29274 (N_29274,N_28101,N_28940);
nor U29275 (N_29275,N_28613,N_28164);
or U29276 (N_29276,N_28148,N_28840);
or U29277 (N_29277,N_28068,N_28461);
and U29278 (N_29278,N_28556,N_28327);
and U29279 (N_29279,N_28930,N_28275);
nor U29280 (N_29280,N_28624,N_28066);
xor U29281 (N_29281,N_28158,N_28841);
nand U29282 (N_29282,N_28848,N_28395);
nand U29283 (N_29283,N_28067,N_28057);
xnor U29284 (N_29284,N_28123,N_28462);
and U29285 (N_29285,N_28436,N_28117);
and U29286 (N_29286,N_28259,N_28901);
and U29287 (N_29287,N_28880,N_28945);
xnor U29288 (N_29288,N_28084,N_28173);
and U29289 (N_29289,N_28920,N_28033);
and U29290 (N_29290,N_28710,N_28663);
nor U29291 (N_29291,N_28204,N_28641);
and U29292 (N_29292,N_28339,N_28865);
nor U29293 (N_29293,N_28298,N_28258);
and U29294 (N_29294,N_28810,N_28035);
nor U29295 (N_29295,N_28620,N_28001);
nand U29296 (N_29296,N_28467,N_28730);
and U29297 (N_29297,N_28143,N_28256);
and U29298 (N_29298,N_28251,N_28342);
and U29299 (N_29299,N_28285,N_28394);
or U29300 (N_29300,N_28454,N_28902);
or U29301 (N_29301,N_28787,N_28282);
xnor U29302 (N_29302,N_28234,N_28254);
or U29303 (N_29303,N_28144,N_28002);
nand U29304 (N_29304,N_28346,N_28111);
and U29305 (N_29305,N_28307,N_28672);
or U29306 (N_29306,N_28139,N_28381);
nor U29307 (N_29307,N_28149,N_28004);
nand U29308 (N_29308,N_28151,N_28958);
nand U29309 (N_29309,N_28864,N_28605);
xor U29310 (N_29310,N_28600,N_28330);
and U29311 (N_29311,N_28759,N_28736);
and U29312 (N_29312,N_28695,N_28691);
nor U29313 (N_29313,N_28223,N_28070);
or U29314 (N_29314,N_28260,N_28410);
or U29315 (N_29315,N_28250,N_28358);
and U29316 (N_29316,N_28506,N_28839);
and U29317 (N_29317,N_28538,N_28969);
nand U29318 (N_29318,N_28690,N_28490);
nand U29319 (N_29319,N_28752,N_28997);
or U29320 (N_29320,N_28792,N_28175);
or U29321 (N_29321,N_28898,N_28397);
or U29322 (N_29322,N_28304,N_28919);
nand U29323 (N_29323,N_28961,N_28982);
and U29324 (N_29324,N_28103,N_28643);
nor U29325 (N_29325,N_28549,N_28380);
and U29326 (N_29326,N_28626,N_28036);
xnor U29327 (N_29327,N_28469,N_28838);
xnor U29328 (N_29328,N_28025,N_28055);
nor U29329 (N_29329,N_28683,N_28347);
nor U29330 (N_29330,N_28897,N_28134);
and U29331 (N_29331,N_28048,N_28451);
and U29332 (N_29332,N_28037,N_28625);
nor U29333 (N_29333,N_28712,N_28703);
nor U29334 (N_29334,N_28485,N_28203);
nand U29335 (N_29335,N_28244,N_28871);
nand U29336 (N_29336,N_28277,N_28868);
or U29337 (N_29337,N_28801,N_28007);
xor U29338 (N_29338,N_28664,N_28344);
and U29339 (N_29339,N_28661,N_28118);
nor U29340 (N_29340,N_28780,N_28953);
nor U29341 (N_29341,N_28005,N_28441);
or U29342 (N_29342,N_28499,N_28310);
or U29343 (N_29343,N_28560,N_28053);
nand U29344 (N_29344,N_28009,N_28987);
nor U29345 (N_29345,N_28708,N_28519);
or U29346 (N_29346,N_28526,N_28121);
xnor U29347 (N_29347,N_28273,N_28614);
or U29348 (N_29348,N_28291,N_28197);
xor U29349 (N_29349,N_28529,N_28951);
and U29350 (N_29350,N_28309,N_28283);
xnor U29351 (N_29351,N_28693,N_28629);
or U29352 (N_29352,N_28916,N_28497);
nand U29353 (N_29353,N_28513,N_28317);
nor U29354 (N_29354,N_28353,N_28533);
nand U29355 (N_29355,N_28230,N_28196);
xor U29356 (N_29356,N_28165,N_28891);
and U29357 (N_29357,N_28371,N_28949);
xnor U29358 (N_29358,N_28333,N_28588);
and U29359 (N_29359,N_28354,N_28419);
and U29360 (N_29360,N_28481,N_28885);
nand U29361 (N_29361,N_28303,N_28131);
or U29362 (N_29362,N_28439,N_28373);
xor U29363 (N_29363,N_28716,N_28700);
nor U29364 (N_29364,N_28832,N_28477);
or U29365 (N_29365,N_28262,N_28579);
or U29366 (N_29366,N_28098,N_28636);
and U29367 (N_29367,N_28073,N_28566);
xor U29368 (N_29368,N_28274,N_28895);
xnor U29369 (N_29369,N_28812,N_28269);
xor U29370 (N_29370,N_28263,N_28622);
nor U29371 (N_29371,N_28903,N_28717);
xnor U29372 (N_29372,N_28830,N_28870);
or U29373 (N_29373,N_28383,N_28112);
and U29374 (N_29374,N_28227,N_28322);
nand U29375 (N_29375,N_28942,N_28719);
nor U29376 (N_29376,N_28202,N_28091);
or U29377 (N_29377,N_28915,N_28646);
xor U29378 (N_29378,N_28470,N_28108);
nor U29379 (N_29379,N_28905,N_28168);
xor U29380 (N_29380,N_28934,N_28032);
or U29381 (N_29381,N_28059,N_28790);
nor U29382 (N_29382,N_28568,N_28109);
and U29383 (N_29383,N_28729,N_28823);
or U29384 (N_29384,N_28302,N_28689);
xor U29385 (N_29385,N_28627,N_28400);
and U29386 (N_29386,N_28331,N_28656);
xor U29387 (N_29387,N_28003,N_28213);
nand U29388 (N_29388,N_28127,N_28157);
xnor U29389 (N_29389,N_28735,N_28120);
or U29390 (N_29390,N_28445,N_28602);
nor U29391 (N_29391,N_28359,N_28246);
and U29392 (N_29392,N_28957,N_28819);
or U29393 (N_29393,N_28518,N_28442);
or U29394 (N_29394,N_28265,N_28199);
nand U29395 (N_29395,N_28286,N_28854);
xor U29396 (N_29396,N_28654,N_28107);
xnor U29397 (N_29397,N_28366,N_28985);
nor U29398 (N_29398,N_28427,N_28874);
and U29399 (N_29399,N_28398,N_28434);
xnor U29400 (N_29400,N_28856,N_28591);
xnor U29401 (N_29401,N_28671,N_28658);
nand U29402 (N_29402,N_28016,N_28686);
or U29403 (N_29403,N_28791,N_28332);
xor U29404 (N_29404,N_28974,N_28496);
or U29405 (N_29405,N_28675,N_28773);
nor U29406 (N_29406,N_28432,N_28799);
or U29407 (N_29407,N_28459,N_28960);
nor U29408 (N_29408,N_28308,N_28356);
nand U29409 (N_29409,N_28563,N_28017);
or U29410 (N_29410,N_28178,N_28833);
nor U29411 (N_29411,N_28607,N_28914);
and U29412 (N_29412,N_28312,N_28160);
xnor U29413 (N_29413,N_28986,N_28795);
and U29414 (N_29414,N_28100,N_28318);
nor U29415 (N_29415,N_28194,N_28884);
nor U29416 (N_29416,N_28647,N_28463);
nor U29417 (N_29417,N_28235,N_28527);
or U29418 (N_29418,N_28998,N_28222);
and U29419 (N_29419,N_28739,N_28074);
and U29420 (N_29420,N_28404,N_28610);
or U29421 (N_29421,N_28668,N_28319);
xor U29422 (N_29422,N_28321,N_28522);
nor U29423 (N_29423,N_28249,N_28290);
or U29424 (N_29424,N_28772,N_28842);
xnor U29425 (N_29425,N_28162,N_28132);
xor U29426 (N_29426,N_28369,N_28858);
and U29427 (N_29427,N_28595,N_28582);
nor U29428 (N_29428,N_28876,N_28508);
xor U29429 (N_29429,N_28287,N_28183);
xnor U29430 (N_29430,N_28236,N_28075);
or U29431 (N_29431,N_28314,N_28894);
and U29432 (N_29432,N_28995,N_28324);
or U29433 (N_29433,N_28429,N_28603);
nand U29434 (N_29434,N_28104,N_28466);
nor U29435 (N_29435,N_28821,N_28926);
xnor U29436 (N_29436,N_28008,N_28013);
nand U29437 (N_29437,N_28753,N_28292);
nand U29438 (N_29438,N_28374,N_28587);
xor U29439 (N_29439,N_28043,N_28946);
or U29440 (N_29440,N_28279,N_28085);
or U29441 (N_29441,N_28154,N_28707);
nand U29442 (N_29442,N_28598,N_28421);
nor U29443 (N_29443,N_28859,N_28415);
and U29444 (N_29444,N_28990,N_28352);
and U29445 (N_29445,N_28879,N_28971);
or U29446 (N_29446,N_28784,N_28449);
nor U29447 (N_29447,N_28367,N_28824);
nand U29448 (N_29448,N_28724,N_28553);
or U29449 (N_29449,N_28530,N_28678);
and U29450 (N_29450,N_28866,N_28783);
and U29451 (N_29451,N_28484,N_28685);
nor U29452 (N_29452,N_28176,N_28831);
nor U29453 (N_29453,N_28450,N_28153);
or U29454 (N_29454,N_28722,N_28520);
nand U29455 (N_29455,N_28102,N_28206);
and U29456 (N_29456,N_28764,N_28446);
or U29457 (N_29457,N_28087,N_28573);
nand U29458 (N_29458,N_28000,N_28912);
nor U29459 (N_29459,N_28713,N_28487);
xor U29460 (N_29460,N_28725,N_28978);
nand U29461 (N_29461,N_28704,N_28798);
nand U29462 (N_29462,N_28938,N_28680);
and U29463 (N_29463,N_28762,N_28904);
xnor U29464 (N_29464,N_28872,N_28240);
and U29465 (N_29465,N_28119,N_28348);
nor U29466 (N_29466,N_28095,N_28498);
xor U29467 (N_29467,N_28300,N_28992);
nand U29468 (N_29468,N_28815,N_28219);
and U29469 (N_29469,N_28950,N_28570);
nor U29470 (N_29470,N_28599,N_28744);
or U29471 (N_29471,N_28126,N_28323);
or U29472 (N_29472,N_28805,N_28435);
or U29473 (N_29473,N_28786,N_28047);
nand U29474 (N_29474,N_28512,N_28847);
nor U29475 (N_29475,N_28072,N_28955);
and U29476 (N_29476,N_28991,N_28738);
nand U29477 (N_29477,N_28097,N_28857);
or U29478 (N_29478,N_28243,N_28021);
xor U29479 (N_29479,N_28051,N_28402);
xnor U29480 (N_29480,N_28802,N_28221);
or U29481 (N_29481,N_28666,N_28150);
or U29482 (N_29482,N_28543,N_28401);
or U29483 (N_29483,N_28679,N_28818);
or U29484 (N_29484,N_28659,N_28836);
or U29485 (N_29485,N_28935,N_28972);
and U29486 (N_29486,N_28060,N_28621);
nand U29487 (N_29487,N_28370,N_28218);
nand U29488 (N_29488,N_28424,N_28630);
or U29489 (N_29489,N_28142,N_28115);
nand U29490 (N_29490,N_28349,N_28586);
xnor U29491 (N_29491,N_28890,N_28140);
xor U29492 (N_29492,N_28718,N_28948);
nand U29493 (N_29493,N_28740,N_28731);
xor U29494 (N_29494,N_28873,N_28418);
and U29495 (N_29495,N_28208,N_28755);
xor U29496 (N_29496,N_28325,N_28299);
nand U29497 (N_29497,N_28617,N_28186);
and U29498 (N_29498,N_28448,N_28855);
nor U29499 (N_29499,N_28372,N_28585);
xor U29500 (N_29500,N_28749,N_28372);
and U29501 (N_29501,N_28539,N_28881);
nor U29502 (N_29502,N_28909,N_28782);
or U29503 (N_29503,N_28643,N_28292);
nand U29504 (N_29504,N_28678,N_28419);
xnor U29505 (N_29505,N_28574,N_28060);
and U29506 (N_29506,N_28622,N_28287);
nand U29507 (N_29507,N_28867,N_28618);
and U29508 (N_29508,N_28299,N_28064);
and U29509 (N_29509,N_28450,N_28877);
xnor U29510 (N_29510,N_28416,N_28349);
and U29511 (N_29511,N_28773,N_28676);
or U29512 (N_29512,N_28684,N_28412);
nand U29513 (N_29513,N_28687,N_28575);
nand U29514 (N_29514,N_28252,N_28162);
xnor U29515 (N_29515,N_28665,N_28911);
xnor U29516 (N_29516,N_28357,N_28631);
and U29517 (N_29517,N_28062,N_28194);
nor U29518 (N_29518,N_28425,N_28848);
or U29519 (N_29519,N_28284,N_28064);
nor U29520 (N_29520,N_28378,N_28967);
and U29521 (N_29521,N_28170,N_28226);
nor U29522 (N_29522,N_28387,N_28273);
nor U29523 (N_29523,N_28195,N_28529);
or U29524 (N_29524,N_28902,N_28357);
nand U29525 (N_29525,N_28869,N_28452);
nor U29526 (N_29526,N_28979,N_28451);
nor U29527 (N_29527,N_28069,N_28784);
and U29528 (N_29528,N_28081,N_28526);
nor U29529 (N_29529,N_28170,N_28364);
nor U29530 (N_29530,N_28652,N_28609);
or U29531 (N_29531,N_28209,N_28724);
or U29532 (N_29532,N_28470,N_28729);
and U29533 (N_29533,N_28765,N_28356);
xor U29534 (N_29534,N_28628,N_28960);
and U29535 (N_29535,N_28040,N_28453);
or U29536 (N_29536,N_28695,N_28276);
xor U29537 (N_29537,N_28818,N_28521);
nand U29538 (N_29538,N_28262,N_28956);
xor U29539 (N_29539,N_28180,N_28205);
nand U29540 (N_29540,N_28875,N_28222);
or U29541 (N_29541,N_28167,N_28176);
and U29542 (N_29542,N_28863,N_28652);
or U29543 (N_29543,N_28230,N_28816);
or U29544 (N_29544,N_28094,N_28843);
nand U29545 (N_29545,N_28729,N_28755);
and U29546 (N_29546,N_28036,N_28866);
or U29547 (N_29547,N_28110,N_28248);
nor U29548 (N_29548,N_28326,N_28126);
or U29549 (N_29549,N_28101,N_28213);
xor U29550 (N_29550,N_28066,N_28612);
nand U29551 (N_29551,N_28094,N_28746);
nor U29552 (N_29552,N_28118,N_28936);
nand U29553 (N_29553,N_28631,N_28714);
nor U29554 (N_29554,N_28059,N_28290);
or U29555 (N_29555,N_28793,N_28705);
and U29556 (N_29556,N_28667,N_28927);
xnor U29557 (N_29557,N_28624,N_28385);
nand U29558 (N_29558,N_28065,N_28838);
and U29559 (N_29559,N_28340,N_28784);
nand U29560 (N_29560,N_28629,N_28786);
nor U29561 (N_29561,N_28900,N_28399);
or U29562 (N_29562,N_28086,N_28213);
xnor U29563 (N_29563,N_28402,N_28154);
nor U29564 (N_29564,N_28133,N_28122);
nand U29565 (N_29565,N_28182,N_28144);
xor U29566 (N_29566,N_28314,N_28626);
and U29567 (N_29567,N_28716,N_28719);
and U29568 (N_29568,N_28094,N_28729);
and U29569 (N_29569,N_28286,N_28709);
and U29570 (N_29570,N_28534,N_28422);
nand U29571 (N_29571,N_28351,N_28564);
nor U29572 (N_29572,N_28696,N_28460);
xnor U29573 (N_29573,N_28924,N_28129);
nand U29574 (N_29574,N_28167,N_28175);
nor U29575 (N_29575,N_28520,N_28261);
nor U29576 (N_29576,N_28282,N_28080);
xnor U29577 (N_29577,N_28947,N_28771);
or U29578 (N_29578,N_28593,N_28072);
or U29579 (N_29579,N_28743,N_28474);
nor U29580 (N_29580,N_28212,N_28944);
nor U29581 (N_29581,N_28631,N_28216);
or U29582 (N_29582,N_28369,N_28972);
nor U29583 (N_29583,N_28402,N_28585);
nand U29584 (N_29584,N_28223,N_28021);
xnor U29585 (N_29585,N_28159,N_28554);
xnor U29586 (N_29586,N_28429,N_28288);
nand U29587 (N_29587,N_28215,N_28294);
and U29588 (N_29588,N_28459,N_28098);
or U29589 (N_29589,N_28073,N_28002);
and U29590 (N_29590,N_28033,N_28441);
nor U29591 (N_29591,N_28793,N_28490);
or U29592 (N_29592,N_28859,N_28243);
or U29593 (N_29593,N_28824,N_28688);
or U29594 (N_29594,N_28296,N_28128);
and U29595 (N_29595,N_28451,N_28582);
or U29596 (N_29596,N_28666,N_28618);
nand U29597 (N_29597,N_28080,N_28126);
and U29598 (N_29598,N_28678,N_28132);
nor U29599 (N_29599,N_28848,N_28627);
and U29600 (N_29600,N_28518,N_28492);
and U29601 (N_29601,N_28561,N_28753);
nor U29602 (N_29602,N_28473,N_28290);
or U29603 (N_29603,N_28338,N_28915);
xor U29604 (N_29604,N_28368,N_28357);
or U29605 (N_29605,N_28365,N_28318);
and U29606 (N_29606,N_28898,N_28454);
and U29607 (N_29607,N_28272,N_28852);
nand U29608 (N_29608,N_28189,N_28787);
nand U29609 (N_29609,N_28782,N_28898);
and U29610 (N_29610,N_28358,N_28054);
and U29611 (N_29611,N_28834,N_28656);
nor U29612 (N_29612,N_28376,N_28672);
nand U29613 (N_29613,N_28426,N_28711);
xor U29614 (N_29614,N_28130,N_28818);
nand U29615 (N_29615,N_28461,N_28382);
and U29616 (N_29616,N_28009,N_28718);
nand U29617 (N_29617,N_28027,N_28641);
nand U29618 (N_29618,N_28450,N_28968);
or U29619 (N_29619,N_28996,N_28616);
or U29620 (N_29620,N_28358,N_28330);
xnor U29621 (N_29621,N_28387,N_28422);
xor U29622 (N_29622,N_28616,N_28343);
and U29623 (N_29623,N_28736,N_28326);
xor U29624 (N_29624,N_28962,N_28252);
nand U29625 (N_29625,N_28301,N_28089);
and U29626 (N_29626,N_28129,N_28416);
nand U29627 (N_29627,N_28845,N_28563);
nand U29628 (N_29628,N_28832,N_28411);
nor U29629 (N_29629,N_28069,N_28527);
nor U29630 (N_29630,N_28878,N_28662);
and U29631 (N_29631,N_28143,N_28426);
and U29632 (N_29632,N_28265,N_28986);
nor U29633 (N_29633,N_28458,N_28111);
xnor U29634 (N_29634,N_28157,N_28844);
and U29635 (N_29635,N_28542,N_28789);
xnor U29636 (N_29636,N_28784,N_28338);
nor U29637 (N_29637,N_28161,N_28968);
nand U29638 (N_29638,N_28562,N_28520);
nor U29639 (N_29639,N_28881,N_28941);
or U29640 (N_29640,N_28968,N_28350);
nor U29641 (N_29641,N_28377,N_28937);
xor U29642 (N_29642,N_28579,N_28399);
nor U29643 (N_29643,N_28082,N_28330);
nor U29644 (N_29644,N_28589,N_28304);
xor U29645 (N_29645,N_28068,N_28095);
and U29646 (N_29646,N_28094,N_28762);
xor U29647 (N_29647,N_28391,N_28201);
nor U29648 (N_29648,N_28706,N_28373);
or U29649 (N_29649,N_28609,N_28249);
xnor U29650 (N_29650,N_28719,N_28479);
nor U29651 (N_29651,N_28522,N_28194);
xnor U29652 (N_29652,N_28475,N_28650);
nand U29653 (N_29653,N_28445,N_28245);
and U29654 (N_29654,N_28200,N_28810);
nor U29655 (N_29655,N_28333,N_28336);
or U29656 (N_29656,N_28551,N_28896);
nand U29657 (N_29657,N_28396,N_28395);
xor U29658 (N_29658,N_28076,N_28336);
nor U29659 (N_29659,N_28204,N_28613);
nand U29660 (N_29660,N_28269,N_28430);
xor U29661 (N_29661,N_28593,N_28474);
or U29662 (N_29662,N_28009,N_28341);
nand U29663 (N_29663,N_28900,N_28649);
and U29664 (N_29664,N_28834,N_28693);
or U29665 (N_29665,N_28129,N_28897);
xnor U29666 (N_29666,N_28719,N_28991);
nand U29667 (N_29667,N_28123,N_28635);
and U29668 (N_29668,N_28335,N_28690);
nand U29669 (N_29669,N_28471,N_28650);
or U29670 (N_29670,N_28544,N_28180);
xor U29671 (N_29671,N_28442,N_28128);
xnor U29672 (N_29672,N_28294,N_28359);
nand U29673 (N_29673,N_28921,N_28708);
xnor U29674 (N_29674,N_28268,N_28357);
or U29675 (N_29675,N_28242,N_28506);
nand U29676 (N_29676,N_28620,N_28964);
or U29677 (N_29677,N_28020,N_28153);
nand U29678 (N_29678,N_28914,N_28515);
nand U29679 (N_29679,N_28762,N_28917);
nand U29680 (N_29680,N_28073,N_28571);
xor U29681 (N_29681,N_28498,N_28436);
xor U29682 (N_29682,N_28161,N_28895);
nand U29683 (N_29683,N_28524,N_28022);
nand U29684 (N_29684,N_28863,N_28682);
xor U29685 (N_29685,N_28154,N_28318);
xor U29686 (N_29686,N_28611,N_28081);
or U29687 (N_29687,N_28941,N_28203);
xor U29688 (N_29688,N_28262,N_28426);
nand U29689 (N_29689,N_28100,N_28493);
nand U29690 (N_29690,N_28371,N_28402);
and U29691 (N_29691,N_28215,N_28257);
nand U29692 (N_29692,N_28169,N_28203);
or U29693 (N_29693,N_28799,N_28040);
nand U29694 (N_29694,N_28914,N_28413);
nand U29695 (N_29695,N_28209,N_28453);
and U29696 (N_29696,N_28964,N_28157);
xor U29697 (N_29697,N_28579,N_28627);
or U29698 (N_29698,N_28348,N_28020);
xor U29699 (N_29699,N_28625,N_28752);
xnor U29700 (N_29700,N_28855,N_28785);
or U29701 (N_29701,N_28872,N_28254);
nand U29702 (N_29702,N_28916,N_28862);
or U29703 (N_29703,N_28214,N_28283);
nor U29704 (N_29704,N_28433,N_28418);
or U29705 (N_29705,N_28252,N_28366);
and U29706 (N_29706,N_28538,N_28013);
nand U29707 (N_29707,N_28640,N_28557);
nor U29708 (N_29708,N_28247,N_28527);
xor U29709 (N_29709,N_28839,N_28362);
nor U29710 (N_29710,N_28702,N_28698);
nor U29711 (N_29711,N_28975,N_28045);
nand U29712 (N_29712,N_28510,N_28972);
xnor U29713 (N_29713,N_28478,N_28528);
nor U29714 (N_29714,N_28233,N_28702);
nand U29715 (N_29715,N_28416,N_28388);
xor U29716 (N_29716,N_28925,N_28288);
nor U29717 (N_29717,N_28541,N_28486);
and U29718 (N_29718,N_28182,N_28824);
or U29719 (N_29719,N_28502,N_28642);
xor U29720 (N_29720,N_28948,N_28730);
nor U29721 (N_29721,N_28458,N_28025);
xor U29722 (N_29722,N_28601,N_28245);
nor U29723 (N_29723,N_28345,N_28309);
xnor U29724 (N_29724,N_28172,N_28510);
or U29725 (N_29725,N_28538,N_28232);
or U29726 (N_29726,N_28148,N_28886);
xnor U29727 (N_29727,N_28771,N_28216);
nor U29728 (N_29728,N_28668,N_28985);
nor U29729 (N_29729,N_28048,N_28725);
and U29730 (N_29730,N_28570,N_28738);
and U29731 (N_29731,N_28767,N_28944);
and U29732 (N_29732,N_28213,N_28359);
nor U29733 (N_29733,N_28089,N_28867);
or U29734 (N_29734,N_28367,N_28280);
and U29735 (N_29735,N_28156,N_28452);
nor U29736 (N_29736,N_28203,N_28609);
or U29737 (N_29737,N_28534,N_28057);
or U29738 (N_29738,N_28679,N_28683);
nor U29739 (N_29739,N_28814,N_28505);
or U29740 (N_29740,N_28713,N_28077);
or U29741 (N_29741,N_28779,N_28937);
and U29742 (N_29742,N_28504,N_28041);
nand U29743 (N_29743,N_28506,N_28980);
xnor U29744 (N_29744,N_28634,N_28178);
xnor U29745 (N_29745,N_28579,N_28926);
xnor U29746 (N_29746,N_28447,N_28449);
xnor U29747 (N_29747,N_28375,N_28203);
and U29748 (N_29748,N_28254,N_28389);
nand U29749 (N_29749,N_28846,N_28219);
nand U29750 (N_29750,N_28962,N_28234);
and U29751 (N_29751,N_28794,N_28609);
and U29752 (N_29752,N_28702,N_28590);
nor U29753 (N_29753,N_28203,N_28283);
or U29754 (N_29754,N_28723,N_28999);
and U29755 (N_29755,N_28411,N_28049);
nor U29756 (N_29756,N_28614,N_28504);
or U29757 (N_29757,N_28941,N_28683);
or U29758 (N_29758,N_28217,N_28306);
or U29759 (N_29759,N_28405,N_28341);
or U29760 (N_29760,N_28073,N_28610);
xnor U29761 (N_29761,N_28652,N_28536);
or U29762 (N_29762,N_28922,N_28879);
nor U29763 (N_29763,N_28835,N_28761);
or U29764 (N_29764,N_28623,N_28532);
nand U29765 (N_29765,N_28937,N_28245);
xnor U29766 (N_29766,N_28294,N_28643);
nand U29767 (N_29767,N_28931,N_28540);
or U29768 (N_29768,N_28245,N_28267);
nand U29769 (N_29769,N_28701,N_28279);
and U29770 (N_29770,N_28350,N_28098);
and U29771 (N_29771,N_28922,N_28691);
nand U29772 (N_29772,N_28554,N_28119);
and U29773 (N_29773,N_28670,N_28240);
xnor U29774 (N_29774,N_28909,N_28104);
or U29775 (N_29775,N_28829,N_28474);
xor U29776 (N_29776,N_28362,N_28417);
or U29777 (N_29777,N_28101,N_28608);
or U29778 (N_29778,N_28499,N_28008);
nand U29779 (N_29779,N_28064,N_28959);
xnor U29780 (N_29780,N_28481,N_28238);
nor U29781 (N_29781,N_28289,N_28603);
nor U29782 (N_29782,N_28265,N_28232);
and U29783 (N_29783,N_28570,N_28963);
nor U29784 (N_29784,N_28242,N_28652);
and U29785 (N_29785,N_28442,N_28011);
and U29786 (N_29786,N_28701,N_28756);
or U29787 (N_29787,N_28374,N_28049);
or U29788 (N_29788,N_28253,N_28248);
and U29789 (N_29789,N_28445,N_28601);
and U29790 (N_29790,N_28955,N_28818);
nor U29791 (N_29791,N_28607,N_28518);
nand U29792 (N_29792,N_28026,N_28813);
nor U29793 (N_29793,N_28698,N_28902);
nand U29794 (N_29794,N_28143,N_28517);
nor U29795 (N_29795,N_28116,N_28291);
xor U29796 (N_29796,N_28616,N_28836);
nand U29797 (N_29797,N_28963,N_28374);
nand U29798 (N_29798,N_28680,N_28724);
xor U29799 (N_29799,N_28914,N_28159);
nand U29800 (N_29800,N_28960,N_28837);
xor U29801 (N_29801,N_28798,N_28905);
and U29802 (N_29802,N_28158,N_28031);
xor U29803 (N_29803,N_28788,N_28464);
xor U29804 (N_29804,N_28908,N_28657);
or U29805 (N_29805,N_28890,N_28044);
nor U29806 (N_29806,N_28894,N_28881);
nand U29807 (N_29807,N_28359,N_28452);
nor U29808 (N_29808,N_28098,N_28795);
or U29809 (N_29809,N_28860,N_28106);
nand U29810 (N_29810,N_28113,N_28230);
or U29811 (N_29811,N_28103,N_28306);
nand U29812 (N_29812,N_28580,N_28131);
or U29813 (N_29813,N_28336,N_28365);
xor U29814 (N_29814,N_28430,N_28196);
nor U29815 (N_29815,N_28881,N_28023);
or U29816 (N_29816,N_28398,N_28411);
or U29817 (N_29817,N_28891,N_28374);
nor U29818 (N_29818,N_28315,N_28868);
xnor U29819 (N_29819,N_28826,N_28305);
or U29820 (N_29820,N_28998,N_28224);
or U29821 (N_29821,N_28644,N_28124);
and U29822 (N_29822,N_28631,N_28000);
nor U29823 (N_29823,N_28275,N_28750);
nand U29824 (N_29824,N_28269,N_28978);
and U29825 (N_29825,N_28284,N_28251);
or U29826 (N_29826,N_28402,N_28291);
or U29827 (N_29827,N_28931,N_28573);
nand U29828 (N_29828,N_28740,N_28586);
or U29829 (N_29829,N_28008,N_28529);
nor U29830 (N_29830,N_28077,N_28715);
nand U29831 (N_29831,N_28555,N_28768);
nand U29832 (N_29832,N_28956,N_28675);
and U29833 (N_29833,N_28335,N_28920);
xnor U29834 (N_29834,N_28858,N_28874);
or U29835 (N_29835,N_28394,N_28703);
or U29836 (N_29836,N_28755,N_28988);
xnor U29837 (N_29837,N_28399,N_28520);
or U29838 (N_29838,N_28915,N_28255);
nor U29839 (N_29839,N_28641,N_28877);
nand U29840 (N_29840,N_28907,N_28456);
xor U29841 (N_29841,N_28409,N_28027);
or U29842 (N_29842,N_28176,N_28924);
and U29843 (N_29843,N_28254,N_28327);
or U29844 (N_29844,N_28006,N_28155);
xnor U29845 (N_29845,N_28349,N_28128);
nor U29846 (N_29846,N_28123,N_28769);
nor U29847 (N_29847,N_28108,N_28615);
xor U29848 (N_29848,N_28916,N_28557);
and U29849 (N_29849,N_28748,N_28980);
nand U29850 (N_29850,N_28891,N_28407);
nand U29851 (N_29851,N_28892,N_28615);
nor U29852 (N_29852,N_28002,N_28062);
nor U29853 (N_29853,N_28480,N_28420);
and U29854 (N_29854,N_28086,N_28663);
nor U29855 (N_29855,N_28436,N_28344);
or U29856 (N_29856,N_28344,N_28615);
xor U29857 (N_29857,N_28749,N_28469);
nand U29858 (N_29858,N_28584,N_28040);
and U29859 (N_29859,N_28403,N_28572);
nor U29860 (N_29860,N_28620,N_28537);
nand U29861 (N_29861,N_28239,N_28052);
nand U29862 (N_29862,N_28985,N_28271);
or U29863 (N_29863,N_28447,N_28147);
nor U29864 (N_29864,N_28164,N_28873);
xnor U29865 (N_29865,N_28016,N_28782);
nand U29866 (N_29866,N_28379,N_28538);
or U29867 (N_29867,N_28434,N_28999);
xnor U29868 (N_29868,N_28324,N_28525);
nand U29869 (N_29869,N_28168,N_28868);
or U29870 (N_29870,N_28658,N_28722);
and U29871 (N_29871,N_28116,N_28616);
or U29872 (N_29872,N_28611,N_28954);
nor U29873 (N_29873,N_28178,N_28126);
nand U29874 (N_29874,N_28140,N_28492);
nor U29875 (N_29875,N_28389,N_28511);
and U29876 (N_29876,N_28994,N_28611);
and U29877 (N_29877,N_28302,N_28168);
and U29878 (N_29878,N_28563,N_28944);
nor U29879 (N_29879,N_28787,N_28490);
and U29880 (N_29880,N_28931,N_28961);
nor U29881 (N_29881,N_28158,N_28162);
nand U29882 (N_29882,N_28563,N_28193);
nand U29883 (N_29883,N_28456,N_28429);
xor U29884 (N_29884,N_28161,N_28438);
nand U29885 (N_29885,N_28181,N_28282);
or U29886 (N_29886,N_28338,N_28984);
or U29887 (N_29887,N_28083,N_28329);
nand U29888 (N_29888,N_28656,N_28693);
nor U29889 (N_29889,N_28974,N_28934);
nand U29890 (N_29890,N_28819,N_28446);
nand U29891 (N_29891,N_28559,N_28672);
nor U29892 (N_29892,N_28072,N_28645);
nand U29893 (N_29893,N_28583,N_28714);
or U29894 (N_29894,N_28182,N_28720);
nand U29895 (N_29895,N_28896,N_28929);
nand U29896 (N_29896,N_28769,N_28413);
nor U29897 (N_29897,N_28842,N_28809);
xnor U29898 (N_29898,N_28809,N_28998);
nand U29899 (N_29899,N_28643,N_28687);
or U29900 (N_29900,N_28818,N_28484);
and U29901 (N_29901,N_28189,N_28481);
nand U29902 (N_29902,N_28563,N_28823);
xor U29903 (N_29903,N_28126,N_28084);
or U29904 (N_29904,N_28383,N_28198);
or U29905 (N_29905,N_28128,N_28952);
or U29906 (N_29906,N_28868,N_28210);
nor U29907 (N_29907,N_28895,N_28233);
nor U29908 (N_29908,N_28093,N_28461);
nand U29909 (N_29909,N_28538,N_28454);
and U29910 (N_29910,N_28190,N_28236);
xor U29911 (N_29911,N_28793,N_28758);
xnor U29912 (N_29912,N_28062,N_28302);
nand U29913 (N_29913,N_28466,N_28431);
and U29914 (N_29914,N_28390,N_28255);
nand U29915 (N_29915,N_28871,N_28707);
nor U29916 (N_29916,N_28063,N_28947);
xor U29917 (N_29917,N_28526,N_28244);
or U29918 (N_29918,N_28481,N_28937);
or U29919 (N_29919,N_28918,N_28248);
or U29920 (N_29920,N_28208,N_28748);
nand U29921 (N_29921,N_28870,N_28805);
or U29922 (N_29922,N_28127,N_28827);
nand U29923 (N_29923,N_28629,N_28375);
xnor U29924 (N_29924,N_28007,N_28419);
nand U29925 (N_29925,N_28879,N_28661);
nand U29926 (N_29926,N_28578,N_28444);
nand U29927 (N_29927,N_28051,N_28816);
or U29928 (N_29928,N_28465,N_28792);
or U29929 (N_29929,N_28444,N_28413);
or U29930 (N_29930,N_28464,N_28129);
nor U29931 (N_29931,N_28936,N_28339);
xnor U29932 (N_29932,N_28050,N_28016);
nor U29933 (N_29933,N_28191,N_28434);
nand U29934 (N_29934,N_28326,N_28797);
and U29935 (N_29935,N_28936,N_28061);
nand U29936 (N_29936,N_28316,N_28356);
and U29937 (N_29937,N_28975,N_28891);
nor U29938 (N_29938,N_28733,N_28308);
nand U29939 (N_29939,N_28448,N_28822);
xnor U29940 (N_29940,N_28400,N_28597);
xnor U29941 (N_29941,N_28078,N_28453);
and U29942 (N_29942,N_28763,N_28914);
xor U29943 (N_29943,N_28329,N_28445);
nor U29944 (N_29944,N_28064,N_28666);
and U29945 (N_29945,N_28699,N_28455);
nand U29946 (N_29946,N_28772,N_28210);
nand U29947 (N_29947,N_28890,N_28249);
nand U29948 (N_29948,N_28524,N_28081);
and U29949 (N_29949,N_28037,N_28732);
or U29950 (N_29950,N_28308,N_28473);
xor U29951 (N_29951,N_28862,N_28439);
or U29952 (N_29952,N_28037,N_28666);
or U29953 (N_29953,N_28206,N_28474);
and U29954 (N_29954,N_28099,N_28874);
nand U29955 (N_29955,N_28626,N_28562);
nand U29956 (N_29956,N_28785,N_28700);
nand U29957 (N_29957,N_28172,N_28114);
nor U29958 (N_29958,N_28964,N_28784);
nor U29959 (N_29959,N_28268,N_28878);
or U29960 (N_29960,N_28712,N_28728);
xnor U29961 (N_29961,N_28196,N_28501);
xor U29962 (N_29962,N_28224,N_28051);
nor U29963 (N_29963,N_28018,N_28920);
nand U29964 (N_29964,N_28584,N_28873);
xnor U29965 (N_29965,N_28655,N_28255);
xor U29966 (N_29966,N_28107,N_28839);
or U29967 (N_29967,N_28673,N_28190);
xor U29968 (N_29968,N_28193,N_28874);
nand U29969 (N_29969,N_28576,N_28259);
xnor U29970 (N_29970,N_28225,N_28968);
nor U29971 (N_29971,N_28291,N_28627);
or U29972 (N_29972,N_28945,N_28613);
xor U29973 (N_29973,N_28862,N_28430);
xnor U29974 (N_29974,N_28591,N_28758);
nor U29975 (N_29975,N_28143,N_28093);
nand U29976 (N_29976,N_28381,N_28587);
nor U29977 (N_29977,N_28582,N_28633);
nor U29978 (N_29978,N_28518,N_28003);
or U29979 (N_29979,N_28512,N_28129);
and U29980 (N_29980,N_28058,N_28302);
xor U29981 (N_29981,N_28561,N_28643);
nand U29982 (N_29982,N_28639,N_28885);
or U29983 (N_29983,N_28447,N_28110);
and U29984 (N_29984,N_28860,N_28866);
nand U29985 (N_29985,N_28986,N_28562);
nor U29986 (N_29986,N_28995,N_28168);
xor U29987 (N_29987,N_28281,N_28517);
xnor U29988 (N_29988,N_28444,N_28498);
or U29989 (N_29989,N_28682,N_28226);
xor U29990 (N_29990,N_28111,N_28548);
or U29991 (N_29991,N_28512,N_28365);
xnor U29992 (N_29992,N_28998,N_28063);
or U29993 (N_29993,N_28559,N_28782);
or U29994 (N_29994,N_28324,N_28659);
xnor U29995 (N_29995,N_28764,N_28746);
xnor U29996 (N_29996,N_28623,N_28667);
and U29997 (N_29997,N_28001,N_28175);
xor U29998 (N_29998,N_28029,N_28419);
and U29999 (N_29999,N_28810,N_28748);
nor U30000 (N_30000,N_29409,N_29921);
nand U30001 (N_30001,N_29764,N_29232);
xnor U30002 (N_30002,N_29662,N_29203);
and U30003 (N_30003,N_29236,N_29710);
or U30004 (N_30004,N_29144,N_29121);
and U30005 (N_30005,N_29931,N_29396);
and U30006 (N_30006,N_29923,N_29102);
and U30007 (N_30007,N_29111,N_29075);
nor U30008 (N_30008,N_29979,N_29344);
or U30009 (N_30009,N_29508,N_29216);
nor U30010 (N_30010,N_29272,N_29847);
and U30011 (N_30011,N_29960,N_29310);
nor U30012 (N_30012,N_29432,N_29224);
xnor U30013 (N_30013,N_29400,N_29909);
nor U30014 (N_30014,N_29407,N_29114);
nand U30015 (N_30015,N_29501,N_29023);
xnor U30016 (N_30016,N_29066,N_29094);
or U30017 (N_30017,N_29564,N_29420);
or U30018 (N_30018,N_29674,N_29273);
and U30019 (N_30019,N_29585,N_29763);
xor U30020 (N_30020,N_29774,N_29520);
nor U30021 (N_30021,N_29324,N_29187);
nor U30022 (N_30022,N_29108,N_29349);
nand U30023 (N_30023,N_29802,N_29255);
xor U30024 (N_30024,N_29748,N_29362);
or U30025 (N_30025,N_29447,N_29715);
nand U30026 (N_30026,N_29575,N_29410);
xor U30027 (N_30027,N_29659,N_29481);
and U30028 (N_30028,N_29222,N_29381);
or U30029 (N_30029,N_29028,N_29772);
nand U30030 (N_30030,N_29598,N_29168);
nand U30031 (N_30031,N_29097,N_29241);
and U30032 (N_30032,N_29178,N_29128);
xor U30033 (N_30033,N_29142,N_29403);
and U30034 (N_30034,N_29237,N_29596);
nand U30035 (N_30035,N_29374,N_29587);
nand U30036 (N_30036,N_29630,N_29424);
xor U30037 (N_30037,N_29051,N_29213);
nor U30038 (N_30038,N_29717,N_29819);
and U30039 (N_30039,N_29716,N_29656);
nor U30040 (N_30040,N_29436,N_29513);
or U30041 (N_30041,N_29820,N_29767);
nor U30042 (N_30042,N_29737,N_29391);
and U30043 (N_30043,N_29570,N_29528);
nand U30044 (N_30044,N_29299,N_29711);
xnor U30045 (N_30045,N_29000,N_29067);
xor U30046 (N_30046,N_29405,N_29679);
nand U30047 (N_30047,N_29597,N_29506);
nand U30048 (N_30048,N_29221,N_29906);
and U30049 (N_30049,N_29437,N_29190);
and U30050 (N_30050,N_29164,N_29101);
or U30051 (N_30051,N_29328,N_29866);
and U30052 (N_30052,N_29929,N_29495);
nand U30053 (N_30053,N_29298,N_29001);
nor U30054 (N_30054,N_29292,N_29683);
or U30055 (N_30055,N_29924,N_29846);
xnor U30056 (N_30056,N_29226,N_29088);
nor U30057 (N_30057,N_29153,N_29617);
nor U30058 (N_30058,N_29208,N_29690);
and U30059 (N_30059,N_29115,N_29078);
or U30060 (N_30060,N_29427,N_29803);
and U30061 (N_30061,N_29070,N_29193);
nand U30062 (N_30062,N_29619,N_29799);
nand U30063 (N_30063,N_29331,N_29395);
nor U30064 (N_30064,N_29635,N_29354);
nor U30065 (N_30065,N_29318,N_29093);
and U30066 (N_30066,N_29859,N_29995);
or U30067 (N_30067,N_29813,N_29548);
xnor U30068 (N_30068,N_29538,N_29179);
xnor U30069 (N_30069,N_29884,N_29608);
nor U30070 (N_30070,N_29430,N_29071);
or U30071 (N_30071,N_29283,N_29138);
nand U30072 (N_30072,N_29282,N_29964);
or U30073 (N_30073,N_29855,N_29275);
xnor U30074 (N_30074,N_29453,N_29245);
xnor U30075 (N_30075,N_29473,N_29456);
and U30076 (N_30076,N_29531,N_29912);
or U30077 (N_30077,N_29810,N_29189);
or U30078 (N_30078,N_29522,N_29346);
or U30079 (N_30079,N_29933,N_29080);
xnor U30080 (N_30080,N_29652,N_29129);
xor U30081 (N_30081,N_29439,N_29512);
and U30082 (N_30082,N_29479,N_29330);
xor U30083 (N_30083,N_29966,N_29347);
xnor U30084 (N_30084,N_29441,N_29239);
xor U30085 (N_30085,N_29691,N_29351);
nand U30086 (N_30086,N_29519,N_29760);
and U30087 (N_30087,N_29042,N_29852);
and U30088 (N_30088,N_29689,N_29712);
xnor U30089 (N_30089,N_29972,N_29758);
and U30090 (N_30090,N_29126,N_29910);
or U30091 (N_30091,N_29687,N_29262);
and U30092 (N_30092,N_29759,N_29254);
and U30093 (N_30093,N_29851,N_29919);
or U30094 (N_30094,N_29735,N_29613);
and U30095 (N_30095,N_29937,N_29918);
xnor U30096 (N_30096,N_29083,N_29697);
nor U30097 (N_30097,N_29326,N_29895);
and U30098 (N_30098,N_29704,N_29151);
xor U30099 (N_30099,N_29584,N_29305);
and U30100 (N_30100,N_29625,N_29804);
or U30101 (N_30101,N_29640,N_29744);
nand U30102 (N_30102,N_29276,N_29798);
and U30103 (N_30103,N_29301,N_29590);
and U30104 (N_30104,N_29337,N_29822);
nand U30105 (N_30105,N_29137,N_29350);
nand U30106 (N_30106,N_29998,N_29100);
xnor U30107 (N_30107,N_29053,N_29206);
nand U30108 (N_30108,N_29369,N_29647);
or U30109 (N_30109,N_29333,N_29302);
xnor U30110 (N_30110,N_29940,N_29387);
and U30111 (N_30111,N_29056,N_29278);
nand U30112 (N_30112,N_29853,N_29844);
and U30113 (N_30113,N_29699,N_29174);
nor U30114 (N_30114,N_29824,N_29365);
and U30115 (N_30115,N_29146,N_29974);
xnor U30116 (N_30116,N_29228,N_29633);
or U30117 (N_30117,N_29818,N_29821);
nor U30118 (N_30118,N_29376,N_29366);
xor U30119 (N_30119,N_29371,N_29729);
nor U30120 (N_30120,N_29665,N_29849);
nand U30121 (N_30121,N_29095,N_29306);
nor U30122 (N_30122,N_29285,N_29728);
xnor U30123 (N_30123,N_29750,N_29487);
xor U30124 (N_30124,N_29762,N_29377);
xor U30125 (N_30125,N_29470,N_29044);
or U30126 (N_30126,N_29279,N_29269);
and U30127 (N_30127,N_29443,N_29181);
xnor U30128 (N_30128,N_29890,N_29594);
nand U30129 (N_30129,N_29010,N_29418);
and U30130 (N_30130,N_29464,N_29989);
nand U30131 (N_30131,N_29110,N_29971);
nor U30132 (N_30132,N_29505,N_29266);
nand U30133 (N_30133,N_29807,N_29314);
and U30134 (N_30134,N_29398,N_29708);
nor U30135 (N_30135,N_29552,N_29719);
or U30136 (N_30136,N_29796,N_29465);
and U30137 (N_30137,N_29503,N_29943);
nor U30138 (N_30138,N_29141,N_29185);
or U30139 (N_30139,N_29877,N_29848);
nand U30140 (N_30140,N_29626,N_29031);
xor U30141 (N_30141,N_29816,N_29104);
nor U30142 (N_30142,N_29364,N_29951);
nor U30143 (N_30143,N_29209,N_29609);
nor U30144 (N_30144,N_29145,N_29671);
and U30145 (N_30145,N_29274,N_29357);
nor U30146 (N_30146,N_29288,N_29198);
and U30147 (N_30147,N_29860,N_29057);
nor U30148 (N_30148,N_29850,N_29593);
or U30149 (N_30149,N_29476,N_29650);
xor U30150 (N_30150,N_29064,N_29021);
or U30151 (N_30151,N_29261,N_29450);
xor U30152 (N_30152,N_29466,N_29657);
xor U30153 (N_30153,N_29646,N_29812);
xnor U30154 (N_30154,N_29707,N_29219);
xnor U30155 (N_30155,N_29233,N_29058);
nor U30156 (N_30156,N_29834,N_29303);
xor U30157 (N_30157,N_29545,N_29361);
xor U30158 (N_30158,N_29170,N_29313);
nand U30159 (N_30159,N_29079,N_29338);
and U30160 (N_30160,N_29257,N_29991);
or U30161 (N_30161,N_29002,N_29060);
and U30162 (N_30162,N_29036,N_29565);
nand U30163 (N_30163,N_29680,N_29211);
and U30164 (N_30164,N_29856,N_29186);
or U30165 (N_30165,N_29461,N_29681);
nor U30166 (N_30166,N_29527,N_29359);
or U30167 (N_30167,N_29876,N_29184);
nand U30168 (N_30168,N_29124,N_29547);
and U30169 (N_30169,N_29891,N_29573);
and U30170 (N_30170,N_29016,N_29908);
nor U30171 (N_30171,N_29325,N_29634);
nand U30172 (N_30172,N_29627,N_29582);
or U30173 (N_30173,N_29014,N_29988);
nor U30174 (N_30174,N_29251,N_29636);
xnor U30175 (N_30175,N_29835,N_29692);
nor U30176 (N_30176,N_29158,N_29823);
or U30177 (N_30177,N_29618,N_29768);
xnor U30178 (N_30178,N_29462,N_29106);
nand U30179 (N_30179,N_29839,N_29382);
xnor U30180 (N_30180,N_29380,N_29591);
or U30181 (N_30181,N_29458,N_29188);
and U30182 (N_30182,N_29030,N_29970);
nor U30183 (N_30183,N_29388,N_29084);
xnor U30184 (N_30184,N_29757,N_29913);
and U30185 (N_30185,N_29831,N_29004);
nor U30186 (N_30186,N_29162,N_29576);
nor U30187 (N_30187,N_29459,N_29342);
nor U30188 (N_30188,N_29862,N_29246);
nand U30189 (N_30189,N_29984,N_29034);
and U30190 (N_30190,N_29235,N_29637);
nand U30191 (N_30191,N_29526,N_29858);
or U30192 (N_30192,N_29800,N_29837);
xor U30193 (N_30193,N_29770,N_29900);
nor U30194 (N_30194,N_29355,N_29392);
xnor U30195 (N_30195,N_29980,N_29752);
xnor U30196 (N_30196,N_29210,N_29502);
and U30197 (N_30197,N_29399,N_29705);
nand U30198 (N_30198,N_29435,N_29007);
nand U30199 (N_30199,N_29358,N_29006);
nor U30200 (N_30200,N_29581,N_29322);
nor U30201 (N_30201,N_29902,N_29069);
nand U30202 (N_30202,N_29082,N_29811);
nor U30203 (N_30203,N_29611,N_29176);
nand U30204 (N_30204,N_29037,N_29947);
and U30205 (N_30205,N_29480,N_29560);
nand U30206 (N_30206,N_29730,N_29589);
or U30207 (N_30207,N_29944,N_29808);
or U30208 (N_30208,N_29726,N_29871);
xnor U30209 (N_30209,N_29309,N_29578);
nor U30210 (N_30210,N_29903,N_29588);
or U30211 (N_30211,N_29277,N_29214);
and U30212 (N_30212,N_29265,N_29063);
nor U30213 (N_30213,N_29996,N_29242);
or U30214 (N_30214,N_29854,N_29732);
and U30215 (N_30215,N_29041,N_29494);
nor U30216 (N_30216,N_29978,N_29655);
nor U30217 (N_30217,N_29651,N_29880);
xnor U30218 (N_30218,N_29826,N_29928);
xor U30219 (N_30219,N_29727,N_29055);
or U30220 (N_30220,N_29167,N_29661);
xnor U30221 (N_30221,N_29562,N_29673);
and U30222 (N_30222,N_29207,N_29696);
or U30223 (N_30223,N_29290,N_29706);
or U30224 (N_30224,N_29892,N_29217);
nand U30225 (N_30225,N_29148,N_29997);
or U30226 (N_30226,N_29434,N_29340);
nand U30227 (N_30227,N_29537,N_29442);
nand U30228 (N_30228,N_29791,N_29348);
xnor U30229 (N_30229,N_29663,N_29356);
or U30230 (N_30230,N_29412,N_29163);
xor U30231 (N_30231,N_29452,N_29676);
xnor U30232 (N_30232,N_29801,N_29054);
or U30233 (N_30233,N_29040,N_29183);
nand U30234 (N_30234,N_29509,N_29092);
nor U30235 (N_30235,N_29507,N_29378);
and U30236 (N_30236,N_29043,N_29857);
nor U30237 (N_30237,N_29927,N_29518);
nor U30238 (N_30238,N_29601,N_29815);
and U30239 (N_30239,N_29047,N_29243);
nor U30240 (N_30240,N_29244,N_29270);
or U30241 (N_30241,N_29402,N_29539);
and U30242 (N_30242,N_29343,N_29334);
and U30243 (N_30243,N_29161,N_29238);
nand U30244 (N_30244,N_29579,N_29113);
xor U30245 (N_30245,N_29032,N_29414);
nand U30246 (N_30246,N_29253,N_29515);
xor U30247 (N_30247,N_29982,N_29052);
and U30248 (N_30248,N_29887,N_29521);
and U30249 (N_30249,N_29878,N_29958);
xor U30250 (N_30250,N_29645,N_29249);
xnor U30251 (N_30251,N_29809,N_29714);
nand U30252 (N_30252,N_29786,N_29499);
or U30253 (N_30253,N_29577,N_29523);
nor U30254 (N_30254,N_29670,N_29199);
and U30255 (N_30255,N_29561,N_29315);
nor U30256 (N_30256,N_29828,N_29467);
or U30257 (N_30257,N_29510,N_29686);
nor U30258 (N_30258,N_29150,N_29999);
xor U30259 (N_30259,N_29899,N_29990);
nand U30260 (N_30260,N_29477,N_29485);
or U30261 (N_30261,N_29742,N_29870);
or U30262 (N_30262,N_29841,N_29894);
or U30263 (N_30263,N_29965,N_29898);
nor U30264 (N_30264,N_29307,N_29907);
and U30265 (N_30265,N_29091,N_29725);
nand U30266 (N_30266,N_29131,N_29781);
nor U30267 (N_30267,N_29949,N_29740);
nand U30268 (N_30268,N_29033,N_29604);
nor U30269 (N_30269,N_29685,N_29486);
or U30270 (N_30270,N_29643,N_29220);
xnor U30271 (N_30271,N_29920,N_29039);
or U30272 (N_30272,N_29879,N_29516);
or U30273 (N_30273,N_29205,N_29905);
nor U30274 (N_30274,N_29155,N_29017);
nand U30275 (N_30275,N_29836,N_29360);
nand U30276 (N_30276,N_29778,N_29574);
and U30277 (N_30277,N_29484,N_29543);
nand U30278 (N_30278,N_29134,N_29780);
nand U30279 (N_30279,N_29688,N_29789);
xor U30280 (N_30280,N_29535,N_29463);
or U30281 (N_30281,N_29621,N_29504);
or U30282 (N_30282,N_29152,N_29336);
xor U30283 (N_30283,N_29015,N_29817);
xor U30284 (N_30284,N_29401,N_29352);
nand U30285 (N_30285,N_29733,N_29829);
and U30286 (N_30286,N_29612,N_29406);
nand U30287 (N_30287,N_29660,N_29747);
nor U30288 (N_30288,N_29250,N_29901);
and U30289 (N_30289,N_29248,N_29620);
nand U30290 (N_30290,N_29022,N_29648);
and U30291 (N_30291,N_29086,N_29160);
and U30292 (N_30292,N_29098,N_29624);
or U30293 (N_30293,N_29975,N_29433);
and U30294 (N_30294,N_29827,N_29335);
nor U30295 (N_30295,N_29460,N_29792);
nor U30296 (N_30296,N_29329,N_29968);
or U30297 (N_30297,N_29379,N_29667);
or U30298 (N_30298,N_29746,N_29976);
or U30299 (N_30299,N_29644,N_29557);
nor U30300 (N_30300,N_29132,N_29474);
nand U30301 (N_30301,N_29428,N_29438);
nand U30302 (N_30302,N_29293,N_29215);
nand U30303 (N_30303,N_29875,N_29109);
nor U30304 (N_30304,N_29986,N_29544);
xnor U30305 (N_30305,N_29073,N_29546);
nand U30306 (N_30306,N_29784,N_29602);
and U30307 (N_30307,N_29606,N_29089);
and U30308 (N_30308,N_29917,N_29166);
or U30309 (N_30309,N_29267,N_29769);
nand U30310 (N_30310,N_29468,N_29204);
nor U30311 (N_30311,N_29953,N_29431);
or U30312 (N_30312,N_29925,N_29195);
and U30313 (N_30313,N_29658,N_29281);
xnor U30314 (N_30314,N_29955,N_29076);
or U30315 (N_30315,N_29311,N_29922);
nor U30316 (N_30316,N_29739,N_29038);
and U30317 (N_30317,N_29223,N_29026);
or U30318 (N_30318,N_29081,N_29191);
or U30319 (N_30319,N_29957,N_29446);
nor U30320 (N_30320,N_29629,N_29771);
xor U30321 (N_30321,N_29316,N_29175);
nor U30322 (N_30322,N_29832,N_29372);
or U30323 (N_30323,N_29120,N_29682);
or U30324 (N_30324,N_29194,N_29616);
nor U30325 (N_30325,N_29904,N_29050);
and U30326 (N_30326,N_29632,N_29698);
nor U30327 (N_30327,N_29230,N_29389);
and U30328 (N_30328,N_29247,N_29312);
xnor U30329 (N_30329,N_29074,N_29814);
or U30330 (N_30330,N_29709,N_29049);
nor U30331 (N_30331,N_29896,N_29469);
xnor U30332 (N_30332,N_29668,N_29099);
xnor U30333 (N_30333,N_29218,N_29926);
or U30334 (N_30334,N_29872,N_29678);
or U30335 (N_30335,N_29046,N_29133);
and U30336 (N_30336,N_29702,N_29173);
nand U30337 (N_30337,N_29795,N_29559);
or U30338 (N_30338,N_29775,N_29946);
nor U30339 (N_30339,N_29289,N_29756);
or U30340 (N_30340,N_29783,N_29787);
xnor U30341 (N_30341,N_29753,N_29993);
or U30342 (N_30342,N_29429,N_29568);
or U30343 (N_30343,N_29411,N_29271);
nand U30344 (N_30344,N_29572,N_29893);
and U30345 (N_30345,N_29096,N_29404);
nand U30346 (N_30346,N_29059,N_29003);
xor U30347 (N_30347,N_29868,N_29765);
xnor U30348 (N_30348,N_29422,N_29229);
nor U30349 (N_30349,N_29669,N_29264);
or U30350 (N_30350,N_29734,N_29553);
nor U30351 (N_30351,N_29182,N_29258);
nor U30352 (N_30352,N_29962,N_29284);
and U30353 (N_30353,N_29840,N_29493);
or U30354 (N_30354,N_29259,N_29451);
or U30355 (N_30355,N_29291,N_29731);
nor U30356 (N_30356,N_29294,N_29534);
xnor U30357 (N_30357,N_29983,N_29319);
nand U30358 (N_30358,N_29024,N_29883);
xor U30359 (N_30359,N_29603,N_29833);
and U30360 (N_30360,N_29845,N_29018);
and U30361 (N_30361,N_29149,N_29751);
nor U30362 (N_30362,N_29642,N_29200);
and U30363 (N_30363,N_29595,N_29754);
nor U30364 (N_30364,N_29062,N_29297);
nand U30365 (N_30365,N_29384,N_29530);
nand U30366 (N_30366,N_29694,N_29788);
xnor U30367 (N_30367,N_29196,N_29571);
nor U30368 (N_30368,N_29440,N_29197);
xnor U30369 (N_30369,N_29779,N_29722);
or U30370 (N_30370,N_29449,N_29136);
and U30371 (N_30371,N_29009,N_29599);
nand U30372 (N_30372,N_29586,N_29454);
and U30373 (N_30373,N_29125,N_29785);
and U30374 (N_30374,N_29280,N_29672);
or U30375 (N_30375,N_29308,N_29304);
xnor U30376 (N_30376,N_29415,N_29533);
and U30377 (N_30377,N_29317,N_29511);
and U30378 (N_30378,N_29421,N_29127);
nand U30379 (N_30379,N_29448,N_29103);
and U30380 (N_30380,N_29367,N_29478);
and U30381 (N_30381,N_29117,N_29939);
and U30382 (N_30382,N_29863,N_29724);
nand U30383 (N_30383,N_29112,N_29386);
nor U30384 (N_30384,N_29061,N_29029);
nand U30385 (N_30385,N_29143,N_29177);
xnor U30386 (N_30386,N_29777,N_29790);
nor U30387 (N_30387,N_29745,N_29268);
or U30388 (N_30388,N_29713,N_29256);
nand U30389 (N_30389,N_29025,N_29390);
and U30390 (N_30390,N_29703,N_29339);
nand U30391 (N_30391,N_29445,N_29171);
nor U30392 (N_30392,N_29628,N_29556);
or U30393 (N_30393,N_29072,N_29130);
or U30394 (N_30394,N_29345,N_29455);
xnor U30395 (N_30395,N_29889,N_29483);
and U30396 (N_30396,N_29723,N_29825);
and U30397 (N_30397,N_29843,N_29550);
and U30398 (N_30398,N_29985,N_29981);
nor U30399 (N_30399,N_29566,N_29934);
or U30400 (N_30400,N_29260,N_29773);
xor U30401 (N_30401,N_29492,N_29373);
or U30402 (N_30402,N_29555,N_29393);
nor U30403 (N_30403,N_29897,N_29695);
or U30404 (N_30404,N_29045,N_29738);
nor U30405 (N_30405,N_29567,N_29419);
xor U30406 (N_30406,N_29558,N_29065);
xor U30407 (N_30407,N_29741,N_29911);
nor U30408 (N_30408,N_29967,N_29416);
nor U30409 (N_30409,N_29491,N_29375);
nor U30410 (N_30410,N_29874,N_29649);
xor U30411 (N_30411,N_29408,N_29225);
nand U30412 (N_30412,N_29529,N_29105);
or U30413 (N_30413,N_29240,N_29180);
or U30414 (N_30414,N_29743,N_29524);
nor U30415 (N_30415,N_29936,N_29135);
and U30416 (N_30416,N_29413,N_29323);
nand U30417 (N_30417,N_29013,N_29631);
or U30418 (N_30418,N_29987,N_29677);
nor U30419 (N_30419,N_29011,N_29157);
nand U30420 (N_30420,N_29118,N_29019);
nor U30421 (N_30421,N_29930,N_29915);
or U30422 (N_30422,N_29623,N_29607);
and U30423 (N_30423,N_29749,N_29948);
or U30424 (N_30424,N_29797,N_29761);
and U30425 (N_30425,N_29363,N_29700);
and U30426 (N_30426,N_29551,N_29532);
and U30427 (N_30427,N_29327,N_29498);
nor U30428 (N_30428,N_29488,N_29638);
or U30429 (N_30429,N_29426,N_29457);
xor U30430 (N_30430,N_29332,N_29782);
xor U30431 (N_30431,N_29489,N_29554);
xor U30432 (N_30432,N_29397,N_29718);
nor U30433 (N_30433,N_29701,N_29385);
and U30434 (N_30434,N_29736,N_29540);
nor U30435 (N_30435,N_29869,N_29615);
nor U30436 (N_30436,N_29838,N_29212);
xor U30437 (N_30437,N_29963,N_29497);
xnor U30438 (N_30438,N_29720,N_29793);
or U30439 (N_30439,N_29942,N_29341);
nor U30440 (N_30440,N_29035,N_29881);
xor U30441 (N_30441,N_29992,N_29012);
and U30442 (N_30442,N_29563,N_29954);
xnor U30443 (N_30443,N_29776,N_29952);
and U30444 (N_30444,N_29592,N_29864);
or U30445 (N_30445,N_29296,N_29549);
xnor U30446 (N_30446,N_29472,N_29156);
and U30447 (N_30447,N_29961,N_29172);
nand U30448 (N_30448,N_29300,N_29471);
or U30449 (N_30449,N_29087,N_29159);
or U30450 (N_30450,N_29542,N_29916);
nor U30451 (N_30451,N_29941,N_29490);
and U30452 (N_30452,N_29865,N_29027);
xnor U30453 (N_30453,N_29295,N_29370);
nand U30454 (N_30454,N_29517,N_29048);
nor U30455 (N_30455,N_29583,N_29614);
and U30456 (N_30456,N_29500,N_29201);
and U30457 (N_30457,N_29580,N_29541);
and U30458 (N_30458,N_29320,N_29423);
nand U30459 (N_30459,N_29202,N_29938);
nor U30460 (N_30460,N_29475,N_29514);
and U30461 (N_30461,N_29861,N_29654);
xnor U30462 (N_30462,N_29885,N_29252);
nand U30463 (N_30463,N_29394,N_29664);
or U30464 (N_30464,N_29231,N_29639);
and U30465 (N_30465,N_29119,N_29482);
xnor U30466 (N_30466,N_29569,N_29417);
nor U30467 (N_30467,N_29994,N_29165);
xor U30468 (N_30468,N_29192,N_29287);
nand U30469 (N_30469,N_29842,N_29977);
xor U30470 (N_30470,N_29122,N_29085);
nand U30471 (N_30471,N_29077,N_29444);
xnor U30472 (N_30472,N_29684,N_29794);
or U30473 (N_30473,N_29068,N_29721);
nor U30474 (N_30474,N_29641,N_29959);
nand U30475 (N_30475,N_29169,N_29286);
and U30476 (N_30476,N_29830,N_29605);
nand U30477 (N_30477,N_29914,N_29116);
xor U30478 (N_30478,N_29935,N_29368);
or U30479 (N_30479,N_29969,N_29263);
or U30480 (N_30480,N_29873,N_29867);
nand U30481 (N_30481,N_29950,N_29154);
nor U30482 (N_30482,N_29806,N_29600);
nand U30483 (N_30483,N_29234,N_29882);
or U30484 (N_30484,N_29107,N_29932);
xnor U30485 (N_30485,N_29622,N_29139);
nor U30486 (N_30486,N_29693,N_29227);
and U30487 (N_30487,N_29805,N_29886);
or U30488 (N_30488,N_29956,N_29140);
and U30489 (N_30489,N_29425,N_29383);
xor U30490 (N_30490,N_29666,N_29766);
nor U30491 (N_30491,N_29353,N_29525);
or U30492 (N_30492,N_29610,N_29147);
nor U30493 (N_30493,N_29675,N_29536);
xor U30494 (N_30494,N_29123,N_29888);
nand U30495 (N_30495,N_29321,N_29755);
and U30496 (N_30496,N_29008,N_29973);
nor U30497 (N_30497,N_29005,N_29090);
or U30498 (N_30498,N_29020,N_29496);
nand U30499 (N_30499,N_29945,N_29653);
nor U30500 (N_30500,N_29561,N_29648);
and U30501 (N_30501,N_29650,N_29319);
nand U30502 (N_30502,N_29091,N_29563);
nand U30503 (N_30503,N_29043,N_29538);
and U30504 (N_30504,N_29188,N_29693);
nand U30505 (N_30505,N_29841,N_29333);
or U30506 (N_30506,N_29287,N_29764);
or U30507 (N_30507,N_29297,N_29063);
and U30508 (N_30508,N_29448,N_29437);
and U30509 (N_30509,N_29653,N_29040);
or U30510 (N_30510,N_29161,N_29200);
xor U30511 (N_30511,N_29363,N_29810);
xor U30512 (N_30512,N_29144,N_29733);
nand U30513 (N_30513,N_29637,N_29639);
nand U30514 (N_30514,N_29075,N_29561);
nor U30515 (N_30515,N_29450,N_29936);
nand U30516 (N_30516,N_29787,N_29820);
nor U30517 (N_30517,N_29643,N_29700);
or U30518 (N_30518,N_29942,N_29601);
nor U30519 (N_30519,N_29156,N_29428);
xor U30520 (N_30520,N_29917,N_29465);
and U30521 (N_30521,N_29499,N_29085);
xnor U30522 (N_30522,N_29712,N_29656);
nor U30523 (N_30523,N_29403,N_29421);
nor U30524 (N_30524,N_29250,N_29096);
xnor U30525 (N_30525,N_29697,N_29018);
and U30526 (N_30526,N_29126,N_29642);
xor U30527 (N_30527,N_29794,N_29485);
nand U30528 (N_30528,N_29396,N_29218);
or U30529 (N_30529,N_29741,N_29509);
or U30530 (N_30530,N_29924,N_29681);
xnor U30531 (N_30531,N_29595,N_29939);
nand U30532 (N_30532,N_29679,N_29915);
or U30533 (N_30533,N_29337,N_29276);
nor U30534 (N_30534,N_29286,N_29609);
xor U30535 (N_30535,N_29917,N_29622);
nor U30536 (N_30536,N_29378,N_29071);
or U30537 (N_30537,N_29471,N_29624);
nand U30538 (N_30538,N_29135,N_29651);
xnor U30539 (N_30539,N_29292,N_29433);
and U30540 (N_30540,N_29734,N_29012);
nor U30541 (N_30541,N_29912,N_29923);
and U30542 (N_30542,N_29917,N_29586);
xor U30543 (N_30543,N_29668,N_29116);
and U30544 (N_30544,N_29489,N_29705);
or U30545 (N_30545,N_29124,N_29505);
nand U30546 (N_30546,N_29320,N_29359);
or U30547 (N_30547,N_29499,N_29854);
nor U30548 (N_30548,N_29406,N_29844);
nor U30549 (N_30549,N_29119,N_29380);
or U30550 (N_30550,N_29890,N_29286);
nand U30551 (N_30551,N_29417,N_29647);
and U30552 (N_30552,N_29248,N_29861);
nand U30553 (N_30553,N_29005,N_29662);
or U30554 (N_30554,N_29453,N_29893);
or U30555 (N_30555,N_29829,N_29757);
and U30556 (N_30556,N_29532,N_29144);
nand U30557 (N_30557,N_29549,N_29080);
nor U30558 (N_30558,N_29299,N_29598);
xnor U30559 (N_30559,N_29525,N_29767);
nand U30560 (N_30560,N_29234,N_29372);
xor U30561 (N_30561,N_29954,N_29045);
nand U30562 (N_30562,N_29102,N_29906);
nor U30563 (N_30563,N_29506,N_29831);
or U30564 (N_30564,N_29513,N_29869);
xor U30565 (N_30565,N_29163,N_29535);
xnor U30566 (N_30566,N_29353,N_29234);
and U30567 (N_30567,N_29975,N_29865);
nor U30568 (N_30568,N_29877,N_29700);
nand U30569 (N_30569,N_29552,N_29586);
xor U30570 (N_30570,N_29945,N_29164);
nor U30571 (N_30571,N_29700,N_29339);
or U30572 (N_30572,N_29436,N_29181);
xnor U30573 (N_30573,N_29478,N_29680);
or U30574 (N_30574,N_29966,N_29655);
xnor U30575 (N_30575,N_29533,N_29274);
nand U30576 (N_30576,N_29973,N_29229);
or U30577 (N_30577,N_29364,N_29341);
nor U30578 (N_30578,N_29015,N_29657);
xor U30579 (N_30579,N_29595,N_29534);
or U30580 (N_30580,N_29177,N_29394);
nand U30581 (N_30581,N_29078,N_29988);
xor U30582 (N_30582,N_29868,N_29906);
nor U30583 (N_30583,N_29727,N_29848);
nor U30584 (N_30584,N_29982,N_29654);
xor U30585 (N_30585,N_29078,N_29319);
xor U30586 (N_30586,N_29516,N_29642);
nand U30587 (N_30587,N_29937,N_29136);
or U30588 (N_30588,N_29895,N_29660);
nor U30589 (N_30589,N_29413,N_29006);
and U30590 (N_30590,N_29048,N_29039);
or U30591 (N_30591,N_29088,N_29351);
xnor U30592 (N_30592,N_29993,N_29142);
and U30593 (N_30593,N_29803,N_29086);
nand U30594 (N_30594,N_29800,N_29050);
nand U30595 (N_30595,N_29825,N_29132);
xnor U30596 (N_30596,N_29047,N_29977);
or U30597 (N_30597,N_29292,N_29247);
nor U30598 (N_30598,N_29562,N_29147);
nand U30599 (N_30599,N_29303,N_29950);
or U30600 (N_30600,N_29108,N_29722);
xor U30601 (N_30601,N_29510,N_29379);
and U30602 (N_30602,N_29191,N_29277);
nand U30603 (N_30603,N_29910,N_29538);
and U30604 (N_30604,N_29594,N_29969);
xnor U30605 (N_30605,N_29416,N_29694);
nor U30606 (N_30606,N_29685,N_29014);
xor U30607 (N_30607,N_29624,N_29706);
nand U30608 (N_30608,N_29441,N_29691);
nor U30609 (N_30609,N_29732,N_29238);
and U30610 (N_30610,N_29138,N_29219);
and U30611 (N_30611,N_29036,N_29228);
xor U30612 (N_30612,N_29014,N_29117);
xor U30613 (N_30613,N_29210,N_29764);
nand U30614 (N_30614,N_29985,N_29448);
nand U30615 (N_30615,N_29271,N_29015);
xnor U30616 (N_30616,N_29131,N_29175);
nor U30617 (N_30617,N_29433,N_29313);
xnor U30618 (N_30618,N_29583,N_29238);
nand U30619 (N_30619,N_29536,N_29726);
xor U30620 (N_30620,N_29962,N_29820);
and U30621 (N_30621,N_29839,N_29582);
nand U30622 (N_30622,N_29031,N_29943);
nand U30623 (N_30623,N_29177,N_29139);
and U30624 (N_30624,N_29925,N_29314);
nor U30625 (N_30625,N_29053,N_29236);
xnor U30626 (N_30626,N_29385,N_29497);
nand U30627 (N_30627,N_29939,N_29771);
and U30628 (N_30628,N_29608,N_29623);
nand U30629 (N_30629,N_29864,N_29055);
nand U30630 (N_30630,N_29852,N_29668);
nand U30631 (N_30631,N_29978,N_29576);
nand U30632 (N_30632,N_29312,N_29845);
xor U30633 (N_30633,N_29132,N_29060);
xnor U30634 (N_30634,N_29694,N_29938);
xnor U30635 (N_30635,N_29824,N_29967);
and U30636 (N_30636,N_29255,N_29249);
nand U30637 (N_30637,N_29804,N_29103);
xor U30638 (N_30638,N_29123,N_29504);
xor U30639 (N_30639,N_29413,N_29044);
or U30640 (N_30640,N_29694,N_29306);
or U30641 (N_30641,N_29683,N_29734);
xor U30642 (N_30642,N_29772,N_29902);
and U30643 (N_30643,N_29373,N_29234);
nor U30644 (N_30644,N_29623,N_29685);
xnor U30645 (N_30645,N_29753,N_29336);
nand U30646 (N_30646,N_29873,N_29465);
nor U30647 (N_30647,N_29705,N_29848);
xnor U30648 (N_30648,N_29547,N_29981);
xnor U30649 (N_30649,N_29953,N_29440);
nor U30650 (N_30650,N_29421,N_29626);
nand U30651 (N_30651,N_29030,N_29768);
nand U30652 (N_30652,N_29067,N_29314);
or U30653 (N_30653,N_29367,N_29258);
and U30654 (N_30654,N_29972,N_29885);
and U30655 (N_30655,N_29360,N_29993);
and U30656 (N_30656,N_29844,N_29122);
nor U30657 (N_30657,N_29847,N_29749);
xor U30658 (N_30658,N_29998,N_29866);
nor U30659 (N_30659,N_29996,N_29431);
or U30660 (N_30660,N_29620,N_29748);
nand U30661 (N_30661,N_29220,N_29804);
nor U30662 (N_30662,N_29567,N_29990);
and U30663 (N_30663,N_29220,N_29802);
nor U30664 (N_30664,N_29305,N_29852);
nor U30665 (N_30665,N_29392,N_29579);
nor U30666 (N_30666,N_29804,N_29360);
and U30667 (N_30667,N_29830,N_29401);
and U30668 (N_30668,N_29901,N_29329);
nand U30669 (N_30669,N_29735,N_29093);
xor U30670 (N_30670,N_29252,N_29175);
nor U30671 (N_30671,N_29026,N_29318);
and U30672 (N_30672,N_29117,N_29400);
and U30673 (N_30673,N_29035,N_29999);
and U30674 (N_30674,N_29211,N_29460);
nor U30675 (N_30675,N_29415,N_29378);
and U30676 (N_30676,N_29675,N_29350);
and U30677 (N_30677,N_29784,N_29418);
and U30678 (N_30678,N_29246,N_29771);
nor U30679 (N_30679,N_29953,N_29107);
nand U30680 (N_30680,N_29363,N_29928);
and U30681 (N_30681,N_29499,N_29051);
nand U30682 (N_30682,N_29362,N_29636);
and U30683 (N_30683,N_29330,N_29265);
xnor U30684 (N_30684,N_29925,N_29266);
nand U30685 (N_30685,N_29196,N_29304);
and U30686 (N_30686,N_29735,N_29064);
xor U30687 (N_30687,N_29981,N_29513);
nand U30688 (N_30688,N_29336,N_29717);
and U30689 (N_30689,N_29576,N_29408);
and U30690 (N_30690,N_29949,N_29257);
xor U30691 (N_30691,N_29209,N_29246);
and U30692 (N_30692,N_29874,N_29556);
xnor U30693 (N_30693,N_29879,N_29092);
or U30694 (N_30694,N_29195,N_29621);
nor U30695 (N_30695,N_29323,N_29474);
nand U30696 (N_30696,N_29680,N_29668);
nand U30697 (N_30697,N_29989,N_29013);
and U30698 (N_30698,N_29370,N_29804);
or U30699 (N_30699,N_29447,N_29321);
or U30700 (N_30700,N_29724,N_29773);
nand U30701 (N_30701,N_29903,N_29509);
xnor U30702 (N_30702,N_29671,N_29786);
nand U30703 (N_30703,N_29601,N_29955);
nor U30704 (N_30704,N_29795,N_29496);
and U30705 (N_30705,N_29228,N_29444);
nor U30706 (N_30706,N_29215,N_29322);
nor U30707 (N_30707,N_29176,N_29060);
xnor U30708 (N_30708,N_29825,N_29638);
nor U30709 (N_30709,N_29652,N_29305);
nor U30710 (N_30710,N_29409,N_29031);
or U30711 (N_30711,N_29722,N_29559);
nand U30712 (N_30712,N_29447,N_29719);
or U30713 (N_30713,N_29243,N_29913);
and U30714 (N_30714,N_29419,N_29960);
xor U30715 (N_30715,N_29966,N_29305);
or U30716 (N_30716,N_29093,N_29987);
xnor U30717 (N_30717,N_29173,N_29890);
or U30718 (N_30718,N_29840,N_29262);
or U30719 (N_30719,N_29328,N_29196);
or U30720 (N_30720,N_29183,N_29618);
nor U30721 (N_30721,N_29410,N_29381);
or U30722 (N_30722,N_29765,N_29545);
or U30723 (N_30723,N_29912,N_29497);
or U30724 (N_30724,N_29194,N_29945);
nor U30725 (N_30725,N_29127,N_29294);
xor U30726 (N_30726,N_29856,N_29839);
nand U30727 (N_30727,N_29879,N_29614);
nand U30728 (N_30728,N_29871,N_29948);
nand U30729 (N_30729,N_29024,N_29380);
nor U30730 (N_30730,N_29753,N_29701);
and U30731 (N_30731,N_29397,N_29524);
nand U30732 (N_30732,N_29013,N_29124);
nand U30733 (N_30733,N_29430,N_29528);
or U30734 (N_30734,N_29454,N_29303);
and U30735 (N_30735,N_29901,N_29125);
nand U30736 (N_30736,N_29534,N_29374);
xor U30737 (N_30737,N_29202,N_29130);
and U30738 (N_30738,N_29533,N_29047);
or U30739 (N_30739,N_29825,N_29457);
xnor U30740 (N_30740,N_29750,N_29119);
and U30741 (N_30741,N_29046,N_29773);
nor U30742 (N_30742,N_29139,N_29050);
nand U30743 (N_30743,N_29287,N_29943);
xor U30744 (N_30744,N_29729,N_29645);
or U30745 (N_30745,N_29277,N_29842);
nor U30746 (N_30746,N_29731,N_29928);
xor U30747 (N_30747,N_29218,N_29555);
nor U30748 (N_30748,N_29354,N_29297);
or U30749 (N_30749,N_29564,N_29184);
nand U30750 (N_30750,N_29381,N_29194);
xnor U30751 (N_30751,N_29708,N_29759);
and U30752 (N_30752,N_29316,N_29751);
nand U30753 (N_30753,N_29477,N_29685);
xor U30754 (N_30754,N_29496,N_29713);
xnor U30755 (N_30755,N_29774,N_29108);
nand U30756 (N_30756,N_29940,N_29464);
nand U30757 (N_30757,N_29230,N_29276);
and U30758 (N_30758,N_29200,N_29669);
or U30759 (N_30759,N_29644,N_29533);
nand U30760 (N_30760,N_29226,N_29970);
nand U30761 (N_30761,N_29166,N_29614);
or U30762 (N_30762,N_29983,N_29575);
or U30763 (N_30763,N_29761,N_29075);
and U30764 (N_30764,N_29535,N_29069);
xnor U30765 (N_30765,N_29859,N_29917);
nor U30766 (N_30766,N_29172,N_29682);
nor U30767 (N_30767,N_29968,N_29337);
nor U30768 (N_30768,N_29952,N_29866);
xnor U30769 (N_30769,N_29949,N_29440);
xor U30770 (N_30770,N_29116,N_29736);
or U30771 (N_30771,N_29806,N_29221);
xor U30772 (N_30772,N_29251,N_29237);
and U30773 (N_30773,N_29798,N_29433);
nand U30774 (N_30774,N_29669,N_29406);
and U30775 (N_30775,N_29444,N_29331);
nand U30776 (N_30776,N_29858,N_29560);
and U30777 (N_30777,N_29482,N_29425);
xor U30778 (N_30778,N_29247,N_29176);
nand U30779 (N_30779,N_29987,N_29277);
xor U30780 (N_30780,N_29604,N_29238);
xor U30781 (N_30781,N_29778,N_29382);
or U30782 (N_30782,N_29808,N_29067);
xor U30783 (N_30783,N_29828,N_29756);
or U30784 (N_30784,N_29386,N_29344);
nand U30785 (N_30785,N_29440,N_29599);
nand U30786 (N_30786,N_29155,N_29139);
and U30787 (N_30787,N_29913,N_29221);
or U30788 (N_30788,N_29559,N_29497);
and U30789 (N_30789,N_29345,N_29259);
and U30790 (N_30790,N_29368,N_29090);
nand U30791 (N_30791,N_29292,N_29925);
and U30792 (N_30792,N_29592,N_29749);
or U30793 (N_30793,N_29234,N_29552);
and U30794 (N_30794,N_29017,N_29425);
or U30795 (N_30795,N_29320,N_29071);
and U30796 (N_30796,N_29044,N_29306);
xnor U30797 (N_30797,N_29555,N_29014);
nor U30798 (N_30798,N_29046,N_29470);
and U30799 (N_30799,N_29566,N_29808);
nand U30800 (N_30800,N_29811,N_29715);
or U30801 (N_30801,N_29904,N_29476);
nand U30802 (N_30802,N_29161,N_29683);
xnor U30803 (N_30803,N_29874,N_29582);
xnor U30804 (N_30804,N_29566,N_29843);
or U30805 (N_30805,N_29250,N_29522);
nor U30806 (N_30806,N_29061,N_29962);
nor U30807 (N_30807,N_29847,N_29981);
nand U30808 (N_30808,N_29575,N_29447);
or U30809 (N_30809,N_29367,N_29989);
nand U30810 (N_30810,N_29868,N_29258);
nor U30811 (N_30811,N_29553,N_29174);
nand U30812 (N_30812,N_29846,N_29754);
or U30813 (N_30813,N_29092,N_29273);
nand U30814 (N_30814,N_29683,N_29556);
nor U30815 (N_30815,N_29489,N_29398);
xor U30816 (N_30816,N_29713,N_29341);
and U30817 (N_30817,N_29486,N_29700);
xnor U30818 (N_30818,N_29311,N_29150);
or U30819 (N_30819,N_29323,N_29714);
nand U30820 (N_30820,N_29703,N_29330);
xnor U30821 (N_30821,N_29816,N_29168);
and U30822 (N_30822,N_29489,N_29651);
nand U30823 (N_30823,N_29362,N_29249);
or U30824 (N_30824,N_29684,N_29820);
xor U30825 (N_30825,N_29181,N_29601);
nand U30826 (N_30826,N_29205,N_29645);
nor U30827 (N_30827,N_29003,N_29813);
or U30828 (N_30828,N_29040,N_29377);
nand U30829 (N_30829,N_29973,N_29416);
and U30830 (N_30830,N_29622,N_29940);
xor U30831 (N_30831,N_29065,N_29505);
or U30832 (N_30832,N_29366,N_29882);
xor U30833 (N_30833,N_29965,N_29880);
or U30834 (N_30834,N_29217,N_29861);
nand U30835 (N_30835,N_29227,N_29182);
or U30836 (N_30836,N_29245,N_29491);
nor U30837 (N_30837,N_29738,N_29047);
nor U30838 (N_30838,N_29417,N_29788);
and U30839 (N_30839,N_29029,N_29912);
nand U30840 (N_30840,N_29272,N_29248);
and U30841 (N_30841,N_29510,N_29895);
xnor U30842 (N_30842,N_29674,N_29711);
nand U30843 (N_30843,N_29014,N_29489);
nand U30844 (N_30844,N_29890,N_29433);
nor U30845 (N_30845,N_29544,N_29509);
and U30846 (N_30846,N_29861,N_29040);
or U30847 (N_30847,N_29463,N_29868);
nor U30848 (N_30848,N_29916,N_29785);
and U30849 (N_30849,N_29973,N_29709);
xor U30850 (N_30850,N_29344,N_29840);
nor U30851 (N_30851,N_29763,N_29228);
or U30852 (N_30852,N_29652,N_29920);
xnor U30853 (N_30853,N_29200,N_29110);
nor U30854 (N_30854,N_29097,N_29900);
or U30855 (N_30855,N_29788,N_29872);
or U30856 (N_30856,N_29439,N_29119);
xor U30857 (N_30857,N_29182,N_29337);
or U30858 (N_30858,N_29460,N_29036);
nor U30859 (N_30859,N_29714,N_29634);
or U30860 (N_30860,N_29284,N_29476);
xor U30861 (N_30861,N_29901,N_29979);
and U30862 (N_30862,N_29397,N_29792);
nand U30863 (N_30863,N_29998,N_29910);
nand U30864 (N_30864,N_29405,N_29959);
nor U30865 (N_30865,N_29483,N_29416);
or U30866 (N_30866,N_29694,N_29799);
or U30867 (N_30867,N_29487,N_29459);
nor U30868 (N_30868,N_29933,N_29614);
nor U30869 (N_30869,N_29813,N_29714);
and U30870 (N_30870,N_29009,N_29681);
nor U30871 (N_30871,N_29149,N_29553);
nor U30872 (N_30872,N_29686,N_29422);
nor U30873 (N_30873,N_29030,N_29048);
and U30874 (N_30874,N_29928,N_29766);
nand U30875 (N_30875,N_29776,N_29947);
xnor U30876 (N_30876,N_29247,N_29366);
nor U30877 (N_30877,N_29407,N_29993);
and U30878 (N_30878,N_29619,N_29657);
nor U30879 (N_30879,N_29524,N_29533);
nor U30880 (N_30880,N_29857,N_29623);
and U30881 (N_30881,N_29816,N_29506);
and U30882 (N_30882,N_29968,N_29433);
or U30883 (N_30883,N_29756,N_29457);
nand U30884 (N_30884,N_29962,N_29551);
or U30885 (N_30885,N_29390,N_29446);
or U30886 (N_30886,N_29255,N_29358);
or U30887 (N_30887,N_29361,N_29993);
nor U30888 (N_30888,N_29748,N_29287);
or U30889 (N_30889,N_29383,N_29377);
xor U30890 (N_30890,N_29456,N_29705);
nor U30891 (N_30891,N_29453,N_29613);
and U30892 (N_30892,N_29839,N_29259);
xnor U30893 (N_30893,N_29246,N_29250);
nand U30894 (N_30894,N_29151,N_29699);
or U30895 (N_30895,N_29150,N_29352);
nor U30896 (N_30896,N_29025,N_29687);
and U30897 (N_30897,N_29608,N_29807);
nand U30898 (N_30898,N_29139,N_29427);
nor U30899 (N_30899,N_29311,N_29020);
nand U30900 (N_30900,N_29803,N_29793);
nor U30901 (N_30901,N_29980,N_29623);
or U30902 (N_30902,N_29542,N_29047);
nor U30903 (N_30903,N_29772,N_29967);
xnor U30904 (N_30904,N_29902,N_29196);
xnor U30905 (N_30905,N_29656,N_29012);
nor U30906 (N_30906,N_29798,N_29139);
and U30907 (N_30907,N_29982,N_29617);
xor U30908 (N_30908,N_29421,N_29508);
and U30909 (N_30909,N_29829,N_29616);
or U30910 (N_30910,N_29026,N_29210);
xor U30911 (N_30911,N_29603,N_29885);
xnor U30912 (N_30912,N_29592,N_29898);
nand U30913 (N_30913,N_29462,N_29195);
nor U30914 (N_30914,N_29811,N_29013);
xor U30915 (N_30915,N_29093,N_29970);
nor U30916 (N_30916,N_29571,N_29138);
nand U30917 (N_30917,N_29604,N_29433);
and U30918 (N_30918,N_29780,N_29684);
nand U30919 (N_30919,N_29634,N_29011);
nor U30920 (N_30920,N_29638,N_29519);
nand U30921 (N_30921,N_29345,N_29603);
xnor U30922 (N_30922,N_29853,N_29027);
or U30923 (N_30923,N_29011,N_29845);
nor U30924 (N_30924,N_29177,N_29560);
nor U30925 (N_30925,N_29885,N_29502);
and U30926 (N_30926,N_29846,N_29048);
nor U30927 (N_30927,N_29423,N_29026);
nor U30928 (N_30928,N_29359,N_29285);
xor U30929 (N_30929,N_29826,N_29154);
or U30930 (N_30930,N_29694,N_29418);
nor U30931 (N_30931,N_29277,N_29910);
or U30932 (N_30932,N_29301,N_29061);
nand U30933 (N_30933,N_29730,N_29970);
xor U30934 (N_30934,N_29208,N_29057);
nand U30935 (N_30935,N_29035,N_29037);
or U30936 (N_30936,N_29919,N_29749);
or U30937 (N_30937,N_29379,N_29481);
xor U30938 (N_30938,N_29349,N_29804);
or U30939 (N_30939,N_29690,N_29127);
nand U30940 (N_30940,N_29702,N_29396);
or U30941 (N_30941,N_29869,N_29483);
or U30942 (N_30942,N_29388,N_29299);
or U30943 (N_30943,N_29952,N_29090);
nor U30944 (N_30944,N_29161,N_29623);
and U30945 (N_30945,N_29902,N_29496);
and U30946 (N_30946,N_29514,N_29030);
and U30947 (N_30947,N_29876,N_29067);
and U30948 (N_30948,N_29195,N_29604);
and U30949 (N_30949,N_29393,N_29772);
or U30950 (N_30950,N_29805,N_29721);
and U30951 (N_30951,N_29616,N_29797);
xnor U30952 (N_30952,N_29600,N_29916);
and U30953 (N_30953,N_29437,N_29893);
xor U30954 (N_30954,N_29318,N_29907);
xor U30955 (N_30955,N_29640,N_29565);
or U30956 (N_30956,N_29544,N_29578);
or U30957 (N_30957,N_29749,N_29068);
or U30958 (N_30958,N_29213,N_29260);
and U30959 (N_30959,N_29549,N_29237);
nor U30960 (N_30960,N_29373,N_29340);
xor U30961 (N_30961,N_29859,N_29008);
xnor U30962 (N_30962,N_29558,N_29691);
nor U30963 (N_30963,N_29909,N_29300);
xor U30964 (N_30964,N_29185,N_29874);
nand U30965 (N_30965,N_29665,N_29463);
nor U30966 (N_30966,N_29167,N_29691);
nand U30967 (N_30967,N_29376,N_29546);
nor U30968 (N_30968,N_29352,N_29749);
or U30969 (N_30969,N_29797,N_29692);
and U30970 (N_30970,N_29985,N_29493);
and U30971 (N_30971,N_29916,N_29951);
nor U30972 (N_30972,N_29005,N_29657);
xor U30973 (N_30973,N_29887,N_29431);
or U30974 (N_30974,N_29170,N_29289);
xor U30975 (N_30975,N_29354,N_29038);
or U30976 (N_30976,N_29572,N_29888);
xor U30977 (N_30977,N_29034,N_29490);
nor U30978 (N_30978,N_29197,N_29895);
nor U30979 (N_30979,N_29516,N_29541);
or U30980 (N_30980,N_29944,N_29948);
or U30981 (N_30981,N_29524,N_29725);
nand U30982 (N_30982,N_29465,N_29425);
nor U30983 (N_30983,N_29975,N_29009);
and U30984 (N_30984,N_29285,N_29641);
and U30985 (N_30985,N_29736,N_29635);
nor U30986 (N_30986,N_29559,N_29277);
or U30987 (N_30987,N_29342,N_29383);
or U30988 (N_30988,N_29268,N_29283);
nor U30989 (N_30989,N_29469,N_29322);
nor U30990 (N_30990,N_29604,N_29053);
and U30991 (N_30991,N_29373,N_29272);
and U30992 (N_30992,N_29541,N_29354);
nor U30993 (N_30993,N_29075,N_29892);
nand U30994 (N_30994,N_29645,N_29383);
nand U30995 (N_30995,N_29453,N_29074);
and U30996 (N_30996,N_29659,N_29742);
nand U30997 (N_30997,N_29011,N_29557);
nor U30998 (N_30998,N_29769,N_29168);
or U30999 (N_30999,N_29292,N_29020);
xor U31000 (N_31000,N_30245,N_30599);
nand U31001 (N_31001,N_30182,N_30088);
nor U31002 (N_31002,N_30218,N_30870);
xor U31003 (N_31003,N_30013,N_30117);
nor U31004 (N_31004,N_30583,N_30416);
nor U31005 (N_31005,N_30615,N_30390);
xor U31006 (N_31006,N_30109,N_30550);
nor U31007 (N_31007,N_30467,N_30370);
nand U31008 (N_31008,N_30662,N_30494);
xor U31009 (N_31009,N_30388,N_30816);
nand U31010 (N_31010,N_30728,N_30696);
nand U31011 (N_31011,N_30092,N_30329);
nand U31012 (N_31012,N_30824,N_30908);
and U31013 (N_31013,N_30246,N_30078);
xor U31014 (N_31014,N_30898,N_30593);
or U31015 (N_31015,N_30429,N_30282);
and U31016 (N_31016,N_30313,N_30353);
nor U31017 (N_31017,N_30845,N_30977);
nor U31018 (N_31018,N_30451,N_30000);
xor U31019 (N_31019,N_30251,N_30236);
nor U31020 (N_31020,N_30255,N_30498);
and U31021 (N_31021,N_30945,N_30697);
and U31022 (N_31022,N_30521,N_30412);
and U31023 (N_31023,N_30985,N_30463);
and U31024 (N_31024,N_30315,N_30764);
or U31025 (N_31025,N_30380,N_30126);
xor U31026 (N_31026,N_30219,N_30719);
nor U31027 (N_31027,N_30374,N_30448);
and U31028 (N_31028,N_30375,N_30886);
nand U31029 (N_31029,N_30426,N_30651);
xor U31030 (N_31030,N_30565,N_30317);
and U31031 (N_31031,N_30130,N_30179);
nor U31032 (N_31032,N_30614,N_30872);
nand U31033 (N_31033,N_30227,N_30865);
or U31034 (N_31034,N_30569,N_30576);
and U31035 (N_31035,N_30685,N_30501);
and U31036 (N_31036,N_30616,N_30938);
nand U31037 (N_31037,N_30570,N_30609);
xor U31038 (N_31038,N_30224,N_30398);
and U31039 (N_31039,N_30488,N_30176);
xnor U31040 (N_31040,N_30237,N_30676);
nand U31041 (N_31041,N_30479,N_30811);
nor U31042 (N_31042,N_30331,N_30554);
nor U31043 (N_31043,N_30699,N_30619);
nor U31044 (N_31044,N_30950,N_30248);
or U31045 (N_31045,N_30392,N_30622);
nor U31046 (N_31046,N_30667,N_30165);
and U31047 (N_31047,N_30956,N_30196);
nor U31048 (N_31048,N_30532,N_30529);
and U31049 (N_31049,N_30447,N_30827);
or U31050 (N_31050,N_30803,N_30613);
nand U31051 (N_31051,N_30597,N_30926);
nand U31052 (N_31052,N_30540,N_30981);
xor U31053 (N_31053,N_30105,N_30516);
xnor U31054 (N_31054,N_30828,N_30156);
and U31055 (N_31055,N_30202,N_30239);
and U31056 (N_31056,N_30914,N_30316);
or U31057 (N_31057,N_30354,N_30743);
or U31058 (N_31058,N_30362,N_30805);
xor U31059 (N_31059,N_30818,N_30393);
or U31060 (N_31060,N_30031,N_30480);
and U31061 (N_31061,N_30919,N_30940);
nor U31062 (N_31062,N_30151,N_30009);
nor U31063 (N_31063,N_30620,N_30855);
and U31064 (N_31064,N_30277,N_30197);
nor U31065 (N_31065,N_30110,N_30044);
and U31066 (N_31066,N_30630,N_30106);
and U31067 (N_31067,N_30976,N_30637);
and U31068 (N_31068,N_30765,N_30600);
or U31069 (N_31069,N_30607,N_30852);
or U31070 (N_31070,N_30234,N_30582);
nor U31071 (N_31071,N_30768,N_30868);
and U31072 (N_31072,N_30233,N_30300);
and U31073 (N_31073,N_30107,N_30829);
xor U31074 (N_31074,N_30999,N_30318);
or U31075 (N_31075,N_30417,N_30832);
or U31076 (N_31076,N_30475,N_30891);
or U31077 (N_31077,N_30876,N_30821);
and U31078 (N_31078,N_30100,N_30345);
nor U31079 (N_31079,N_30559,N_30884);
nor U31080 (N_31080,N_30113,N_30680);
xnor U31081 (N_31081,N_30528,N_30762);
and U31082 (N_31082,N_30677,N_30720);
and U31083 (N_31083,N_30035,N_30076);
and U31084 (N_31084,N_30123,N_30575);
nor U31085 (N_31085,N_30268,N_30466);
and U31086 (N_31086,N_30850,N_30312);
nand U31087 (N_31087,N_30026,N_30885);
nand U31088 (N_31088,N_30483,N_30936);
and U31089 (N_31089,N_30840,N_30589);
nor U31090 (N_31090,N_30860,N_30703);
and U31091 (N_31091,N_30311,N_30003);
nand U31092 (N_31092,N_30937,N_30671);
nor U31093 (N_31093,N_30546,N_30799);
xor U31094 (N_31094,N_30695,N_30511);
or U31095 (N_31095,N_30681,N_30208);
nor U31096 (N_31096,N_30309,N_30889);
nand U31097 (N_31097,N_30906,N_30658);
nand U31098 (N_31098,N_30191,N_30733);
xor U31099 (N_31099,N_30396,N_30557);
or U31100 (N_31100,N_30931,N_30160);
and U31101 (N_31101,N_30204,N_30709);
nor U31102 (N_31102,N_30661,N_30486);
or U31103 (N_31103,N_30297,N_30863);
and U31104 (N_31104,N_30518,N_30669);
or U31105 (N_31105,N_30675,N_30826);
xnor U31106 (N_31106,N_30545,N_30017);
nand U31107 (N_31107,N_30663,N_30339);
nor U31108 (N_31108,N_30952,N_30064);
nand U31109 (N_31109,N_30562,N_30415);
nor U31110 (N_31110,N_30602,N_30049);
or U31111 (N_31111,N_30686,N_30955);
nor U31112 (N_31112,N_30817,N_30115);
or U31113 (N_31113,N_30376,N_30961);
and U31114 (N_31114,N_30453,N_30842);
or U31115 (N_31115,N_30556,N_30118);
nor U31116 (N_31116,N_30144,N_30445);
xnor U31117 (N_31117,N_30913,N_30971);
nor U31118 (N_31118,N_30834,N_30158);
and U31119 (N_31119,N_30778,N_30385);
nor U31120 (N_31120,N_30982,N_30427);
nor U31121 (N_31121,N_30298,N_30425);
or U31122 (N_31122,N_30611,N_30257);
nor U31123 (N_31123,N_30332,N_30809);
nand U31124 (N_31124,N_30075,N_30420);
xor U31125 (N_31125,N_30779,N_30223);
nand U31126 (N_31126,N_30294,N_30063);
xor U31127 (N_31127,N_30129,N_30469);
nor U31128 (N_31128,N_30405,N_30624);
or U31129 (N_31129,N_30621,N_30207);
nand U31130 (N_31130,N_30683,N_30735);
nor U31131 (N_31131,N_30154,N_30142);
and U31132 (N_31132,N_30638,N_30867);
xor U31133 (N_31133,N_30359,N_30992);
or U31134 (N_31134,N_30900,N_30749);
or U31135 (N_31135,N_30175,N_30640);
or U31136 (N_31136,N_30355,N_30526);
nor U31137 (N_31137,N_30969,N_30032);
and U31138 (N_31138,N_30149,N_30260);
nor U31139 (N_31139,N_30065,N_30929);
nand U31140 (N_31140,N_30979,N_30904);
xnor U31141 (N_31141,N_30171,N_30520);
xnor U31142 (N_31142,N_30679,N_30966);
nand U31143 (N_31143,N_30334,N_30738);
and U31144 (N_31144,N_30098,N_30962);
xnor U31145 (N_31145,N_30783,N_30150);
xnor U31146 (N_31146,N_30361,N_30153);
and U31147 (N_31147,N_30543,N_30323);
or U31148 (N_31148,N_30691,N_30281);
and U31149 (N_31149,N_30839,N_30465);
xor U31150 (N_31150,N_30083,N_30776);
nor U31151 (N_31151,N_30563,N_30019);
xnor U31152 (N_31152,N_30972,N_30786);
xor U31153 (N_31153,N_30653,N_30866);
and U31154 (N_31154,N_30259,N_30220);
and U31155 (N_31155,N_30287,N_30437);
nor U31156 (N_31156,N_30174,N_30434);
nor U31157 (N_31157,N_30721,N_30717);
nor U31158 (N_31158,N_30538,N_30435);
nand U31159 (N_31159,N_30849,N_30090);
nor U31160 (N_31160,N_30221,N_30641);
and U31161 (N_31161,N_30184,N_30773);
or U31162 (N_31162,N_30310,N_30124);
xor U31163 (N_31163,N_30784,N_30005);
and U31164 (N_31164,N_30292,N_30580);
nor U31165 (N_31165,N_30070,N_30188);
or U31166 (N_31166,N_30632,N_30833);
nor U31167 (N_31167,N_30490,N_30140);
and U31168 (N_31168,N_30099,N_30045);
xnor U31169 (N_31169,N_30284,N_30957);
and U31170 (N_31170,N_30102,N_30760);
xnor U31171 (N_31171,N_30209,N_30499);
and U31172 (N_31172,N_30054,N_30590);
xnor U31173 (N_31173,N_30432,N_30302);
or U31174 (N_31174,N_30723,N_30710);
nand U31175 (N_31175,N_30892,N_30431);
or U31176 (N_31176,N_30715,N_30880);
nand U31177 (N_31177,N_30649,N_30414);
and U31178 (N_31178,N_30103,N_30455);
xor U31179 (N_31179,N_30605,N_30594);
nand U31180 (N_31180,N_30496,N_30306);
xnor U31181 (N_31181,N_30497,N_30513);
xnor U31182 (N_31182,N_30491,N_30023);
nor U31183 (N_31183,N_30947,N_30672);
nand U31184 (N_31184,N_30056,N_30128);
and U31185 (N_31185,N_30617,N_30271);
nand U31186 (N_31186,N_30010,N_30213);
nand U31187 (N_31187,N_30895,N_30835);
or U31188 (N_31188,N_30507,N_30327);
and U31189 (N_31189,N_30322,N_30958);
xor U31190 (N_31190,N_30047,N_30544);
nor U31191 (N_31191,N_30745,N_30980);
nor U31192 (N_31192,N_30069,N_30456);
xor U31193 (N_31193,N_30888,N_30305);
nand U31194 (N_31194,N_30934,N_30942);
or U31195 (N_31195,N_30403,N_30091);
xor U31196 (N_31196,N_30567,N_30192);
and U31197 (N_31197,N_30481,N_30584);
and U31198 (N_31198,N_30383,N_30674);
and U31199 (N_31199,N_30771,N_30943);
nand U31200 (N_31200,N_30350,N_30579);
xnor U31201 (N_31201,N_30748,N_30214);
nor U31202 (N_31202,N_30378,N_30231);
xnor U31203 (N_31203,N_30249,N_30235);
xor U31204 (N_31204,N_30813,N_30039);
and U31205 (N_31205,N_30907,N_30304);
nor U31206 (N_31206,N_30785,N_30788);
or U31207 (N_31207,N_30635,N_30727);
or U31208 (N_31208,N_30731,N_30462);
nand U31209 (N_31209,N_30874,N_30363);
nand U31210 (N_31210,N_30858,N_30360);
or U31211 (N_31211,N_30276,N_30280);
and U31212 (N_31212,N_30804,N_30066);
nor U31213 (N_31213,N_30470,N_30984);
nand U31214 (N_31214,N_30753,N_30903);
xnor U31215 (N_31215,N_30911,N_30650);
nor U31216 (N_31216,N_30657,N_30407);
or U31217 (N_31217,N_30111,N_30705);
nand U31218 (N_31218,N_30780,N_30012);
nand U31219 (N_31219,N_30542,N_30485);
or U31220 (N_31220,N_30052,N_30033);
or U31221 (N_31221,N_30143,N_30022);
xor U31222 (N_31222,N_30133,N_30071);
nor U31223 (N_31223,N_30801,N_30206);
nand U31224 (N_31224,N_30229,N_30324);
nor U31225 (N_31225,N_30744,N_30458);
nand U31226 (N_31226,N_30505,N_30761);
and U31227 (N_31227,N_30264,N_30881);
xor U31228 (N_31228,N_30851,N_30319);
nor U31229 (N_31229,N_30732,N_30147);
and U31230 (N_31230,N_30541,N_30132);
xnor U31231 (N_31231,N_30061,N_30746);
xor U31232 (N_31232,N_30928,N_30391);
nand U31233 (N_31233,N_30262,N_30401);
or U31234 (N_31234,N_30419,N_30564);
or U31235 (N_31235,N_30062,N_30410);
xnor U31236 (N_31236,N_30772,N_30949);
or U31237 (N_31237,N_30433,N_30986);
or U31238 (N_31238,N_30509,N_30095);
and U31239 (N_31239,N_30702,N_30228);
nor U31240 (N_31240,N_30493,N_30181);
nor U31241 (N_31241,N_30163,N_30665);
or U31242 (N_31242,N_30423,N_30578);
and U31243 (N_31243,N_30792,N_30708);
or U31244 (N_31244,N_30660,N_30814);
xor U31245 (N_31245,N_30112,N_30517);
or U31246 (N_31246,N_30856,N_30591);
or U31247 (N_31247,N_30688,N_30604);
xnor U31248 (N_31248,N_30468,N_30240);
xnor U31249 (N_31249,N_30755,N_30379);
or U31250 (N_31250,N_30596,N_30524);
xor U31251 (N_31251,N_30395,N_30975);
xnor U31252 (N_31252,N_30386,N_30384);
nor U31253 (N_31253,N_30289,N_30222);
nand U31254 (N_31254,N_30381,N_30758);
or U31255 (N_31255,N_30629,N_30647);
and U31256 (N_31256,N_30838,N_30910);
nor U31257 (N_31257,N_30241,N_30137);
nor U31258 (N_31258,N_30377,N_30750);
or U31259 (N_31259,N_30861,N_30178);
nor U31260 (N_31260,N_30689,N_30549);
or U31261 (N_31261,N_30534,N_30085);
nor U31262 (N_31262,N_30766,N_30057);
or U31263 (N_31263,N_30759,N_30418);
nor U31264 (N_31264,N_30368,N_30014);
nor U31265 (N_31265,N_30996,N_30016);
xor U31266 (N_31266,N_30279,N_30612);
or U31267 (N_31267,N_30642,N_30742);
nor U31268 (N_31268,N_30210,N_30527);
nor U31269 (N_31269,N_30333,N_30897);
nor U31270 (N_31270,N_30648,N_30185);
nor U31271 (N_31271,N_30547,N_30096);
nor U31272 (N_31272,N_30963,N_30476);
xnor U31273 (N_31273,N_30998,N_30916);
xor U31274 (N_31274,N_30119,N_30021);
or U31275 (N_31275,N_30243,N_30537);
and U31276 (N_31276,N_30654,N_30440);
nor U31277 (N_31277,N_30751,N_30552);
nand U31278 (N_31278,N_30295,N_30242);
xnor U31279 (N_31279,N_30330,N_30757);
and U31280 (N_31280,N_30905,N_30443);
or U31281 (N_31281,N_30893,N_30436);
or U31282 (N_31282,N_30274,N_30389);
xor U31283 (N_31283,N_30625,N_30121);
nor U31284 (N_31284,N_30195,N_30299);
nand U31285 (N_31285,N_30519,N_30970);
or U31286 (N_31286,N_30424,N_30040);
xnor U31287 (N_31287,N_30168,N_30215);
nor U31288 (N_31288,N_30180,N_30571);
nand U31289 (N_31289,N_30225,N_30734);
or U31290 (N_31290,N_30588,N_30633);
nand U31291 (N_31291,N_30079,N_30566);
and U31292 (N_31292,N_30442,N_30533);
or U31293 (N_31293,N_30741,N_30203);
and U31294 (N_31294,N_30046,N_30523);
and U31295 (N_31295,N_30560,N_30756);
or U31296 (N_31296,N_30474,N_30967);
nand U31297 (N_31297,N_30795,N_30120);
or U31298 (N_31298,N_30628,N_30166);
or U31299 (N_31299,N_30530,N_30877);
and U31300 (N_31300,N_30053,N_30639);
nand U31301 (N_31301,N_30670,N_30067);
nand U31302 (N_31302,N_30230,N_30349);
and U31303 (N_31303,N_30673,N_30244);
xnor U31304 (N_31304,N_30011,N_30328);
xor U31305 (N_31305,N_30901,N_30921);
and U31306 (N_31306,N_30636,N_30161);
nor U31307 (N_31307,N_30266,N_30170);
or U31308 (N_31308,N_30946,N_30351);
xor U31309 (N_31309,N_30413,N_30058);
and U31310 (N_31310,N_30608,N_30232);
or U31311 (N_31311,N_30555,N_30995);
and U31312 (N_31312,N_30652,N_30815);
nor U31313 (N_31313,N_30592,N_30878);
xor U31314 (N_31314,N_30348,N_30767);
nand U31315 (N_31315,N_30344,N_30770);
nor U31316 (N_31316,N_30347,N_30270);
and U31317 (N_31317,N_30890,N_30836);
or U31318 (N_31318,N_30645,N_30598);
xnor U31319 (N_31319,N_30960,N_30793);
nand U31320 (N_31320,N_30912,N_30918);
xor U31321 (N_31321,N_30250,N_30183);
or U31322 (N_31322,N_30714,N_30358);
nand U31323 (N_31323,N_30082,N_30807);
and U31324 (N_31324,N_30138,N_30774);
and U31325 (N_31325,N_30135,N_30293);
and U31326 (N_31326,N_30428,N_30101);
or U31327 (N_31327,N_30626,N_30382);
or U31328 (N_31328,N_30932,N_30190);
xor U31329 (N_31329,N_30997,N_30296);
xor U31330 (N_31330,N_30189,N_30968);
or U31331 (N_31331,N_30460,N_30782);
nor U31332 (N_31332,N_30114,N_30978);
nor U31333 (N_31333,N_30864,N_30366);
xor U31334 (N_31334,N_30337,N_30531);
and U31335 (N_31335,N_30343,N_30558);
or U31336 (N_31336,N_30253,N_30777);
and U31337 (N_31337,N_30577,N_30217);
and U31338 (N_31338,N_30325,N_30726);
nor U31339 (N_31339,N_30167,N_30790);
or U31340 (N_31340,N_30059,N_30164);
and U31341 (N_31341,N_30627,N_30973);
nand U31342 (N_31342,N_30983,N_30902);
and U31343 (N_31343,N_30216,N_30707);
nand U31344 (N_31344,N_30145,N_30736);
or U31345 (N_31345,N_30682,N_30352);
and U31346 (N_31346,N_30646,N_30015);
nor U31347 (N_31347,N_30941,N_30944);
nor U31348 (N_31348,N_30853,N_30915);
and U31349 (N_31349,N_30369,N_30152);
xor U31350 (N_31350,N_30535,N_30198);
xnor U31351 (N_31351,N_30029,N_30643);
nand U31352 (N_31352,N_30514,N_30825);
nor U31353 (N_31353,N_30724,N_30283);
xor U31354 (N_31354,N_30201,N_30326);
or U31355 (N_31355,N_30806,N_30737);
or U31356 (N_31356,N_30684,N_30042);
nor U31357 (N_31357,N_30678,N_30991);
nand U31358 (N_31358,N_30854,N_30848);
nand U31359 (N_31359,N_30357,N_30716);
nor U31360 (N_31360,N_30291,N_30730);
xnor U31361 (N_31361,N_30887,N_30857);
nand U31362 (N_31362,N_30252,N_30974);
or U31363 (N_31363,N_30822,N_30051);
xnor U31364 (N_31364,N_30038,N_30879);
or U31365 (N_31365,N_30037,N_30964);
nand U31366 (N_31366,N_30173,N_30800);
nor U31367 (N_31367,N_30587,N_30787);
xnor U31368 (N_31368,N_30585,N_30859);
nor U31369 (N_31369,N_30084,N_30211);
nand U31370 (N_31370,N_30953,N_30692);
nor U31371 (N_31371,N_30894,N_30698);
and U31372 (N_31372,N_30553,N_30406);
xnor U31373 (N_31373,N_30595,N_30018);
nand U31374 (N_31374,N_30471,N_30338);
nand U31375 (N_31375,N_30080,N_30157);
and U31376 (N_31376,N_30796,N_30439);
nand U31377 (N_31377,N_30551,N_30446);
nand U31378 (N_31378,N_30186,N_30548);
nand U31379 (N_31379,N_30116,N_30454);
or U31380 (N_31380,N_30200,N_30263);
and U31381 (N_31381,N_30089,N_30506);
xor U31382 (N_31382,N_30797,N_30572);
nor U31383 (N_31383,N_30808,N_30581);
xnor U31384 (N_31384,N_30896,N_30830);
or U31385 (N_31385,N_30254,N_30093);
nand U31386 (N_31386,N_30314,N_30993);
or U31387 (N_31387,N_30586,N_30387);
or U31388 (N_31388,N_30482,N_30108);
nand U31389 (N_31389,N_30162,N_30837);
nor U31390 (N_31390,N_30372,N_30024);
xor U31391 (N_31391,N_30286,N_30288);
xnor U31392 (N_31392,N_30875,N_30141);
or U31393 (N_31393,N_30030,N_30364);
or U31394 (N_31394,N_30989,N_30273);
or U31395 (N_31395,N_30452,N_30290);
or U31396 (N_31396,N_30341,N_30873);
xnor U31397 (N_31397,N_30810,N_30712);
xnor U31398 (N_31398,N_30843,N_30644);
nor U31399 (N_31399,N_30094,N_30267);
or U31400 (N_31400,N_30134,N_30438);
xor U31401 (N_31401,N_30367,N_30373);
nor U31402 (N_31402,N_30489,N_30948);
and U31403 (N_31403,N_30238,N_30097);
nand U31404 (N_31404,N_30336,N_30146);
or U31405 (N_31405,N_30515,N_30034);
nor U31406 (N_31406,N_30508,N_30711);
nor U31407 (N_31407,N_30307,N_30930);
xor U31408 (N_31408,N_30073,N_30394);
xnor U31409 (N_31409,N_30927,N_30275);
nand U31410 (N_31410,N_30573,N_30457);
and U31411 (N_31411,N_30127,N_30177);
or U31412 (N_31412,N_30869,N_30951);
nand U31413 (N_31413,N_30994,N_30704);
nand U31414 (N_31414,N_30408,N_30959);
and U31415 (N_31415,N_30603,N_30001);
nand U31416 (N_31416,N_30008,N_30002);
or U31417 (N_31417,N_30340,N_30444);
xor U31418 (N_31418,N_30402,N_30502);
nor U31419 (N_31419,N_30072,N_30522);
and U31420 (N_31420,N_30725,N_30812);
xnor U31421 (N_31421,N_30285,N_30713);
nand U31422 (N_31422,N_30028,N_30988);
nand U31423 (N_31423,N_30449,N_30871);
or U31424 (N_31424,N_30618,N_30122);
or U31425 (N_31425,N_30495,N_30265);
or U31426 (N_31426,N_30775,N_30823);
or U31427 (N_31427,N_30409,N_30461);
or U31428 (N_31428,N_30939,N_30882);
and U31429 (N_31429,N_30321,N_30909);
nand U31430 (N_31430,N_30050,N_30729);
nand U31431 (N_31431,N_30272,N_30631);
xnor U31432 (N_31432,N_30077,N_30020);
or U31433 (N_31433,N_30346,N_30668);
xnor U31434 (N_31434,N_30987,N_30159);
xnor U31435 (N_31435,N_30819,N_30718);
nor U31436 (N_31436,N_30802,N_30139);
nand U31437 (N_31437,N_30539,N_30536);
or U31438 (N_31438,N_30763,N_30278);
or U31439 (N_31439,N_30068,N_30430);
xor U31440 (N_31440,N_30212,N_30883);
xnor U31441 (N_31441,N_30193,N_30954);
or U31442 (N_31442,N_30694,N_30256);
xnor U31443 (N_31443,N_30831,N_30990);
nor U31444 (N_31444,N_30404,N_30512);
or U31445 (N_31445,N_30935,N_30769);
or U31446 (N_31446,N_30187,N_30478);
xor U31447 (N_31447,N_30269,N_30747);
and U31448 (N_31448,N_30397,N_30798);
and U31449 (N_31449,N_30226,N_30081);
or U31450 (N_31450,N_30862,N_30687);
xnor U31451 (N_31451,N_30477,N_30504);
and U31452 (N_31452,N_30342,N_30706);
nor U31453 (N_31453,N_30791,N_30087);
xnor U31454 (N_31454,N_30301,N_30664);
xor U31455 (N_31455,N_30693,N_30303);
xnor U31456 (N_31456,N_30666,N_30104);
nand U31457 (N_31457,N_30459,N_30060);
or U31458 (N_31458,N_30933,N_30450);
xnor U31459 (N_31459,N_30754,N_30048);
or U31460 (N_31460,N_30917,N_30036);
xnor U31461 (N_31461,N_30841,N_30623);
nand U31462 (N_31462,N_30172,N_30335);
nor U31463 (N_31463,N_30155,N_30525);
or U31464 (N_31464,N_30441,N_30422);
xor U31465 (N_31465,N_30131,N_30574);
and U31466 (N_31466,N_30924,N_30820);
or U31467 (N_31467,N_30086,N_30473);
or U31468 (N_31468,N_30258,N_30421);
and U31469 (N_31469,N_30794,N_30371);
or U31470 (N_31470,N_30399,N_30148);
and U31471 (N_31471,N_30055,N_30846);
nand U31472 (N_31472,N_30027,N_30472);
nand U31473 (N_31473,N_30847,N_30043);
nand U31474 (N_31474,N_30510,N_30606);
and U31475 (N_31475,N_30923,N_30247);
nand U31476 (N_31476,N_30041,N_30965);
or U31477 (N_31477,N_30356,N_30655);
xnor U31478 (N_31478,N_30503,N_30136);
nand U31479 (N_31479,N_30925,N_30125);
or U31480 (N_31480,N_30205,N_30601);
nand U31481 (N_31481,N_30740,N_30025);
nand U31482 (N_31482,N_30659,N_30261);
nor U31483 (N_31483,N_30700,N_30484);
nand U31484 (N_31484,N_30690,N_30610);
nand U31485 (N_31485,N_30492,N_30789);
xor U31486 (N_31486,N_30701,N_30568);
or U31487 (N_31487,N_30400,N_30007);
xnor U31488 (N_31488,N_30752,N_30844);
nand U31489 (N_31489,N_30464,N_30781);
and U31490 (N_31490,N_30920,N_30169);
and U31491 (N_31491,N_30320,N_30365);
or U31492 (N_31492,N_30074,N_30561);
or U31493 (N_31493,N_30656,N_30500);
or U31494 (N_31494,N_30006,N_30199);
nor U31495 (N_31495,N_30411,N_30739);
and U31496 (N_31496,N_30194,N_30899);
or U31497 (N_31497,N_30004,N_30722);
or U31498 (N_31498,N_30487,N_30922);
nor U31499 (N_31499,N_30308,N_30634);
and U31500 (N_31500,N_30368,N_30580);
xnor U31501 (N_31501,N_30234,N_30938);
and U31502 (N_31502,N_30261,N_30159);
xnor U31503 (N_31503,N_30669,N_30729);
nor U31504 (N_31504,N_30436,N_30330);
and U31505 (N_31505,N_30920,N_30749);
nor U31506 (N_31506,N_30716,N_30360);
nor U31507 (N_31507,N_30702,N_30977);
or U31508 (N_31508,N_30667,N_30594);
nor U31509 (N_31509,N_30110,N_30922);
nor U31510 (N_31510,N_30470,N_30983);
nor U31511 (N_31511,N_30235,N_30078);
nand U31512 (N_31512,N_30196,N_30522);
and U31513 (N_31513,N_30134,N_30351);
or U31514 (N_31514,N_30645,N_30422);
nor U31515 (N_31515,N_30866,N_30617);
xnor U31516 (N_31516,N_30242,N_30315);
or U31517 (N_31517,N_30422,N_30444);
xor U31518 (N_31518,N_30419,N_30524);
or U31519 (N_31519,N_30441,N_30148);
nand U31520 (N_31520,N_30317,N_30328);
and U31521 (N_31521,N_30682,N_30884);
nor U31522 (N_31522,N_30571,N_30592);
xor U31523 (N_31523,N_30377,N_30230);
and U31524 (N_31524,N_30106,N_30964);
xor U31525 (N_31525,N_30199,N_30291);
xnor U31526 (N_31526,N_30924,N_30054);
nor U31527 (N_31527,N_30458,N_30123);
xnor U31528 (N_31528,N_30728,N_30874);
and U31529 (N_31529,N_30236,N_30506);
nand U31530 (N_31530,N_30653,N_30417);
nor U31531 (N_31531,N_30947,N_30466);
nand U31532 (N_31532,N_30584,N_30553);
nand U31533 (N_31533,N_30973,N_30561);
xnor U31534 (N_31534,N_30539,N_30413);
and U31535 (N_31535,N_30648,N_30562);
nor U31536 (N_31536,N_30916,N_30011);
or U31537 (N_31537,N_30485,N_30673);
nand U31538 (N_31538,N_30532,N_30156);
or U31539 (N_31539,N_30324,N_30802);
or U31540 (N_31540,N_30884,N_30025);
and U31541 (N_31541,N_30467,N_30289);
nor U31542 (N_31542,N_30191,N_30549);
or U31543 (N_31543,N_30744,N_30552);
xnor U31544 (N_31544,N_30597,N_30136);
and U31545 (N_31545,N_30851,N_30842);
or U31546 (N_31546,N_30432,N_30940);
or U31547 (N_31547,N_30807,N_30869);
or U31548 (N_31548,N_30255,N_30880);
nor U31549 (N_31549,N_30944,N_30934);
nor U31550 (N_31550,N_30073,N_30100);
nand U31551 (N_31551,N_30799,N_30388);
or U31552 (N_31552,N_30232,N_30854);
or U31553 (N_31553,N_30512,N_30013);
nor U31554 (N_31554,N_30798,N_30364);
nor U31555 (N_31555,N_30594,N_30051);
xor U31556 (N_31556,N_30939,N_30339);
nand U31557 (N_31557,N_30944,N_30412);
or U31558 (N_31558,N_30793,N_30843);
or U31559 (N_31559,N_30495,N_30021);
and U31560 (N_31560,N_30291,N_30153);
and U31561 (N_31561,N_30420,N_30558);
nor U31562 (N_31562,N_30003,N_30805);
and U31563 (N_31563,N_30464,N_30140);
or U31564 (N_31564,N_30278,N_30513);
or U31565 (N_31565,N_30613,N_30526);
nand U31566 (N_31566,N_30280,N_30438);
nor U31567 (N_31567,N_30504,N_30869);
xor U31568 (N_31568,N_30714,N_30481);
xnor U31569 (N_31569,N_30813,N_30485);
nor U31570 (N_31570,N_30083,N_30922);
or U31571 (N_31571,N_30463,N_30565);
xnor U31572 (N_31572,N_30786,N_30370);
nor U31573 (N_31573,N_30544,N_30188);
xor U31574 (N_31574,N_30903,N_30702);
nor U31575 (N_31575,N_30220,N_30864);
or U31576 (N_31576,N_30094,N_30527);
or U31577 (N_31577,N_30497,N_30334);
nor U31578 (N_31578,N_30388,N_30789);
and U31579 (N_31579,N_30698,N_30833);
nand U31580 (N_31580,N_30068,N_30538);
and U31581 (N_31581,N_30367,N_30362);
or U31582 (N_31582,N_30392,N_30760);
nor U31583 (N_31583,N_30503,N_30740);
and U31584 (N_31584,N_30068,N_30977);
and U31585 (N_31585,N_30146,N_30053);
nand U31586 (N_31586,N_30703,N_30434);
nor U31587 (N_31587,N_30454,N_30113);
nor U31588 (N_31588,N_30078,N_30167);
nand U31589 (N_31589,N_30365,N_30108);
xor U31590 (N_31590,N_30471,N_30609);
nor U31591 (N_31591,N_30302,N_30318);
xor U31592 (N_31592,N_30077,N_30846);
xnor U31593 (N_31593,N_30518,N_30100);
xnor U31594 (N_31594,N_30184,N_30916);
or U31595 (N_31595,N_30591,N_30217);
nand U31596 (N_31596,N_30614,N_30195);
or U31597 (N_31597,N_30584,N_30430);
nand U31598 (N_31598,N_30342,N_30851);
nor U31599 (N_31599,N_30861,N_30846);
nand U31600 (N_31600,N_30502,N_30037);
or U31601 (N_31601,N_30848,N_30549);
nor U31602 (N_31602,N_30495,N_30504);
nor U31603 (N_31603,N_30095,N_30126);
xor U31604 (N_31604,N_30221,N_30750);
or U31605 (N_31605,N_30254,N_30097);
nor U31606 (N_31606,N_30942,N_30494);
nor U31607 (N_31607,N_30567,N_30782);
xor U31608 (N_31608,N_30846,N_30373);
and U31609 (N_31609,N_30945,N_30143);
nor U31610 (N_31610,N_30811,N_30266);
or U31611 (N_31611,N_30139,N_30996);
and U31612 (N_31612,N_30131,N_30135);
nand U31613 (N_31613,N_30765,N_30206);
nand U31614 (N_31614,N_30900,N_30184);
nand U31615 (N_31615,N_30165,N_30597);
xnor U31616 (N_31616,N_30059,N_30721);
xor U31617 (N_31617,N_30158,N_30770);
nor U31618 (N_31618,N_30795,N_30755);
or U31619 (N_31619,N_30617,N_30413);
xnor U31620 (N_31620,N_30026,N_30568);
or U31621 (N_31621,N_30002,N_30479);
and U31622 (N_31622,N_30040,N_30521);
xnor U31623 (N_31623,N_30499,N_30084);
and U31624 (N_31624,N_30686,N_30508);
nor U31625 (N_31625,N_30824,N_30660);
nand U31626 (N_31626,N_30103,N_30936);
or U31627 (N_31627,N_30346,N_30953);
nor U31628 (N_31628,N_30279,N_30540);
nor U31629 (N_31629,N_30839,N_30666);
nor U31630 (N_31630,N_30207,N_30529);
or U31631 (N_31631,N_30019,N_30403);
nand U31632 (N_31632,N_30019,N_30789);
nand U31633 (N_31633,N_30913,N_30321);
or U31634 (N_31634,N_30806,N_30964);
xnor U31635 (N_31635,N_30946,N_30978);
or U31636 (N_31636,N_30887,N_30645);
nor U31637 (N_31637,N_30295,N_30855);
nor U31638 (N_31638,N_30489,N_30203);
nor U31639 (N_31639,N_30812,N_30621);
xnor U31640 (N_31640,N_30859,N_30474);
nand U31641 (N_31641,N_30489,N_30276);
or U31642 (N_31642,N_30928,N_30725);
nor U31643 (N_31643,N_30754,N_30322);
and U31644 (N_31644,N_30506,N_30782);
or U31645 (N_31645,N_30089,N_30031);
nor U31646 (N_31646,N_30507,N_30512);
nor U31647 (N_31647,N_30258,N_30559);
xnor U31648 (N_31648,N_30210,N_30362);
or U31649 (N_31649,N_30825,N_30000);
and U31650 (N_31650,N_30444,N_30907);
nand U31651 (N_31651,N_30125,N_30892);
or U31652 (N_31652,N_30181,N_30324);
nor U31653 (N_31653,N_30673,N_30460);
or U31654 (N_31654,N_30025,N_30519);
xnor U31655 (N_31655,N_30526,N_30192);
nand U31656 (N_31656,N_30293,N_30022);
nor U31657 (N_31657,N_30117,N_30183);
xor U31658 (N_31658,N_30722,N_30855);
nand U31659 (N_31659,N_30853,N_30845);
xor U31660 (N_31660,N_30906,N_30005);
nand U31661 (N_31661,N_30633,N_30216);
xnor U31662 (N_31662,N_30837,N_30801);
nor U31663 (N_31663,N_30939,N_30160);
nand U31664 (N_31664,N_30867,N_30620);
nor U31665 (N_31665,N_30005,N_30723);
and U31666 (N_31666,N_30546,N_30653);
or U31667 (N_31667,N_30865,N_30534);
or U31668 (N_31668,N_30325,N_30412);
xnor U31669 (N_31669,N_30804,N_30241);
xnor U31670 (N_31670,N_30935,N_30399);
nand U31671 (N_31671,N_30305,N_30135);
and U31672 (N_31672,N_30192,N_30267);
nand U31673 (N_31673,N_30225,N_30582);
and U31674 (N_31674,N_30800,N_30407);
and U31675 (N_31675,N_30787,N_30260);
nand U31676 (N_31676,N_30834,N_30000);
and U31677 (N_31677,N_30657,N_30628);
or U31678 (N_31678,N_30194,N_30087);
nor U31679 (N_31679,N_30088,N_30179);
xor U31680 (N_31680,N_30155,N_30173);
nand U31681 (N_31681,N_30887,N_30509);
nor U31682 (N_31682,N_30416,N_30975);
and U31683 (N_31683,N_30216,N_30945);
xor U31684 (N_31684,N_30236,N_30203);
or U31685 (N_31685,N_30339,N_30392);
and U31686 (N_31686,N_30277,N_30097);
nand U31687 (N_31687,N_30987,N_30477);
xor U31688 (N_31688,N_30553,N_30291);
and U31689 (N_31689,N_30734,N_30883);
xor U31690 (N_31690,N_30603,N_30837);
and U31691 (N_31691,N_30032,N_30737);
and U31692 (N_31692,N_30151,N_30673);
or U31693 (N_31693,N_30460,N_30848);
xor U31694 (N_31694,N_30875,N_30712);
xnor U31695 (N_31695,N_30014,N_30029);
and U31696 (N_31696,N_30183,N_30047);
and U31697 (N_31697,N_30780,N_30598);
and U31698 (N_31698,N_30561,N_30049);
xnor U31699 (N_31699,N_30270,N_30715);
nand U31700 (N_31700,N_30544,N_30225);
or U31701 (N_31701,N_30392,N_30074);
and U31702 (N_31702,N_30678,N_30523);
xnor U31703 (N_31703,N_30186,N_30347);
nand U31704 (N_31704,N_30445,N_30616);
and U31705 (N_31705,N_30505,N_30515);
and U31706 (N_31706,N_30965,N_30172);
or U31707 (N_31707,N_30337,N_30142);
and U31708 (N_31708,N_30867,N_30930);
nand U31709 (N_31709,N_30121,N_30349);
nor U31710 (N_31710,N_30187,N_30367);
nand U31711 (N_31711,N_30508,N_30154);
nand U31712 (N_31712,N_30407,N_30372);
xor U31713 (N_31713,N_30208,N_30192);
or U31714 (N_31714,N_30326,N_30174);
xor U31715 (N_31715,N_30698,N_30766);
or U31716 (N_31716,N_30371,N_30402);
nor U31717 (N_31717,N_30033,N_30926);
xnor U31718 (N_31718,N_30132,N_30452);
nor U31719 (N_31719,N_30854,N_30820);
xnor U31720 (N_31720,N_30104,N_30405);
nand U31721 (N_31721,N_30057,N_30054);
xor U31722 (N_31722,N_30952,N_30630);
nand U31723 (N_31723,N_30853,N_30033);
and U31724 (N_31724,N_30130,N_30705);
and U31725 (N_31725,N_30605,N_30651);
and U31726 (N_31726,N_30830,N_30753);
xnor U31727 (N_31727,N_30630,N_30282);
xor U31728 (N_31728,N_30467,N_30458);
xor U31729 (N_31729,N_30600,N_30429);
nor U31730 (N_31730,N_30911,N_30439);
nand U31731 (N_31731,N_30073,N_30108);
and U31732 (N_31732,N_30176,N_30141);
nor U31733 (N_31733,N_30610,N_30966);
and U31734 (N_31734,N_30059,N_30397);
nor U31735 (N_31735,N_30008,N_30554);
xnor U31736 (N_31736,N_30212,N_30116);
xor U31737 (N_31737,N_30955,N_30131);
xnor U31738 (N_31738,N_30622,N_30903);
xnor U31739 (N_31739,N_30879,N_30911);
or U31740 (N_31740,N_30380,N_30672);
and U31741 (N_31741,N_30945,N_30544);
xor U31742 (N_31742,N_30779,N_30257);
nor U31743 (N_31743,N_30951,N_30492);
nor U31744 (N_31744,N_30870,N_30617);
xnor U31745 (N_31745,N_30252,N_30255);
nand U31746 (N_31746,N_30018,N_30824);
or U31747 (N_31747,N_30285,N_30907);
nor U31748 (N_31748,N_30573,N_30529);
nor U31749 (N_31749,N_30793,N_30508);
or U31750 (N_31750,N_30814,N_30413);
xnor U31751 (N_31751,N_30815,N_30256);
nor U31752 (N_31752,N_30399,N_30120);
nand U31753 (N_31753,N_30087,N_30085);
or U31754 (N_31754,N_30237,N_30996);
nor U31755 (N_31755,N_30490,N_30537);
nor U31756 (N_31756,N_30314,N_30770);
and U31757 (N_31757,N_30291,N_30126);
nor U31758 (N_31758,N_30617,N_30616);
or U31759 (N_31759,N_30692,N_30939);
nor U31760 (N_31760,N_30740,N_30012);
xor U31761 (N_31761,N_30101,N_30872);
or U31762 (N_31762,N_30720,N_30243);
nor U31763 (N_31763,N_30863,N_30372);
and U31764 (N_31764,N_30801,N_30487);
or U31765 (N_31765,N_30803,N_30191);
or U31766 (N_31766,N_30547,N_30891);
and U31767 (N_31767,N_30924,N_30650);
nor U31768 (N_31768,N_30027,N_30299);
nor U31769 (N_31769,N_30623,N_30982);
xor U31770 (N_31770,N_30067,N_30429);
or U31771 (N_31771,N_30982,N_30576);
xnor U31772 (N_31772,N_30323,N_30405);
or U31773 (N_31773,N_30540,N_30281);
nor U31774 (N_31774,N_30888,N_30894);
and U31775 (N_31775,N_30888,N_30495);
nor U31776 (N_31776,N_30270,N_30820);
nor U31777 (N_31777,N_30687,N_30031);
nand U31778 (N_31778,N_30369,N_30093);
nand U31779 (N_31779,N_30435,N_30348);
or U31780 (N_31780,N_30859,N_30084);
nand U31781 (N_31781,N_30120,N_30291);
or U31782 (N_31782,N_30919,N_30668);
or U31783 (N_31783,N_30199,N_30727);
nor U31784 (N_31784,N_30216,N_30593);
or U31785 (N_31785,N_30139,N_30462);
and U31786 (N_31786,N_30358,N_30373);
nor U31787 (N_31787,N_30162,N_30226);
and U31788 (N_31788,N_30376,N_30636);
or U31789 (N_31789,N_30124,N_30216);
xor U31790 (N_31790,N_30535,N_30846);
nand U31791 (N_31791,N_30511,N_30909);
nand U31792 (N_31792,N_30116,N_30774);
or U31793 (N_31793,N_30669,N_30307);
or U31794 (N_31794,N_30273,N_30025);
and U31795 (N_31795,N_30814,N_30437);
or U31796 (N_31796,N_30057,N_30168);
nor U31797 (N_31797,N_30776,N_30298);
nor U31798 (N_31798,N_30690,N_30146);
or U31799 (N_31799,N_30321,N_30080);
nand U31800 (N_31800,N_30121,N_30482);
and U31801 (N_31801,N_30277,N_30419);
and U31802 (N_31802,N_30225,N_30547);
nand U31803 (N_31803,N_30309,N_30835);
and U31804 (N_31804,N_30119,N_30063);
and U31805 (N_31805,N_30808,N_30150);
xnor U31806 (N_31806,N_30050,N_30516);
or U31807 (N_31807,N_30062,N_30476);
xnor U31808 (N_31808,N_30227,N_30792);
nor U31809 (N_31809,N_30400,N_30344);
nand U31810 (N_31810,N_30076,N_30819);
xor U31811 (N_31811,N_30777,N_30594);
and U31812 (N_31812,N_30458,N_30616);
and U31813 (N_31813,N_30512,N_30901);
nor U31814 (N_31814,N_30184,N_30458);
nor U31815 (N_31815,N_30423,N_30249);
xnor U31816 (N_31816,N_30711,N_30618);
or U31817 (N_31817,N_30184,N_30451);
nor U31818 (N_31818,N_30910,N_30263);
xor U31819 (N_31819,N_30925,N_30055);
and U31820 (N_31820,N_30926,N_30823);
and U31821 (N_31821,N_30554,N_30066);
and U31822 (N_31822,N_30267,N_30954);
or U31823 (N_31823,N_30119,N_30023);
nor U31824 (N_31824,N_30829,N_30195);
xnor U31825 (N_31825,N_30807,N_30286);
xnor U31826 (N_31826,N_30284,N_30596);
or U31827 (N_31827,N_30448,N_30194);
or U31828 (N_31828,N_30949,N_30613);
nor U31829 (N_31829,N_30949,N_30945);
or U31830 (N_31830,N_30908,N_30393);
and U31831 (N_31831,N_30950,N_30490);
nor U31832 (N_31832,N_30706,N_30200);
or U31833 (N_31833,N_30884,N_30243);
or U31834 (N_31834,N_30297,N_30381);
nor U31835 (N_31835,N_30761,N_30399);
nand U31836 (N_31836,N_30836,N_30444);
or U31837 (N_31837,N_30083,N_30021);
or U31838 (N_31838,N_30985,N_30522);
nand U31839 (N_31839,N_30461,N_30787);
nand U31840 (N_31840,N_30844,N_30308);
nor U31841 (N_31841,N_30061,N_30976);
xnor U31842 (N_31842,N_30598,N_30431);
nor U31843 (N_31843,N_30716,N_30959);
nor U31844 (N_31844,N_30205,N_30866);
nor U31845 (N_31845,N_30932,N_30688);
or U31846 (N_31846,N_30479,N_30065);
nand U31847 (N_31847,N_30147,N_30740);
and U31848 (N_31848,N_30064,N_30447);
or U31849 (N_31849,N_30800,N_30824);
xnor U31850 (N_31850,N_30995,N_30998);
nor U31851 (N_31851,N_30752,N_30450);
nor U31852 (N_31852,N_30792,N_30768);
nand U31853 (N_31853,N_30598,N_30050);
or U31854 (N_31854,N_30311,N_30114);
nand U31855 (N_31855,N_30932,N_30097);
or U31856 (N_31856,N_30863,N_30238);
or U31857 (N_31857,N_30277,N_30266);
nor U31858 (N_31858,N_30477,N_30760);
or U31859 (N_31859,N_30971,N_30369);
or U31860 (N_31860,N_30312,N_30521);
nor U31861 (N_31861,N_30185,N_30272);
nand U31862 (N_31862,N_30477,N_30476);
and U31863 (N_31863,N_30568,N_30105);
nand U31864 (N_31864,N_30504,N_30806);
nor U31865 (N_31865,N_30586,N_30154);
nor U31866 (N_31866,N_30990,N_30596);
nor U31867 (N_31867,N_30579,N_30689);
and U31868 (N_31868,N_30464,N_30338);
nor U31869 (N_31869,N_30269,N_30489);
nor U31870 (N_31870,N_30589,N_30012);
xor U31871 (N_31871,N_30902,N_30133);
xor U31872 (N_31872,N_30018,N_30482);
xnor U31873 (N_31873,N_30018,N_30232);
xor U31874 (N_31874,N_30248,N_30457);
or U31875 (N_31875,N_30388,N_30925);
and U31876 (N_31876,N_30897,N_30455);
nand U31877 (N_31877,N_30545,N_30152);
and U31878 (N_31878,N_30338,N_30734);
nand U31879 (N_31879,N_30316,N_30343);
and U31880 (N_31880,N_30617,N_30912);
nor U31881 (N_31881,N_30117,N_30104);
or U31882 (N_31882,N_30240,N_30059);
nand U31883 (N_31883,N_30194,N_30376);
or U31884 (N_31884,N_30835,N_30522);
nand U31885 (N_31885,N_30986,N_30319);
or U31886 (N_31886,N_30931,N_30303);
xnor U31887 (N_31887,N_30142,N_30357);
xnor U31888 (N_31888,N_30258,N_30961);
or U31889 (N_31889,N_30577,N_30325);
xor U31890 (N_31890,N_30815,N_30098);
xnor U31891 (N_31891,N_30331,N_30684);
nand U31892 (N_31892,N_30866,N_30095);
or U31893 (N_31893,N_30607,N_30099);
and U31894 (N_31894,N_30714,N_30287);
or U31895 (N_31895,N_30752,N_30062);
or U31896 (N_31896,N_30241,N_30430);
and U31897 (N_31897,N_30040,N_30651);
or U31898 (N_31898,N_30082,N_30471);
xnor U31899 (N_31899,N_30302,N_30891);
xnor U31900 (N_31900,N_30281,N_30539);
xor U31901 (N_31901,N_30735,N_30324);
nand U31902 (N_31902,N_30785,N_30578);
nor U31903 (N_31903,N_30384,N_30976);
nand U31904 (N_31904,N_30660,N_30955);
nand U31905 (N_31905,N_30405,N_30056);
and U31906 (N_31906,N_30770,N_30596);
nor U31907 (N_31907,N_30866,N_30818);
or U31908 (N_31908,N_30234,N_30152);
or U31909 (N_31909,N_30124,N_30683);
nor U31910 (N_31910,N_30864,N_30486);
and U31911 (N_31911,N_30466,N_30267);
and U31912 (N_31912,N_30163,N_30136);
or U31913 (N_31913,N_30423,N_30547);
or U31914 (N_31914,N_30199,N_30798);
or U31915 (N_31915,N_30188,N_30644);
nor U31916 (N_31916,N_30018,N_30669);
nor U31917 (N_31917,N_30450,N_30871);
xor U31918 (N_31918,N_30632,N_30012);
xnor U31919 (N_31919,N_30187,N_30789);
nor U31920 (N_31920,N_30882,N_30413);
xor U31921 (N_31921,N_30536,N_30640);
or U31922 (N_31922,N_30553,N_30634);
nor U31923 (N_31923,N_30693,N_30290);
and U31924 (N_31924,N_30573,N_30626);
nand U31925 (N_31925,N_30067,N_30305);
xnor U31926 (N_31926,N_30253,N_30476);
xor U31927 (N_31927,N_30855,N_30289);
and U31928 (N_31928,N_30821,N_30888);
xnor U31929 (N_31929,N_30744,N_30835);
nand U31930 (N_31930,N_30244,N_30198);
and U31931 (N_31931,N_30670,N_30351);
and U31932 (N_31932,N_30712,N_30621);
and U31933 (N_31933,N_30070,N_30752);
and U31934 (N_31934,N_30123,N_30465);
or U31935 (N_31935,N_30429,N_30952);
and U31936 (N_31936,N_30013,N_30583);
nand U31937 (N_31937,N_30255,N_30488);
or U31938 (N_31938,N_30230,N_30829);
nand U31939 (N_31939,N_30177,N_30077);
nor U31940 (N_31940,N_30889,N_30126);
and U31941 (N_31941,N_30092,N_30199);
xor U31942 (N_31942,N_30791,N_30046);
nand U31943 (N_31943,N_30901,N_30989);
nor U31944 (N_31944,N_30340,N_30509);
xnor U31945 (N_31945,N_30080,N_30548);
nand U31946 (N_31946,N_30479,N_30723);
and U31947 (N_31947,N_30445,N_30542);
xnor U31948 (N_31948,N_30921,N_30143);
or U31949 (N_31949,N_30208,N_30377);
nor U31950 (N_31950,N_30287,N_30985);
nor U31951 (N_31951,N_30751,N_30429);
nand U31952 (N_31952,N_30851,N_30640);
or U31953 (N_31953,N_30104,N_30360);
nand U31954 (N_31954,N_30820,N_30795);
xor U31955 (N_31955,N_30981,N_30832);
nor U31956 (N_31956,N_30329,N_30440);
nand U31957 (N_31957,N_30960,N_30248);
or U31958 (N_31958,N_30824,N_30003);
nand U31959 (N_31959,N_30675,N_30530);
nor U31960 (N_31960,N_30842,N_30896);
nor U31961 (N_31961,N_30060,N_30092);
and U31962 (N_31962,N_30016,N_30318);
nand U31963 (N_31963,N_30491,N_30391);
nand U31964 (N_31964,N_30670,N_30715);
and U31965 (N_31965,N_30438,N_30524);
nand U31966 (N_31966,N_30531,N_30278);
and U31967 (N_31967,N_30852,N_30888);
nor U31968 (N_31968,N_30318,N_30059);
and U31969 (N_31969,N_30433,N_30010);
nand U31970 (N_31970,N_30776,N_30764);
nor U31971 (N_31971,N_30484,N_30504);
xnor U31972 (N_31972,N_30313,N_30640);
nor U31973 (N_31973,N_30180,N_30281);
xnor U31974 (N_31974,N_30799,N_30341);
or U31975 (N_31975,N_30396,N_30159);
and U31976 (N_31976,N_30725,N_30280);
or U31977 (N_31977,N_30173,N_30649);
xnor U31978 (N_31978,N_30031,N_30959);
nand U31979 (N_31979,N_30507,N_30911);
and U31980 (N_31980,N_30494,N_30023);
xor U31981 (N_31981,N_30858,N_30719);
nand U31982 (N_31982,N_30768,N_30787);
xor U31983 (N_31983,N_30528,N_30285);
or U31984 (N_31984,N_30407,N_30727);
xor U31985 (N_31985,N_30274,N_30266);
xor U31986 (N_31986,N_30997,N_30038);
nor U31987 (N_31987,N_30437,N_30766);
nand U31988 (N_31988,N_30434,N_30701);
and U31989 (N_31989,N_30724,N_30870);
nand U31990 (N_31990,N_30270,N_30173);
nor U31991 (N_31991,N_30040,N_30101);
and U31992 (N_31992,N_30026,N_30116);
nand U31993 (N_31993,N_30224,N_30981);
nand U31994 (N_31994,N_30027,N_30781);
xor U31995 (N_31995,N_30384,N_30989);
nand U31996 (N_31996,N_30642,N_30750);
and U31997 (N_31997,N_30393,N_30046);
xnor U31998 (N_31998,N_30555,N_30853);
or U31999 (N_31999,N_30445,N_30276);
or U32000 (N_32000,N_31451,N_31112);
nor U32001 (N_32001,N_31904,N_31897);
xnor U32002 (N_32002,N_31801,N_31173);
and U32003 (N_32003,N_31729,N_31001);
and U32004 (N_32004,N_31760,N_31289);
xnor U32005 (N_32005,N_31363,N_31196);
xnor U32006 (N_32006,N_31641,N_31181);
and U32007 (N_32007,N_31975,N_31156);
nand U32008 (N_32008,N_31361,N_31479);
nand U32009 (N_32009,N_31371,N_31403);
nor U32010 (N_32010,N_31531,N_31901);
and U32011 (N_32011,N_31033,N_31638);
xor U32012 (N_32012,N_31567,N_31958);
nand U32013 (N_32013,N_31459,N_31551);
and U32014 (N_32014,N_31094,N_31581);
nand U32015 (N_32015,N_31832,N_31034);
and U32016 (N_32016,N_31983,N_31994);
or U32017 (N_32017,N_31322,N_31616);
xnor U32018 (N_32018,N_31954,N_31596);
xnor U32019 (N_32019,N_31464,N_31239);
nor U32020 (N_32020,N_31389,N_31853);
nand U32021 (N_32021,N_31758,N_31810);
or U32022 (N_32022,N_31797,N_31323);
or U32023 (N_32023,N_31227,N_31827);
and U32024 (N_32024,N_31053,N_31846);
or U32025 (N_32025,N_31183,N_31896);
nor U32026 (N_32026,N_31730,N_31973);
nor U32027 (N_32027,N_31413,N_31829);
xor U32028 (N_32028,N_31334,N_31948);
or U32029 (N_32029,N_31280,N_31978);
and U32030 (N_32030,N_31905,N_31169);
nor U32031 (N_32031,N_31397,N_31633);
nor U32032 (N_32032,N_31436,N_31842);
or U32033 (N_32033,N_31400,N_31944);
or U32034 (N_32034,N_31935,N_31252);
xor U32035 (N_32035,N_31009,N_31737);
and U32036 (N_32036,N_31606,N_31131);
and U32037 (N_32037,N_31898,N_31279);
nor U32038 (N_32038,N_31664,N_31051);
and U32039 (N_32039,N_31063,N_31221);
nand U32040 (N_32040,N_31226,N_31177);
nand U32041 (N_32041,N_31611,N_31467);
and U32042 (N_32042,N_31534,N_31979);
or U32043 (N_32043,N_31881,N_31912);
or U32044 (N_32044,N_31012,N_31122);
nand U32045 (N_32045,N_31207,N_31791);
and U32046 (N_32046,N_31320,N_31027);
or U32047 (N_32047,N_31779,N_31355);
nor U32048 (N_32048,N_31845,N_31340);
or U32049 (N_32049,N_31670,N_31483);
nor U32050 (N_32050,N_31811,N_31894);
nand U32051 (N_32051,N_31293,N_31563);
or U32052 (N_32052,N_31546,N_31667);
xor U32053 (N_32053,N_31775,N_31380);
and U32054 (N_32054,N_31578,N_31420);
and U32055 (N_32055,N_31088,N_31060);
xnor U32056 (N_32056,N_31594,N_31140);
nor U32057 (N_32057,N_31374,N_31536);
nor U32058 (N_32058,N_31931,N_31520);
nand U32059 (N_32059,N_31532,N_31964);
nand U32060 (N_32060,N_31158,N_31786);
or U32061 (N_32061,N_31042,N_31178);
or U32062 (N_32062,N_31584,N_31657);
xor U32063 (N_32063,N_31615,N_31794);
and U32064 (N_32064,N_31602,N_31268);
and U32065 (N_32065,N_31351,N_31133);
nor U32066 (N_32066,N_31702,N_31992);
xor U32067 (N_32067,N_31834,N_31650);
nand U32068 (N_32068,N_31461,N_31151);
or U32069 (N_32069,N_31127,N_31362);
xor U32070 (N_32070,N_31301,N_31428);
or U32071 (N_32071,N_31022,N_31540);
or U32072 (N_32072,N_31463,N_31785);
nand U32073 (N_32073,N_31206,N_31020);
nor U32074 (N_32074,N_31422,N_31684);
or U32075 (N_32075,N_31035,N_31683);
nor U32076 (N_32076,N_31561,N_31315);
and U32077 (N_32077,N_31365,N_31445);
nand U32078 (N_32078,N_31082,N_31883);
nand U32079 (N_32079,N_31195,N_31701);
nand U32080 (N_32080,N_31241,N_31704);
nand U32081 (N_32081,N_31333,N_31840);
or U32082 (N_32082,N_31346,N_31266);
xor U32083 (N_32083,N_31887,N_31052);
xor U32084 (N_32084,N_31432,N_31854);
nor U32085 (N_32085,N_31861,N_31774);
or U32086 (N_32086,N_31273,N_31435);
nand U32087 (N_32087,N_31076,N_31538);
nand U32088 (N_32088,N_31449,N_31286);
xor U32089 (N_32089,N_31360,N_31695);
xor U32090 (N_32090,N_31607,N_31850);
nor U32091 (N_32091,N_31314,N_31145);
nand U32092 (N_32092,N_31216,N_31645);
and U32093 (N_32093,N_31044,N_31822);
or U32094 (N_32094,N_31613,N_31788);
nand U32095 (N_32095,N_31185,N_31799);
xnor U32096 (N_32096,N_31516,N_31671);
and U32097 (N_32097,N_31477,N_31240);
nand U32098 (N_32098,N_31608,N_31056);
and U32099 (N_32099,N_31751,N_31620);
xnor U32100 (N_32100,N_31324,N_31424);
nor U32101 (N_32101,N_31356,N_31587);
nand U32102 (N_32102,N_31752,N_31621);
xnor U32103 (N_32103,N_31798,N_31271);
xnor U32104 (N_32104,N_31238,N_31625);
xor U32105 (N_32105,N_31098,N_31844);
xor U32106 (N_32106,N_31640,N_31599);
nand U32107 (N_32107,N_31685,N_31163);
or U32108 (N_32108,N_31568,N_31366);
nand U32109 (N_32109,N_31580,N_31182);
and U32110 (N_32110,N_31984,N_31203);
or U32111 (N_32111,N_31655,N_31624);
nor U32112 (N_32112,N_31600,N_31336);
nand U32113 (N_32113,N_31038,N_31610);
nand U32114 (N_32114,N_31288,N_31265);
nor U32115 (N_32115,N_31705,N_31263);
or U32116 (N_32116,N_31512,N_31833);
nand U32117 (N_32117,N_31628,N_31865);
nor U32118 (N_32118,N_31899,N_31426);
and U32119 (N_32119,N_31824,N_31807);
or U32120 (N_32120,N_31116,N_31444);
xor U32121 (N_32121,N_31858,N_31443);
xnor U32122 (N_32122,N_31826,N_31966);
and U32123 (N_32123,N_31511,N_31915);
and U32124 (N_32124,N_31668,N_31062);
xnor U32125 (N_32125,N_31500,N_31588);
nor U32126 (N_32126,N_31418,N_31805);
xor U32127 (N_32127,N_31302,N_31951);
and U32128 (N_32128,N_31651,N_31728);
or U32129 (N_32129,N_31055,N_31697);
xnor U32130 (N_32130,N_31254,N_31859);
xnor U32131 (N_32131,N_31184,N_31072);
nand U32132 (N_32132,N_31687,N_31851);
xor U32133 (N_32133,N_31748,N_31485);
and U32134 (N_32134,N_31727,N_31490);
nand U32135 (N_32135,N_31732,N_31455);
or U32136 (N_32136,N_31764,N_31554);
xor U32137 (N_32137,N_31117,N_31576);
xor U32138 (N_32138,N_31714,N_31011);
nor U32139 (N_32139,N_31803,N_31558);
nor U32140 (N_32140,N_31662,N_31390);
or U32141 (N_32141,N_31812,N_31553);
or U32142 (N_32142,N_31202,N_31749);
nand U32143 (N_32143,N_31077,N_31916);
xor U32144 (N_32144,N_31497,N_31820);
and U32145 (N_32145,N_31115,N_31802);
nor U32146 (N_32146,N_31108,N_31719);
xor U32147 (N_32147,N_31157,N_31547);
and U32148 (N_32148,N_31943,N_31016);
or U32149 (N_32149,N_31379,N_31257);
or U32150 (N_32150,N_31080,N_31929);
nor U32151 (N_32151,N_31880,N_31849);
xnor U32152 (N_32152,N_31586,N_31574);
or U32153 (N_32153,N_31715,N_31046);
and U32154 (N_32154,N_31643,N_31223);
and U32155 (N_32155,N_31783,N_31126);
or U32156 (N_32156,N_31562,N_31735);
or U32157 (N_32157,N_31677,N_31014);
xor U32158 (N_32158,N_31959,N_31109);
xor U32159 (N_32159,N_31407,N_31470);
xnor U32160 (N_32160,N_31676,N_31637);
and U32161 (N_32161,N_31468,N_31523);
or U32162 (N_32162,N_31316,N_31731);
and U32163 (N_32163,N_31101,N_31498);
or U32164 (N_32164,N_31245,N_31300);
nand U32165 (N_32165,N_31525,N_31047);
and U32166 (N_32166,N_31328,N_31617);
and U32167 (N_32167,N_31548,N_31416);
and U32168 (N_32168,N_31137,N_31394);
and U32169 (N_32169,N_31879,N_31246);
xnor U32170 (N_32170,N_31491,N_31770);
nand U32171 (N_32171,N_31527,N_31373);
nand U32172 (N_32172,N_31890,N_31214);
and U32173 (N_32173,N_31125,N_31260);
nor U32174 (N_32174,N_31440,N_31255);
nand U32175 (N_32175,N_31437,N_31644);
nor U32176 (N_32176,N_31068,N_31800);
xor U32177 (N_32177,N_31040,N_31065);
and U32178 (N_32178,N_31544,N_31556);
or U32179 (N_32179,N_31739,N_31968);
nand U32180 (N_32180,N_31867,N_31130);
or U32181 (N_32181,N_31384,N_31589);
nand U32182 (N_32182,N_31989,N_31093);
or U32183 (N_32183,N_31388,N_31933);
nor U32184 (N_32184,N_31176,N_31004);
and U32185 (N_32185,N_31285,N_31318);
xor U32186 (N_32186,N_31796,N_31233);
nor U32187 (N_32187,N_31926,N_31903);
and U32188 (N_32188,N_31224,N_31253);
and U32189 (N_32189,N_31090,N_31306);
nor U32190 (N_32190,N_31187,N_31745);
or U32191 (N_32191,N_31308,N_31514);
or U32192 (N_32192,N_31136,N_31746);
and U32193 (N_32193,N_31790,N_31338);
nand U32194 (N_32194,N_31993,N_31290);
or U32195 (N_32195,N_31383,N_31283);
nand U32196 (N_32196,N_31160,N_31331);
and U32197 (N_32197,N_31595,N_31629);
xnor U32198 (N_32198,N_31287,N_31194);
or U32199 (N_32199,N_31930,N_31393);
and U32200 (N_32200,N_31692,N_31956);
xnor U32201 (N_32201,N_31504,N_31965);
or U32202 (N_32202,N_31906,N_31953);
or U32203 (N_32203,N_31612,N_31067);
xor U32204 (N_32204,N_31674,N_31635);
nor U32205 (N_32205,N_31381,N_31937);
nand U32206 (N_32206,N_31541,N_31878);
or U32207 (N_32207,N_31804,N_31493);
or U32208 (N_32208,N_31352,N_31741);
nor U32209 (N_32209,N_31032,N_31866);
nand U32210 (N_32210,N_31335,N_31086);
xnor U32211 (N_32211,N_31707,N_31663);
or U32212 (N_32212,N_31010,N_31089);
nand U32213 (N_32213,N_31962,N_31756);
nand U32214 (N_32214,N_31700,N_31609);
nor U32215 (N_32215,N_31847,N_31092);
nor U32216 (N_32216,N_31682,N_31874);
nand U32217 (N_32217,N_31367,N_31294);
and U32218 (N_32218,N_31515,N_31138);
nand U32219 (N_32219,N_31069,N_31917);
nor U32220 (N_32220,N_31496,N_31876);
nand U32221 (N_32221,N_31278,N_31703);
nor U32222 (N_32222,N_31050,N_31311);
nor U32223 (N_32223,N_31484,N_31210);
nor U32224 (N_32224,N_31593,N_31292);
nor U32225 (N_32225,N_31186,N_31572);
or U32226 (N_32226,N_31166,N_31114);
or U32227 (N_32227,N_31919,N_31066);
nand U32228 (N_32228,N_31354,N_31539);
xor U32229 (N_32229,N_31597,N_31763);
and U32230 (N_32230,N_31559,N_31211);
nor U32231 (N_32231,N_31344,N_31911);
or U32232 (N_32232,N_31319,N_31345);
nor U32233 (N_32233,N_31141,N_31139);
xnor U32234 (N_32234,N_31711,N_31402);
nand U32235 (N_32235,N_31773,N_31873);
or U32236 (N_32236,N_31699,N_31401);
or U32237 (N_32237,N_31134,N_31781);
nand U32238 (N_32238,N_31936,N_31005);
and U32239 (N_32239,N_31924,N_31408);
or U32240 (N_32240,N_31619,N_31395);
xnor U32241 (N_32241,N_31870,N_31232);
and U32242 (N_32242,N_31678,N_31605);
nand U32243 (N_32243,N_31375,N_31332);
nor U32244 (N_32244,N_31037,N_31149);
or U32245 (N_32245,N_31144,N_31575);
nand U32246 (N_32246,N_31771,N_31425);
nor U32247 (N_32247,N_31941,N_31099);
and U32248 (N_32248,N_31601,N_31350);
nor U32249 (N_32249,N_31660,N_31618);
nand U32250 (N_32250,N_31049,N_31018);
or U32251 (N_32251,N_31446,N_31891);
nor U32252 (N_32252,N_31236,N_31565);
xor U32253 (N_32253,N_31008,N_31955);
and U32254 (N_32254,N_31475,N_31398);
nor U32255 (N_32255,N_31421,N_31517);
nand U32256 (N_32256,N_31342,N_31368);
or U32257 (N_32257,N_31220,N_31521);
nand U32258 (N_32258,N_31075,N_31995);
nor U32259 (N_32259,N_31852,N_31990);
or U32260 (N_32260,N_31998,N_31113);
nand U32261 (N_32261,N_31478,N_31922);
nand U32262 (N_32262,N_31305,N_31209);
nand U32263 (N_32263,N_31495,N_31839);
xor U32264 (N_32264,N_31923,N_31469);
nand U32265 (N_32265,N_31769,N_31171);
xnor U32266 (N_32266,N_31698,N_31070);
and U32267 (N_32267,N_31025,N_31213);
nor U32268 (N_32268,N_31466,N_31843);
xnor U32269 (N_32269,N_31501,N_31458);
nand U32270 (N_32270,N_31877,N_31604);
xnor U32271 (N_32271,N_31806,N_31084);
nand U32272 (N_32272,N_31048,N_31198);
and U32273 (N_32273,N_31622,N_31471);
nand U32274 (N_32274,N_31079,N_31019);
nand U32275 (N_32275,N_31369,N_31439);
nand U32276 (N_32276,N_31681,N_31128);
xor U32277 (N_32277,N_31623,N_31603);
nand U32278 (N_32278,N_31180,N_31808);
xor U32279 (N_32279,N_31399,N_31585);
xor U32280 (N_32280,N_31480,N_31441);
or U32281 (N_32281,N_31487,N_31768);
xnor U32282 (N_32282,N_31339,N_31091);
or U32283 (N_32283,N_31583,N_31230);
xnor U32284 (N_32284,N_31672,N_31100);
and U32285 (N_32285,N_31474,N_31343);
and U32286 (N_32286,N_31448,N_31789);
nor U32287 (N_32287,N_31248,N_31148);
and U32288 (N_32288,N_31353,N_31337);
or U32289 (N_32289,N_31256,N_31892);
nor U32290 (N_32290,N_31460,N_31205);
nor U32291 (N_32291,N_31885,N_31999);
and U32292 (N_32292,N_31653,N_31918);
nor U32293 (N_32293,N_31696,N_31564);
or U32294 (N_32294,N_31242,N_31074);
nand U32295 (N_32295,N_31431,N_31039);
and U32296 (N_32296,N_31809,N_31957);
nor U32297 (N_32297,N_31864,N_31064);
and U32298 (N_32298,N_31244,N_31105);
nand U32299 (N_32299,N_31712,N_31251);
and U32300 (N_32300,N_31900,N_31329);
nand U32301 (N_32301,N_31427,N_31188);
nand U32302 (N_32302,N_31762,N_31147);
and U32303 (N_32303,N_31830,N_31942);
and U32304 (N_32304,N_31269,N_31723);
and U32305 (N_32305,N_31190,N_31502);
and U32306 (N_32306,N_31738,N_31003);
xnor U32307 (N_32307,N_31888,N_31433);
and U32308 (N_32308,N_31325,N_31831);
nand U32309 (N_32309,N_31073,N_31893);
or U32310 (N_32310,N_31454,N_31974);
and U32311 (N_32311,N_31518,N_31658);
or U32312 (N_32312,N_31875,N_31818);
and U32313 (N_32313,N_31987,N_31192);
xnor U32314 (N_32314,N_31218,N_31028);
nand U32315 (N_32315,N_31920,N_31243);
and U32316 (N_32316,N_31921,N_31225);
and U32317 (N_32317,N_31489,N_31412);
nand U32318 (N_32318,N_31526,N_31259);
xnor U32319 (N_32319,N_31364,N_31882);
or U32320 (N_32320,N_31952,N_31309);
xnor U32321 (N_32321,N_31519,N_31823);
nand U32322 (N_32322,N_31270,N_31405);
or U32323 (N_32323,N_31197,N_31659);
and U32324 (N_32324,N_31646,N_31571);
or U32325 (N_32325,N_31652,N_31792);
nand U32326 (N_32326,N_31036,N_31761);
nor U32327 (N_32327,N_31940,N_31939);
and U32328 (N_32328,N_31825,N_31235);
and U32329 (N_32329,N_31041,N_31642);
xor U32330 (N_32330,N_31175,N_31179);
xnor U32331 (N_32331,N_31472,N_31152);
xnor U32332 (N_32332,N_31647,N_31945);
and U32333 (N_32333,N_31733,N_31299);
nand U32334 (N_32334,N_31102,N_31950);
and U32335 (N_32335,N_31780,N_31330);
nand U32336 (N_32336,N_31111,N_31988);
nand U32337 (N_32337,N_31766,N_31215);
and U32338 (N_32338,N_31910,N_31162);
xnor U32339 (N_32339,N_31784,N_31550);
nand U32340 (N_32340,N_31423,N_31560);
xnor U32341 (N_32341,N_31121,N_31058);
nor U32342 (N_32342,N_31376,N_31656);
or U32343 (N_32343,N_31972,N_31669);
nor U32344 (N_32344,N_31598,N_31303);
nand U32345 (N_32345,N_31410,N_31262);
nand U32346 (N_32346,N_31537,N_31726);
or U32347 (N_32347,N_31636,N_31476);
nand U32348 (N_32348,N_31078,N_31895);
nand U32349 (N_32349,N_31317,N_31710);
nand U32350 (N_32350,N_31409,N_31632);
xnor U32351 (N_32351,N_31247,N_31872);
xnor U32352 (N_32352,N_31626,N_31396);
and U32353 (N_32353,N_31986,N_31757);
or U32354 (N_32354,N_31026,N_31778);
and U32355 (N_32355,N_31776,N_31661);
or U32356 (N_32356,N_31835,N_31297);
nor U32357 (N_32357,N_31414,N_31524);
xor U32358 (N_32358,N_31284,N_31530);
and U32359 (N_32359,N_31411,N_31848);
and U32360 (N_32360,N_31577,N_31997);
and U32361 (N_32361,N_31155,N_31680);
and U32362 (N_32362,N_31694,N_31347);
or U32363 (N_32363,N_31579,N_31170);
nand U32364 (N_32364,N_31691,N_31782);
nor U32365 (N_32365,N_31506,N_31816);
or U32366 (N_32366,N_31960,N_31724);
and U32367 (N_32367,N_31884,N_31391);
nand U32368 (N_32368,N_31429,N_31281);
or U32369 (N_32369,N_31573,N_31120);
xor U32370 (N_32370,N_31015,N_31907);
and U32371 (N_32371,N_31725,N_31119);
nor U32372 (N_32372,N_31902,N_31002);
or U32373 (N_32373,N_31234,N_31971);
or U32374 (N_32374,N_31718,N_31570);
nor U32375 (N_32375,N_31963,N_31860);
xor U32376 (N_32376,N_31191,N_31529);
nor U32377 (N_32377,N_31510,N_31021);
and U32378 (N_32378,N_31296,N_31688);
nor U32379 (N_32379,N_31291,N_31857);
or U32380 (N_32380,N_31406,N_31321);
nand U32381 (N_32381,N_31648,N_31542);
and U32382 (N_32382,N_31980,N_31666);
and U32383 (N_32383,N_31819,N_31313);
xnor U32384 (N_32384,N_31693,N_31482);
xor U32385 (N_32385,N_31499,N_31465);
xnor U32386 (N_32386,N_31535,N_31552);
nor U32387 (N_32387,N_31507,N_31675);
and U32388 (N_32388,N_31889,N_31492);
nand U32389 (N_32389,N_31934,N_31392);
xor U32390 (N_32390,N_31654,N_31000);
nand U32391 (N_32391,N_31932,N_31359);
or U32392 (N_32392,N_31310,N_31208);
or U32393 (N_32393,N_31634,N_31085);
or U32394 (N_32394,N_31167,N_31708);
or U32395 (N_32395,N_31689,N_31153);
xnor U32396 (N_32396,N_31341,N_31985);
and U32397 (N_32397,N_31118,N_31837);
and U32398 (N_32398,N_31417,N_31777);
xor U32399 (N_32399,N_31276,N_31795);
nand U32400 (N_32400,N_31555,N_31862);
or U32401 (N_32401,N_31753,N_31868);
and U32402 (N_32402,N_31017,N_31106);
and U32403 (N_32403,N_31097,N_31249);
nor U32404 (N_32404,N_31057,N_31045);
nor U32405 (N_32405,N_31582,N_31107);
nor U32406 (N_32406,N_31061,N_31772);
xnor U32407 (N_32407,N_31592,N_31528);
nor U32408 (N_32408,N_31456,N_31168);
or U32409 (N_32409,N_31630,N_31307);
nor U32410 (N_32410,N_31434,N_31631);
and U32411 (N_32411,N_31023,N_31457);
xor U32412 (N_32412,N_31508,N_31522);
nand U32413 (N_32413,N_31913,N_31081);
nand U32414 (N_32414,N_31327,N_31679);
or U32415 (N_32415,N_31549,N_31229);
nor U32416 (N_32416,N_31452,N_31349);
nor U32417 (N_32417,N_31787,N_31473);
and U32418 (N_32418,N_31566,N_31029);
nor U32419 (N_32419,N_31231,N_31071);
or U32420 (N_32420,N_31754,N_31513);
nor U32421 (N_32421,N_31744,N_31386);
and U32422 (N_32422,N_31970,N_31649);
nand U32423 (N_32423,N_31981,N_31357);
or U32424 (N_32424,N_31007,N_31836);
nand U32425 (N_32425,N_31264,N_31043);
xnor U32426 (N_32426,N_31404,N_31488);
nand U32427 (N_32427,N_31569,N_31372);
and U32428 (N_32428,N_31982,N_31886);
xor U32429 (N_32429,N_31871,N_31274);
nand U32430 (N_32430,N_31450,N_31172);
or U32431 (N_32431,N_31298,N_31031);
nand U32432 (N_32432,N_31201,N_31348);
nand U32433 (N_32433,N_31486,N_31096);
nand U32434 (N_32434,N_31419,N_31736);
nand U32435 (N_32435,N_31557,N_31146);
or U32436 (N_32436,N_31841,N_31104);
and U32437 (N_32437,N_31765,N_31716);
or U32438 (N_32438,N_31509,N_31481);
xor U32439 (N_32439,N_31747,N_31415);
nor U32440 (N_32440,N_31665,N_31838);
and U32441 (N_32441,N_31438,N_31969);
nand U32442 (N_32442,N_31947,N_31909);
xnor U32443 (N_32443,N_31750,N_31855);
and U32444 (N_32444,N_31272,N_31275);
nor U32445 (N_32445,N_31755,N_31869);
or U32446 (N_32446,N_31154,N_31124);
nand U32447 (N_32447,N_31150,N_31237);
and U32448 (N_32448,N_31219,N_31713);
nor U32449 (N_32449,N_31813,N_31721);
nor U32450 (N_32450,N_31949,N_31142);
nor U32451 (N_32451,N_31991,N_31013);
and U32452 (N_32452,N_31250,N_31793);
nor U32453 (N_32453,N_31159,N_31814);
and U32454 (N_32454,N_31908,N_31914);
and U32455 (N_32455,N_31453,N_31590);
xnor U32456 (N_32456,N_31382,N_31006);
and U32457 (N_32457,N_31815,N_31204);
and U32458 (N_32458,N_31996,N_31129);
nand U32459 (N_32459,N_31686,N_31030);
nand U32460 (N_32460,N_31087,N_31828);
xor U32461 (N_32461,N_31734,N_31165);
nand U32462 (N_32462,N_31024,N_31863);
nand U32463 (N_32463,N_31326,N_31946);
nand U32464 (N_32464,N_31967,N_31817);
nand U32465 (N_32465,N_31927,N_31282);
and U32466 (N_32466,N_31174,N_31673);
nand U32467 (N_32467,N_31494,N_31200);
and U32468 (N_32468,N_31387,N_31358);
or U32469 (N_32469,N_31742,N_31977);
xor U32470 (N_32470,N_31132,N_31312);
or U32471 (N_32471,N_31503,N_31161);
or U32472 (N_32472,N_31543,N_31743);
and U32473 (N_32473,N_31709,N_31103);
nand U32474 (N_32474,N_31447,N_31639);
or U32475 (N_32475,N_31261,N_31222);
nand U32476 (N_32476,N_31267,N_31545);
and U32477 (N_32477,N_31083,N_31759);
nor U32478 (N_32478,N_31110,N_31189);
and U32479 (N_32479,N_31143,N_31533);
or U32480 (N_32480,N_31370,N_31123);
and U32481 (N_32481,N_31193,N_31385);
xor U32482 (N_32482,N_31304,N_31706);
nor U32483 (N_32483,N_31722,N_31442);
or U32484 (N_32484,N_31462,N_31217);
nand U32485 (N_32485,N_31135,N_31054);
nor U32486 (N_32486,N_31591,N_31627);
nand U32487 (N_32487,N_31976,N_31767);
nor U32488 (N_32488,N_31925,N_31821);
nor U32489 (N_32489,N_31258,N_31212);
nand U32490 (N_32490,N_31228,N_31961);
and U32491 (N_32491,N_31717,N_31377);
or U32492 (N_32492,N_31277,N_31295);
xnor U32493 (N_32493,N_31505,N_31690);
nand U32494 (N_32494,N_31928,N_31430);
or U32495 (N_32495,N_31378,N_31614);
or U32496 (N_32496,N_31059,N_31856);
and U32497 (N_32497,N_31199,N_31095);
nand U32498 (N_32498,N_31740,N_31164);
and U32499 (N_32499,N_31938,N_31720);
or U32500 (N_32500,N_31368,N_31121);
and U32501 (N_32501,N_31840,N_31760);
nor U32502 (N_32502,N_31577,N_31283);
nor U32503 (N_32503,N_31125,N_31870);
nand U32504 (N_32504,N_31641,N_31772);
and U32505 (N_32505,N_31530,N_31351);
and U32506 (N_32506,N_31181,N_31057);
xor U32507 (N_32507,N_31291,N_31859);
xnor U32508 (N_32508,N_31094,N_31184);
xor U32509 (N_32509,N_31625,N_31189);
or U32510 (N_32510,N_31987,N_31230);
xnor U32511 (N_32511,N_31581,N_31725);
and U32512 (N_32512,N_31989,N_31326);
or U32513 (N_32513,N_31685,N_31258);
or U32514 (N_32514,N_31884,N_31394);
nor U32515 (N_32515,N_31750,N_31601);
nand U32516 (N_32516,N_31113,N_31506);
nor U32517 (N_32517,N_31357,N_31238);
and U32518 (N_32518,N_31637,N_31730);
xnor U32519 (N_32519,N_31911,N_31940);
nand U32520 (N_32520,N_31415,N_31351);
xnor U32521 (N_32521,N_31824,N_31247);
and U32522 (N_32522,N_31594,N_31639);
and U32523 (N_32523,N_31296,N_31397);
nand U32524 (N_32524,N_31303,N_31910);
or U32525 (N_32525,N_31634,N_31475);
nor U32526 (N_32526,N_31367,N_31147);
or U32527 (N_32527,N_31834,N_31664);
nor U32528 (N_32528,N_31948,N_31692);
nand U32529 (N_32529,N_31749,N_31704);
xnor U32530 (N_32530,N_31930,N_31281);
xor U32531 (N_32531,N_31294,N_31642);
xor U32532 (N_32532,N_31000,N_31402);
xor U32533 (N_32533,N_31230,N_31569);
nor U32534 (N_32534,N_31701,N_31228);
and U32535 (N_32535,N_31969,N_31925);
and U32536 (N_32536,N_31653,N_31640);
or U32537 (N_32537,N_31793,N_31655);
nand U32538 (N_32538,N_31319,N_31535);
or U32539 (N_32539,N_31558,N_31324);
and U32540 (N_32540,N_31068,N_31458);
xor U32541 (N_32541,N_31327,N_31888);
or U32542 (N_32542,N_31378,N_31846);
nor U32543 (N_32543,N_31184,N_31297);
and U32544 (N_32544,N_31133,N_31140);
nor U32545 (N_32545,N_31646,N_31860);
xor U32546 (N_32546,N_31133,N_31979);
xnor U32547 (N_32547,N_31007,N_31543);
nand U32548 (N_32548,N_31339,N_31086);
or U32549 (N_32549,N_31241,N_31556);
and U32550 (N_32550,N_31405,N_31366);
xor U32551 (N_32551,N_31395,N_31627);
nor U32552 (N_32552,N_31801,N_31119);
nand U32553 (N_32553,N_31070,N_31910);
and U32554 (N_32554,N_31958,N_31722);
and U32555 (N_32555,N_31031,N_31049);
nor U32556 (N_32556,N_31430,N_31470);
nor U32557 (N_32557,N_31295,N_31153);
nand U32558 (N_32558,N_31623,N_31048);
nor U32559 (N_32559,N_31325,N_31102);
or U32560 (N_32560,N_31599,N_31970);
or U32561 (N_32561,N_31605,N_31912);
nor U32562 (N_32562,N_31636,N_31944);
nand U32563 (N_32563,N_31783,N_31319);
nand U32564 (N_32564,N_31275,N_31493);
or U32565 (N_32565,N_31810,N_31096);
xor U32566 (N_32566,N_31505,N_31991);
and U32567 (N_32567,N_31203,N_31012);
and U32568 (N_32568,N_31191,N_31007);
or U32569 (N_32569,N_31466,N_31062);
xnor U32570 (N_32570,N_31548,N_31299);
xnor U32571 (N_32571,N_31389,N_31331);
nand U32572 (N_32572,N_31053,N_31136);
xnor U32573 (N_32573,N_31469,N_31001);
or U32574 (N_32574,N_31415,N_31853);
nor U32575 (N_32575,N_31838,N_31553);
and U32576 (N_32576,N_31873,N_31917);
and U32577 (N_32577,N_31784,N_31491);
and U32578 (N_32578,N_31165,N_31151);
nor U32579 (N_32579,N_31715,N_31680);
and U32580 (N_32580,N_31290,N_31306);
nor U32581 (N_32581,N_31946,N_31425);
xnor U32582 (N_32582,N_31420,N_31755);
or U32583 (N_32583,N_31426,N_31282);
and U32584 (N_32584,N_31809,N_31221);
nand U32585 (N_32585,N_31757,N_31600);
or U32586 (N_32586,N_31893,N_31756);
xor U32587 (N_32587,N_31895,N_31928);
or U32588 (N_32588,N_31308,N_31536);
or U32589 (N_32589,N_31505,N_31206);
or U32590 (N_32590,N_31504,N_31880);
xor U32591 (N_32591,N_31968,N_31707);
or U32592 (N_32592,N_31390,N_31400);
or U32593 (N_32593,N_31985,N_31009);
and U32594 (N_32594,N_31436,N_31008);
and U32595 (N_32595,N_31655,N_31370);
or U32596 (N_32596,N_31751,N_31314);
xor U32597 (N_32597,N_31160,N_31078);
and U32598 (N_32598,N_31650,N_31238);
nor U32599 (N_32599,N_31971,N_31372);
xor U32600 (N_32600,N_31896,N_31590);
nor U32601 (N_32601,N_31616,N_31912);
or U32602 (N_32602,N_31523,N_31832);
nand U32603 (N_32603,N_31953,N_31303);
nor U32604 (N_32604,N_31183,N_31671);
or U32605 (N_32605,N_31833,N_31725);
xor U32606 (N_32606,N_31869,N_31837);
or U32607 (N_32607,N_31283,N_31190);
and U32608 (N_32608,N_31320,N_31364);
xor U32609 (N_32609,N_31325,N_31388);
nor U32610 (N_32610,N_31788,N_31440);
xor U32611 (N_32611,N_31852,N_31475);
nor U32612 (N_32612,N_31715,N_31481);
nand U32613 (N_32613,N_31593,N_31637);
xnor U32614 (N_32614,N_31231,N_31953);
and U32615 (N_32615,N_31679,N_31012);
nand U32616 (N_32616,N_31033,N_31529);
nand U32617 (N_32617,N_31968,N_31586);
or U32618 (N_32618,N_31878,N_31884);
xor U32619 (N_32619,N_31536,N_31270);
nor U32620 (N_32620,N_31514,N_31830);
nand U32621 (N_32621,N_31110,N_31748);
nand U32622 (N_32622,N_31560,N_31528);
nor U32623 (N_32623,N_31474,N_31451);
nand U32624 (N_32624,N_31483,N_31369);
nand U32625 (N_32625,N_31435,N_31976);
nand U32626 (N_32626,N_31134,N_31153);
nand U32627 (N_32627,N_31267,N_31542);
or U32628 (N_32628,N_31522,N_31303);
xnor U32629 (N_32629,N_31504,N_31282);
or U32630 (N_32630,N_31011,N_31190);
nand U32631 (N_32631,N_31545,N_31305);
xnor U32632 (N_32632,N_31587,N_31179);
nand U32633 (N_32633,N_31787,N_31700);
nand U32634 (N_32634,N_31896,N_31676);
nand U32635 (N_32635,N_31558,N_31202);
and U32636 (N_32636,N_31723,N_31484);
nor U32637 (N_32637,N_31972,N_31913);
and U32638 (N_32638,N_31512,N_31522);
nor U32639 (N_32639,N_31448,N_31466);
nor U32640 (N_32640,N_31585,N_31287);
or U32641 (N_32641,N_31510,N_31255);
and U32642 (N_32642,N_31771,N_31332);
nor U32643 (N_32643,N_31335,N_31248);
nor U32644 (N_32644,N_31129,N_31225);
nor U32645 (N_32645,N_31713,N_31674);
nand U32646 (N_32646,N_31750,N_31403);
xor U32647 (N_32647,N_31092,N_31180);
xnor U32648 (N_32648,N_31876,N_31372);
xor U32649 (N_32649,N_31623,N_31137);
nand U32650 (N_32650,N_31347,N_31510);
nor U32651 (N_32651,N_31102,N_31688);
or U32652 (N_32652,N_31221,N_31609);
xor U32653 (N_32653,N_31353,N_31948);
and U32654 (N_32654,N_31192,N_31196);
nor U32655 (N_32655,N_31643,N_31863);
and U32656 (N_32656,N_31436,N_31467);
or U32657 (N_32657,N_31767,N_31731);
nor U32658 (N_32658,N_31353,N_31476);
nor U32659 (N_32659,N_31313,N_31295);
xnor U32660 (N_32660,N_31653,N_31383);
nor U32661 (N_32661,N_31500,N_31364);
and U32662 (N_32662,N_31423,N_31378);
or U32663 (N_32663,N_31171,N_31184);
or U32664 (N_32664,N_31407,N_31142);
xor U32665 (N_32665,N_31691,N_31747);
xnor U32666 (N_32666,N_31149,N_31212);
xor U32667 (N_32667,N_31655,N_31481);
and U32668 (N_32668,N_31787,N_31803);
nor U32669 (N_32669,N_31236,N_31605);
and U32670 (N_32670,N_31412,N_31049);
nand U32671 (N_32671,N_31758,N_31095);
or U32672 (N_32672,N_31753,N_31553);
and U32673 (N_32673,N_31903,N_31914);
and U32674 (N_32674,N_31493,N_31487);
nand U32675 (N_32675,N_31246,N_31249);
nand U32676 (N_32676,N_31139,N_31784);
nor U32677 (N_32677,N_31408,N_31566);
nor U32678 (N_32678,N_31224,N_31791);
or U32679 (N_32679,N_31146,N_31196);
and U32680 (N_32680,N_31722,N_31702);
xnor U32681 (N_32681,N_31048,N_31214);
and U32682 (N_32682,N_31200,N_31725);
nand U32683 (N_32683,N_31614,N_31831);
and U32684 (N_32684,N_31228,N_31604);
nor U32685 (N_32685,N_31713,N_31656);
nor U32686 (N_32686,N_31181,N_31100);
and U32687 (N_32687,N_31889,N_31074);
and U32688 (N_32688,N_31739,N_31839);
nor U32689 (N_32689,N_31912,N_31693);
and U32690 (N_32690,N_31438,N_31234);
or U32691 (N_32691,N_31363,N_31805);
nand U32692 (N_32692,N_31484,N_31892);
nand U32693 (N_32693,N_31357,N_31112);
xnor U32694 (N_32694,N_31728,N_31249);
and U32695 (N_32695,N_31317,N_31327);
nand U32696 (N_32696,N_31603,N_31631);
nor U32697 (N_32697,N_31015,N_31805);
and U32698 (N_32698,N_31082,N_31131);
xor U32699 (N_32699,N_31962,N_31177);
xnor U32700 (N_32700,N_31272,N_31321);
xor U32701 (N_32701,N_31407,N_31222);
or U32702 (N_32702,N_31132,N_31811);
nand U32703 (N_32703,N_31049,N_31298);
or U32704 (N_32704,N_31692,N_31413);
nor U32705 (N_32705,N_31238,N_31837);
nor U32706 (N_32706,N_31573,N_31306);
and U32707 (N_32707,N_31829,N_31920);
xnor U32708 (N_32708,N_31393,N_31715);
nor U32709 (N_32709,N_31233,N_31094);
and U32710 (N_32710,N_31844,N_31696);
nand U32711 (N_32711,N_31382,N_31196);
or U32712 (N_32712,N_31606,N_31937);
xor U32713 (N_32713,N_31649,N_31358);
nor U32714 (N_32714,N_31460,N_31254);
nand U32715 (N_32715,N_31085,N_31331);
nand U32716 (N_32716,N_31393,N_31899);
and U32717 (N_32717,N_31869,N_31661);
nor U32718 (N_32718,N_31222,N_31553);
or U32719 (N_32719,N_31284,N_31027);
nor U32720 (N_32720,N_31839,N_31351);
xnor U32721 (N_32721,N_31367,N_31675);
or U32722 (N_32722,N_31485,N_31800);
or U32723 (N_32723,N_31281,N_31026);
and U32724 (N_32724,N_31500,N_31819);
xnor U32725 (N_32725,N_31936,N_31329);
xor U32726 (N_32726,N_31677,N_31168);
xor U32727 (N_32727,N_31795,N_31755);
or U32728 (N_32728,N_31437,N_31511);
xor U32729 (N_32729,N_31181,N_31739);
xnor U32730 (N_32730,N_31985,N_31767);
nand U32731 (N_32731,N_31288,N_31970);
or U32732 (N_32732,N_31142,N_31924);
xor U32733 (N_32733,N_31976,N_31481);
nand U32734 (N_32734,N_31306,N_31044);
xor U32735 (N_32735,N_31051,N_31457);
or U32736 (N_32736,N_31012,N_31746);
or U32737 (N_32737,N_31115,N_31388);
xnor U32738 (N_32738,N_31544,N_31023);
or U32739 (N_32739,N_31988,N_31445);
or U32740 (N_32740,N_31967,N_31102);
nor U32741 (N_32741,N_31613,N_31111);
nand U32742 (N_32742,N_31868,N_31065);
and U32743 (N_32743,N_31290,N_31446);
or U32744 (N_32744,N_31039,N_31837);
or U32745 (N_32745,N_31937,N_31967);
nor U32746 (N_32746,N_31516,N_31710);
nor U32747 (N_32747,N_31797,N_31642);
and U32748 (N_32748,N_31341,N_31587);
nor U32749 (N_32749,N_31828,N_31219);
and U32750 (N_32750,N_31170,N_31118);
nor U32751 (N_32751,N_31394,N_31266);
or U32752 (N_32752,N_31018,N_31169);
or U32753 (N_32753,N_31551,N_31495);
and U32754 (N_32754,N_31642,N_31367);
nand U32755 (N_32755,N_31549,N_31801);
and U32756 (N_32756,N_31517,N_31262);
or U32757 (N_32757,N_31630,N_31132);
nand U32758 (N_32758,N_31191,N_31919);
nand U32759 (N_32759,N_31829,N_31772);
nand U32760 (N_32760,N_31319,N_31045);
xor U32761 (N_32761,N_31254,N_31915);
and U32762 (N_32762,N_31826,N_31863);
or U32763 (N_32763,N_31914,N_31122);
or U32764 (N_32764,N_31142,N_31324);
or U32765 (N_32765,N_31613,N_31384);
xor U32766 (N_32766,N_31122,N_31700);
xnor U32767 (N_32767,N_31016,N_31163);
nand U32768 (N_32768,N_31263,N_31081);
and U32769 (N_32769,N_31514,N_31747);
and U32770 (N_32770,N_31474,N_31829);
nor U32771 (N_32771,N_31222,N_31436);
nand U32772 (N_32772,N_31789,N_31174);
nor U32773 (N_32773,N_31472,N_31330);
xor U32774 (N_32774,N_31753,N_31878);
and U32775 (N_32775,N_31516,N_31674);
and U32776 (N_32776,N_31086,N_31551);
nor U32777 (N_32777,N_31091,N_31003);
nand U32778 (N_32778,N_31795,N_31308);
or U32779 (N_32779,N_31991,N_31713);
and U32780 (N_32780,N_31658,N_31226);
or U32781 (N_32781,N_31073,N_31300);
xnor U32782 (N_32782,N_31236,N_31331);
or U32783 (N_32783,N_31071,N_31353);
and U32784 (N_32784,N_31473,N_31642);
or U32785 (N_32785,N_31729,N_31332);
or U32786 (N_32786,N_31907,N_31871);
and U32787 (N_32787,N_31690,N_31926);
nor U32788 (N_32788,N_31041,N_31375);
xor U32789 (N_32789,N_31962,N_31689);
nor U32790 (N_32790,N_31053,N_31968);
xnor U32791 (N_32791,N_31163,N_31890);
nand U32792 (N_32792,N_31770,N_31683);
xor U32793 (N_32793,N_31112,N_31554);
nand U32794 (N_32794,N_31047,N_31101);
nand U32795 (N_32795,N_31060,N_31630);
or U32796 (N_32796,N_31204,N_31206);
xnor U32797 (N_32797,N_31108,N_31863);
xor U32798 (N_32798,N_31186,N_31203);
or U32799 (N_32799,N_31448,N_31833);
xnor U32800 (N_32800,N_31245,N_31529);
nand U32801 (N_32801,N_31368,N_31236);
and U32802 (N_32802,N_31236,N_31748);
and U32803 (N_32803,N_31261,N_31088);
or U32804 (N_32804,N_31206,N_31351);
nand U32805 (N_32805,N_31492,N_31844);
or U32806 (N_32806,N_31821,N_31935);
nand U32807 (N_32807,N_31076,N_31418);
nor U32808 (N_32808,N_31305,N_31649);
xor U32809 (N_32809,N_31733,N_31322);
or U32810 (N_32810,N_31912,N_31860);
nand U32811 (N_32811,N_31072,N_31065);
xor U32812 (N_32812,N_31440,N_31946);
or U32813 (N_32813,N_31973,N_31392);
nand U32814 (N_32814,N_31318,N_31957);
nand U32815 (N_32815,N_31764,N_31788);
nor U32816 (N_32816,N_31425,N_31791);
or U32817 (N_32817,N_31013,N_31607);
nor U32818 (N_32818,N_31843,N_31944);
nor U32819 (N_32819,N_31850,N_31522);
nor U32820 (N_32820,N_31632,N_31468);
or U32821 (N_32821,N_31337,N_31513);
xnor U32822 (N_32822,N_31162,N_31286);
and U32823 (N_32823,N_31773,N_31095);
and U32824 (N_32824,N_31855,N_31265);
and U32825 (N_32825,N_31979,N_31271);
xnor U32826 (N_32826,N_31613,N_31869);
nor U32827 (N_32827,N_31823,N_31341);
nand U32828 (N_32828,N_31765,N_31791);
and U32829 (N_32829,N_31213,N_31998);
or U32830 (N_32830,N_31538,N_31010);
nor U32831 (N_32831,N_31044,N_31996);
or U32832 (N_32832,N_31487,N_31034);
nor U32833 (N_32833,N_31800,N_31974);
xnor U32834 (N_32834,N_31683,N_31305);
or U32835 (N_32835,N_31598,N_31761);
or U32836 (N_32836,N_31200,N_31105);
nand U32837 (N_32837,N_31299,N_31114);
nor U32838 (N_32838,N_31669,N_31114);
nand U32839 (N_32839,N_31834,N_31901);
nand U32840 (N_32840,N_31073,N_31102);
xor U32841 (N_32841,N_31048,N_31774);
xor U32842 (N_32842,N_31090,N_31581);
nand U32843 (N_32843,N_31250,N_31670);
nor U32844 (N_32844,N_31845,N_31211);
or U32845 (N_32845,N_31066,N_31314);
and U32846 (N_32846,N_31902,N_31867);
xnor U32847 (N_32847,N_31351,N_31552);
nor U32848 (N_32848,N_31000,N_31806);
xor U32849 (N_32849,N_31494,N_31401);
nor U32850 (N_32850,N_31178,N_31847);
xor U32851 (N_32851,N_31790,N_31936);
and U32852 (N_32852,N_31118,N_31381);
and U32853 (N_32853,N_31969,N_31911);
and U32854 (N_32854,N_31001,N_31396);
nor U32855 (N_32855,N_31029,N_31089);
xnor U32856 (N_32856,N_31640,N_31702);
or U32857 (N_32857,N_31045,N_31996);
or U32858 (N_32858,N_31924,N_31842);
nor U32859 (N_32859,N_31849,N_31235);
or U32860 (N_32860,N_31698,N_31262);
and U32861 (N_32861,N_31147,N_31004);
nand U32862 (N_32862,N_31068,N_31568);
or U32863 (N_32863,N_31126,N_31086);
xor U32864 (N_32864,N_31307,N_31188);
and U32865 (N_32865,N_31740,N_31473);
xnor U32866 (N_32866,N_31204,N_31656);
and U32867 (N_32867,N_31624,N_31733);
nand U32868 (N_32868,N_31458,N_31534);
nor U32869 (N_32869,N_31539,N_31124);
nand U32870 (N_32870,N_31844,N_31550);
nor U32871 (N_32871,N_31853,N_31031);
and U32872 (N_32872,N_31772,N_31664);
nor U32873 (N_32873,N_31872,N_31663);
nor U32874 (N_32874,N_31383,N_31470);
xnor U32875 (N_32875,N_31351,N_31962);
nand U32876 (N_32876,N_31279,N_31664);
nor U32877 (N_32877,N_31808,N_31489);
xnor U32878 (N_32878,N_31112,N_31995);
nor U32879 (N_32879,N_31183,N_31141);
xnor U32880 (N_32880,N_31750,N_31509);
and U32881 (N_32881,N_31869,N_31680);
xor U32882 (N_32882,N_31406,N_31455);
nor U32883 (N_32883,N_31035,N_31463);
or U32884 (N_32884,N_31524,N_31707);
and U32885 (N_32885,N_31956,N_31203);
xnor U32886 (N_32886,N_31752,N_31472);
nor U32887 (N_32887,N_31510,N_31214);
xnor U32888 (N_32888,N_31144,N_31906);
xnor U32889 (N_32889,N_31368,N_31041);
and U32890 (N_32890,N_31313,N_31244);
nor U32891 (N_32891,N_31202,N_31594);
nor U32892 (N_32892,N_31477,N_31052);
xnor U32893 (N_32893,N_31305,N_31504);
nand U32894 (N_32894,N_31846,N_31616);
nand U32895 (N_32895,N_31413,N_31630);
nand U32896 (N_32896,N_31891,N_31527);
and U32897 (N_32897,N_31736,N_31011);
or U32898 (N_32898,N_31289,N_31857);
and U32899 (N_32899,N_31945,N_31757);
nand U32900 (N_32900,N_31921,N_31044);
xor U32901 (N_32901,N_31409,N_31002);
or U32902 (N_32902,N_31918,N_31045);
or U32903 (N_32903,N_31715,N_31928);
nor U32904 (N_32904,N_31070,N_31151);
and U32905 (N_32905,N_31302,N_31646);
or U32906 (N_32906,N_31678,N_31649);
xnor U32907 (N_32907,N_31000,N_31261);
xor U32908 (N_32908,N_31356,N_31202);
and U32909 (N_32909,N_31838,N_31769);
and U32910 (N_32910,N_31883,N_31241);
nor U32911 (N_32911,N_31958,N_31867);
or U32912 (N_32912,N_31811,N_31688);
or U32913 (N_32913,N_31209,N_31541);
and U32914 (N_32914,N_31105,N_31263);
xnor U32915 (N_32915,N_31125,N_31009);
or U32916 (N_32916,N_31263,N_31944);
and U32917 (N_32917,N_31318,N_31798);
nor U32918 (N_32918,N_31765,N_31867);
xnor U32919 (N_32919,N_31458,N_31758);
nand U32920 (N_32920,N_31186,N_31512);
nor U32921 (N_32921,N_31150,N_31186);
nand U32922 (N_32922,N_31541,N_31355);
nand U32923 (N_32923,N_31255,N_31756);
xnor U32924 (N_32924,N_31394,N_31372);
or U32925 (N_32925,N_31979,N_31424);
nand U32926 (N_32926,N_31119,N_31780);
and U32927 (N_32927,N_31277,N_31413);
and U32928 (N_32928,N_31515,N_31852);
nand U32929 (N_32929,N_31358,N_31006);
nor U32930 (N_32930,N_31345,N_31160);
nor U32931 (N_32931,N_31262,N_31929);
and U32932 (N_32932,N_31542,N_31407);
or U32933 (N_32933,N_31591,N_31022);
and U32934 (N_32934,N_31164,N_31823);
nor U32935 (N_32935,N_31887,N_31662);
xnor U32936 (N_32936,N_31880,N_31072);
xnor U32937 (N_32937,N_31633,N_31110);
and U32938 (N_32938,N_31924,N_31991);
and U32939 (N_32939,N_31062,N_31061);
and U32940 (N_32940,N_31784,N_31002);
xnor U32941 (N_32941,N_31722,N_31593);
nand U32942 (N_32942,N_31512,N_31070);
or U32943 (N_32943,N_31500,N_31417);
xor U32944 (N_32944,N_31868,N_31261);
nor U32945 (N_32945,N_31896,N_31032);
or U32946 (N_32946,N_31361,N_31020);
nor U32947 (N_32947,N_31281,N_31266);
nor U32948 (N_32948,N_31705,N_31461);
xnor U32949 (N_32949,N_31300,N_31074);
xor U32950 (N_32950,N_31050,N_31573);
nor U32951 (N_32951,N_31851,N_31986);
nor U32952 (N_32952,N_31376,N_31927);
nor U32953 (N_32953,N_31536,N_31843);
and U32954 (N_32954,N_31984,N_31590);
xnor U32955 (N_32955,N_31531,N_31856);
or U32956 (N_32956,N_31534,N_31841);
nand U32957 (N_32957,N_31009,N_31657);
nand U32958 (N_32958,N_31871,N_31873);
nand U32959 (N_32959,N_31799,N_31719);
and U32960 (N_32960,N_31197,N_31305);
nand U32961 (N_32961,N_31407,N_31615);
nor U32962 (N_32962,N_31994,N_31943);
nand U32963 (N_32963,N_31031,N_31939);
and U32964 (N_32964,N_31221,N_31662);
or U32965 (N_32965,N_31222,N_31354);
and U32966 (N_32966,N_31088,N_31469);
nand U32967 (N_32967,N_31971,N_31862);
nor U32968 (N_32968,N_31483,N_31717);
xor U32969 (N_32969,N_31424,N_31113);
xnor U32970 (N_32970,N_31672,N_31590);
xnor U32971 (N_32971,N_31588,N_31172);
nand U32972 (N_32972,N_31389,N_31064);
and U32973 (N_32973,N_31774,N_31937);
xnor U32974 (N_32974,N_31076,N_31319);
and U32975 (N_32975,N_31268,N_31073);
xor U32976 (N_32976,N_31580,N_31796);
and U32977 (N_32977,N_31227,N_31071);
xor U32978 (N_32978,N_31190,N_31487);
nand U32979 (N_32979,N_31372,N_31004);
xnor U32980 (N_32980,N_31718,N_31299);
nor U32981 (N_32981,N_31559,N_31965);
and U32982 (N_32982,N_31459,N_31617);
and U32983 (N_32983,N_31110,N_31622);
nand U32984 (N_32984,N_31245,N_31849);
and U32985 (N_32985,N_31241,N_31383);
nor U32986 (N_32986,N_31594,N_31167);
or U32987 (N_32987,N_31302,N_31501);
or U32988 (N_32988,N_31785,N_31172);
nor U32989 (N_32989,N_31688,N_31166);
or U32990 (N_32990,N_31587,N_31852);
and U32991 (N_32991,N_31651,N_31733);
and U32992 (N_32992,N_31881,N_31884);
nand U32993 (N_32993,N_31151,N_31162);
or U32994 (N_32994,N_31815,N_31355);
or U32995 (N_32995,N_31703,N_31911);
and U32996 (N_32996,N_31231,N_31957);
or U32997 (N_32997,N_31584,N_31850);
xnor U32998 (N_32998,N_31891,N_31668);
and U32999 (N_32999,N_31129,N_31621);
nand U33000 (N_33000,N_32197,N_32574);
nor U33001 (N_33001,N_32837,N_32713);
and U33002 (N_33002,N_32024,N_32431);
nor U33003 (N_33003,N_32471,N_32691);
or U33004 (N_33004,N_32988,N_32060);
nand U33005 (N_33005,N_32482,N_32853);
nor U33006 (N_33006,N_32188,N_32229);
xor U33007 (N_33007,N_32566,N_32783);
nor U33008 (N_33008,N_32746,N_32932);
xnor U33009 (N_33009,N_32429,N_32308);
xor U33010 (N_33010,N_32523,N_32138);
or U33011 (N_33011,N_32495,N_32982);
or U33012 (N_33012,N_32112,N_32362);
nor U33013 (N_33013,N_32442,N_32305);
and U33014 (N_33014,N_32347,N_32017);
or U33015 (N_33015,N_32407,N_32217);
or U33016 (N_33016,N_32199,N_32022);
nand U33017 (N_33017,N_32789,N_32264);
and U33018 (N_33018,N_32425,N_32408);
xor U33019 (N_33019,N_32587,N_32351);
nor U33020 (N_33020,N_32326,N_32657);
nor U33021 (N_33021,N_32702,N_32526);
xnor U33022 (N_33022,N_32121,N_32033);
nand U33023 (N_33023,N_32763,N_32277);
xnor U33024 (N_33024,N_32677,N_32740);
nor U33025 (N_33025,N_32851,N_32933);
nor U33026 (N_33026,N_32039,N_32714);
and U33027 (N_33027,N_32070,N_32293);
nor U33028 (N_33028,N_32300,N_32899);
nor U33029 (N_33029,N_32370,N_32669);
xnor U33030 (N_33030,N_32272,N_32075);
nor U33031 (N_33031,N_32211,N_32614);
nand U33032 (N_33032,N_32536,N_32306);
xnor U33033 (N_33033,N_32001,N_32196);
nor U33034 (N_33034,N_32828,N_32884);
nand U33035 (N_33035,N_32808,N_32765);
nor U33036 (N_33036,N_32413,N_32575);
nor U33037 (N_33037,N_32236,N_32115);
or U33038 (N_33038,N_32053,N_32498);
and U33039 (N_33039,N_32318,N_32662);
and U33040 (N_33040,N_32984,N_32462);
xor U33041 (N_33041,N_32269,N_32481);
nor U33042 (N_33042,N_32220,N_32928);
nand U33043 (N_33043,N_32667,N_32364);
nand U33044 (N_33044,N_32080,N_32924);
nor U33045 (N_33045,N_32049,N_32720);
xor U33046 (N_33046,N_32971,N_32164);
nand U33047 (N_33047,N_32023,N_32289);
nand U33048 (N_33048,N_32965,N_32005);
nand U33049 (N_33049,N_32866,N_32156);
nor U33050 (N_33050,N_32317,N_32360);
nor U33051 (N_33051,N_32799,N_32281);
or U33052 (N_33052,N_32215,N_32962);
nor U33053 (N_33053,N_32203,N_32478);
and U33054 (N_33054,N_32245,N_32149);
nor U33055 (N_33055,N_32037,N_32622);
nor U33056 (N_33056,N_32592,N_32371);
xor U33057 (N_33057,N_32675,N_32985);
and U33058 (N_33058,N_32943,N_32313);
or U33059 (N_33059,N_32180,N_32729);
nand U33060 (N_33060,N_32441,N_32346);
or U33061 (N_33061,N_32190,N_32081);
nand U33062 (N_33062,N_32865,N_32448);
or U33063 (N_33063,N_32843,N_32086);
nor U33064 (N_33064,N_32282,N_32824);
nor U33065 (N_33065,N_32268,N_32493);
nand U33066 (N_33066,N_32440,N_32076);
xor U33067 (N_33067,N_32189,N_32959);
nor U33068 (N_33068,N_32650,N_32434);
nand U33069 (N_33069,N_32455,N_32626);
nor U33070 (N_33070,N_32106,N_32003);
and U33071 (N_33071,N_32820,N_32031);
nand U33072 (N_33072,N_32607,N_32627);
or U33073 (N_33073,N_32420,N_32500);
or U33074 (N_33074,N_32689,N_32375);
nor U33075 (N_33075,N_32134,N_32176);
nand U33076 (N_33076,N_32548,N_32841);
nand U33077 (N_33077,N_32946,N_32116);
nand U33078 (N_33078,N_32635,N_32571);
nand U33079 (N_33079,N_32887,N_32530);
nor U33080 (N_33080,N_32251,N_32972);
and U33081 (N_33081,N_32382,N_32775);
or U33082 (N_33082,N_32405,N_32496);
or U33083 (N_33083,N_32288,N_32485);
nand U33084 (N_33084,N_32201,N_32873);
xnor U33085 (N_33085,N_32468,N_32761);
or U33086 (N_33086,N_32903,N_32432);
nor U33087 (N_33087,N_32367,N_32557);
nor U33088 (N_33088,N_32867,N_32334);
nand U33089 (N_33089,N_32718,N_32999);
nor U33090 (N_33090,N_32803,N_32815);
nor U33091 (N_33091,N_32111,N_32414);
nand U33092 (N_33092,N_32400,N_32386);
nor U33093 (N_33093,N_32886,N_32205);
nand U33094 (N_33094,N_32206,N_32531);
and U33095 (N_33095,N_32396,N_32067);
and U33096 (N_33096,N_32731,N_32410);
nand U33097 (N_33097,N_32983,N_32778);
or U33098 (N_33098,N_32178,N_32036);
xnor U33099 (N_33099,N_32030,N_32917);
and U33100 (N_33100,N_32320,N_32467);
and U33101 (N_33101,N_32093,N_32255);
nor U33102 (N_33102,N_32920,N_32350);
nand U33103 (N_33103,N_32144,N_32257);
nand U33104 (N_33104,N_32921,N_32950);
and U33105 (N_33105,N_32435,N_32054);
nand U33106 (N_33106,N_32072,N_32006);
nor U33107 (N_33107,N_32788,N_32826);
nand U33108 (N_33108,N_32524,N_32751);
and U33109 (N_33109,N_32916,N_32831);
or U33110 (N_33110,N_32135,N_32995);
nand U33111 (N_33111,N_32918,N_32732);
and U33112 (N_33112,N_32028,N_32249);
xnor U33113 (N_33113,N_32380,N_32658);
and U33114 (N_33114,N_32940,N_32609);
nand U33115 (N_33115,N_32838,N_32353);
nand U33116 (N_33116,N_32167,N_32114);
and U33117 (N_33117,N_32143,N_32693);
and U33118 (N_33118,N_32007,N_32673);
or U33119 (N_33119,N_32891,N_32861);
and U33120 (N_33120,N_32155,N_32449);
or U33121 (N_33121,N_32337,N_32146);
or U33122 (N_33122,N_32046,N_32295);
xnor U33123 (N_33123,N_32221,N_32395);
nor U33124 (N_33124,N_32951,N_32686);
or U33125 (N_33125,N_32543,N_32428);
or U33126 (N_33126,N_32094,N_32291);
xor U33127 (N_33127,N_32562,N_32653);
or U33128 (N_33128,N_32676,N_32058);
nor U33129 (N_33129,N_32503,N_32707);
and U33130 (N_33130,N_32508,N_32847);
and U33131 (N_33131,N_32942,N_32085);
nand U33132 (N_33132,N_32564,N_32792);
or U33133 (N_33133,N_32252,N_32097);
and U33134 (N_33134,N_32666,N_32781);
xor U33135 (N_33135,N_32889,N_32758);
and U33136 (N_33136,N_32931,N_32234);
or U33137 (N_33137,N_32577,N_32324);
and U33138 (N_33138,N_32749,N_32734);
nand U33139 (N_33139,N_32628,N_32404);
xor U33140 (N_33140,N_32911,N_32358);
nand U33141 (N_33141,N_32491,N_32095);
xnor U33142 (N_33142,N_32338,N_32898);
nand U33143 (N_33143,N_32172,N_32356);
or U33144 (N_33144,N_32430,N_32256);
nand U33145 (N_33145,N_32807,N_32872);
and U33146 (N_33146,N_32954,N_32542);
nand U33147 (N_33147,N_32796,N_32907);
or U33148 (N_33148,N_32992,N_32618);
nand U33149 (N_33149,N_32230,N_32701);
nand U33150 (N_33150,N_32363,N_32671);
nand U33151 (N_33151,N_32977,N_32079);
xnor U33152 (N_33152,N_32549,N_32239);
nor U33153 (N_33153,N_32640,N_32705);
nor U33154 (N_33154,N_32848,N_32069);
xor U33155 (N_33155,N_32605,N_32219);
and U33156 (N_33156,N_32736,N_32868);
nor U33157 (N_33157,N_32223,N_32665);
xnor U33158 (N_33158,N_32596,N_32050);
xor U33159 (N_33159,N_32525,N_32451);
and U33160 (N_33160,N_32019,N_32238);
or U33161 (N_33161,N_32142,N_32610);
xnor U33162 (N_33162,N_32539,N_32532);
or U33163 (N_33163,N_32439,N_32949);
nand U33164 (N_33164,N_32603,N_32325);
or U33165 (N_33165,N_32846,N_32029);
or U33166 (N_33166,N_32699,N_32329);
or U33167 (N_33167,N_32963,N_32926);
and U33168 (N_33168,N_32032,N_32569);
nand U33169 (N_33169,N_32266,N_32585);
nand U33170 (N_33170,N_32099,N_32715);
xor U33171 (N_33171,N_32927,N_32730);
or U33172 (N_33172,N_32941,N_32104);
xnor U33173 (N_33173,N_32208,N_32506);
nand U33174 (N_33174,N_32579,N_32727);
and U33175 (N_33175,N_32819,N_32157);
nor U33176 (N_33176,N_32896,N_32975);
nor U33177 (N_33177,N_32688,N_32647);
xnor U33178 (N_33178,N_32009,N_32960);
and U33179 (N_33179,N_32581,N_32348);
xor U33180 (N_33180,N_32991,N_32993);
or U33181 (N_33181,N_32475,N_32381);
or U33182 (N_33182,N_32922,N_32047);
nor U33183 (N_33183,N_32314,N_32604);
xnor U33184 (N_33184,N_32473,N_32694);
xor U33185 (N_33185,N_32162,N_32725);
nor U33186 (N_33186,N_32845,N_32588);
and U33187 (N_33187,N_32644,N_32589);
nor U33188 (N_33188,N_32110,N_32515);
nand U33189 (N_33189,N_32421,N_32674);
nand U33190 (N_33190,N_32745,N_32417);
xor U33191 (N_33191,N_32335,N_32177);
and U33192 (N_33192,N_32136,N_32849);
nand U33193 (N_33193,N_32710,N_32790);
xor U33194 (N_33194,N_32812,N_32833);
nand U33195 (N_33195,N_32042,N_32565);
xnor U33196 (N_33196,N_32297,N_32186);
nand U33197 (N_33197,N_32519,N_32860);
nor U33198 (N_33198,N_32641,N_32222);
xnor U33199 (N_33199,N_32038,N_32064);
nand U33200 (N_33200,N_32100,N_32169);
or U33201 (N_33201,N_32474,N_32411);
and U33202 (N_33202,N_32298,N_32881);
nand U33203 (N_33203,N_32192,N_32102);
and U33204 (N_33204,N_32012,N_32472);
nor U33205 (N_33205,N_32590,N_32956);
nand U33206 (N_33206,N_32128,N_32020);
and U33207 (N_33207,N_32782,N_32418);
xnor U33208 (N_33208,N_32900,N_32398);
or U33209 (N_33209,N_32355,N_32332);
and U33210 (N_33210,N_32213,N_32857);
nor U33211 (N_33211,N_32385,N_32952);
or U33212 (N_33212,N_32810,N_32466);
xor U33213 (N_33213,N_32476,N_32057);
xor U33214 (N_33214,N_32646,N_32243);
nand U33215 (N_33215,N_32384,N_32158);
or U33216 (N_33216,N_32880,N_32994);
or U33217 (N_33217,N_32773,N_32232);
nor U33218 (N_33218,N_32859,N_32179);
or U33219 (N_33219,N_32556,N_32161);
nor U33220 (N_33220,N_32250,N_32387);
nor U33221 (N_33221,N_32690,N_32901);
xor U33222 (N_33222,N_32550,N_32580);
nand U33223 (N_33223,N_32762,N_32620);
xnor U33224 (N_33224,N_32538,N_32593);
nor U33225 (N_33225,N_32632,N_32154);
nand U33226 (N_33226,N_32415,N_32748);
nor U33227 (N_33227,N_32814,N_32913);
nor U33228 (N_33228,N_32310,N_32754);
nand U33229 (N_33229,N_32235,N_32888);
or U33230 (N_33230,N_32349,N_32997);
xor U33231 (N_33231,N_32505,N_32487);
xor U33232 (N_33232,N_32105,N_32004);
xnor U33233 (N_33233,N_32263,N_32809);
xor U33234 (N_33234,N_32541,N_32254);
xor U33235 (N_33235,N_32312,N_32021);
nand U33236 (N_33236,N_32262,N_32122);
nand U33237 (N_33237,N_32444,N_32551);
nor U33238 (N_33238,N_32366,N_32150);
or U33239 (N_33239,N_32096,N_32141);
and U33240 (N_33240,N_32433,N_32759);
nor U33241 (N_33241,N_32996,N_32168);
and U33242 (N_33242,N_32267,N_32611);
nand U33243 (N_33243,N_32450,N_32802);
nor U33244 (N_33244,N_32120,N_32805);
nor U33245 (N_33245,N_32777,N_32737);
nand U33246 (N_33246,N_32661,N_32704);
nand U33247 (N_33247,N_32247,N_32642);
nor U33248 (N_33248,N_32461,N_32212);
nor U33249 (N_33249,N_32744,N_32533);
and U33250 (N_33250,N_32711,N_32124);
and U33251 (N_33251,N_32406,N_32108);
or U33252 (N_33252,N_32345,N_32813);
or U33253 (N_33253,N_32753,N_32739);
or U33254 (N_33254,N_32774,N_32035);
nor U33255 (N_33255,N_32659,N_32507);
or U33256 (N_33256,N_32275,N_32591);
and U33257 (N_33257,N_32629,N_32490);
xnor U33258 (N_33258,N_32027,N_32521);
and U33259 (N_33259,N_32204,N_32460);
and U33260 (N_33260,N_32193,N_32552);
xor U33261 (N_33261,N_32595,N_32957);
nand U33262 (N_33262,N_32131,N_32504);
xnor U33263 (N_33263,N_32925,N_32352);
xnor U33264 (N_33264,N_32163,N_32682);
nand U33265 (N_33265,N_32173,N_32651);
nand U33266 (N_33266,N_32559,N_32426);
xor U33267 (N_33267,N_32553,N_32311);
xor U33268 (N_33268,N_32379,N_32098);
and U33269 (N_33269,N_32445,N_32091);
nor U33270 (N_33270,N_32258,N_32750);
or U33271 (N_33271,N_32517,N_32403);
and U33272 (N_33272,N_32283,N_32130);
xor U33273 (N_33273,N_32637,N_32228);
and U33274 (N_33274,N_32409,N_32512);
nor U33275 (N_33275,N_32897,N_32459);
nor U33276 (N_33276,N_32735,N_32225);
xnor U33277 (N_33277,N_32365,N_32852);
and U33278 (N_33278,N_32113,N_32265);
xor U33279 (N_33279,N_32546,N_32002);
or U33280 (N_33280,N_32246,N_32437);
nand U33281 (N_33281,N_32516,N_32339);
or U33282 (N_33282,N_32465,N_32499);
nand U33283 (N_33283,N_32034,N_32502);
nand U33284 (N_33284,N_32638,N_32087);
nor U33285 (N_33285,N_32066,N_32547);
nor U33286 (N_33286,N_32331,N_32798);
nor U33287 (N_33287,N_32818,N_32680);
and U33288 (N_33288,N_32890,N_32484);
nand U33289 (N_33289,N_32107,N_32520);
xnor U33290 (N_33290,N_32578,N_32025);
nor U33291 (N_33291,N_32301,N_32078);
xnor U33292 (N_33292,N_32801,N_32989);
nor U33293 (N_33293,N_32719,N_32576);
nand U33294 (N_33294,N_32606,N_32752);
nor U33295 (N_33295,N_32117,N_32287);
xnor U33296 (N_33296,N_32560,N_32392);
nand U33297 (N_33297,N_32393,N_32863);
nand U33298 (N_33298,N_32529,N_32043);
nor U33299 (N_33299,N_32194,N_32563);
or U33300 (N_33300,N_32929,N_32584);
xor U33301 (N_33301,N_32717,N_32870);
or U33302 (N_33302,N_32464,N_32955);
xor U33303 (N_33303,N_32290,N_32200);
nor U33304 (N_33304,N_32074,N_32817);
or U33305 (N_33305,N_32486,N_32935);
or U33306 (N_33306,N_32261,N_32373);
xnor U33307 (N_33307,N_32118,N_32684);
and U33308 (N_33308,N_32132,N_32660);
nand U33309 (N_33309,N_32769,N_32741);
nand U33310 (N_33310,N_32510,N_32259);
or U33311 (N_33311,N_32296,N_32764);
nor U33312 (N_33312,N_32315,N_32617);
xor U33313 (N_33313,N_32242,N_32766);
nand U33314 (N_33314,N_32767,N_32388);
and U33315 (N_33315,N_32902,N_32904);
xnor U33316 (N_33316,N_32497,N_32816);
or U33317 (N_33317,N_32885,N_32906);
nand U33318 (N_33318,N_32453,N_32438);
xor U33319 (N_33319,N_32757,N_32015);
or U33320 (N_33320,N_32077,N_32480);
and U33321 (N_33321,N_32248,N_32323);
and U33322 (N_33322,N_32534,N_32998);
xnor U33323 (N_33323,N_32390,N_32152);
or U33324 (N_33324,N_32554,N_32555);
nand U33325 (N_33325,N_32760,N_32600);
xor U33326 (N_33326,N_32260,N_32509);
or U33327 (N_33327,N_32276,N_32939);
or U33328 (N_33328,N_32830,N_32883);
nand U33329 (N_33329,N_32171,N_32655);
and U33330 (N_33330,N_32597,N_32974);
xnor U33331 (N_33331,N_32174,N_32160);
nor U33332 (N_33332,N_32703,N_32964);
and U33333 (N_33333,N_32780,N_32724);
nand U33334 (N_33334,N_32126,N_32842);
xnor U33335 (N_33335,N_32274,N_32436);
nor U33336 (N_33336,N_32327,N_32092);
xor U33337 (N_33337,N_32527,N_32309);
nand U33338 (N_33338,N_32083,N_32018);
nand U33339 (N_33339,N_32089,N_32583);
xnor U33340 (N_33340,N_32090,N_32864);
nand U33341 (N_33341,N_32071,N_32947);
and U33342 (N_33342,N_32771,N_32619);
xor U33343 (N_33343,N_32470,N_32513);
nor U33344 (N_33344,N_32494,N_32755);
nor U33345 (N_33345,N_32936,N_32695);
nand U33346 (N_33346,N_32582,N_32728);
nand U33347 (N_33347,N_32643,N_32664);
and U33348 (N_33348,N_32244,N_32151);
and U33349 (N_33349,N_32391,N_32785);
xor U33350 (N_33350,N_32008,N_32422);
xnor U33351 (N_33351,N_32065,N_32051);
xor U33352 (N_33352,N_32616,N_32594);
or U33353 (N_33353,N_32811,N_32227);
nor U33354 (N_33354,N_32923,N_32284);
xnor U33355 (N_33355,N_32374,N_32967);
nand U33356 (N_33356,N_32446,N_32402);
nor U33357 (N_33357,N_32834,N_32458);
nor U33358 (N_33358,N_32825,N_32109);
xnor U33359 (N_33359,N_32010,N_32401);
nor U33360 (N_33360,N_32148,N_32698);
nand U33361 (N_33361,N_32361,N_32056);
or U33362 (N_33362,N_32185,N_32804);
nand U33363 (N_33363,N_32854,N_32787);
or U33364 (N_33364,N_32681,N_32061);
xor U33365 (N_33365,N_32654,N_32633);
nand U33366 (N_33366,N_32139,N_32195);
or U33367 (N_33367,N_32127,N_32561);
nor U33368 (N_33368,N_32958,N_32978);
nor U33369 (N_33369,N_32285,N_32631);
xnor U33370 (N_33370,N_32342,N_32806);
nor U33371 (N_33371,N_32545,N_32145);
nand U33372 (N_33372,N_32303,N_32014);
xor U33373 (N_33373,N_32937,N_32776);
and U33374 (N_33374,N_32218,N_32454);
and U33375 (N_33375,N_32125,N_32210);
nor U33376 (N_33376,N_32747,N_32424);
or U33377 (N_33377,N_32101,N_32469);
or U33378 (N_33378,N_32452,N_32416);
or U33379 (N_33379,N_32599,N_32930);
xnor U33380 (N_33380,N_32912,N_32568);
and U33381 (N_33381,N_32011,N_32123);
xnor U33382 (N_33382,N_32772,N_32700);
xor U33383 (N_33383,N_32624,N_32489);
nor U33384 (N_33384,N_32456,N_32844);
or U33385 (N_33385,N_32419,N_32336);
or U33386 (N_33386,N_32687,N_32307);
or U33387 (N_33387,N_32187,N_32668);
xor U33388 (N_33388,N_32797,N_32910);
xnor U33389 (N_33389,N_32165,N_32829);
nand U33390 (N_33390,N_32447,N_32961);
nor U33391 (N_33391,N_32770,N_32905);
and U33392 (N_33392,N_32823,N_32586);
nand U33393 (N_33393,N_32322,N_32501);
or U33394 (N_33394,N_32882,N_32793);
nor U33395 (N_33395,N_32966,N_32540);
nand U33396 (N_33396,N_32721,N_32827);
nand U33397 (N_33397,N_32679,N_32708);
xor U33398 (N_33398,N_32625,N_32376);
nor U33399 (N_33399,N_32483,N_32723);
nand U33400 (N_33400,N_32119,N_32822);
nand U33401 (N_33401,N_32394,N_32986);
xnor U33402 (N_33402,N_32184,N_32639);
or U33403 (N_33403,N_32202,N_32621);
or U33404 (N_33404,N_32084,N_32040);
nor U33405 (N_33405,N_32207,N_32492);
or U33406 (N_33406,N_32514,N_32427);
or U33407 (N_33407,N_32649,N_32722);
or U33408 (N_33408,N_32328,N_32378);
or U33409 (N_33409,N_32858,N_32648);
or U33410 (N_33410,N_32292,N_32878);
nor U33411 (N_33411,N_32241,N_32976);
xnor U33412 (N_33412,N_32794,N_32636);
xnor U33413 (N_33413,N_32055,N_32981);
xnor U33414 (N_33414,N_32894,N_32457);
nand U33415 (N_33415,N_32000,N_32558);
nor U33416 (N_33416,N_32048,N_32052);
and U33417 (N_33417,N_32953,N_32062);
xor U33418 (N_33418,N_32175,N_32987);
xnor U33419 (N_33419,N_32535,N_32567);
or U33420 (N_33420,N_32615,N_32608);
and U33421 (N_33421,N_32874,N_32879);
and U33422 (N_33422,N_32572,N_32970);
or U33423 (N_33423,N_32423,N_32214);
nor U33424 (N_33424,N_32333,N_32279);
or U33425 (N_33425,N_32573,N_32463);
xnor U33426 (N_33426,N_32663,N_32270);
or U33427 (N_33427,N_32341,N_32630);
nand U33428 (N_33428,N_32672,N_32877);
or U33429 (N_33429,N_32656,N_32862);
xnor U33430 (N_33430,N_32836,N_32181);
nor U33431 (N_33431,N_32738,N_32915);
nand U33432 (N_33432,N_32231,N_32839);
and U33433 (N_33433,N_32224,N_32733);
xnor U33434 (N_33434,N_32613,N_32909);
and U33435 (N_33435,N_32990,N_32948);
xor U33436 (N_33436,N_32372,N_32602);
xnor U33437 (N_33437,N_32895,N_32712);
or U33438 (N_33438,N_32980,N_32412);
or U33439 (N_33439,N_32893,N_32368);
or U33440 (N_33440,N_32330,N_32237);
nor U33441 (N_33441,N_32013,N_32399);
or U33442 (N_33442,N_32742,N_32026);
and U33443 (N_33443,N_32129,N_32875);
nand U33444 (N_33444,N_32319,N_32488);
nor U33445 (N_33445,N_32286,N_32377);
xnor U33446 (N_33446,N_32103,N_32479);
xor U33447 (N_33447,N_32945,N_32354);
or U33448 (N_33448,N_32938,N_32968);
xnor U33449 (N_33449,N_32045,N_32850);
or U33450 (N_33450,N_32278,N_32344);
xnor U33451 (N_33451,N_32088,N_32073);
nor U33452 (N_33452,N_32357,N_32183);
and U33453 (N_33453,N_32063,N_32209);
nand U33454 (N_33454,N_32159,N_32343);
and U33455 (N_33455,N_32598,N_32233);
or U33456 (N_33456,N_32709,N_32316);
xor U33457 (N_33457,N_32716,N_32198);
xor U33458 (N_33458,N_32869,N_32059);
and U33459 (N_33459,N_32795,N_32170);
and U33460 (N_33460,N_32756,N_32443);
and U33461 (N_33461,N_32253,N_32645);
nor U33462 (N_33462,N_32147,N_32768);
nor U33463 (N_33463,N_32182,N_32685);
and U33464 (N_33464,N_32601,N_32835);
xnor U33465 (N_33465,N_32068,N_32697);
nand U33466 (N_33466,N_32216,N_32840);
nand U33467 (N_33467,N_32166,N_32226);
xnor U33468 (N_33468,N_32280,N_32137);
and U33469 (N_33469,N_32871,N_32240);
xor U33470 (N_33470,N_32389,N_32786);
nand U33471 (N_33471,N_32570,N_32696);
and U33472 (N_33472,N_32477,N_32294);
xnor U33473 (N_33473,N_32271,N_32979);
or U33474 (N_33474,N_32133,N_32973);
xor U33475 (N_33475,N_32041,N_32383);
or U33476 (N_33476,N_32726,N_32914);
or U33477 (N_33477,N_32800,N_32016);
nor U33478 (N_33478,N_32856,N_32544);
nor U33479 (N_33479,N_32528,N_32743);
nand U33480 (N_33480,N_32369,N_32397);
xor U33481 (N_33481,N_32340,N_32623);
nand U33482 (N_33482,N_32082,N_32321);
xnor U33483 (N_33483,N_32140,N_32359);
or U33484 (N_33484,N_32934,N_32304);
nand U33485 (N_33485,N_32302,N_32299);
or U33486 (N_33486,N_32876,N_32537);
nor U33487 (N_33487,N_32791,N_32779);
nand U33488 (N_33488,N_32273,N_32678);
nand U33489 (N_33489,N_32153,N_32908);
and U33490 (N_33490,N_32855,N_32683);
or U33491 (N_33491,N_32670,N_32919);
xor U33492 (N_33492,N_32044,N_32522);
and U33493 (N_33493,N_32518,N_32969);
xnor U33494 (N_33494,N_32892,N_32706);
and U33495 (N_33495,N_32784,N_32191);
nand U33496 (N_33496,N_32511,N_32634);
xnor U33497 (N_33497,N_32692,N_32652);
xnor U33498 (N_33498,N_32821,N_32944);
or U33499 (N_33499,N_32832,N_32612);
nand U33500 (N_33500,N_32963,N_32882);
xor U33501 (N_33501,N_32350,N_32834);
and U33502 (N_33502,N_32821,N_32933);
nor U33503 (N_33503,N_32631,N_32577);
and U33504 (N_33504,N_32253,N_32546);
or U33505 (N_33505,N_32971,N_32123);
nor U33506 (N_33506,N_32795,N_32378);
or U33507 (N_33507,N_32817,N_32704);
nor U33508 (N_33508,N_32654,N_32897);
nor U33509 (N_33509,N_32461,N_32947);
nand U33510 (N_33510,N_32893,N_32477);
nand U33511 (N_33511,N_32706,N_32248);
xor U33512 (N_33512,N_32080,N_32150);
nor U33513 (N_33513,N_32570,N_32981);
nand U33514 (N_33514,N_32470,N_32118);
or U33515 (N_33515,N_32536,N_32041);
or U33516 (N_33516,N_32649,N_32516);
nand U33517 (N_33517,N_32095,N_32654);
or U33518 (N_33518,N_32254,N_32909);
xor U33519 (N_33519,N_32702,N_32780);
nor U33520 (N_33520,N_32987,N_32233);
nor U33521 (N_33521,N_32023,N_32824);
or U33522 (N_33522,N_32721,N_32577);
nor U33523 (N_33523,N_32327,N_32896);
xor U33524 (N_33524,N_32723,N_32529);
and U33525 (N_33525,N_32134,N_32156);
nand U33526 (N_33526,N_32889,N_32981);
nor U33527 (N_33527,N_32198,N_32903);
nor U33528 (N_33528,N_32731,N_32426);
xnor U33529 (N_33529,N_32070,N_32399);
and U33530 (N_33530,N_32681,N_32606);
xnor U33531 (N_33531,N_32532,N_32013);
and U33532 (N_33532,N_32810,N_32412);
nor U33533 (N_33533,N_32244,N_32525);
and U33534 (N_33534,N_32898,N_32243);
nor U33535 (N_33535,N_32890,N_32038);
and U33536 (N_33536,N_32579,N_32485);
xnor U33537 (N_33537,N_32093,N_32983);
nor U33538 (N_33538,N_32928,N_32274);
and U33539 (N_33539,N_32707,N_32897);
nand U33540 (N_33540,N_32771,N_32156);
nand U33541 (N_33541,N_32796,N_32661);
nand U33542 (N_33542,N_32413,N_32381);
and U33543 (N_33543,N_32012,N_32631);
nor U33544 (N_33544,N_32052,N_32070);
nand U33545 (N_33545,N_32261,N_32331);
and U33546 (N_33546,N_32777,N_32739);
or U33547 (N_33547,N_32535,N_32821);
or U33548 (N_33548,N_32658,N_32969);
nor U33549 (N_33549,N_32047,N_32868);
nand U33550 (N_33550,N_32740,N_32988);
and U33551 (N_33551,N_32306,N_32478);
and U33552 (N_33552,N_32146,N_32069);
and U33553 (N_33553,N_32374,N_32902);
and U33554 (N_33554,N_32497,N_32951);
xnor U33555 (N_33555,N_32477,N_32591);
or U33556 (N_33556,N_32782,N_32928);
xnor U33557 (N_33557,N_32563,N_32138);
xnor U33558 (N_33558,N_32115,N_32449);
or U33559 (N_33559,N_32757,N_32551);
xnor U33560 (N_33560,N_32081,N_32181);
xnor U33561 (N_33561,N_32495,N_32903);
nand U33562 (N_33562,N_32283,N_32476);
or U33563 (N_33563,N_32984,N_32920);
and U33564 (N_33564,N_32658,N_32403);
xnor U33565 (N_33565,N_32120,N_32992);
nand U33566 (N_33566,N_32793,N_32985);
nor U33567 (N_33567,N_32304,N_32155);
xor U33568 (N_33568,N_32175,N_32895);
and U33569 (N_33569,N_32362,N_32759);
nor U33570 (N_33570,N_32711,N_32338);
nand U33571 (N_33571,N_32640,N_32817);
and U33572 (N_33572,N_32641,N_32879);
xor U33573 (N_33573,N_32965,N_32443);
and U33574 (N_33574,N_32597,N_32342);
nand U33575 (N_33575,N_32166,N_32273);
and U33576 (N_33576,N_32576,N_32725);
or U33577 (N_33577,N_32149,N_32903);
and U33578 (N_33578,N_32927,N_32375);
and U33579 (N_33579,N_32147,N_32540);
and U33580 (N_33580,N_32852,N_32105);
and U33581 (N_33581,N_32744,N_32347);
xor U33582 (N_33582,N_32878,N_32686);
xor U33583 (N_33583,N_32050,N_32786);
and U33584 (N_33584,N_32929,N_32663);
or U33585 (N_33585,N_32982,N_32828);
and U33586 (N_33586,N_32079,N_32817);
or U33587 (N_33587,N_32263,N_32782);
and U33588 (N_33588,N_32546,N_32583);
xnor U33589 (N_33589,N_32810,N_32657);
xnor U33590 (N_33590,N_32235,N_32195);
xor U33591 (N_33591,N_32229,N_32416);
nand U33592 (N_33592,N_32329,N_32855);
nor U33593 (N_33593,N_32041,N_32193);
or U33594 (N_33594,N_32181,N_32678);
and U33595 (N_33595,N_32652,N_32376);
nand U33596 (N_33596,N_32960,N_32264);
nand U33597 (N_33597,N_32245,N_32891);
xor U33598 (N_33598,N_32928,N_32852);
or U33599 (N_33599,N_32604,N_32211);
nor U33600 (N_33600,N_32541,N_32190);
nand U33601 (N_33601,N_32481,N_32952);
nor U33602 (N_33602,N_32742,N_32532);
nor U33603 (N_33603,N_32240,N_32622);
nor U33604 (N_33604,N_32450,N_32007);
and U33605 (N_33605,N_32019,N_32128);
xor U33606 (N_33606,N_32719,N_32637);
nand U33607 (N_33607,N_32795,N_32004);
xor U33608 (N_33608,N_32307,N_32674);
and U33609 (N_33609,N_32368,N_32116);
or U33610 (N_33610,N_32234,N_32797);
and U33611 (N_33611,N_32823,N_32843);
xor U33612 (N_33612,N_32431,N_32194);
nor U33613 (N_33613,N_32715,N_32633);
nand U33614 (N_33614,N_32985,N_32483);
and U33615 (N_33615,N_32062,N_32170);
and U33616 (N_33616,N_32853,N_32711);
and U33617 (N_33617,N_32558,N_32094);
xnor U33618 (N_33618,N_32647,N_32158);
xor U33619 (N_33619,N_32459,N_32946);
xnor U33620 (N_33620,N_32207,N_32614);
nand U33621 (N_33621,N_32034,N_32714);
nor U33622 (N_33622,N_32179,N_32959);
xor U33623 (N_33623,N_32633,N_32854);
xor U33624 (N_33624,N_32156,N_32516);
xnor U33625 (N_33625,N_32592,N_32057);
and U33626 (N_33626,N_32494,N_32974);
xnor U33627 (N_33627,N_32151,N_32088);
nor U33628 (N_33628,N_32690,N_32626);
xnor U33629 (N_33629,N_32054,N_32585);
and U33630 (N_33630,N_32185,N_32229);
or U33631 (N_33631,N_32988,N_32631);
or U33632 (N_33632,N_32185,N_32624);
nand U33633 (N_33633,N_32943,N_32676);
xnor U33634 (N_33634,N_32339,N_32736);
nand U33635 (N_33635,N_32775,N_32588);
or U33636 (N_33636,N_32054,N_32607);
or U33637 (N_33637,N_32307,N_32165);
nand U33638 (N_33638,N_32176,N_32747);
xnor U33639 (N_33639,N_32577,N_32064);
and U33640 (N_33640,N_32800,N_32333);
nand U33641 (N_33641,N_32608,N_32857);
and U33642 (N_33642,N_32182,N_32839);
nand U33643 (N_33643,N_32966,N_32004);
nand U33644 (N_33644,N_32099,N_32059);
or U33645 (N_33645,N_32832,N_32672);
xnor U33646 (N_33646,N_32862,N_32966);
and U33647 (N_33647,N_32305,N_32120);
or U33648 (N_33648,N_32021,N_32336);
xnor U33649 (N_33649,N_32568,N_32893);
and U33650 (N_33650,N_32344,N_32942);
nor U33651 (N_33651,N_32534,N_32266);
and U33652 (N_33652,N_32133,N_32901);
or U33653 (N_33653,N_32836,N_32747);
xor U33654 (N_33654,N_32309,N_32933);
nor U33655 (N_33655,N_32537,N_32237);
xor U33656 (N_33656,N_32193,N_32314);
and U33657 (N_33657,N_32884,N_32981);
nand U33658 (N_33658,N_32982,N_32133);
nor U33659 (N_33659,N_32461,N_32590);
nand U33660 (N_33660,N_32370,N_32007);
nor U33661 (N_33661,N_32729,N_32659);
or U33662 (N_33662,N_32715,N_32616);
and U33663 (N_33663,N_32587,N_32043);
xor U33664 (N_33664,N_32817,N_32270);
or U33665 (N_33665,N_32929,N_32137);
xnor U33666 (N_33666,N_32679,N_32189);
and U33667 (N_33667,N_32798,N_32522);
and U33668 (N_33668,N_32180,N_32054);
xnor U33669 (N_33669,N_32070,N_32475);
and U33670 (N_33670,N_32323,N_32048);
xor U33671 (N_33671,N_32969,N_32060);
nor U33672 (N_33672,N_32065,N_32761);
xor U33673 (N_33673,N_32142,N_32039);
and U33674 (N_33674,N_32726,N_32214);
xor U33675 (N_33675,N_32004,N_32463);
and U33676 (N_33676,N_32912,N_32804);
nor U33677 (N_33677,N_32734,N_32206);
nor U33678 (N_33678,N_32001,N_32529);
nand U33679 (N_33679,N_32912,N_32462);
xnor U33680 (N_33680,N_32912,N_32776);
and U33681 (N_33681,N_32965,N_32926);
and U33682 (N_33682,N_32973,N_32152);
xnor U33683 (N_33683,N_32805,N_32453);
xor U33684 (N_33684,N_32196,N_32992);
xnor U33685 (N_33685,N_32827,N_32236);
or U33686 (N_33686,N_32043,N_32450);
xnor U33687 (N_33687,N_32463,N_32191);
or U33688 (N_33688,N_32019,N_32852);
nor U33689 (N_33689,N_32621,N_32417);
and U33690 (N_33690,N_32758,N_32789);
and U33691 (N_33691,N_32581,N_32908);
xor U33692 (N_33692,N_32373,N_32082);
nand U33693 (N_33693,N_32227,N_32098);
or U33694 (N_33694,N_32790,N_32250);
xor U33695 (N_33695,N_32060,N_32430);
nor U33696 (N_33696,N_32289,N_32368);
or U33697 (N_33697,N_32297,N_32500);
xor U33698 (N_33698,N_32987,N_32060);
nor U33699 (N_33699,N_32330,N_32636);
nand U33700 (N_33700,N_32759,N_32944);
nand U33701 (N_33701,N_32406,N_32177);
or U33702 (N_33702,N_32778,N_32519);
or U33703 (N_33703,N_32359,N_32342);
or U33704 (N_33704,N_32931,N_32301);
or U33705 (N_33705,N_32959,N_32300);
xor U33706 (N_33706,N_32283,N_32360);
xor U33707 (N_33707,N_32587,N_32290);
xnor U33708 (N_33708,N_32960,N_32104);
nand U33709 (N_33709,N_32959,N_32068);
or U33710 (N_33710,N_32130,N_32372);
nand U33711 (N_33711,N_32624,N_32432);
nand U33712 (N_33712,N_32807,N_32425);
or U33713 (N_33713,N_32588,N_32598);
nor U33714 (N_33714,N_32277,N_32439);
xor U33715 (N_33715,N_32401,N_32648);
and U33716 (N_33716,N_32039,N_32032);
nand U33717 (N_33717,N_32729,N_32885);
or U33718 (N_33718,N_32015,N_32643);
or U33719 (N_33719,N_32424,N_32425);
xor U33720 (N_33720,N_32428,N_32330);
or U33721 (N_33721,N_32397,N_32686);
and U33722 (N_33722,N_32785,N_32187);
and U33723 (N_33723,N_32707,N_32649);
and U33724 (N_33724,N_32626,N_32854);
or U33725 (N_33725,N_32441,N_32189);
or U33726 (N_33726,N_32929,N_32421);
or U33727 (N_33727,N_32103,N_32738);
nor U33728 (N_33728,N_32591,N_32071);
and U33729 (N_33729,N_32586,N_32410);
nand U33730 (N_33730,N_32508,N_32891);
nand U33731 (N_33731,N_32540,N_32971);
nand U33732 (N_33732,N_32950,N_32881);
xnor U33733 (N_33733,N_32046,N_32132);
nor U33734 (N_33734,N_32290,N_32397);
xor U33735 (N_33735,N_32253,N_32651);
or U33736 (N_33736,N_32304,N_32803);
and U33737 (N_33737,N_32295,N_32433);
nand U33738 (N_33738,N_32075,N_32507);
nor U33739 (N_33739,N_32026,N_32291);
nor U33740 (N_33740,N_32364,N_32024);
xor U33741 (N_33741,N_32965,N_32922);
nand U33742 (N_33742,N_32300,N_32689);
or U33743 (N_33743,N_32615,N_32944);
nor U33744 (N_33744,N_32764,N_32829);
xnor U33745 (N_33745,N_32699,N_32377);
nor U33746 (N_33746,N_32738,N_32374);
nand U33747 (N_33747,N_32923,N_32617);
xnor U33748 (N_33748,N_32269,N_32761);
xor U33749 (N_33749,N_32223,N_32405);
or U33750 (N_33750,N_32802,N_32953);
xnor U33751 (N_33751,N_32094,N_32937);
and U33752 (N_33752,N_32174,N_32711);
and U33753 (N_33753,N_32139,N_32569);
and U33754 (N_33754,N_32524,N_32909);
or U33755 (N_33755,N_32281,N_32304);
nor U33756 (N_33756,N_32083,N_32632);
and U33757 (N_33757,N_32538,N_32796);
nand U33758 (N_33758,N_32849,N_32755);
xnor U33759 (N_33759,N_32566,N_32886);
or U33760 (N_33760,N_32408,N_32870);
xor U33761 (N_33761,N_32639,N_32562);
or U33762 (N_33762,N_32359,N_32263);
xnor U33763 (N_33763,N_32994,N_32570);
xnor U33764 (N_33764,N_32824,N_32529);
or U33765 (N_33765,N_32366,N_32461);
nand U33766 (N_33766,N_32495,N_32588);
nand U33767 (N_33767,N_32162,N_32749);
and U33768 (N_33768,N_32739,N_32414);
and U33769 (N_33769,N_32510,N_32084);
and U33770 (N_33770,N_32526,N_32654);
xor U33771 (N_33771,N_32221,N_32467);
and U33772 (N_33772,N_32717,N_32624);
nor U33773 (N_33773,N_32073,N_32353);
nand U33774 (N_33774,N_32355,N_32671);
xnor U33775 (N_33775,N_32739,N_32160);
nor U33776 (N_33776,N_32410,N_32371);
xnor U33777 (N_33777,N_32551,N_32827);
or U33778 (N_33778,N_32602,N_32257);
nand U33779 (N_33779,N_32040,N_32707);
nor U33780 (N_33780,N_32565,N_32854);
and U33781 (N_33781,N_32605,N_32898);
or U33782 (N_33782,N_32851,N_32001);
nand U33783 (N_33783,N_32259,N_32880);
nand U33784 (N_33784,N_32073,N_32523);
nand U33785 (N_33785,N_32988,N_32724);
or U33786 (N_33786,N_32740,N_32219);
and U33787 (N_33787,N_32416,N_32260);
nor U33788 (N_33788,N_32319,N_32469);
xor U33789 (N_33789,N_32826,N_32819);
and U33790 (N_33790,N_32817,N_32964);
xnor U33791 (N_33791,N_32445,N_32800);
xor U33792 (N_33792,N_32245,N_32631);
nand U33793 (N_33793,N_32444,N_32011);
nand U33794 (N_33794,N_32570,N_32333);
or U33795 (N_33795,N_32094,N_32193);
nor U33796 (N_33796,N_32587,N_32317);
nor U33797 (N_33797,N_32730,N_32330);
nand U33798 (N_33798,N_32716,N_32279);
xor U33799 (N_33799,N_32197,N_32732);
nand U33800 (N_33800,N_32964,N_32913);
xnor U33801 (N_33801,N_32742,N_32710);
nor U33802 (N_33802,N_32398,N_32502);
or U33803 (N_33803,N_32777,N_32107);
xnor U33804 (N_33804,N_32269,N_32497);
xor U33805 (N_33805,N_32007,N_32883);
nand U33806 (N_33806,N_32635,N_32201);
nand U33807 (N_33807,N_32408,N_32004);
or U33808 (N_33808,N_32669,N_32148);
nor U33809 (N_33809,N_32543,N_32424);
or U33810 (N_33810,N_32248,N_32945);
nand U33811 (N_33811,N_32157,N_32679);
or U33812 (N_33812,N_32646,N_32557);
xor U33813 (N_33813,N_32700,N_32066);
nand U33814 (N_33814,N_32323,N_32774);
xnor U33815 (N_33815,N_32848,N_32862);
nor U33816 (N_33816,N_32295,N_32132);
nor U33817 (N_33817,N_32828,N_32090);
and U33818 (N_33818,N_32570,N_32562);
xnor U33819 (N_33819,N_32700,N_32338);
or U33820 (N_33820,N_32943,N_32521);
and U33821 (N_33821,N_32086,N_32169);
nor U33822 (N_33822,N_32864,N_32495);
and U33823 (N_33823,N_32757,N_32059);
or U33824 (N_33824,N_32720,N_32998);
nor U33825 (N_33825,N_32808,N_32608);
and U33826 (N_33826,N_32254,N_32982);
xor U33827 (N_33827,N_32994,N_32396);
nand U33828 (N_33828,N_32602,N_32778);
nand U33829 (N_33829,N_32570,N_32453);
nand U33830 (N_33830,N_32283,N_32273);
or U33831 (N_33831,N_32695,N_32985);
and U33832 (N_33832,N_32696,N_32410);
nand U33833 (N_33833,N_32158,N_32342);
nand U33834 (N_33834,N_32122,N_32960);
or U33835 (N_33835,N_32768,N_32259);
nand U33836 (N_33836,N_32406,N_32759);
nor U33837 (N_33837,N_32196,N_32603);
nand U33838 (N_33838,N_32087,N_32184);
and U33839 (N_33839,N_32525,N_32963);
and U33840 (N_33840,N_32852,N_32079);
or U33841 (N_33841,N_32406,N_32407);
nor U33842 (N_33842,N_32901,N_32402);
nor U33843 (N_33843,N_32399,N_32695);
nor U33844 (N_33844,N_32141,N_32304);
nor U33845 (N_33845,N_32027,N_32280);
or U33846 (N_33846,N_32264,N_32155);
xor U33847 (N_33847,N_32211,N_32057);
xnor U33848 (N_33848,N_32115,N_32451);
nor U33849 (N_33849,N_32738,N_32994);
nand U33850 (N_33850,N_32241,N_32424);
xor U33851 (N_33851,N_32271,N_32343);
nand U33852 (N_33852,N_32457,N_32706);
nand U33853 (N_33853,N_32408,N_32571);
or U33854 (N_33854,N_32513,N_32186);
or U33855 (N_33855,N_32800,N_32458);
xor U33856 (N_33856,N_32925,N_32177);
nor U33857 (N_33857,N_32993,N_32274);
or U33858 (N_33858,N_32180,N_32922);
xor U33859 (N_33859,N_32774,N_32027);
and U33860 (N_33860,N_32210,N_32247);
and U33861 (N_33861,N_32243,N_32009);
xnor U33862 (N_33862,N_32622,N_32720);
and U33863 (N_33863,N_32668,N_32576);
xnor U33864 (N_33864,N_32311,N_32259);
or U33865 (N_33865,N_32279,N_32135);
xnor U33866 (N_33866,N_32358,N_32631);
nand U33867 (N_33867,N_32417,N_32897);
nand U33868 (N_33868,N_32314,N_32896);
or U33869 (N_33869,N_32302,N_32660);
nand U33870 (N_33870,N_32331,N_32829);
nor U33871 (N_33871,N_32606,N_32380);
nor U33872 (N_33872,N_32074,N_32192);
or U33873 (N_33873,N_32992,N_32743);
xnor U33874 (N_33874,N_32889,N_32123);
or U33875 (N_33875,N_32652,N_32325);
and U33876 (N_33876,N_32658,N_32360);
nor U33877 (N_33877,N_32066,N_32031);
nor U33878 (N_33878,N_32309,N_32500);
xnor U33879 (N_33879,N_32738,N_32569);
and U33880 (N_33880,N_32130,N_32588);
and U33881 (N_33881,N_32785,N_32472);
and U33882 (N_33882,N_32012,N_32086);
xnor U33883 (N_33883,N_32669,N_32845);
nand U33884 (N_33884,N_32041,N_32164);
nand U33885 (N_33885,N_32061,N_32526);
or U33886 (N_33886,N_32033,N_32507);
xor U33887 (N_33887,N_32203,N_32989);
and U33888 (N_33888,N_32978,N_32755);
nand U33889 (N_33889,N_32424,N_32510);
or U33890 (N_33890,N_32897,N_32644);
nor U33891 (N_33891,N_32320,N_32913);
and U33892 (N_33892,N_32895,N_32308);
nor U33893 (N_33893,N_32990,N_32047);
or U33894 (N_33894,N_32664,N_32750);
xnor U33895 (N_33895,N_32411,N_32286);
and U33896 (N_33896,N_32069,N_32804);
nor U33897 (N_33897,N_32767,N_32216);
or U33898 (N_33898,N_32096,N_32519);
nor U33899 (N_33899,N_32300,N_32807);
or U33900 (N_33900,N_32439,N_32950);
and U33901 (N_33901,N_32760,N_32005);
nand U33902 (N_33902,N_32224,N_32766);
nand U33903 (N_33903,N_32406,N_32615);
nor U33904 (N_33904,N_32729,N_32649);
xor U33905 (N_33905,N_32757,N_32690);
nor U33906 (N_33906,N_32968,N_32964);
nand U33907 (N_33907,N_32322,N_32268);
nand U33908 (N_33908,N_32858,N_32758);
nand U33909 (N_33909,N_32286,N_32991);
and U33910 (N_33910,N_32630,N_32891);
nor U33911 (N_33911,N_32251,N_32838);
and U33912 (N_33912,N_32105,N_32287);
nor U33913 (N_33913,N_32856,N_32129);
xnor U33914 (N_33914,N_32071,N_32868);
xor U33915 (N_33915,N_32564,N_32703);
or U33916 (N_33916,N_32025,N_32814);
and U33917 (N_33917,N_32339,N_32165);
and U33918 (N_33918,N_32327,N_32782);
or U33919 (N_33919,N_32383,N_32205);
xnor U33920 (N_33920,N_32572,N_32125);
nor U33921 (N_33921,N_32536,N_32387);
and U33922 (N_33922,N_32763,N_32940);
and U33923 (N_33923,N_32634,N_32885);
nor U33924 (N_33924,N_32062,N_32400);
nor U33925 (N_33925,N_32357,N_32005);
and U33926 (N_33926,N_32318,N_32955);
nand U33927 (N_33927,N_32500,N_32539);
nand U33928 (N_33928,N_32510,N_32715);
nor U33929 (N_33929,N_32232,N_32492);
nor U33930 (N_33930,N_32796,N_32481);
and U33931 (N_33931,N_32382,N_32708);
nand U33932 (N_33932,N_32860,N_32513);
nor U33933 (N_33933,N_32572,N_32936);
xnor U33934 (N_33934,N_32418,N_32389);
or U33935 (N_33935,N_32079,N_32844);
xnor U33936 (N_33936,N_32476,N_32360);
nor U33937 (N_33937,N_32616,N_32216);
and U33938 (N_33938,N_32420,N_32196);
and U33939 (N_33939,N_32879,N_32498);
or U33940 (N_33940,N_32853,N_32315);
or U33941 (N_33941,N_32087,N_32709);
nor U33942 (N_33942,N_32004,N_32213);
and U33943 (N_33943,N_32216,N_32523);
and U33944 (N_33944,N_32416,N_32034);
or U33945 (N_33945,N_32669,N_32497);
xor U33946 (N_33946,N_32779,N_32352);
or U33947 (N_33947,N_32567,N_32362);
or U33948 (N_33948,N_32057,N_32849);
nor U33949 (N_33949,N_32403,N_32822);
xnor U33950 (N_33950,N_32803,N_32988);
nor U33951 (N_33951,N_32405,N_32698);
and U33952 (N_33952,N_32245,N_32868);
nand U33953 (N_33953,N_32471,N_32543);
xnor U33954 (N_33954,N_32681,N_32648);
and U33955 (N_33955,N_32353,N_32946);
xor U33956 (N_33956,N_32150,N_32712);
xnor U33957 (N_33957,N_32712,N_32597);
nand U33958 (N_33958,N_32289,N_32814);
nor U33959 (N_33959,N_32610,N_32660);
and U33960 (N_33960,N_32851,N_32444);
or U33961 (N_33961,N_32667,N_32974);
nand U33962 (N_33962,N_32494,N_32108);
nor U33963 (N_33963,N_32410,N_32160);
xor U33964 (N_33964,N_32506,N_32360);
nor U33965 (N_33965,N_32923,N_32084);
xor U33966 (N_33966,N_32861,N_32025);
nor U33967 (N_33967,N_32622,N_32935);
nor U33968 (N_33968,N_32571,N_32657);
nand U33969 (N_33969,N_32109,N_32454);
and U33970 (N_33970,N_32937,N_32389);
nor U33971 (N_33971,N_32048,N_32784);
nor U33972 (N_33972,N_32562,N_32797);
nand U33973 (N_33973,N_32829,N_32125);
and U33974 (N_33974,N_32397,N_32612);
and U33975 (N_33975,N_32548,N_32835);
or U33976 (N_33976,N_32412,N_32489);
xnor U33977 (N_33977,N_32706,N_32427);
nor U33978 (N_33978,N_32918,N_32661);
and U33979 (N_33979,N_32831,N_32817);
nor U33980 (N_33980,N_32167,N_32853);
xnor U33981 (N_33981,N_32643,N_32238);
nand U33982 (N_33982,N_32479,N_32171);
or U33983 (N_33983,N_32105,N_32129);
nand U33984 (N_33984,N_32348,N_32843);
xnor U33985 (N_33985,N_32731,N_32734);
and U33986 (N_33986,N_32256,N_32901);
nand U33987 (N_33987,N_32050,N_32325);
and U33988 (N_33988,N_32874,N_32027);
xor U33989 (N_33989,N_32952,N_32120);
and U33990 (N_33990,N_32756,N_32841);
xnor U33991 (N_33991,N_32867,N_32030);
xor U33992 (N_33992,N_32272,N_32441);
nand U33993 (N_33993,N_32486,N_32537);
nor U33994 (N_33994,N_32526,N_32635);
nor U33995 (N_33995,N_32960,N_32925);
xnor U33996 (N_33996,N_32962,N_32642);
nand U33997 (N_33997,N_32614,N_32212);
and U33998 (N_33998,N_32700,N_32388);
xnor U33999 (N_33999,N_32721,N_32355);
or U34000 (N_34000,N_33959,N_33036);
xnor U34001 (N_34001,N_33958,N_33520);
and U34002 (N_34002,N_33667,N_33688);
nand U34003 (N_34003,N_33917,N_33945);
and U34004 (N_34004,N_33042,N_33185);
xnor U34005 (N_34005,N_33724,N_33478);
nand U34006 (N_34006,N_33481,N_33912);
or U34007 (N_34007,N_33795,N_33980);
nand U34008 (N_34008,N_33691,N_33549);
nor U34009 (N_34009,N_33944,N_33129);
nor U34010 (N_34010,N_33551,N_33940);
nand U34011 (N_34011,N_33321,N_33438);
nand U34012 (N_34012,N_33843,N_33697);
or U34013 (N_34013,N_33661,N_33953);
and U34014 (N_34014,N_33493,N_33911);
nor U34015 (N_34015,N_33647,N_33238);
and U34016 (N_34016,N_33791,N_33543);
nand U34017 (N_34017,N_33556,N_33573);
xor U34018 (N_34018,N_33487,N_33417);
nand U34019 (N_34019,N_33152,N_33369);
nor U34020 (N_34020,N_33637,N_33390);
and U34021 (N_34021,N_33279,N_33705);
xnor U34022 (N_34022,N_33222,N_33502);
nor U34023 (N_34023,N_33995,N_33351);
and U34024 (N_34024,N_33357,N_33726);
nor U34025 (N_34025,N_33905,N_33656);
and U34026 (N_34026,N_33847,N_33579);
xnor U34027 (N_34027,N_33160,N_33437);
nand U34028 (N_34028,N_33739,N_33400);
xor U34029 (N_34029,N_33224,N_33327);
nand U34030 (N_34030,N_33654,N_33055);
or U34031 (N_34031,N_33054,N_33641);
nand U34032 (N_34032,N_33996,N_33646);
or U34033 (N_34033,N_33028,N_33061);
and U34034 (N_34034,N_33069,N_33193);
and U34035 (N_34035,N_33132,N_33283);
and U34036 (N_34036,N_33013,N_33367);
nor U34037 (N_34037,N_33976,N_33902);
or U34038 (N_34038,N_33602,N_33049);
nor U34039 (N_34039,N_33232,N_33931);
nand U34040 (N_34040,N_33259,N_33806);
or U34041 (N_34041,N_33308,N_33883);
nor U34042 (N_34042,N_33348,N_33865);
nor U34043 (N_34043,N_33825,N_33627);
or U34044 (N_34044,N_33001,N_33058);
and U34045 (N_34045,N_33457,N_33335);
xnor U34046 (N_34046,N_33267,N_33601);
nand U34047 (N_34047,N_33532,N_33972);
nor U34048 (N_34048,N_33141,N_33153);
nand U34049 (N_34049,N_33639,N_33422);
nor U34050 (N_34050,N_33057,N_33219);
nand U34051 (N_34051,N_33137,N_33799);
xor U34052 (N_34052,N_33901,N_33146);
or U34053 (N_34053,N_33459,N_33398);
or U34054 (N_34054,N_33827,N_33067);
nor U34055 (N_34055,N_33625,N_33612);
or U34056 (N_34056,N_33519,N_33017);
nor U34057 (N_34057,N_33112,N_33251);
xor U34058 (N_34058,N_33288,N_33529);
nor U34059 (N_34059,N_33712,N_33167);
and U34060 (N_34060,N_33758,N_33298);
or U34061 (N_34061,N_33109,N_33614);
nand U34062 (N_34062,N_33033,N_33361);
nor U34063 (N_34063,N_33441,N_33266);
and U34064 (N_34064,N_33908,N_33040);
or U34065 (N_34065,N_33622,N_33087);
nor U34066 (N_34066,N_33031,N_33411);
nor U34067 (N_34067,N_33164,N_33515);
and U34068 (N_34068,N_33766,N_33926);
and U34069 (N_34069,N_33938,N_33347);
nand U34070 (N_34070,N_33702,N_33096);
or U34071 (N_34071,N_33964,N_33518);
and U34072 (N_34072,N_33056,N_33870);
or U34073 (N_34073,N_33135,N_33690);
nand U34074 (N_34074,N_33730,N_33858);
and U34075 (N_34075,N_33815,N_33787);
and U34076 (N_34076,N_33019,N_33133);
nand U34077 (N_34077,N_33854,N_33504);
nor U34078 (N_34078,N_33618,N_33273);
and U34079 (N_34079,N_33919,N_33672);
and U34080 (N_34080,N_33605,N_33254);
or U34081 (N_34081,N_33371,N_33820);
xnor U34082 (N_34082,N_33342,N_33247);
or U34083 (N_34083,N_33760,N_33391);
xnor U34084 (N_34084,N_33047,N_33203);
nand U34085 (N_34085,N_33703,N_33158);
nor U34086 (N_34086,N_33184,N_33068);
or U34087 (N_34087,N_33215,N_33468);
or U34088 (N_34088,N_33349,N_33638);
and U34089 (N_34089,N_33377,N_33981);
nor U34090 (N_34090,N_33150,N_33440);
nor U34091 (N_34091,N_33966,N_33253);
and U34092 (N_34092,N_33101,N_33256);
nand U34093 (N_34093,N_33530,N_33053);
nand U34094 (N_34094,N_33894,N_33838);
or U34095 (N_34095,N_33803,N_33707);
or U34096 (N_34096,N_33380,N_33754);
and U34097 (N_34097,N_33269,N_33932);
or U34098 (N_34098,N_33145,N_33263);
or U34099 (N_34099,N_33234,N_33379);
and U34100 (N_34100,N_33116,N_33781);
nor U34101 (N_34101,N_33965,N_33542);
nand U34102 (N_34102,N_33951,N_33334);
or U34103 (N_34103,N_33075,N_33466);
or U34104 (N_34104,N_33686,N_33824);
and U34105 (N_34105,N_33546,N_33372);
xnor U34106 (N_34106,N_33503,N_33793);
or U34107 (N_34107,N_33078,N_33217);
nor U34108 (N_34108,N_33406,N_33859);
xnor U34109 (N_34109,N_33114,N_33500);
xnor U34110 (N_34110,N_33695,N_33428);
and U34111 (N_34111,N_33170,N_33201);
and U34112 (N_34112,N_33626,N_33678);
nor U34113 (N_34113,N_33063,N_33378);
or U34114 (N_34114,N_33252,N_33445);
and U34115 (N_34115,N_33734,N_33942);
and U34116 (N_34116,N_33018,N_33986);
nor U34117 (N_34117,N_33125,N_33420);
nor U34118 (N_34118,N_33014,N_33143);
and U34119 (N_34119,N_33607,N_33552);
or U34120 (N_34120,N_33444,N_33740);
and U34121 (N_34121,N_33590,N_33257);
or U34122 (N_34122,N_33842,N_33363);
or U34123 (N_34123,N_33623,N_33002);
or U34124 (N_34124,N_33861,N_33448);
or U34125 (N_34125,N_33709,N_33665);
and U34126 (N_34126,N_33452,N_33316);
nor U34127 (N_34127,N_33241,N_33844);
and U34128 (N_34128,N_33093,N_33589);
or U34129 (N_34129,N_33421,N_33115);
and U34130 (N_34130,N_33855,N_33370);
xor U34131 (N_34131,N_33020,N_33818);
and U34132 (N_34132,N_33717,N_33175);
xor U34133 (N_34133,N_33154,N_33299);
nor U34134 (N_34134,N_33302,N_33447);
nand U34135 (N_34135,N_33650,N_33489);
nand U34136 (N_34136,N_33325,N_33933);
or U34137 (N_34137,N_33710,N_33197);
nor U34138 (N_34138,N_33648,N_33821);
xor U34139 (N_34139,N_33867,N_33628);
nor U34140 (N_34140,N_33236,N_33742);
xnor U34141 (N_34141,N_33807,N_33248);
xor U34142 (N_34142,N_33041,N_33523);
nor U34143 (N_34143,N_33609,N_33365);
nand U34144 (N_34144,N_33169,N_33122);
or U34145 (N_34145,N_33220,N_33786);
nand U34146 (N_34146,N_33613,N_33830);
or U34147 (N_34147,N_33458,N_33831);
nor U34148 (N_34148,N_33097,N_33282);
or U34149 (N_34149,N_33578,N_33330);
xor U34150 (N_34150,N_33679,N_33011);
and U34151 (N_34151,N_33998,N_33025);
xnor U34152 (N_34152,N_33209,N_33584);
and U34153 (N_34153,N_33508,N_33591);
nor U34154 (N_34154,N_33166,N_33183);
nand U34155 (N_34155,N_33410,N_33255);
xnor U34156 (N_34156,N_33872,N_33762);
nor U34157 (N_34157,N_33332,N_33425);
and U34158 (N_34158,N_33599,N_33923);
and U34159 (N_34159,N_33927,N_33239);
nor U34160 (N_34160,N_33967,N_33585);
or U34161 (N_34161,N_33675,N_33176);
or U34162 (N_34162,N_33687,N_33943);
xnor U34163 (N_34163,N_33443,N_33271);
or U34164 (N_34164,N_33205,N_33937);
nand U34165 (N_34165,N_33403,N_33700);
xnor U34166 (N_34166,N_33840,N_33513);
xnor U34167 (N_34167,N_33208,N_33317);
xnor U34168 (N_34168,N_33890,N_33524);
nor U34169 (N_34169,N_33083,N_33533);
nand U34170 (N_34170,N_33566,N_33670);
nor U34171 (N_34171,N_33326,N_33381);
and U34172 (N_34172,N_33027,N_33461);
xor U34173 (N_34173,N_33889,N_33262);
and U34174 (N_34174,N_33356,N_33906);
and U34175 (N_34175,N_33582,N_33849);
nor U34176 (N_34176,N_33698,N_33879);
xnor U34177 (N_34177,N_33449,N_33021);
nand U34178 (N_34178,N_33322,N_33435);
nand U34179 (N_34179,N_33065,N_33505);
or U34180 (N_34180,N_33388,N_33539);
nand U34181 (N_34181,N_33303,N_33396);
nor U34182 (N_34182,N_33869,N_33721);
xor U34183 (N_34183,N_33059,N_33072);
or U34184 (N_34184,N_33290,N_33352);
nor U34185 (N_34185,N_33727,N_33113);
nand U34186 (N_34186,N_33293,N_33716);
nor U34187 (N_34187,N_33752,N_33473);
nor U34188 (N_34188,N_33106,N_33202);
xnor U34189 (N_34189,N_33817,N_33231);
nor U34190 (N_34190,N_33948,N_33856);
or U34191 (N_34191,N_33026,N_33774);
nand U34192 (N_34192,N_33694,N_33392);
nor U34193 (N_34193,N_33947,N_33264);
nand U34194 (N_34194,N_33200,N_33887);
nand U34195 (N_34195,N_33826,N_33431);
nand U34196 (N_34196,N_33358,N_33659);
nand U34197 (N_34197,N_33198,N_33778);
xnor U34198 (N_34198,N_33402,N_33460);
nand U34199 (N_34199,N_33767,N_33472);
and U34200 (N_34200,N_33527,N_33603);
and U34201 (N_34201,N_33009,N_33899);
and U34202 (N_34202,N_33066,N_33593);
nand U34203 (N_34203,N_33975,N_33029);
nor U34204 (N_34204,N_33822,N_33353);
and U34205 (N_34205,N_33368,N_33857);
or U34206 (N_34206,N_33194,N_33492);
nand U34207 (N_34207,N_33880,N_33233);
nand U34208 (N_34208,N_33569,N_33914);
xor U34209 (N_34209,N_33973,N_33415);
xnor U34210 (N_34210,N_33120,N_33761);
or U34211 (N_34211,N_33676,N_33276);
nor U34212 (N_34212,N_33540,N_33376);
nand U34213 (N_34213,N_33913,N_33465);
nor U34214 (N_34214,N_33517,N_33711);
nor U34215 (N_34215,N_33571,N_33155);
and U34216 (N_34216,N_33086,N_33790);
xnor U34217 (N_34217,N_33871,N_33414);
and U34218 (N_34218,N_33074,N_33588);
nand U34219 (N_34219,N_33346,N_33993);
nand U34220 (N_34220,N_33689,N_33983);
nor U34221 (N_34221,N_33521,N_33497);
nor U34222 (N_34222,N_33151,N_33181);
nor U34223 (N_34223,N_33768,N_33512);
xor U34224 (N_34224,N_33038,N_33832);
or U34225 (N_34225,N_33792,N_33280);
nand U34226 (N_34226,N_33863,N_33952);
xnor U34227 (N_34227,N_33925,N_33785);
xor U34228 (N_34228,N_33470,N_33836);
nor U34229 (N_34229,N_33541,N_33079);
xor U34230 (N_34230,N_33910,N_33544);
or U34231 (N_34231,N_33681,N_33624);
and U34232 (N_34232,N_33749,N_33596);
nor U34233 (N_34233,N_33763,N_33801);
nor U34234 (N_34234,N_33499,N_33629);
nor U34235 (N_34235,N_33265,N_33204);
nand U34236 (N_34236,N_33634,N_33606);
and U34237 (N_34237,N_33528,N_33394);
nor U34238 (N_34238,N_33977,N_33393);
or U34239 (N_34239,N_33076,N_33139);
xnor U34240 (N_34240,N_33008,N_33907);
nand U34241 (N_34241,N_33426,N_33619);
or U34242 (N_34242,N_33103,N_33315);
and U34243 (N_34243,N_33773,N_33463);
and U34244 (N_34244,N_33180,N_33099);
and U34245 (N_34245,N_33554,N_33216);
xnor U34246 (N_34246,N_33851,N_33868);
or U34247 (N_34247,N_33475,N_33359);
or U34248 (N_34248,N_33604,N_33731);
xnor U34249 (N_34249,N_33553,N_33000);
and U34250 (N_34250,N_33568,N_33617);
nor U34251 (N_34251,N_33455,N_33732);
xor U34252 (N_34252,N_33214,N_33783);
and U34253 (N_34253,N_33957,N_33587);
xnor U34254 (N_34254,N_33765,N_33451);
xnor U34255 (N_34255,N_33156,N_33312);
and U34256 (N_34256,N_33495,N_33892);
xor U34257 (N_34257,N_33003,N_33319);
nor U34258 (N_34258,N_33649,N_33534);
or U34259 (N_34259,N_33506,N_33804);
nor U34260 (N_34260,N_33294,N_33477);
nand U34261 (N_34261,N_33416,N_33608);
xor U34262 (N_34262,N_33121,N_33989);
nor U34263 (N_34263,N_33131,N_33467);
and U34264 (N_34264,N_33991,N_33071);
nand U34265 (N_34265,N_33275,N_33077);
or U34266 (N_34266,N_33800,N_33979);
nor U34267 (N_34267,N_33389,N_33755);
xor U34268 (N_34268,N_33080,N_33757);
xor U34269 (N_34269,N_33187,N_33736);
nand U34270 (N_34270,N_33984,N_33704);
and U34271 (N_34271,N_33545,N_33130);
xnor U34272 (N_34272,N_33227,N_33482);
or U34273 (N_34273,N_33360,N_33597);
nor U34274 (N_34274,N_33811,N_33576);
nand U34275 (N_34275,N_33918,N_33620);
nand U34276 (N_34276,N_33124,N_33935);
and U34277 (N_34277,N_33882,N_33666);
nor U34278 (N_34278,N_33301,N_33404);
nand U34279 (N_34279,N_33873,N_33138);
nand U34280 (N_34280,N_33016,N_33829);
or U34281 (N_34281,N_33561,N_33343);
or U34282 (N_34282,N_33024,N_33237);
nand U34283 (N_34283,N_33484,N_33307);
nor U34284 (N_34284,N_33229,N_33772);
or U34285 (N_34285,N_33660,N_33538);
xor U34286 (N_34286,N_33841,N_33043);
nor U34287 (N_34287,N_33364,N_33718);
and U34288 (N_34288,N_33782,N_33268);
or U34289 (N_34289,N_33722,N_33305);
nand U34290 (N_34290,N_33725,N_33412);
nor U34291 (N_34291,N_33581,N_33699);
xor U34292 (N_34292,N_33751,N_33719);
nand U34293 (N_34293,N_33329,N_33728);
nor U34294 (N_34294,N_33488,N_33595);
or U34295 (N_34295,N_33397,N_33249);
nand U34296 (N_34296,N_33149,N_33577);
nor U34297 (N_34297,N_33373,N_33118);
and U34298 (N_34298,N_33759,N_33833);
xnor U34299 (N_34299,N_33985,N_33970);
nor U34300 (N_34300,N_33992,N_33994);
or U34301 (N_34301,N_33206,N_33875);
xor U34302 (N_34302,N_33794,N_33924);
nand U34303 (N_34303,N_33640,N_33630);
nand U34304 (N_34304,N_33693,N_33771);
nor U34305 (N_34305,N_33982,N_33453);
nand U34306 (N_34306,N_33474,N_33936);
or U34307 (N_34307,N_33548,N_33564);
and U34308 (N_34308,N_33098,N_33123);
nand U34309 (N_34309,N_33107,N_33070);
nor U34310 (N_34310,N_33344,N_33600);
nand U34311 (N_34311,N_33246,N_33583);
nand U34312 (N_34312,N_33295,N_33310);
nand U34313 (N_34313,N_33738,N_33030);
xnor U34314 (N_34314,N_33320,N_33188);
and U34315 (N_34315,N_33105,N_33845);
nor U34316 (N_34316,N_33955,N_33696);
and U34317 (N_34317,N_33157,N_33386);
nor U34318 (N_34318,N_33337,N_33277);
xnor U34319 (N_34319,N_33651,N_33611);
xor U34320 (N_34320,N_33483,N_33598);
and U34321 (N_34321,N_33621,N_33091);
or U34322 (N_34322,N_33401,N_33789);
or U34323 (N_34323,N_33090,N_33685);
or U34324 (N_34324,N_33888,N_33062);
or U34325 (N_34325,N_33557,N_33374);
or U34326 (N_34326,N_33189,N_33427);
or U34327 (N_34327,N_33382,N_33172);
and U34328 (N_34328,N_33903,N_33929);
and U34329 (N_34329,N_33244,N_33633);
nand U34330 (N_34330,N_33173,N_33708);
xnor U34331 (N_34331,N_33430,N_33559);
or U34332 (N_34332,N_33978,N_33195);
nor U34333 (N_34333,N_33338,N_33490);
nor U34334 (N_34334,N_33741,N_33210);
nand U34335 (N_34335,N_33436,N_33594);
and U34336 (N_34336,N_33769,N_33405);
xnor U34337 (N_34337,N_33498,N_33387);
xnor U34338 (N_34338,N_33044,N_33142);
and U34339 (N_34339,N_33941,N_33345);
xor U34340 (N_34340,N_33684,N_33272);
nand U34341 (N_34341,N_33802,N_33297);
nor U34342 (N_34342,N_33092,N_33285);
or U34343 (N_34343,N_33969,N_33567);
xor U34344 (N_34344,N_33218,N_33039);
nand U34345 (N_34345,N_33615,N_33161);
or U34346 (N_34346,N_33653,N_33525);
nor U34347 (N_34347,N_33260,N_33850);
and U34348 (N_34348,N_33207,N_33102);
xor U34349 (N_34349,N_33796,N_33954);
and U34350 (N_34350,N_33399,N_33987);
nand U34351 (N_34351,N_33341,N_33439);
and U34352 (N_34352,N_33962,N_33834);
and U34353 (N_34353,N_33891,N_33007);
or U34354 (N_34354,N_33284,N_33968);
or U34355 (N_34355,N_33126,N_33896);
or U34356 (N_34356,N_33258,N_33570);
and U34357 (N_34357,N_33798,N_33922);
nor U34358 (N_34358,N_33306,N_33963);
nand U34359 (N_34359,N_33419,N_33339);
or U34360 (N_34360,N_33333,N_33464);
or U34361 (N_34361,N_33846,N_33119);
xor U34362 (N_34362,N_33961,N_33848);
xnor U34363 (N_34363,N_33706,N_33291);
xnor U34364 (N_34364,N_33336,N_33535);
nand U34365 (N_34365,N_33034,N_33035);
xor U34366 (N_34366,N_33934,N_33323);
and U34367 (N_34367,N_33111,N_33720);
nand U34368 (N_34368,N_33230,N_33494);
and U34369 (N_34369,N_33108,N_33226);
or U34370 (N_34370,N_33324,N_33876);
nor U34371 (N_34371,N_33228,N_33997);
nor U34372 (N_34372,N_33900,N_33878);
xnor U34373 (N_34373,N_33159,N_33574);
and U34374 (N_34374,N_33864,N_33723);
nor U34375 (N_34375,N_33182,N_33839);
nor U34376 (N_34376,N_33171,N_33866);
and U34377 (N_34377,N_33300,N_33395);
xor U34378 (N_34378,N_33211,N_33434);
nand U34379 (N_34379,N_33562,N_33898);
nor U34380 (N_34380,N_33212,N_33432);
xnor U34381 (N_34381,N_33668,N_33015);
or U34382 (N_34382,N_33930,N_33278);
and U34383 (N_34383,N_33743,N_33663);
xnor U34384 (N_34384,N_33221,N_33809);
xor U34385 (N_34385,N_33558,N_33823);
xnor U34386 (N_34386,N_33261,N_33309);
nand U34387 (N_34387,N_33877,N_33565);
or U34388 (N_34388,N_33296,N_33196);
xnor U34389 (N_34389,N_33433,N_33897);
or U34390 (N_34390,N_33814,N_33988);
nand U34391 (N_34391,N_33516,N_33446);
nor U34392 (N_34392,N_33136,N_33714);
nor U34393 (N_34393,N_33127,N_33311);
nand U34394 (N_34394,N_33148,N_33128);
nand U34395 (N_34395,N_33852,N_33046);
nand U34396 (N_34396,N_33162,N_33423);
and U34397 (N_34397,N_33191,N_33168);
nor U34398 (N_34398,N_33550,N_33163);
and U34399 (N_34399,N_33971,N_33895);
xor U34400 (N_34400,N_33045,N_33756);
nor U34401 (N_34401,N_33413,N_33281);
or U34402 (N_34402,N_33536,N_33424);
nand U34403 (N_34403,N_33701,N_33085);
nand U34404 (N_34404,N_33526,N_33064);
nor U34405 (N_34405,N_33733,N_33745);
or U34406 (N_34406,N_33586,N_33592);
or U34407 (N_34407,N_33511,N_33853);
nand U34408 (N_34408,N_33784,N_33885);
or U34409 (N_34409,N_33580,N_33383);
and U34410 (N_34410,N_33480,N_33134);
nor U34411 (N_34411,N_33764,N_33713);
or U34412 (N_34412,N_33921,N_33920);
or U34413 (N_34413,N_33174,N_33682);
xnor U34414 (N_34414,N_33022,N_33671);
nand U34415 (N_34415,N_33616,N_33645);
xor U34416 (N_34416,N_33737,N_33032);
or U34417 (N_34417,N_33192,N_33813);
nor U34418 (N_34418,N_33355,N_33362);
or U34419 (N_34419,N_33939,N_33644);
or U34420 (N_34420,N_33735,N_33753);
xnor U34421 (N_34421,N_33006,N_33575);
and U34422 (N_34422,N_33313,N_33089);
nor U34423 (N_34423,N_33631,N_33023);
or U34424 (N_34424,N_33050,N_33409);
nand U34425 (N_34425,N_33746,N_33304);
nand U34426 (N_34426,N_33479,N_33110);
or U34427 (N_34427,N_33144,N_33531);
xor U34428 (N_34428,N_33274,N_33104);
or U34429 (N_34429,N_33496,N_33328);
nand U34430 (N_34430,N_33956,N_33081);
xor U34431 (N_34431,N_33779,N_33454);
xor U34432 (N_34432,N_33915,N_33744);
nor U34433 (N_34433,N_33366,N_33094);
and U34434 (N_34434,N_33407,N_33904);
or U34435 (N_34435,N_33178,N_33893);
xor U34436 (N_34436,N_33747,N_33340);
and U34437 (N_34437,N_33632,N_33916);
or U34438 (N_34438,N_33292,N_33331);
nor U34439 (N_34439,N_33010,N_33471);
xor U34440 (N_34440,N_33729,N_33837);
and U34441 (N_34441,N_33664,N_33385);
nand U34442 (N_34442,N_33828,N_33776);
and U34443 (N_34443,N_33485,N_33770);
nor U34444 (N_34444,N_33657,N_33286);
nand U34445 (N_34445,N_33117,N_33507);
nor U34446 (N_34446,N_33450,N_33673);
xor U34447 (N_34447,N_33186,N_33537);
xor U34448 (N_34448,N_33060,N_33004);
and U34449 (N_34449,N_33881,N_33350);
nor U34450 (N_34450,N_33949,N_33147);
xor U34451 (N_34451,N_33509,N_33812);
or U34452 (N_34452,N_33456,N_33950);
or U34453 (N_34453,N_33270,N_33384);
or U34454 (N_34454,N_33354,N_33037);
or U34455 (N_34455,N_33810,N_33674);
and U34456 (N_34456,N_33662,N_33788);
or U34457 (N_34457,N_33652,N_33669);
nor U34458 (N_34458,N_33177,N_33469);
xnor U34459 (N_34459,N_33692,N_33715);
nor U34460 (N_34460,N_33860,N_33874);
nor U34461 (N_34461,N_33642,N_33240);
nand U34462 (N_34462,N_33835,N_33658);
and U34463 (N_34463,N_33572,N_33677);
or U34464 (N_34464,N_33095,N_33190);
or U34465 (N_34465,N_33225,N_33418);
or U34466 (N_34466,N_33082,N_33408);
or U34467 (N_34467,N_33242,N_33928);
and U34468 (N_34468,N_33635,N_33052);
nor U34469 (N_34469,N_33250,N_33862);
nand U34470 (N_34470,N_33213,N_33816);
or U34471 (N_34471,N_33073,N_33797);
and U34472 (N_34472,N_33289,N_33990);
xnor U34473 (N_34473,N_33501,N_33375);
and U34474 (N_34474,N_33775,N_33808);
xor U34475 (N_34475,N_33819,N_33522);
nand U34476 (N_34476,N_33223,N_33610);
and U34477 (N_34477,N_33442,N_33683);
nor U34478 (N_34478,N_33563,N_33510);
xnor U34479 (N_34479,N_33748,N_33486);
and U34480 (N_34480,N_33051,N_33088);
and U34481 (N_34481,N_33462,N_33100);
and U34482 (N_34482,N_33560,N_33974);
xor U34483 (N_34483,N_33780,N_33960);
nand U34484 (N_34484,N_33005,N_33314);
or U34485 (N_34485,N_33243,N_33179);
nor U34486 (N_34486,N_33680,N_33245);
xor U34487 (N_34487,N_33048,N_33084);
nand U34488 (N_34488,N_33012,N_33884);
nor U34489 (N_34489,N_33235,N_33547);
nand U34490 (N_34490,N_33140,N_33318);
nor U34491 (N_34491,N_33429,N_33655);
nor U34492 (N_34492,N_33777,N_33886);
nor U34493 (N_34493,N_33999,N_33555);
or U34494 (N_34494,N_33491,N_33514);
and U34495 (N_34495,N_33805,N_33636);
nor U34496 (N_34496,N_33909,N_33643);
nor U34497 (N_34497,N_33476,N_33750);
xnor U34498 (N_34498,N_33199,N_33165);
or U34499 (N_34499,N_33946,N_33287);
nor U34500 (N_34500,N_33799,N_33822);
xor U34501 (N_34501,N_33711,N_33537);
or U34502 (N_34502,N_33050,N_33059);
and U34503 (N_34503,N_33617,N_33792);
nor U34504 (N_34504,N_33009,N_33719);
nor U34505 (N_34505,N_33913,N_33513);
nor U34506 (N_34506,N_33566,N_33415);
and U34507 (N_34507,N_33313,N_33703);
nor U34508 (N_34508,N_33994,N_33418);
and U34509 (N_34509,N_33389,N_33705);
xor U34510 (N_34510,N_33986,N_33634);
and U34511 (N_34511,N_33138,N_33022);
or U34512 (N_34512,N_33841,N_33151);
nand U34513 (N_34513,N_33440,N_33364);
nand U34514 (N_34514,N_33750,N_33145);
or U34515 (N_34515,N_33297,N_33927);
xnor U34516 (N_34516,N_33477,N_33228);
nand U34517 (N_34517,N_33566,N_33758);
or U34518 (N_34518,N_33342,N_33459);
xnor U34519 (N_34519,N_33139,N_33015);
or U34520 (N_34520,N_33941,N_33971);
or U34521 (N_34521,N_33973,N_33535);
xnor U34522 (N_34522,N_33412,N_33526);
xnor U34523 (N_34523,N_33525,N_33481);
and U34524 (N_34524,N_33351,N_33085);
xnor U34525 (N_34525,N_33464,N_33947);
xnor U34526 (N_34526,N_33809,N_33334);
nor U34527 (N_34527,N_33061,N_33573);
nor U34528 (N_34528,N_33899,N_33449);
and U34529 (N_34529,N_33917,N_33162);
nand U34530 (N_34530,N_33175,N_33942);
and U34531 (N_34531,N_33689,N_33164);
and U34532 (N_34532,N_33312,N_33894);
xnor U34533 (N_34533,N_33674,N_33974);
nor U34534 (N_34534,N_33700,N_33068);
nand U34535 (N_34535,N_33852,N_33510);
nand U34536 (N_34536,N_33122,N_33304);
and U34537 (N_34537,N_33047,N_33287);
xor U34538 (N_34538,N_33811,N_33365);
and U34539 (N_34539,N_33542,N_33759);
nor U34540 (N_34540,N_33469,N_33880);
xnor U34541 (N_34541,N_33321,N_33505);
nor U34542 (N_34542,N_33955,N_33916);
or U34543 (N_34543,N_33936,N_33013);
nor U34544 (N_34544,N_33653,N_33483);
or U34545 (N_34545,N_33894,N_33564);
and U34546 (N_34546,N_33527,N_33909);
or U34547 (N_34547,N_33890,N_33995);
and U34548 (N_34548,N_33678,N_33081);
and U34549 (N_34549,N_33961,N_33860);
or U34550 (N_34550,N_33281,N_33468);
or U34551 (N_34551,N_33420,N_33297);
nand U34552 (N_34552,N_33191,N_33279);
nor U34553 (N_34553,N_33315,N_33764);
or U34554 (N_34554,N_33948,N_33262);
nor U34555 (N_34555,N_33760,N_33942);
or U34556 (N_34556,N_33654,N_33613);
xnor U34557 (N_34557,N_33118,N_33969);
nor U34558 (N_34558,N_33251,N_33029);
xnor U34559 (N_34559,N_33663,N_33027);
xor U34560 (N_34560,N_33613,N_33479);
or U34561 (N_34561,N_33326,N_33247);
and U34562 (N_34562,N_33441,N_33140);
or U34563 (N_34563,N_33516,N_33570);
nand U34564 (N_34564,N_33109,N_33626);
nand U34565 (N_34565,N_33541,N_33882);
or U34566 (N_34566,N_33238,N_33147);
and U34567 (N_34567,N_33921,N_33775);
xnor U34568 (N_34568,N_33765,N_33994);
or U34569 (N_34569,N_33791,N_33146);
nand U34570 (N_34570,N_33635,N_33509);
nor U34571 (N_34571,N_33726,N_33408);
nand U34572 (N_34572,N_33946,N_33107);
or U34573 (N_34573,N_33801,N_33766);
xor U34574 (N_34574,N_33583,N_33517);
or U34575 (N_34575,N_33694,N_33661);
or U34576 (N_34576,N_33702,N_33549);
nand U34577 (N_34577,N_33024,N_33277);
nor U34578 (N_34578,N_33571,N_33284);
xor U34579 (N_34579,N_33041,N_33883);
nor U34580 (N_34580,N_33979,N_33993);
nand U34581 (N_34581,N_33707,N_33676);
nand U34582 (N_34582,N_33521,N_33441);
xor U34583 (N_34583,N_33608,N_33816);
and U34584 (N_34584,N_33344,N_33156);
nor U34585 (N_34585,N_33675,N_33657);
nand U34586 (N_34586,N_33484,N_33077);
and U34587 (N_34587,N_33141,N_33749);
or U34588 (N_34588,N_33441,N_33226);
or U34589 (N_34589,N_33745,N_33884);
nand U34590 (N_34590,N_33774,N_33645);
nor U34591 (N_34591,N_33151,N_33818);
nand U34592 (N_34592,N_33947,N_33876);
nor U34593 (N_34593,N_33980,N_33649);
xnor U34594 (N_34594,N_33628,N_33833);
nor U34595 (N_34595,N_33997,N_33606);
nand U34596 (N_34596,N_33900,N_33712);
nor U34597 (N_34597,N_33396,N_33103);
nor U34598 (N_34598,N_33878,N_33820);
xor U34599 (N_34599,N_33111,N_33742);
or U34600 (N_34600,N_33882,N_33652);
or U34601 (N_34601,N_33869,N_33933);
or U34602 (N_34602,N_33849,N_33533);
and U34603 (N_34603,N_33468,N_33220);
and U34604 (N_34604,N_33496,N_33727);
or U34605 (N_34605,N_33127,N_33882);
or U34606 (N_34606,N_33496,N_33697);
and U34607 (N_34607,N_33874,N_33322);
nor U34608 (N_34608,N_33764,N_33460);
nand U34609 (N_34609,N_33602,N_33215);
nor U34610 (N_34610,N_33712,N_33033);
nor U34611 (N_34611,N_33384,N_33521);
xor U34612 (N_34612,N_33544,N_33474);
xnor U34613 (N_34613,N_33471,N_33783);
nor U34614 (N_34614,N_33744,N_33125);
nand U34615 (N_34615,N_33996,N_33417);
and U34616 (N_34616,N_33705,N_33874);
and U34617 (N_34617,N_33703,N_33782);
xor U34618 (N_34618,N_33614,N_33576);
and U34619 (N_34619,N_33627,N_33132);
or U34620 (N_34620,N_33275,N_33586);
nand U34621 (N_34621,N_33568,N_33268);
and U34622 (N_34622,N_33723,N_33438);
xor U34623 (N_34623,N_33329,N_33536);
or U34624 (N_34624,N_33539,N_33306);
nor U34625 (N_34625,N_33577,N_33177);
nand U34626 (N_34626,N_33940,N_33042);
or U34627 (N_34627,N_33562,N_33603);
xnor U34628 (N_34628,N_33911,N_33821);
or U34629 (N_34629,N_33877,N_33748);
xor U34630 (N_34630,N_33323,N_33288);
xor U34631 (N_34631,N_33367,N_33855);
or U34632 (N_34632,N_33086,N_33297);
and U34633 (N_34633,N_33880,N_33885);
xnor U34634 (N_34634,N_33516,N_33979);
nand U34635 (N_34635,N_33678,N_33122);
nor U34636 (N_34636,N_33754,N_33895);
xnor U34637 (N_34637,N_33867,N_33812);
nand U34638 (N_34638,N_33933,N_33179);
nand U34639 (N_34639,N_33647,N_33414);
nor U34640 (N_34640,N_33991,N_33593);
nand U34641 (N_34641,N_33256,N_33369);
and U34642 (N_34642,N_33615,N_33488);
nor U34643 (N_34643,N_33834,N_33028);
nand U34644 (N_34644,N_33768,N_33944);
nand U34645 (N_34645,N_33453,N_33359);
xnor U34646 (N_34646,N_33232,N_33140);
nor U34647 (N_34647,N_33791,N_33745);
nand U34648 (N_34648,N_33433,N_33350);
nor U34649 (N_34649,N_33781,N_33578);
and U34650 (N_34650,N_33245,N_33515);
and U34651 (N_34651,N_33095,N_33073);
or U34652 (N_34652,N_33822,N_33725);
and U34653 (N_34653,N_33073,N_33725);
nor U34654 (N_34654,N_33474,N_33561);
nor U34655 (N_34655,N_33364,N_33050);
or U34656 (N_34656,N_33308,N_33021);
nand U34657 (N_34657,N_33616,N_33367);
and U34658 (N_34658,N_33497,N_33820);
nand U34659 (N_34659,N_33496,N_33575);
or U34660 (N_34660,N_33162,N_33594);
xor U34661 (N_34661,N_33639,N_33684);
or U34662 (N_34662,N_33599,N_33535);
nand U34663 (N_34663,N_33302,N_33889);
and U34664 (N_34664,N_33697,N_33860);
nand U34665 (N_34665,N_33056,N_33328);
nor U34666 (N_34666,N_33658,N_33153);
and U34667 (N_34667,N_33315,N_33071);
or U34668 (N_34668,N_33032,N_33468);
xnor U34669 (N_34669,N_33564,N_33288);
and U34670 (N_34670,N_33077,N_33201);
xor U34671 (N_34671,N_33344,N_33214);
and U34672 (N_34672,N_33961,N_33834);
xnor U34673 (N_34673,N_33331,N_33934);
xor U34674 (N_34674,N_33777,N_33795);
nor U34675 (N_34675,N_33469,N_33107);
xnor U34676 (N_34676,N_33693,N_33762);
nand U34677 (N_34677,N_33142,N_33581);
xnor U34678 (N_34678,N_33963,N_33308);
xor U34679 (N_34679,N_33341,N_33281);
xnor U34680 (N_34680,N_33763,N_33984);
nand U34681 (N_34681,N_33773,N_33059);
nor U34682 (N_34682,N_33269,N_33999);
nand U34683 (N_34683,N_33669,N_33912);
nor U34684 (N_34684,N_33050,N_33213);
and U34685 (N_34685,N_33789,N_33660);
xor U34686 (N_34686,N_33604,N_33117);
xor U34687 (N_34687,N_33601,N_33254);
or U34688 (N_34688,N_33608,N_33924);
xor U34689 (N_34689,N_33336,N_33500);
nor U34690 (N_34690,N_33224,N_33240);
or U34691 (N_34691,N_33380,N_33955);
nand U34692 (N_34692,N_33763,N_33061);
nand U34693 (N_34693,N_33336,N_33141);
and U34694 (N_34694,N_33242,N_33815);
nor U34695 (N_34695,N_33993,N_33696);
xor U34696 (N_34696,N_33173,N_33850);
xnor U34697 (N_34697,N_33201,N_33425);
nand U34698 (N_34698,N_33294,N_33718);
and U34699 (N_34699,N_33943,N_33386);
and U34700 (N_34700,N_33384,N_33708);
or U34701 (N_34701,N_33887,N_33880);
and U34702 (N_34702,N_33438,N_33458);
and U34703 (N_34703,N_33850,N_33317);
nor U34704 (N_34704,N_33121,N_33022);
xnor U34705 (N_34705,N_33536,N_33082);
or U34706 (N_34706,N_33809,N_33330);
nor U34707 (N_34707,N_33428,N_33730);
nand U34708 (N_34708,N_33093,N_33885);
and U34709 (N_34709,N_33998,N_33644);
nand U34710 (N_34710,N_33408,N_33115);
nor U34711 (N_34711,N_33765,N_33008);
and U34712 (N_34712,N_33101,N_33316);
nand U34713 (N_34713,N_33087,N_33173);
xnor U34714 (N_34714,N_33950,N_33874);
nand U34715 (N_34715,N_33512,N_33550);
nor U34716 (N_34716,N_33775,N_33679);
and U34717 (N_34717,N_33067,N_33662);
nand U34718 (N_34718,N_33016,N_33167);
or U34719 (N_34719,N_33750,N_33692);
or U34720 (N_34720,N_33303,N_33221);
xor U34721 (N_34721,N_33264,N_33665);
nor U34722 (N_34722,N_33874,N_33697);
xor U34723 (N_34723,N_33454,N_33531);
nand U34724 (N_34724,N_33590,N_33583);
nand U34725 (N_34725,N_33763,N_33872);
nand U34726 (N_34726,N_33318,N_33834);
or U34727 (N_34727,N_33946,N_33770);
and U34728 (N_34728,N_33648,N_33299);
or U34729 (N_34729,N_33004,N_33744);
or U34730 (N_34730,N_33623,N_33287);
or U34731 (N_34731,N_33880,N_33939);
and U34732 (N_34732,N_33226,N_33286);
and U34733 (N_34733,N_33122,N_33280);
xnor U34734 (N_34734,N_33442,N_33997);
nor U34735 (N_34735,N_33753,N_33042);
and U34736 (N_34736,N_33343,N_33927);
nand U34737 (N_34737,N_33660,N_33834);
and U34738 (N_34738,N_33769,N_33058);
xor U34739 (N_34739,N_33614,N_33117);
or U34740 (N_34740,N_33393,N_33159);
or U34741 (N_34741,N_33842,N_33900);
xnor U34742 (N_34742,N_33945,N_33585);
and U34743 (N_34743,N_33457,N_33815);
and U34744 (N_34744,N_33605,N_33207);
nand U34745 (N_34745,N_33497,N_33484);
nand U34746 (N_34746,N_33477,N_33241);
and U34747 (N_34747,N_33968,N_33053);
xnor U34748 (N_34748,N_33661,N_33806);
or U34749 (N_34749,N_33276,N_33895);
nand U34750 (N_34750,N_33934,N_33727);
and U34751 (N_34751,N_33578,N_33422);
and U34752 (N_34752,N_33458,N_33489);
and U34753 (N_34753,N_33386,N_33878);
or U34754 (N_34754,N_33480,N_33565);
nor U34755 (N_34755,N_33571,N_33679);
nand U34756 (N_34756,N_33328,N_33318);
nand U34757 (N_34757,N_33704,N_33483);
nand U34758 (N_34758,N_33258,N_33906);
xnor U34759 (N_34759,N_33931,N_33117);
nor U34760 (N_34760,N_33774,N_33821);
or U34761 (N_34761,N_33668,N_33766);
xor U34762 (N_34762,N_33299,N_33079);
nand U34763 (N_34763,N_33674,N_33682);
xnor U34764 (N_34764,N_33017,N_33975);
and U34765 (N_34765,N_33238,N_33339);
and U34766 (N_34766,N_33695,N_33635);
and U34767 (N_34767,N_33639,N_33786);
or U34768 (N_34768,N_33985,N_33466);
and U34769 (N_34769,N_33829,N_33906);
and U34770 (N_34770,N_33079,N_33289);
xnor U34771 (N_34771,N_33311,N_33239);
xor U34772 (N_34772,N_33758,N_33382);
nand U34773 (N_34773,N_33228,N_33756);
xor U34774 (N_34774,N_33878,N_33021);
or U34775 (N_34775,N_33259,N_33987);
and U34776 (N_34776,N_33024,N_33687);
nor U34777 (N_34777,N_33835,N_33958);
nand U34778 (N_34778,N_33462,N_33918);
or U34779 (N_34779,N_33542,N_33809);
xor U34780 (N_34780,N_33221,N_33896);
nor U34781 (N_34781,N_33157,N_33956);
or U34782 (N_34782,N_33364,N_33791);
nand U34783 (N_34783,N_33315,N_33954);
nand U34784 (N_34784,N_33846,N_33302);
nor U34785 (N_34785,N_33076,N_33176);
nor U34786 (N_34786,N_33365,N_33013);
or U34787 (N_34787,N_33661,N_33531);
or U34788 (N_34788,N_33865,N_33951);
nand U34789 (N_34789,N_33690,N_33313);
and U34790 (N_34790,N_33391,N_33993);
nand U34791 (N_34791,N_33333,N_33431);
nand U34792 (N_34792,N_33782,N_33269);
xor U34793 (N_34793,N_33941,N_33896);
nor U34794 (N_34794,N_33089,N_33886);
nand U34795 (N_34795,N_33492,N_33289);
or U34796 (N_34796,N_33314,N_33086);
and U34797 (N_34797,N_33733,N_33301);
and U34798 (N_34798,N_33018,N_33799);
xnor U34799 (N_34799,N_33705,N_33019);
and U34800 (N_34800,N_33011,N_33867);
nor U34801 (N_34801,N_33411,N_33488);
or U34802 (N_34802,N_33749,N_33582);
xnor U34803 (N_34803,N_33038,N_33840);
nor U34804 (N_34804,N_33008,N_33992);
or U34805 (N_34805,N_33711,N_33362);
nor U34806 (N_34806,N_33900,N_33750);
and U34807 (N_34807,N_33169,N_33568);
xor U34808 (N_34808,N_33338,N_33854);
or U34809 (N_34809,N_33968,N_33980);
and U34810 (N_34810,N_33701,N_33841);
or U34811 (N_34811,N_33507,N_33842);
xor U34812 (N_34812,N_33017,N_33661);
nand U34813 (N_34813,N_33301,N_33960);
or U34814 (N_34814,N_33321,N_33205);
and U34815 (N_34815,N_33002,N_33376);
nor U34816 (N_34816,N_33792,N_33225);
nor U34817 (N_34817,N_33077,N_33836);
xor U34818 (N_34818,N_33800,N_33205);
or U34819 (N_34819,N_33707,N_33645);
nand U34820 (N_34820,N_33575,N_33941);
nor U34821 (N_34821,N_33023,N_33757);
and U34822 (N_34822,N_33514,N_33098);
nor U34823 (N_34823,N_33656,N_33820);
nand U34824 (N_34824,N_33797,N_33400);
and U34825 (N_34825,N_33124,N_33876);
and U34826 (N_34826,N_33616,N_33691);
or U34827 (N_34827,N_33238,N_33424);
nand U34828 (N_34828,N_33125,N_33721);
nand U34829 (N_34829,N_33777,N_33184);
nor U34830 (N_34830,N_33767,N_33214);
nand U34831 (N_34831,N_33885,N_33072);
and U34832 (N_34832,N_33913,N_33042);
xnor U34833 (N_34833,N_33052,N_33004);
or U34834 (N_34834,N_33086,N_33474);
or U34835 (N_34835,N_33730,N_33962);
or U34836 (N_34836,N_33795,N_33375);
xor U34837 (N_34837,N_33099,N_33027);
nor U34838 (N_34838,N_33613,N_33193);
nor U34839 (N_34839,N_33097,N_33119);
nand U34840 (N_34840,N_33658,N_33654);
or U34841 (N_34841,N_33495,N_33705);
nand U34842 (N_34842,N_33114,N_33673);
xnor U34843 (N_34843,N_33101,N_33679);
and U34844 (N_34844,N_33464,N_33846);
or U34845 (N_34845,N_33280,N_33050);
xnor U34846 (N_34846,N_33458,N_33350);
or U34847 (N_34847,N_33382,N_33281);
xor U34848 (N_34848,N_33599,N_33897);
or U34849 (N_34849,N_33298,N_33180);
xnor U34850 (N_34850,N_33593,N_33474);
xnor U34851 (N_34851,N_33269,N_33859);
and U34852 (N_34852,N_33864,N_33395);
or U34853 (N_34853,N_33055,N_33898);
or U34854 (N_34854,N_33204,N_33692);
and U34855 (N_34855,N_33160,N_33992);
and U34856 (N_34856,N_33032,N_33883);
nand U34857 (N_34857,N_33580,N_33040);
or U34858 (N_34858,N_33086,N_33340);
nand U34859 (N_34859,N_33938,N_33368);
and U34860 (N_34860,N_33505,N_33157);
xnor U34861 (N_34861,N_33951,N_33963);
or U34862 (N_34862,N_33151,N_33995);
xor U34863 (N_34863,N_33741,N_33756);
nand U34864 (N_34864,N_33110,N_33455);
or U34865 (N_34865,N_33090,N_33864);
nand U34866 (N_34866,N_33108,N_33100);
nor U34867 (N_34867,N_33178,N_33815);
xnor U34868 (N_34868,N_33125,N_33404);
or U34869 (N_34869,N_33462,N_33639);
and U34870 (N_34870,N_33449,N_33067);
xnor U34871 (N_34871,N_33280,N_33009);
xnor U34872 (N_34872,N_33655,N_33618);
and U34873 (N_34873,N_33056,N_33658);
or U34874 (N_34874,N_33611,N_33850);
nor U34875 (N_34875,N_33814,N_33240);
nand U34876 (N_34876,N_33422,N_33380);
or U34877 (N_34877,N_33966,N_33648);
nand U34878 (N_34878,N_33451,N_33620);
xnor U34879 (N_34879,N_33307,N_33857);
and U34880 (N_34880,N_33535,N_33685);
xor U34881 (N_34881,N_33766,N_33081);
nand U34882 (N_34882,N_33668,N_33498);
and U34883 (N_34883,N_33221,N_33983);
xor U34884 (N_34884,N_33709,N_33913);
nor U34885 (N_34885,N_33160,N_33383);
nor U34886 (N_34886,N_33019,N_33139);
xor U34887 (N_34887,N_33232,N_33392);
xnor U34888 (N_34888,N_33982,N_33050);
and U34889 (N_34889,N_33826,N_33469);
and U34890 (N_34890,N_33722,N_33242);
and U34891 (N_34891,N_33294,N_33540);
or U34892 (N_34892,N_33081,N_33069);
nand U34893 (N_34893,N_33992,N_33183);
nor U34894 (N_34894,N_33635,N_33938);
xnor U34895 (N_34895,N_33926,N_33880);
xnor U34896 (N_34896,N_33402,N_33886);
or U34897 (N_34897,N_33524,N_33201);
nand U34898 (N_34898,N_33377,N_33695);
nand U34899 (N_34899,N_33976,N_33249);
and U34900 (N_34900,N_33937,N_33925);
nor U34901 (N_34901,N_33959,N_33151);
nand U34902 (N_34902,N_33115,N_33217);
nand U34903 (N_34903,N_33887,N_33806);
or U34904 (N_34904,N_33236,N_33080);
nand U34905 (N_34905,N_33898,N_33147);
or U34906 (N_34906,N_33637,N_33801);
or U34907 (N_34907,N_33868,N_33025);
xnor U34908 (N_34908,N_33445,N_33298);
and U34909 (N_34909,N_33167,N_33374);
and U34910 (N_34910,N_33810,N_33499);
nand U34911 (N_34911,N_33311,N_33713);
nand U34912 (N_34912,N_33789,N_33597);
and U34913 (N_34913,N_33314,N_33623);
nor U34914 (N_34914,N_33547,N_33924);
nor U34915 (N_34915,N_33632,N_33082);
and U34916 (N_34916,N_33295,N_33961);
or U34917 (N_34917,N_33804,N_33238);
nand U34918 (N_34918,N_33198,N_33378);
nor U34919 (N_34919,N_33174,N_33185);
xor U34920 (N_34920,N_33746,N_33799);
or U34921 (N_34921,N_33110,N_33736);
nand U34922 (N_34922,N_33141,N_33748);
or U34923 (N_34923,N_33232,N_33176);
nand U34924 (N_34924,N_33320,N_33305);
nand U34925 (N_34925,N_33593,N_33623);
xnor U34926 (N_34926,N_33975,N_33840);
xnor U34927 (N_34927,N_33812,N_33841);
nand U34928 (N_34928,N_33512,N_33765);
and U34929 (N_34929,N_33957,N_33061);
nor U34930 (N_34930,N_33993,N_33781);
xnor U34931 (N_34931,N_33137,N_33836);
and U34932 (N_34932,N_33562,N_33043);
nor U34933 (N_34933,N_33929,N_33277);
nor U34934 (N_34934,N_33449,N_33705);
and U34935 (N_34935,N_33046,N_33257);
and U34936 (N_34936,N_33351,N_33847);
or U34937 (N_34937,N_33665,N_33818);
xor U34938 (N_34938,N_33079,N_33624);
and U34939 (N_34939,N_33825,N_33333);
nand U34940 (N_34940,N_33685,N_33433);
nor U34941 (N_34941,N_33620,N_33159);
and U34942 (N_34942,N_33451,N_33983);
xor U34943 (N_34943,N_33160,N_33613);
nor U34944 (N_34944,N_33768,N_33918);
xnor U34945 (N_34945,N_33955,N_33570);
or U34946 (N_34946,N_33707,N_33000);
and U34947 (N_34947,N_33890,N_33341);
xor U34948 (N_34948,N_33007,N_33211);
nand U34949 (N_34949,N_33544,N_33156);
or U34950 (N_34950,N_33906,N_33230);
xor U34951 (N_34951,N_33568,N_33092);
and U34952 (N_34952,N_33995,N_33208);
nor U34953 (N_34953,N_33947,N_33440);
or U34954 (N_34954,N_33218,N_33597);
nor U34955 (N_34955,N_33750,N_33776);
nor U34956 (N_34956,N_33059,N_33080);
nand U34957 (N_34957,N_33081,N_33537);
nand U34958 (N_34958,N_33482,N_33986);
and U34959 (N_34959,N_33937,N_33763);
or U34960 (N_34960,N_33182,N_33987);
and U34961 (N_34961,N_33333,N_33318);
xnor U34962 (N_34962,N_33783,N_33525);
nor U34963 (N_34963,N_33345,N_33615);
and U34964 (N_34964,N_33271,N_33551);
nand U34965 (N_34965,N_33281,N_33368);
xor U34966 (N_34966,N_33213,N_33942);
and U34967 (N_34967,N_33746,N_33777);
and U34968 (N_34968,N_33801,N_33884);
xnor U34969 (N_34969,N_33016,N_33918);
nand U34970 (N_34970,N_33910,N_33909);
nand U34971 (N_34971,N_33894,N_33895);
nand U34972 (N_34972,N_33853,N_33009);
nor U34973 (N_34973,N_33519,N_33553);
xor U34974 (N_34974,N_33731,N_33507);
nand U34975 (N_34975,N_33112,N_33124);
and U34976 (N_34976,N_33174,N_33563);
and U34977 (N_34977,N_33678,N_33038);
or U34978 (N_34978,N_33452,N_33758);
or U34979 (N_34979,N_33979,N_33694);
and U34980 (N_34980,N_33727,N_33665);
and U34981 (N_34981,N_33950,N_33812);
or U34982 (N_34982,N_33381,N_33528);
or U34983 (N_34983,N_33137,N_33774);
nand U34984 (N_34984,N_33980,N_33207);
xor U34985 (N_34985,N_33216,N_33932);
and U34986 (N_34986,N_33522,N_33026);
and U34987 (N_34987,N_33646,N_33904);
nor U34988 (N_34988,N_33665,N_33109);
nand U34989 (N_34989,N_33881,N_33858);
xnor U34990 (N_34990,N_33723,N_33453);
xnor U34991 (N_34991,N_33114,N_33630);
nand U34992 (N_34992,N_33015,N_33338);
nor U34993 (N_34993,N_33437,N_33318);
nor U34994 (N_34994,N_33106,N_33824);
xnor U34995 (N_34995,N_33548,N_33618);
and U34996 (N_34996,N_33570,N_33501);
or U34997 (N_34997,N_33609,N_33124);
and U34998 (N_34998,N_33326,N_33525);
nand U34999 (N_34999,N_33587,N_33498);
nor U35000 (N_35000,N_34680,N_34064);
nand U35001 (N_35001,N_34016,N_34158);
xnor U35002 (N_35002,N_34115,N_34171);
or U35003 (N_35003,N_34869,N_34394);
nand U35004 (N_35004,N_34276,N_34445);
or U35005 (N_35005,N_34474,N_34047);
and U35006 (N_35006,N_34997,N_34086);
and U35007 (N_35007,N_34591,N_34592);
or U35008 (N_35008,N_34184,N_34325);
nor U35009 (N_35009,N_34254,N_34930);
or U35010 (N_35010,N_34863,N_34439);
nor U35011 (N_35011,N_34471,N_34765);
xnor U35012 (N_35012,N_34023,N_34759);
nor U35013 (N_35013,N_34854,N_34101);
nor U35014 (N_35014,N_34665,N_34488);
nand U35015 (N_35015,N_34646,N_34326);
nand U35016 (N_35016,N_34905,N_34727);
nand U35017 (N_35017,N_34752,N_34927);
nand U35018 (N_35018,N_34786,N_34923);
nand U35019 (N_35019,N_34845,N_34437);
and U35020 (N_35020,N_34622,N_34203);
nor U35021 (N_35021,N_34972,N_34459);
and U35022 (N_35022,N_34550,N_34684);
and U35023 (N_35023,N_34220,N_34539);
and U35024 (N_35024,N_34698,N_34682);
xnor U35025 (N_35025,N_34559,N_34771);
and U35026 (N_35026,N_34837,N_34195);
and U35027 (N_35027,N_34371,N_34004);
and U35028 (N_35028,N_34781,N_34238);
or U35029 (N_35029,N_34027,N_34348);
or U35030 (N_35030,N_34758,N_34129);
or U35031 (N_35031,N_34624,N_34926);
or U35032 (N_35032,N_34636,N_34260);
or U35033 (N_35033,N_34971,N_34921);
and U35034 (N_35034,N_34545,N_34832);
nor U35035 (N_35035,N_34168,N_34777);
xor U35036 (N_35036,N_34312,N_34172);
and U35037 (N_35037,N_34491,N_34204);
or U35038 (N_35038,N_34618,N_34750);
xnor U35039 (N_35039,N_34511,N_34537);
or U35040 (N_35040,N_34892,N_34187);
and U35041 (N_35041,N_34249,N_34661);
xnor U35042 (N_35042,N_34035,N_34141);
and U35043 (N_35043,N_34749,N_34008);
nand U35044 (N_35044,N_34753,N_34933);
nand U35045 (N_35045,N_34526,N_34484);
or U35046 (N_35046,N_34370,N_34907);
nor U35047 (N_35047,N_34599,N_34029);
nand U35048 (N_35048,N_34876,N_34039);
and U35049 (N_35049,N_34958,N_34495);
and U35050 (N_35050,N_34843,N_34882);
and U35051 (N_35051,N_34784,N_34945);
or U35052 (N_35052,N_34766,N_34337);
xor U35053 (N_35053,N_34896,N_34134);
xor U35054 (N_35054,N_34691,N_34557);
nor U35055 (N_35055,N_34475,N_34149);
xor U35056 (N_35056,N_34621,N_34946);
nor U35057 (N_35057,N_34009,N_34292);
and U35058 (N_35058,N_34351,N_34272);
or U35059 (N_35059,N_34441,N_34556);
nand U35060 (N_35060,N_34055,N_34365);
or U35061 (N_35061,N_34660,N_34476);
or U35062 (N_35062,N_34431,N_34800);
nor U35063 (N_35063,N_34306,N_34755);
or U35064 (N_35064,N_34740,N_34797);
nand U35065 (N_35065,N_34320,N_34030);
xnor U35066 (N_35066,N_34173,N_34938);
nand U35067 (N_35067,N_34779,N_34527);
xor U35068 (N_35068,N_34226,N_34572);
or U35069 (N_35069,N_34121,N_34018);
nand U35070 (N_35070,N_34335,N_34770);
xnor U35071 (N_35071,N_34117,N_34970);
nand U35072 (N_35072,N_34595,N_34332);
nor U35073 (N_35073,N_34396,N_34935);
nor U35074 (N_35074,N_34066,N_34073);
and U35075 (N_35075,N_34163,N_34726);
nor U35076 (N_35076,N_34225,N_34780);
nor U35077 (N_35077,N_34688,N_34872);
nand U35078 (N_35078,N_34369,N_34707);
nor U35079 (N_35079,N_34553,N_34323);
and U35080 (N_35080,N_34552,N_34918);
nand U35081 (N_35081,N_34915,N_34356);
and U35082 (N_35082,N_34668,N_34314);
and U35083 (N_35083,N_34640,N_34216);
and U35084 (N_35084,N_34625,N_34290);
nor U35085 (N_35085,N_34060,N_34307);
xor U35086 (N_35086,N_34222,N_34014);
nor U35087 (N_35087,N_34864,N_34390);
xor U35088 (N_35088,N_34404,N_34637);
and U35089 (N_35089,N_34453,N_34783);
xnor U35090 (N_35090,N_34514,N_34531);
nand U35091 (N_35091,N_34152,N_34499);
or U35092 (N_35092,N_34182,N_34889);
or U35093 (N_35093,N_34528,N_34577);
or U35094 (N_35094,N_34062,N_34135);
nor U35095 (N_35095,N_34022,N_34125);
xnor U35096 (N_35096,N_34413,N_34457);
or U35097 (N_35097,N_34075,N_34300);
nand U35098 (N_35098,N_34996,N_34099);
xnor U35099 (N_35099,N_34520,N_34201);
xnor U35100 (N_35100,N_34833,N_34639);
or U35101 (N_35101,N_34380,N_34130);
nor U35102 (N_35102,N_34309,N_34798);
nand U35103 (N_35103,N_34360,N_34011);
and U35104 (N_35104,N_34106,N_34259);
and U35105 (N_35105,N_34724,N_34664);
xor U35106 (N_35106,N_34339,N_34068);
nor U35107 (N_35107,N_34477,N_34188);
or U35108 (N_35108,N_34078,N_34811);
xnor U35109 (N_35109,N_34825,N_34675);
nand U35110 (N_35110,N_34283,N_34578);
xor U35111 (N_35111,N_34033,N_34223);
and U35112 (N_35112,N_34534,N_34709);
nor U35113 (N_35113,N_34217,N_34012);
and U35114 (N_35114,N_34028,N_34983);
nor U35115 (N_35115,N_34100,N_34059);
nor U35116 (N_35116,N_34543,N_34447);
and U35117 (N_35117,N_34388,N_34436);
nand U35118 (N_35118,N_34560,N_34213);
or U35119 (N_35119,N_34420,N_34993);
xnor U35120 (N_35120,N_34190,N_34296);
or U35121 (N_35121,N_34063,N_34076);
or U35122 (N_35122,N_34812,N_34735);
xnor U35123 (N_35123,N_34347,N_34738);
or U35124 (N_35124,N_34775,N_34629);
nor U35125 (N_35125,N_34576,N_34362);
nor U35126 (N_35126,N_34040,N_34888);
and U35127 (N_35127,N_34287,N_34105);
and U35128 (N_35128,N_34359,N_34044);
and U35129 (N_35129,N_34991,N_34391);
xnor U35130 (N_35130,N_34914,N_34401);
nand U35131 (N_35131,N_34443,N_34089);
and U35132 (N_35132,N_34823,N_34649);
nand U35133 (N_35133,N_34252,N_34703);
or U35134 (N_35134,N_34403,N_34103);
and U35135 (N_35135,N_34170,N_34179);
xor U35136 (N_35136,N_34953,N_34840);
nor U35137 (N_35137,N_34248,N_34286);
or U35138 (N_35138,N_34334,N_34400);
xor U35139 (N_35139,N_34198,N_34432);
or U35140 (N_35140,N_34712,N_34763);
nand U35141 (N_35141,N_34246,N_34697);
nand U35142 (N_35142,N_34271,N_34229);
nor U35143 (N_35143,N_34670,N_34126);
and U35144 (N_35144,N_34674,N_34270);
nor U35145 (N_35145,N_34166,N_34005);
xnor U35146 (N_35146,N_34808,N_34265);
nor U35147 (N_35147,N_34257,N_34718);
and U35148 (N_35148,N_34042,N_34731);
or U35149 (N_35149,N_34962,N_34212);
or U35150 (N_35150,N_34316,N_34087);
nor U35151 (N_35151,N_34581,N_34666);
nand U35152 (N_35152,N_34155,N_34357);
and U35153 (N_35153,N_34449,N_34289);
nor U35154 (N_35154,N_34717,N_34116);
nand U35155 (N_35155,N_34333,N_34500);
nor U35156 (N_35156,N_34136,N_34795);
and U35157 (N_35157,N_34451,N_34153);
nor U35158 (N_35158,N_34767,N_34679);
nand U35159 (N_35159,N_34659,N_34151);
nor U35160 (N_35160,N_34501,N_34279);
and U35161 (N_35161,N_34446,N_34722);
nand U35162 (N_35162,N_34275,N_34548);
nand U35163 (N_35163,N_34414,N_34482);
and U35164 (N_35164,N_34327,N_34853);
and U35165 (N_35165,N_34744,N_34769);
or U35166 (N_35166,N_34866,N_34821);
xnor U35167 (N_35167,N_34025,N_34603);
and U35168 (N_35168,N_34774,N_34980);
nand U35169 (N_35169,N_34429,N_34920);
xnor U35170 (N_35170,N_34588,N_34317);
xor U35171 (N_35171,N_34716,N_34486);
or U35172 (N_35172,N_34694,N_34992);
nand U35173 (N_35173,N_34407,N_34515);
and U35174 (N_35174,N_34937,N_34194);
nand U35175 (N_35175,N_34813,N_34579);
or U35176 (N_35176,N_34378,N_34313);
nand U35177 (N_35177,N_34858,N_34990);
or U35178 (N_35178,N_34344,N_34143);
nor U35179 (N_35179,N_34234,N_34667);
or U35180 (N_35180,N_34051,N_34352);
or U35181 (N_35181,N_34886,N_34002);
and U35182 (N_35182,N_34240,N_34412);
or U35183 (N_35183,N_34540,N_34341);
and U35184 (N_35184,N_34302,N_34139);
nor U35185 (N_35185,N_34608,N_34549);
nand U35186 (N_35186,N_34093,N_34473);
and U35187 (N_35187,N_34934,N_34031);
nand U35188 (N_35188,N_34806,N_34834);
or U35189 (N_35189,N_34176,N_34338);
or U35190 (N_35190,N_34050,N_34433);
nor U35191 (N_35191,N_34000,N_34623);
nand U35192 (N_35192,N_34802,N_34109);
or U35193 (N_35193,N_34868,N_34428);
or U35194 (N_35194,N_34999,N_34746);
xor U35195 (N_35195,N_34734,N_34444);
nand U35196 (N_35196,N_34605,N_34138);
nor U35197 (N_35197,N_34650,N_34175);
and U35198 (N_35198,N_34430,N_34742);
nor U35199 (N_35199,N_34601,N_34232);
nand U35200 (N_35200,N_34288,N_34828);
nand U35201 (N_35201,N_34424,N_34416);
nor U35202 (N_35202,N_34693,N_34221);
xnor U35203 (N_35203,N_34386,N_34901);
xnor U35204 (N_35204,N_34277,N_34110);
nand U35205 (N_35205,N_34522,N_34523);
or U35206 (N_35206,N_34810,N_34494);
or U35207 (N_35207,N_34835,N_34793);
or U35208 (N_35208,N_34354,N_34974);
or U35209 (N_35209,N_34897,N_34911);
and U35210 (N_35210,N_34342,N_34676);
xnor U35211 (N_35211,N_34924,N_34525);
nand U35212 (N_35212,N_34367,N_34045);
nand U35213 (N_35213,N_34585,N_34931);
nor U35214 (N_35214,N_34161,N_34733);
xnor U35215 (N_35215,N_34502,N_34114);
and U35216 (N_35216,N_34468,N_34957);
or U35217 (N_35217,N_34487,N_34049);
nand U35218 (N_35218,N_34651,N_34298);
nor U35219 (N_35219,N_34399,N_34162);
and U35220 (N_35220,N_34455,N_34328);
nor U35221 (N_35221,N_34434,N_34303);
nor U35222 (N_35222,N_34202,N_34778);
xor U35223 (N_35223,N_34695,N_34479);
xnor U35224 (N_35224,N_34794,N_34336);
and U35225 (N_35225,N_34977,N_34311);
nor U35226 (N_35226,N_34376,N_34242);
nor U35227 (N_35227,N_34418,N_34575);
or U35228 (N_35228,N_34205,N_34791);
nor U35229 (N_35229,N_34614,N_34003);
nand U35230 (N_35230,N_34379,N_34186);
or U35231 (N_35231,N_34681,N_34224);
nand U35232 (N_35232,N_34554,N_34566);
nand U35233 (N_35233,N_34615,N_34529);
or U35234 (N_35234,N_34177,N_34903);
and U35235 (N_35235,N_34253,N_34739);
nand U35236 (N_35236,N_34839,N_34278);
xor U35237 (N_35237,N_34538,N_34017);
or U35238 (N_35238,N_34616,N_34638);
and U35239 (N_35239,N_34867,N_34088);
or U35240 (N_35240,N_34510,N_34409);
and U35241 (N_35241,N_34112,N_34206);
nand U35242 (N_35242,N_34816,N_34850);
or U35243 (N_35243,N_34015,N_34363);
nor U35244 (N_35244,N_34984,N_34826);
xor U35245 (N_35245,N_34330,N_34448);
xor U35246 (N_35246,N_34497,N_34207);
and U35247 (N_35247,N_34824,N_34587);
nor U35248 (N_35248,N_34366,N_34174);
xor U35249 (N_35249,N_34541,N_34393);
nand U35250 (N_35250,N_34561,N_34193);
and U35251 (N_35251,N_34569,N_34095);
nand U35252 (N_35252,N_34757,N_34438);
nor U35253 (N_35253,N_34489,N_34090);
nand U35254 (N_35254,N_34730,N_34619);
and U35255 (N_35255,N_34788,N_34013);
xor U35256 (N_35256,N_34879,N_34966);
xnor U35257 (N_35257,N_34452,N_34836);
xor U35258 (N_35258,N_34120,N_34975);
nor U35259 (N_35259,N_34498,N_34237);
nor U35260 (N_35260,N_34273,N_34567);
xor U35261 (N_35261,N_34656,N_34041);
nor U35262 (N_35262,N_34963,N_34805);
and U35263 (N_35263,N_34415,N_34633);
nand U35264 (N_35264,N_34925,N_34199);
or U35265 (N_35265,N_34644,N_34936);
and U35266 (N_35266,N_34111,N_34720);
nand U35267 (N_35267,N_34916,N_34465);
nand U35268 (N_35268,N_34210,N_34819);
xnor U35269 (N_35269,N_34729,N_34654);
nand U35270 (N_35270,N_34589,N_34208);
or U35271 (N_35271,N_34372,N_34862);
and U35272 (N_35272,N_34301,N_34949);
nor U35273 (N_35273,N_34227,N_34532);
nand U35274 (N_35274,N_34282,N_34425);
nand U35275 (N_35275,N_34061,N_34492);
or U35276 (N_35276,N_34702,N_34546);
nand U35277 (N_35277,N_34382,N_34353);
xnor U35278 (N_35278,N_34961,N_34214);
xor U35279 (N_35279,N_34760,N_34450);
xnor U35280 (N_35280,N_34374,N_34939);
or U35281 (N_35281,N_34381,N_34846);
nor U35282 (N_35282,N_34512,N_34435);
nand U35283 (N_35283,N_34950,N_34524);
nor U35284 (N_35284,N_34427,N_34102);
nand U35285 (N_35285,N_34671,N_34917);
or U35286 (N_35286,N_34887,N_34036);
nand U35287 (N_35287,N_34809,N_34375);
nor U35288 (N_35288,N_34085,N_34861);
xnor U35289 (N_35289,N_34197,N_34144);
nand U35290 (N_35290,N_34267,N_34988);
or U35291 (N_35291,N_34948,N_34714);
xor U35292 (N_35292,N_34235,N_34507);
xnor U35293 (N_35293,N_34324,N_34606);
nor U35294 (N_35294,N_34628,N_34870);
xnor U35295 (N_35295,N_34642,N_34973);
and U35296 (N_35296,N_34250,N_34598);
or U35297 (N_35297,N_34683,N_34987);
nor U35298 (N_35298,N_34142,N_34461);
or U35299 (N_35299,N_34231,N_34890);
and U35300 (N_35300,N_34191,N_34304);
and U35301 (N_35301,N_34140,N_34426);
or U35302 (N_35302,N_34124,N_34701);
nor U35303 (N_35303,N_34299,N_34728);
nor U35304 (N_35304,N_34536,N_34322);
and U35305 (N_35305,N_34402,N_34180);
and U35306 (N_35306,N_34083,N_34266);
nor U35307 (N_35307,N_34831,N_34590);
nor U35308 (N_35308,N_34119,N_34183);
and U35309 (N_35309,N_34137,N_34613);
xor U35310 (N_35310,N_34908,N_34768);
xnor U35311 (N_35311,N_34704,N_34294);
xor U35312 (N_35312,N_34192,N_34956);
and U35313 (N_35313,N_34293,N_34065);
and U35314 (N_35314,N_34251,N_34519);
nand U35315 (N_35315,N_34421,N_34885);
nand U35316 (N_35316,N_34094,N_34133);
nor U35317 (N_35317,N_34384,N_34032);
or U35318 (N_35318,N_34493,N_34932);
nor U35319 (N_35319,N_34269,N_34620);
xor U35320 (N_35320,N_34849,N_34851);
and U35321 (N_35321,N_34228,N_34626);
or U35322 (N_35322,N_34842,N_34838);
or U35323 (N_35323,N_34690,N_34215);
or U35324 (N_35324,N_34721,N_34280);
nor U35325 (N_35325,N_34969,N_34108);
and U35326 (N_35326,N_34700,N_34264);
nand U35327 (N_35327,N_34263,N_34178);
nand U35328 (N_35328,N_34736,N_34057);
xor U35329 (N_35329,N_34167,N_34219);
xor U35330 (N_35330,N_34368,N_34555);
xnor U35331 (N_35331,N_34422,N_34982);
or U35332 (N_35332,N_34995,N_34669);
xnor U35333 (N_35333,N_34239,N_34685);
and U35334 (N_35334,N_34773,N_34570);
nand U35335 (N_35335,N_34829,N_34258);
nand U35336 (N_35336,N_34052,N_34308);
nor U35337 (N_35337,N_34211,N_34077);
nor U35338 (N_35338,N_34848,N_34860);
or U35339 (N_35339,N_34634,N_34818);
xor U35340 (N_35340,N_34072,N_34127);
nor U35341 (N_35341,N_34978,N_34558);
xnor U35342 (N_35342,N_34145,N_34241);
nand U35343 (N_35343,N_34817,N_34852);
or U35344 (N_35344,N_34274,N_34516);
nor U35345 (N_35345,N_34648,N_34686);
nor U35346 (N_35346,N_34247,N_34196);
or U35347 (N_35347,N_34392,N_34010);
nor U35348 (N_35348,N_34535,N_34678);
and U35349 (N_35349,N_34218,N_34967);
nand U35350 (N_35350,N_34513,N_34097);
xor U35351 (N_35351,N_34460,N_34245);
xnor U35352 (N_35352,N_34884,N_34079);
and U35353 (N_35353,N_34456,N_34132);
nor U35354 (N_35354,N_34944,N_34723);
or U35355 (N_35355,N_34844,N_34454);
and U35356 (N_35356,N_34785,N_34019);
or U35357 (N_35357,N_34408,N_34804);
nor U35358 (N_35358,N_34562,N_34377);
nand U35359 (N_35359,N_34909,N_34713);
nor U35360 (N_35360,N_34244,N_34796);
or U35361 (N_35361,N_34792,N_34913);
nor U35362 (N_35362,N_34627,N_34893);
xnor U35363 (N_35363,N_34912,N_34910);
and U35364 (N_35364,N_34998,N_34941);
xnor U35365 (N_35365,N_34715,N_34297);
nor U35366 (N_35366,N_34877,N_34521);
and U35367 (N_35367,N_34689,N_34647);
or U35368 (N_35368,N_34255,N_34157);
nor U35369 (N_35369,N_34243,N_34530);
nand U35370 (N_35370,N_34054,N_34349);
nand U35371 (N_35371,N_34256,N_34483);
and U35372 (N_35372,N_34319,N_34960);
and U35373 (N_35373,N_34955,N_34582);
nand U35374 (N_35374,N_34803,N_34021);
xnor U35375 (N_35375,N_34883,N_34128);
nand U35376 (N_35376,N_34747,N_34919);
xnor U35377 (N_35377,N_34165,N_34026);
and U35378 (N_35378,N_34906,N_34827);
or U35379 (N_35379,N_34355,N_34951);
xor U35380 (N_35380,N_34902,N_34894);
nor U35381 (N_35381,N_34706,N_34586);
xor U35382 (N_35382,N_34001,N_34904);
nor U35383 (N_35383,N_34071,N_34985);
or U35384 (N_35384,N_34472,N_34899);
xnor U35385 (N_35385,N_34122,N_34604);
nor U35386 (N_35386,N_34478,N_34708);
nand U35387 (N_35387,N_34573,N_34508);
and U35388 (N_35388,N_34631,N_34593);
nor U35389 (N_35389,N_34547,N_34741);
xnor U35390 (N_35390,N_34209,N_34859);
or U35391 (N_35391,N_34754,N_34976);
nand U35392 (N_35392,N_34600,N_34262);
nor U35393 (N_35393,N_34470,N_34189);
and U35394 (N_35394,N_34373,N_34979);
or U35395 (N_35395,N_34799,N_34981);
nand U35396 (N_35396,N_34159,N_34096);
nor U35397 (N_35397,N_34156,N_34350);
nor U35398 (N_35398,N_34080,N_34696);
and U35399 (N_35399,N_34321,N_34505);
nor U35400 (N_35400,N_34481,N_34565);
nand U35401 (N_35401,N_34285,N_34891);
nor U35402 (N_35402,N_34672,N_34580);
and U35403 (N_35403,N_34947,N_34284);
or U35404 (N_35404,N_34964,N_34563);
or U35405 (N_35405,N_34787,N_34857);
and U35406 (N_35406,N_34607,N_34801);
and U35407 (N_35407,N_34395,N_34150);
or U35408 (N_35408,N_34632,N_34346);
and U35409 (N_35409,N_34480,N_34281);
xor U35410 (N_35410,N_34994,N_34574);
nor U35411 (N_35411,N_34082,N_34942);
and U35412 (N_35412,N_34411,N_34692);
xnor U35413 (N_35413,N_34789,N_34725);
xor U35414 (N_35414,N_34389,N_34007);
and U35415 (N_35415,N_34236,N_34815);
xnor U35416 (N_35416,N_34410,N_34464);
or U35417 (N_35417,N_34874,N_34034);
and U35418 (N_35418,N_34687,N_34113);
nor U35419 (N_35419,N_34310,N_34533);
xnor U35420 (N_35420,N_34385,N_34131);
nand U35421 (N_35421,N_34544,N_34856);
and U35422 (N_35422,N_34053,N_34705);
nand U35423 (N_35423,N_34814,N_34645);
and U35424 (N_35424,N_34871,N_34020);
nor U35425 (N_35425,N_34084,N_34596);
or U35426 (N_35426,N_34611,N_34602);
xnor U35427 (N_35427,N_34610,N_34551);
nand U35428 (N_35428,N_34875,N_34658);
and U35429 (N_35429,N_34417,N_34074);
and U35430 (N_35430,N_34807,N_34069);
nand U35431 (N_35431,N_34748,N_34663);
xor U35432 (N_35432,N_34361,N_34469);
xor U35433 (N_35433,N_34822,N_34617);
xnor U35434 (N_35434,N_34635,N_34081);
nand U35435 (N_35435,N_34764,N_34268);
and U35436 (N_35436,N_34710,N_34181);
and U35437 (N_35437,N_34761,N_34387);
nand U35438 (N_35438,N_34677,N_34340);
and U35439 (N_35439,N_34657,N_34878);
xnor U35440 (N_35440,N_34169,N_34952);
and U35441 (N_35441,N_34873,N_34318);
and U35442 (N_35442,N_34772,N_34440);
or U35443 (N_35443,N_34732,N_34230);
xnor U35444 (N_35444,N_34584,N_34107);
or U35445 (N_35445,N_34364,N_34467);
and U35446 (N_35446,N_34024,N_34643);
xnor U35447 (N_35447,N_34820,N_34331);
and U35448 (N_35448,N_34092,N_34517);
or U35449 (N_35449,N_34895,N_34123);
xor U35450 (N_35450,N_34406,N_34583);
xor U35451 (N_35451,N_34048,N_34782);
or U35452 (N_35452,N_34067,N_34405);
and U35453 (N_35453,N_34751,N_34006);
xor U35454 (N_35454,N_34959,N_34641);
or U35455 (N_35455,N_34880,N_34419);
nand U35456 (N_35456,N_34058,N_34295);
nand U35457 (N_35457,N_34164,N_34423);
and U35458 (N_35458,N_34518,N_34898);
or U35459 (N_35459,N_34954,N_34329);
nand U35460 (N_35460,N_34929,N_34743);
or U35461 (N_35461,N_34496,N_34790);
xor U35462 (N_35462,N_34200,N_34711);
or U35463 (N_35463,N_34989,N_34506);
and U35464 (N_35464,N_34699,N_34485);
xnor U35465 (N_35465,N_34397,N_34291);
and U35466 (N_35466,N_34841,N_34847);
and U35467 (N_35467,N_34233,N_34185);
xnor U35468 (N_35468,N_34719,N_34865);
xor U35469 (N_35469,N_34564,N_34398);
or U35470 (N_35470,N_34542,N_34043);
nand U35471 (N_35471,N_34148,N_34745);
and U35472 (N_35472,N_34922,N_34940);
nor U35473 (N_35473,N_34466,N_34383);
and U35474 (N_35474,N_34652,N_34965);
xnor U35475 (N_35475,N_34928,N_34756);
or U35476 (N_35476,N_34830,N_34630);
nand U35477 (N_35477,N_34463,N_34056);
nand U35478 (N_35478,N_34038,N_34261);
nor U35479 (N_35479,N_34662,N_34146);
nand U35480 (N_35480,N_34881,N_34943);
or U35481 (N_35481,N_34358,N_34315);
xnor U35482 (N_35482,N_34855,N_34509);
nand U35483 (N_35483,N_34762,N_34490);
nand U35484 (N_35484,N_34046,N_34968);
nor U35485 (N_35485,N_34504,N_34037);
and U35486 (N_35486,N_34442,N_34655);
nand U35487 (N_35487,N_34462,N_34160);
nor U35488 (N_35488,N_34070,N_34594);
nor U35489 (N_35489,N_34458,N_34147);
nor U35490 (N_35490,N_34737,N_34568);
nor U35491 (N_35491,N_34118,N_34305);
nand U35492 (N_35492,N_34098,N_34612);
nor U35493 (N_35493,N_34609,N_34673);
nor U35494 (N_35494,N_34503,N_34343);
or U35495 (N_35495,N_34104,N_34571);
or U35496 (N_35496,N_34653,N_34900);
and U35497 (N_35497,N_34986,N_34091);
and U35498 (N_35498,N_34597,N_34154);
nand U35499 (N_35499,N_34776,N_34345);
or U35500 (N_35500,N_34574,N_34580);
xor U35501 (N_35501,N_34635,N_34510);
or U35502 (N_35502,N_34069,N_34854);
and U35503 (N_35503,N_34181,N_34405);
xnor U35504 (N_35504,N_34635,N_34646);
or U35505 (N_35505,N_34213,N_34427);
nand U35506 (N_35506,N_34558,N_34617);
and U35507 (N_35507,N_34790,N_34387);
or U35508 (N_35508,N_34820,N_34180);
nor U35509 (N_35509,N_34405,N_34772);
or U35510 (N_35510,N_34054,N_34360);
xor U35511 (N_35511,N_34930,N_34113);
and U35512 (N_35512,N_34963,N_34276);
nor U35513 (N_35513,N_34574,N_34736);
xnor U35514 (N_35514,N_34820,N_34989);
xor U35515 (N_35515,N_34704,N_34754);
and U35516 (N_35516,N_34322,N_34836);
or U35517 (N_35517,N_34584,N_34860);
xnor U35518 (N_35518,N_34787,N_34083);
nand U35519 (N_35519,N_34595,N_34453);
nor U35520 (N_35520,N_34287,N_34450);
or U35521 (N_35521,N_34195,N_34646);
nor U35522 (N_35522,N_34396,N_34093);
or U35523 (N_35523,N_34321,N_34622);
and U35524 (N_35524,N_34499,N_34562);
and U35525 (N_35525,N_34630,N_34133);
or U35526 (N_35526,N_34719,N_34057);
or U35527 (N_35527,N_34309,N_34844);
nand U35528 (N_35528,N_34298,N_34417);
or U35529 (N_35529,N_34866,N_34397);
nor U35530 (N_35530,N_34709,N_34970);
nand U35531 (N_35531,N_34036,N_34971);
and U35532 (N_35532,N_34166,N_34104);
nand U35533 (N_35533,N_34255,N_34085);
xor U35534 (N_35534,N_34037,N_34820);
nand U35535 (N_35535,N_34163,N_34740);
xnor U35536 (N_35536,N_34482,N_34400);
xnor U35537 (N_35537,N_34876,N_34721);
or U35538 (N_35538,N_34495,N_34572);
and U35539 (N_35539,N_34463,N_34364);
xor U35540 (N_35540,N_34325,N_34748);
xnor U35541 (N_35541,N_34170,N_34618);
nor U35542 (N_35542,N_34825,N_34641);
xnor U35543 (N_35543,N_34549,N_34508);
or U35544 (N_35544,N_34734,N_34599);
or U35545 (N_35545,N_34952,N_34721);
and U35546 (N_35546,N_34916,N_34941);
nor U35547 (N_35547,N_34829,N_34814);
and U35548 (N_35548,N_34195,N_34577);
or U35549 (N_35549,N_34810,N_34713);
and U35550 (N_35550,N_34614,N_34679);
or U35551 (N_35551,N_34265,N_34244);
or U35552 (N_35552,N_34814,N_34298);
xnor U35553 (N_35553,N_34561,N_34147);
and U35554 (N_35554,N_34363,N_34531);
or U35555 (N_35555,N_34883,N_34736);
and U35556 (N_35556,N_34715,N_34170);
xnor U35557 (N_35557,N_34974,N_34589);
nand U35558 (N_35558,N_34370,N_34794);
xor U35559 (N_35559,N_34735,N_34948);
or U35560 (N_35560,N_34577,N_34720);
or U35561 (N_35561,N_34031,N_34549);
or U35562 (N_35562,N_34394,N_34315);
or U35563 (N_35563,N_34383,N_34434);
nor U35564 (N_35564,N_34854,N_34922);
xnor U35565 (N_35565,N_34019,N_34928);
and U35566 (N_35566,N_34310,N_34724);
or U35567 (N_35567,N_34696,N_34538);
nor U35568 (N_35568,N_34925,N_34809);
xnor U35569 (N_35569,N_34778,N_34699);
xnor U35570 (N_35570,N_34021,N_34952);
or U35571 (N_35571,N_34320,N_34726);
or U35572 (N_35572,N_34061,N_34044);
nand U35573 (N_35573,N_34732,N_34728);
nand U35574 (N_35574,N_34709,N_34634);
and U35575 (N_35575,N_34194,N_34189);
xnor U35576 (N_35576,N_34007,N_34768);
nand U35577 (N_35577,N_34561,N_34189);
and U35578 (N_35578,N_34010,N_34787);
and U35579 (N_35579,N_34025,N_34132);
nand U35580 (N_35580,N_34393,N_34669);
or U35581 (N_35581,N_34792,N_34261);
nor U35582 (N_35582,N_34013,N_34266);
nor U35583 (N_35583,N_34980,N_34634);
or U35584 (N_35584,N_34681,N_34961);
or U35585 (N_35585,N_34991,N_34406);
nor U35586 (N_35586,N_34191,N_34892);
nand U35587 (N_35587,N_34854,N_34450);
xor U35588 (N_35588,N_34632,N_34024);
xor U35589 (N_35589,N_34032,N_34580);
nand U35590 (N_35590,N_34285,N_34102);
and U35591 (N_35591,N_34955,N_34072);
nor U35592 (N_35592,N_34375,N_34251);
and U35593 (N_35593,N_34266,N_34461);
xnor U35594 (N_35594,N_34652,N_34230);
and U35595 (N_35595,N_34382,N_34838);
or U35596 (N_35596,N_34776,N_34820);
nor U35597 (N_35597,N_34536,N_34361);
nor U35598 (N_35598,N_34435,N_34394);
nand U35599 (N_35599,N_34366,N_34315);
nand U35600 (N_35600,N_34504,N_34515);
nand U35601 (N_35601,N_34117,N_34177);
nor U35602 (N_35602,N_34573,N_34101);
xnor U35603 (N_35603,N_34500,N_34429);
nor U35604 (N_35604,N_34582,N_34519);
nor U35605 (N_35605,N_34876,N_34409);
and U35606 (N_35606,N_34542,N_34402);
nand U35607 (N_35607,N_34954,N_34743);
nand U35608 (N_35608,N_34314,N_34630);
or U35609 (N_35609,N_34875,N_34305);
nor U35610 (N_35610,N_34236,N_34984);
nand U35611 (N_35611,N_34247,N_34725);
and U35612 (N_35612,N_34085,N_34776);
and U35613 (N_35613,N_34598,N_34931);
nand U35614 (N_35614,N_34999,N_34418);
and U35615 (N_35615,N_34817,N_34381);
xnor U35616 (N_35616,N_34910,N_34150);
and U35617 (N_35617,N_34956,N_34885);
xor U35618 (N_35618,N_34734,N_34155);
or U35619 (N_35619,N_34923,N_34620);
nand U35620 (N_35620,N_34610,N_34384);
nor U35621 (N_35621,N_34515,N_34324);
or U35622 (N_35622,N_34136,N_34061);
and U35623 (N_35623,N_34801,N_34819);
xnor U35624 (N_35624,N_34078,N_34112);
and U35625 (N_35625,N_34792,N_34326);
or U35626 (N_35626,N_34029,N_34741);
nor U35627 (N_35627,N_34494,N_34570);
nand U35628 (N_35628,N_34640,N_34234);
nand U35629 (N_35629,N_34419,N_34223);
or U35630 (N_35630,N_34902,N_34713);
nand U35631 (N_35631,N_34653,N_34301);
or U35632 (N_35632,N_34929,N_34573);
or U35633 (N_35633,N_34431,N_34563);
and U35634 (N_35634,N_34245,N_34474);
xor U35635 (N_35635,N_34965,N_34873);
nand U35636 (N_35636,N_34355,N_34455);
nand U35637 (N_35637,N_34244,N_34874);
or U35638 (N_35638,N_34872,N_34236);
nor U35639 (N_35639,N_34203,N_34041);
nor U35640 (N_35640,N_34447,N_34646);
nor U35641 (N_35641,N_34354,N_34186);
or U35642 (N_35642,N_34829,N_34635);
nor U35643 (N_35643,N_34580,N_34262);
nand U35644 (N_35644,N_34358,N_34325);
xnor U35645 (N_35645,N_34116,N_34968);
or U35646 (N_35646,N_34829,N_34563);
or U35647 (N_35647,N_34966,N_34618);
nand U35648 (N_35648,N_34303,N_34889);
nand U35649 (N_35649,N_34971,N_34825);
nor U35650 (N_35650,N_34460,N_34006);
or U35651 (N_35651,N_34405,N_34607);
nand U35652 (N_35652,N_34390,N_34290);
and U35653 (N_35653,N_34395,N_34860);
or U35654 (N_35654,N_34547,N_34705);
xnor U35655 (N_35655,N_34985,N_34166);
and U35656 (N_35656,N_34430,N_34739);
and U35657 (N_35657,N_34643,N_34963);
and U35658 (N_35658,N_34676,N_34814);
nor U35659 (N_35659,N_34773,N_34981);
and U35660 (N_35660,N_34626,N_34402);
xnor U35661 (N_35661,N_34468,N_34686);
xor U35662 (N_35662,N_34062,N_34463);
xor U35663 (N_35663,N_34426,N_34298);
xor U35664 (N_35664,N_34288,N_34595);
xor U35665 (N_35665,N_34461,N_34753);
and U35666 (N_35666,N_34177,N_34164);
nand U35667 (N_35667,N_34805,N_34309);
and U35668 (N_35668,N_34915,N_34500);
and U35669 (N_35669,N_34873,N_34004);
nand U35670 (N_35670,N_34725,N_34121);
or U35671 (N_35671,N_34124,N_34047);
and U35672 (N_35672,N_34167,N_34614);
xor U35673 (N_35673,N_34001,N_34079);
and U35674 (N_35674,N_34456,N_34530);
nand U35675 (N_35675,N_34000,N_34708);
xnor U35676 (N_35676,N_34827,N_34847);
or U35677 (N_35677,N_34314,N_34586);
nor U35678 (N_35678,N_34813,N_34470);
and U35679 (N_35679,N_34555,N_34985);
and U35680 (N_35680,N_34847,N_34724);
and U35681 (N_35681,N_34557,N_34911);
nand U35682 (N_35682,N_34084,N_34691);
or U35683 (N_35683,N_34578,N_34108);
or U35684 (N_35684,N_34798,N_34853);
nor U35685 (N_35685,N_34350,N_34950);
nand U35686 (N_35686,N_34059,N_34647);
xor U35687 (N_35687,N_34171,N_34545);
xor U35688 (N_35688,N_34804,N_34861);
nor U35689 (N_35689,N_34570,N_34873);
nor U35690 (N_35690,N_34106,N_34627);
nand U35691 (N_35691,N_34563,N_34386);
xor U35692 (N_35692,N_34181,N_34009);
nand U35693 (N_35693,N_34267,N_34233);
nor U35694 (N_35694,N_34494,N_34223);
or U35695 (N_35695,N_34882,N_34484);
or U35696 (N_35696,N_34788,N_34604);
nand U35697 (N_35697,N_34247,N_34793);
and U35698 (N_35698,N_34477,N_34575);
nor U35699 (N_35699,N_34251,N_34282);
and U35700 (N_35700,N_34925,N_34354);
nor U35701 (N_35701,N_34840,N_34870);
nor U35702 (N_35702,N_34549,N_34423);
nand U35703 (N_35703,N_34706,N_34599);
or U35704 (N_35704,N_34000,N_34118);
xor U35705 (N_35705,N_34106,N_34954);
and U35706 (N_35706,N_34594,N_34496);
nor U35707 (N_35707,N_34346,N_34653);
or U35708 (N_35708,N_34088,N_34253);
or U35709 (N_35709,N_34098,N_34173);
nor U35710 (N_35710,N_34626,N_34271);
and U35711 (N_35711,N_34495,N_34887);
and U35712 (N_35712,N_34861,N_34751);
nand U35713 (N_35713,N_34979,N_34870);
nor U35714 (N_35714,N_34111,N_34274);
nor U35715 (N_35715,N_34399,N_34512);
nor U35716 (N_35716,N_34675,N_34192);
or U35717 (N_35717,N_34753,N_34098);
or U35718 (N_35718,N_34754,N_34707);
nand U35719 (N_35719,N_34755,N_34041);
nor U35720 (N_35720,N_34799,N_34721);
nor U35721 (N_35721,N_34485,N_34042);
or U35722 (N_35722,N_34888,N_34597);
nor U35723 (N_35723,N_34356,N_34436);
nand U35724 (N_35724,N_34591,N_34759);
nor U35725 (N_35725,N_34913,N_34147);
or U35726 (N_35726,N_34518,N_34992);
nor U35727 (N_35727,N_34383,N_34993);
nor U35728 (N_35728,N_34262,N_34271);
nand U35729 (N_35729,N_34304,N_34096);
nor U35730 (N_35730,N_34425,N_34142);
nand U35731 (N_35731,N_34123,N_34235);
and U35732 (N_35732,N_34279,N_34699);
and U35733 (N_35733,N_34869,N_34114);
and U35734 (N_35734,N_34623,N_34929);
and U35735 (N_35735,N_34011,N_34434);
or U35736 (N_35736,N_34526,N_34146);
nor U35737 (N_35737,N_34438,N_34168);
and U35738 (N_35738,N_34954,N_34968);
and U35739 (N_35739,N_34060,N_34269);
xnor U35740 (N_35740,N_34341,N_34778);
xor U35741 (N_35741,N_34434,N_34734);
and U35742 (N_35742,N_34083,N_34856);
nor U35743 (N_35743,N_34372,N_34681);
and U35744 (N_35744,N_34434,N_34420);
nor U35745 (N_35745,N_34722,N_34066);
and U35746 (N_35746,N_34128,N_34691);
xnor U35747 (N_35747,N_34675,N_34625);
xor U35748 (N_35748,N_34091,N_34747);
or U35749 (N_35749,N_34957,N_34521);
nand U35750 (N_35750,N_34607,N_34170);
and U35751 (N_35751,N_34077,N_34923);
xnor U35752 (N_35752,N_34193,N_34933);
nor U35753 (N_35753,N_34726,N_34060);
and U35754 (N_35754,N_34443,N_34322);
or U35755 (N_35755,N_34498,N_34789);
nor U35756 (N_35756,N_34634,N_34292);
or U35757 (N_35757,N_34959,N_34590);
nand U35758 (N_35758,N_34469,N_34378);
or U35759 (N_35759,N_34727,N_34993);
and U35760 (N_35760,N_34111,N_34222);
nand U35761 (N_35761,N_34520,N_34907);
xnor U35762 (N_35762,N_34087,N_34436);
xnor U35763 (N_35763,N_34325,N_34028);
or U35764 (N_35764,N_34301,N_34084);
or U35765 (N_35765,N_34563,N_34989);
xnor U35766 (N_35766,N_34690,N_34902);
or U35767 (N_35767,N_34394,N_34928);
nor U35768 (N_35768,N_34863,N_34666);
or U35769 (N_35769,N_34984,N_34686);
nor U35770 (N_35770,N_34152,N_34716);
xor U35771 (N_35771,N_34238,N_34925);
or U35772 (N_35772,N_34987,N_34087);
nand U35773 (N_35773,N_34378,N_34744);
nand U35774 (N_35774,N_34856,N_34589);
xor U35775 (N_35775,N_34584,N_34926);
nor U35776 (N_35776,N_34042,N_34300);
nor U35777 (N_35777,N_34407,N_34761);
and U35778 (N_35778,N_34282,N_34792);
xnor U35779 (N_35779,N_34713,N_34354);
nor U35780 (N_35780,N_34279,N_34959);
and U35781 (N_35781,N_34820,N_34182);
or U35782 (N_35782,N_34740,N_34677);
and U35783 (N_35783,N_34222,N_34269);
or U35784 (N_35784,N_34562,N_34180);
nand U35785 (N_35785,N_34884,N_34133);
or U35786 (N_35786,N_34935,N_34163);
nand U35787 (N_35787,N_34129,N_34839);
or U35788 (N_35788,N_34011,N_34883);
xor U35789 (N_35789,N_34029,N_34023);
and U35790 (N_35790,N_34825,N_34094);
nor U35791 (N_35791,N_34937,N_34085);
xnor U35792 (N_35792,N_34292,N_34989);
or U35793 (N_35793,N_34723,N_34476);
and U35794 (N_35794,N_34889,N_34933);
and U35795 (N_35795,N_34855,N_34801);
or U35796 (N_35796,N_34714,N_34603);
nor U35797 (N_35797,N_34625,N_34365);
xor U35798 (N_35798,N_34230,N_34492);
nor U35799 (N_35799,N_34546,N_34107);
nor U35800 (N_35800,N_34457,N_34666);
nand U35801 (N_35801,N_34647,N_34959);
or U35802 (N_35802,N_34272,N_34243);
xnor U35803 (N_35803,N_34147,N_34937);
and U35804 (N_35804,N_34656,N_34464);
or U35805 (N_35805,N_34145,N_34032);
and U35806 (N_35806,N_34691,N_34558);
nand U35807 (N_35807,N_34204,N_34028);
and U35808 (N_35808,N_34218,N_34541);
nor U35809 (N_35809,N_34102,N_34563);
nand U35810 (N_35810,N_34782,N_34336);
or U35811 (N_35811,N_34526,N_34073);
or U35812 (N_35812,N_34028,N_34663);
and U35813 (N_35813,N_34484,N_34530);
nand U35814 (N_35814,N_34546,N_34418);
and U35815 (N_35815,N_34297,N_34106);
and U35816 (N_35816,N_34237,N_34426);
and U35817 (N_35817,N_34234,N_34831);
nand U35818 (N_35818,N_34110,N_34709);
nor U35819 (N_35819,N_34007,N_34764);
nand U35820 (N_35820,N_34934,N_34339);
xor U35821 (N_35821,N_34137,N_34790);
or U35822 (N_35822,N_34833,N_34836);
nor U35823 (N_35823,N_34962,N_34209);
xnor U35824 (N_35824,N_34021,N_34343);
nand U35825 (N_35825,N_34641,N_34924);
nand U35826 (N_35826,N_34204,N_34338);
or U35827 (N_35827,N_34311,N_34025);
nand U35828 (N_35828,N_34680,N_34869);
nor U35829 (N_35829,N_34461,N_34819);
nor U35830 (N_35830,N_34325,N_34634);
nand U35831 (N_35831,N_34583,N_34992);
nand U35832 (N_35832,N_34629,N_34204);
or U35833 (N_35833,N_34936,N_34885);
or U35834 (N_35834,N_34114,N_34588);
nand U35835 (N_35835,N_34347,N_34956);
or U35836 (N_35836,N_34639,N_34437);
xor U35837 (N_35837,N_34629,N_34220);
nand U35838 (N_35838,N_34183,N_34434);
nand U35839 (N_35839,N_34556,N_34974);
nand U35840 (N_35840,N_34590,N_34106);
xnor U35841 (N_35841,N_34382,N_34215);
nand U35842 (N_35842,N_34251,N_34087);
nand U35843 (N_35843,N_34242,N_34988);
nor U35844 (N_35844,N_34516,N_34561);
and U35845 (N_35845,N_34455,N_34963);
and U35846 (N_35846,N_34233,N_34510);
or U35847 (N_35847,N_34406,N_34327);
or U35848 (N_35848,N_34089,N_34034);
nand U35849 (N_35849,N_34057,N_34462);
nand U35850 (N_35850,N_34785,N_34557);
and U35851 (N_35851,N_34497,N_34291);
or U35852 (N_35852,N_34289,N_34323);
xnor U35853 (N_35853,N_34064,N_34116);
and U35854 (N_35854,N_34254,N_34935);
xnor U35855 (N_35855,N_34519,N_34765);
and U35856 (N_35856,N_34978,N_34231);
xnor U35857 (N_35857,N_34484,N_34390);
or U35858 (N_35858,N_34331,N_34510);
or U35859 (N_35859,N_34024,N_34502);
nor U35860 (N_35860,N_34509,N_34295);
or U35861 (N_35861,N_34177,N_34634);
nand U35862 (N_35862,N_34051,N_34271);
or U35863 (N_35863,N_34128,N_34790);
nand U35864 (N_35864,N_34368,N_34201);
and U35865 (N_35865,N_34371,N_34128);
nor U35866 (N_35866,N_34867,N_34336);
and U35867 (N_35867,N_34916,N_34416);
or U35868 (N_35868,N_34976,N_34045);
nand U35869 (N_35869,N_34492,N_34085);
nand U35870 (N_35870,N_34688,N_34297);
or U35871 (N_35871,N_34019,N_34820);
and U35872 (N_35872,N_34465,N_34173);
nand U35873 (N_35873,N_34878,N_34970);
nor U35874 (N_35874,N_34858,N_34451);
nor U35875 (N_35875,N_34300,N_34185);
nor U35876 (N_35876,N_34342,N_34321);
and U35877 (N_35877,N_34426,N_34689);
nor U35878 (N_35878,N_34612,N_34509);
or U35879 (N_35879,N_34698,N_34477);
xor U35880 (N_35880,N_34103,N_34440);
or U35881 (N_35881,N_34399,N_34258);
nor U35882 (N_35882,N_34814,N_34779);
xnor U35883 (N_35883,N_34233,N_34040);
and U35884 (N_35884,N_34360,N_34091);
nand U35885 (N_35885,N_34979,N_34467);
or U35886 (N_35886,N_34021,N_34123);
nand U35887 (N_35887,N_34195,N_34149);
nand U35888 (N_35888,N_34821,N_34681);
nand U35889 (N_35889,N_34451,N_34674);
nor U35890 (N_35890,N_34917,N_34827);
or U35891 (N_35891,N_34009,N_34560);
nand U35892 (N_35892,N_34265,N_34471);
xnor U35893 (N_35893,N_34326,N_34457);
or U35894 (N_35894,N_34908,N_34913);
xnor U35895 (N_35895,N_34799,N_34962);
or U35896 (N_35896,N_34597,N_34645);
nand U35897 (N_35897,N_34785,N_34987);
nand U35898 (N_35898,N_34283,N_34282);
or U35899 (N_35899,N_34482,N_34292);
nand U35900 (N_35900,N_34249,N_34030);
nand U35901 (N_35901,N_34074,N_34361);
nand U35902 (N_35902,N_34741,N_34203);
or U35903 (N_35903,N_34201,N_34497);
xor U35904 (N_35904,N_34128,N_34846);
nor U35905 (N_35905,N_34333,N_34071);
nand U35906 (N_35906,N_34400,N_34782);
nand U35907 (N_35907,N_34854,N_34967);
nor U35908 (N_35908,N_34283,N_34193);
nand U35909 (N_35909,N_34012,N_34902);
or U35910 (N_35910,N_34223,N_34653);
nand U35911 (N_35911,N_34181,N_34016);
or U35912 (N_35912,N_34730,N_34671);
xor U35913 (N_35913,N_34359,N_34528);
and U35914 (N_35914,N_34063,N_34065);
and U35915 (N_35915,N_34534,N_34040);
xor U35916 (N_35916,N_34940,N_34139);
nor U35917 (N_35917,N_34264,N_34300);
nand U35918 (N_35918,N_34142,N_34857);
and U35919 (N_35919,N_34831,N_34550);
nor U35920 (N_35920,N_34423,N_34032);
nor U35921 (N_35921,N_34007,N_34513);
nand U35922 (N_35922,N_34140,N_34505);
nor U35923 (N_35923,N_34236,N_34341);
nand U35924 (N_35924,N_34685,N_34286);
nor U35925 (N_35925,N_34117,N_34968);
and U35926 (N_35926,N_34521,N_34229);
and U35927 (N_35927,N_34938,N_34927);
and U35928 (N_35928,N_34790,N_34404);
nand U35929 (N_35929,N_34408,N_34034);
nor U35930 (N_35930,N_34347,N_34875);
xor U35931 (N_35931,N_34648,N_34685);
nand U35932 (N_35932,N_34173,N_34292);
nand U35933 (N_35933,N_34546,N_34419);
nand U35934 (N_35934,N_34351,N_34647);
xnor U35935 (N_35935,N_34391,N_34193);
or U35936 (N_35936,N_34285,N_34163);
xnor U35937 (N_35937,N_34534,N_34876);
xnor U35938 (N_35938,N_34359,N_34221);
nor U35939 (N_35939,N_34667,N_34996);
nand U35940 (N_35940,N_34673,N_34975);
xnor U35941 (N_35941,N_34120,N_34706);
nor U35942 (N_35942,N_34942,N_34002);
xnor U35943 (N_35943,N_34582,N_34296);
xnor U35944 (N_35944,N_34798,N_34165);
and U35945 (N_35945,N_34266,N_34732);
xnor U35946 (N_35946,N_34540,N_34862);
or U35947 (N_35947,N_34224,N_34343);
or U35948 (N_35948,N_34739,N_34462);
xor U35949 (N_35949,N_34429,N_34487);
and U35950 (N_35950,N_34852,N_34339);
nand U35951 (N_35951,N_34620,N_34601);
nor U35952 (N_35952,N_34588,N_34304);
xnor U35953 (N_35953,N_34403,N_34425);
and U35954 (N_35954,N_34262,N_34627);
nor U35955 (N_35955,N_34083,N_34311);
nor U35956 (N_35956,N_34726,N_34951);
and U35957 (N_35957,N_34191,N_34153);
or U35958 (N_35958,N_34375,N_34817);
and U35959 (N_35959,N_34052,N_34984);
nor U35960 (N_35960,N_34360,N_34508);
nor U35961 (N_35961,N_34684,N_34362);
nor U35962 (N_35962,N_34624,N_34982);
nand U35963 (N_35963,N_34157,N_34338);
nand U35964 (N_35964,N_34712,N_34104);
or U35965 (N_35965,N_34973,N_34136);
and U35966 (N_35966,N_34790,N_34785);
or U35967 (N_35967,N_34374,N_34322);
and U35968 (N_35968,N_34435,N_34668);
nand U35969 (N_35969,N_34445,N_34698);
nor U35970 (N_35970,N_34631,N_34242);
or U35971 (N_35971,N_34382,N_34272);
nor U35972 (N_35972,N_34534,N_34411);
nand U35973 (N_35973,N_34252,N_34163);
nor U35974 (N_35974,N_34605,N_34883);
or U35975 (N_35975,N_34432,N_34659);
nand U35976 (N_35976,N_34424,N_34759);
nor U35977 (N_35977,N_34864,N_34730);
xor U35978 (N_35978,N_34428,N_34951);
and U35979 (N_35979,N_34846,N_34611);
xor U35980 (N_35980,N_34841,N_34395);
nand U35981 (N_35981,N_34548,N_34801);
or U35982 (N_35982,N_34602,N_34737);
nand U35983 (N_35983,N_34177,N_34956);
nand U35984 (N_35984,N_34651,N_34322);
and U35985 (N_35985,N_34751,N_34788);
nand U35986 (N_35986,N_34492,N_34203);
or U35987 (N_35987,N_34997,N_34506);
or U35988 (N_35988,N_34183,N_34437);
or U35989 (N_35989,N_34028,N_34754);
nor U35990 (N_35990,N_34809,N_34669);
and U35991 (N_35991,N_34431,N_34955);
xnor U35992 (N_35992,N_34094,N_34637);
nand U35993 (N_35993,N_34952,N_34230);
xor U35994 (N_35994,N_34924,N_34727);
and U35995 (N_35995,N_34673,N_34375);
or U35996 (N_35996,N_34943,N_34415);
xor U35997 (N_35997,N_34945,N_34016);
nor U35998 (N_35998,N_34466,N_34916);
or U35999 (N_35999,N_34619,N_34051);
or U36000 (N_36000,N_35671,N_35912);
and U36001 (N_36001,N_35449,N_35651);
and U36002 (N_36002,N_35828,N_35756);
nand U36003 (N_36003,N_35321,N_35084);
nor U36004 (N_36004,N_35182,N_35240);
nor U36005 (N_36005,N_35626,N_35409);
xor U36006 (N_36006,N_35832,N_35101);
nand U36007 (N_36007,N_35502,N_35247);
or U36008 (N_36008,N_35676,N_35166);
nand U36009 (N_36009,N_35578,N_35752);
or U36010 (N_36010,N_35083,N_35538);
nor U36011 (N_36011,N_35356,N_35929);
xnor U36012 (N_36012,N_35076,N_35318);
or U36013 (N_36013,N_35085,N_35117);
and U36014 (N_36014,N_35373,N_35993);
or U36015 (N_36015,N_35333,N_35021);
xor U36016 (N_36016,N_35557,N_35797);
nor U36017 (N_36017,N_35881,N_35453);
xnor U36018 (N_36018,N_35906,N_35656);
and U36019 (N_36019,N_35150,N_35174);
and U36020 (N_36020,N_35282,N_35505);
and U36021 (N_36021,N_35307,N_35000);
and U36022 (N_36022,N_35404,N_35056);
nor U36023 (N_36023,N_35726,N_35209);
nand U36024 (N_36024,N_35919,N_35283);
nor U36025 (N_36025,N_35062,N_35996);
nand U36026 (N_36026,N_35067,N_35214);
xor U36027 (N_36027,N_35904,N_35415);
nand U36028 (N_36028,N_35312,N_35138);
and U36029 (N_36029,N_35611,N_35025);
nand U36030 (N_36030,N_35670,N_35364);
nand U36031 (N_36031,N_35794,N_35679);
and U36032 (N_36032,N_35571,N_35770);
and U36033 (N_36033,N_35090,N_35535);
nor U36034 (N_36034,N_35091,N_35457);
or U36035 (N_36035,N_35329,N_35494);
xor U36036 (N_36036,N_35274,N_35830);
xnor U36037 (N_36037,N_35099,N_35965);
xor U36038 (N_36038,N_35521,N_35545);
or U36039 (N_36039,N_35880,N_35028);
nor U36040 (N_36040,N_35530,N_35582);
and U36041 (N_36041,N_35336,N_35779);
xor U36042 (N_36042,N_35745,N_35501);
nor U36043 (N_36043,N_35314,N_35115);
nand U36044 (N_36044,N_35600,N_35735);
or U36045 (N_36045,N_35599,N_35682);
nor U36046 (N_36046,N_35562,N_35456);
nor U36047 (N_36047,N_35143,N_35662);
or U36048 (N_36048,N_35232,N_35548);
and U36049 (N_36049,N_35528,N_35660);
and U36050 (N_36050,N_35144,N_35591);
nor U36051 (N_36051,N_35402,N_35430);
nor U36052 (N_36052,N_35332,N_35434);
nand U36053 (N_36053,N_35316,N_35390);
xor U36054 (N_36054,N_35771,N_35086);
nand U36055 (N_36055,N_35211,N_35948);
xor U36056 (N_36056,N_35933,N_35720);
xor U36057 (N_36057,N_35026,N_35495);
xor U36058 (N_36058,N_35552,N_35903);
or U36059 (N_36059,N_35053,N_35196);
xnor U36060 (N_36060,N_35672,N_35173);
or U36061 (N_36061,N_35969,N_35864);
or U36062 (N_36062,N_35338,N_35098);
nand U36063 (N_36063,N_35841,N_35048);
and U36064 (N_36064,N_35829,N_35259);
or U36065 (N_36065,N_35280,N_35825);
nor U36066 (N_36066,N_35287,N_35382);
or U36067 (N_36067,N_35536,N_35376);
xnor U36068 (N_36068,N_35069,N_35826);
nand U36069 (N_36069,N_35616,N_35399);
xnor U36070 (N_36070,N_35709,N_35315);
xnor U36071 (N_36071,N_35947,N_35408);
and U36072 (N_36072,N_35435,N_35856);
nor U36073 (N_36073,N_35303,N_35849);
or U36074 (N_36074,N_35284,N_35928);
or U36075 (N_36075,N_35313,N_35732);
and U36076 (N_36076,N_35576,N_35942);
nor U36077 (N_36077,N_35954,N_35890);
xnor U36078 (N_36078,N_35967,N_35210);
nor U36079 (N_36079,N_35386,N_35328);
or U36080 (N_36080,N_35568,N_35186);
xor U36081 (N_36081,N_35717,N_35116);
xor U36082 (N_36082,N_35515,N_35573);
and U36083 (N_36083,N_35847,N_35747);
or U36084 (N_36084,N_35995,N_35853);
xor U36085 (N_36085,N_35987,N_35788);
and U36086 (N_36086,N_35234,N_35131);
and U36087 (N_36087,N_35029,N_35020);
and U36088 (N_36088,N_35251,N_35135);
or U36089 (N_36089,N_35127,N_35882);
xor U36090 (N_36090,N_35989,N_35913);
nor U36091 (N_36091,N_35721,N_35862);
and U36092 (N_36092,N_35191,N_35613);
nor U36093 (N_36093,N_35711,N_35347);
xor U36094 (N_36094,N_35877,N_35057);
and U36095 (N_36095,N_35815,N_35510);
nor U36096 (N_36096,N_35664,N_35237);
and U36097 (N_36097,N_35041,N_35524);
and U36098 (N_36098,N_35963,N_35052);
nand U36099 (N_36099,N_35397,N_35661);
nor U36100 (N_36100,N_35908,N_35991);
or U36101 (N_36101,N_35139,N_35132);
or U36102 (N_36102,N_35629,N_35035);
xnor U36103 (N_36103,N_35219,N_35221);
and U36104 (N_36104,N_35990,N_35097);
nor U36105 (N_36105,N_35750,N_35407);
or U36106 (N_36106,N_35394,N_35270);
and U36107 (N_36107,N_35520,N_35128);
xor U36108 (N_36108,N_35612,N_35032);
xnor U36109 (N_36109,N_35644,N_35622);
nand U36110 (N_36110,N_35901,N_35044);
and U36111 (N_36111,N_35839,N_35134);
xor U36112 (N_36112,N_35248,N_35137);
nand U36113 (N_36113,N_35759,N_35066);
nor U36114 (N_36114,N_35850,N_35125);
xnor U36115 (N_36115,N_35767,N_35869);
nor U36116 (N_36116,N_35961,N_35884);
nor U36117 (N_36117,N_35840,N_35631);
or U36118 (N_36118,N_35722,N_35206);
nand U36119 (N_36119,N_35061,N_35851);
or U36120 (N_36120,N_35891,N_35606);
nor U36121 (N_36121,N_35045,N_35590);
nor U36122 (N_36122,N_35075,N_35485);
nor U36123 (N_36123,N_35204,N_35027);
or U36124 (N_36124,N_35892,N_35741);
nand U36125 (N_36125,N_35413,N_35843);
nor U36126 (N_36126,N_35202,N_35439);
or U36127 (N_36127,N_35162,N_35569);
xor U36128 (N_36128,N_35030,N_35320);
or U36129 (N_36129,N_35130,N_35774);
xnor U36130 (N_36130,N_35384,N_35179);
nand U36131 (N_36131,N_35738,N_35419);
xor U36132 (N_36132,N_35441,N_35959);
and U36133 (N_36133,N_35362,N_35970);
and U36134 (N_36134,N_35063,N_35498);
nor U36135 (N_36135,N_35658,N_35366);
xor U36136 (N_36136,N_35950,N_35807);
and U36137 (N_36137,N_35700,N_35277);
nand U36138 (N_36138,N_35295,N_35380);
nand U36139 (N_36139,N_35769,N_35411);
and U36140 (N_36140,N_35563,N_35178);
and U36141 (N_36141,N_35955,N_35418);
and U36142 (N_36142,N_35523,N_35089);
nand U36143 (N_36143,N_35454,N_35565);
nor U36144 (N_36144,N_35760,N_35707);
or U36145 (N_36145,N_35768,N_35058);
nor U36146 (N_36146,N_35688,N_35713);
nor U36147 (N_36147,N_35640,N_35647);
nand U36148 (N_36148,N_35633,N_35715);
and U36149 (N_36149,N_35653,N_35118);
xnor U36150 (N_36150,N_35164,N_35425);
and U36151 (N_36151,N_35437,N_35823);
and U36152 (N_36152,N_35152,N_35648);
or U36153 (N_36153,N_35790,N_35155);
and U36154 (N_36154,N_35059,N_35055);
nand U36155 (N_36155,N_35281,N_35291);
and U36156 (N_36156,N_35911,N_35801);
xor U36157 (N_36157,N_35226,N_35780);
nand U36158 (N_36158,N_35577,N_35699);
nor U36159 (N_36159,N_35141,N_35817);
xnor U36160 (N_36160,N_35852,N_35541);
or U36161 (N_36161,N_35123,N_35938);
xor U36162 (N_36162,N_35215,N_35657);
nor U36163 (N_36163,N_35529,N_35039);
xor U36164 (N_36164,N_35249,N_35385);
nor U36165 (N_36165,N_35940,N_35533);
nand U36166 (N_36166,N_35263,N_35952);
nor U36167 (N_36167,N_35188,N_35345);
nor U36168 (N_36168,N_35575,N_35836);
nand U36169 (N_36169,N_35806,N_35939);
and U36170 (N_36170,N_35690,N_35739);
or U36171 (N_36171,N_35875,N_35354);
nand U36172 (N_36172,N_35496,N_35238);
xor U36173 (N_36173,N_35513,N_35918);
xor U36174 (N_36174,N_35398,N_35532);
xnor U36175 (N_36175,N_35983,N_35956);
nor U36176 (N_36176,N_35223,N_35558);
or U36177 (N_36177,N_35669,N_35924);
and U36178 (N_36178,N_35006,N_35725);
or U36179 (N_36179,N_35213,N_35714);
and U36180 (N_36180,N_35073,N_35728);
xnor U36181 (N_36181,N_35666,N_35325);
and U36182 (N_36182,N_35848,N_35698);
nor U36183 (N_36183,N_35466,N_35033);
xor U36184 (N_36184,N_35620,N_35153);
nand U36185 (N_36185,N_35710,N_35391);
nor U36186 (N_36186,N_35289,N_35412);
nand U36187 (N_36187,N_35842,N_35811);
and U36188 (N_36188,N_35833,N_35361);
xnor U36189 (N_36189,N_35465,N_35450);
xnor U36190 (N_36190,N_35685,N_35821);
and U36191 (N_36191,N_35550,N_35646);
nor U36192 (N_36192,N_35190,N_35812);
and U36193 (N_36193,N_35865,N_35471);
xnor U36194 (N_36194,N_35697,N_35224);
or U36195 (N_36195,N_35844,N_35203);
nor U36196 (N_36196,N_35427,N_35317);
or U36197 (N_36197,N_35497,N_35870);
xor U36198 (N_36198,N_35013,N_35043);
or U36199 (N_36199,N_35945,N_35899);
nand U36200 (N_36200,N_35922,N_35478);
and U36201 (N_36201,N_35953,N_35677);
nor U36202 (N_36202,N_35740,N_35334);
xor U36203 (N_36203,N_35617,N_35252);
nand U36204 (N_36204,N_35424,N_35159);
xnor U36205 (N_36205,N_35151,N_35476);
xnor U36206 (N_36206,N_35936,N_35477);
and U36207 (N_36207,N_35293,N_35292);
nor U36208 (N_36208,N_35860,N_35507);
or U36209 (N_36209,N_35448,N_35786);
and U36210 (N_36210,N_35587,N_35614);
xor U36211 (N_36211,N_35262,N_35019);
nand U36212 (N_36212,N_35663,N_35369);
xnor U36213 (N_36213,N_35623,N_35866);
nand U36214 (N_36214,N_35094,N_35193);
nand U36215 (N_36215,N_35349,N_35440);
nor U36216 (N_36216,N_35584,N_35250);
xnor U36217 (N_36217,N_35265,N_35119);
xor U36218 (N_36218,N_35944,N_35683);
or U36219 (N_36219,N_35773,N_35642);
nand U36220 (N_36220,N_35235,N_35170);
or U36221 (N_36221,N_35375,N_35181);
or U36222 (N_36222,N_35225,N_35493);
or U36223 (N_36223,N_35500,N_35158);
nand U36224 (N_36224,N_35136,N_35286);
nor U36225 (N_36225,N_35167,N_35042);
xor U36226 (N_36226,N_35988,N_35298);
xnor U36227 (N_36227,N_35005,N_35087);
nand U36228 (N_36228,N_35619,N_35464);
nor U36229 (N_36229,N_35808,N_35346);
and U36230 (N_36230,N_35517,N_35652);
xor U36231 (N_36231,N_35926,N_35737);
or U36232 (N_36232,N_35161,N_35288);
and U36233 (N_36233,N_35992,N_35570);
or U36234 (N_36234,N_35560,N_35207);
and U36235 (N_36235,N_35932,N_35696);
nor U36236 (N_36236,N_35896,N_35960);
or U36237 (N_36237,N_35290,N_35650);
nor U36238 (N_36238,N_35754,N_35104);
nor U36239 (N_36239,N_35330,N_35074);
xor U36240 (N_36240,N_35574,N_35596);
nand U36241 (N_36241,N_35719,N_35949);
or U36242 (N_36242,N_35300,N_35145);
and U36243 (N_36243,N_35986,N_35387);
nor U36244 (N_36244,N_35337,N_35004);
nor U36245 (N_36245,N_35475,N_35902);
xnor U36246 (N_36246,N_35879,N_35302);
nor U36247 (N_36247,N_35031,N_35327);
nand U36248 (N_36248,N_35508,N_35766);
and U36249 (N_36249,N_35294,N_35267);
and U36250 (N_36250,N_35659,N_35064);
nand U36251 (N_36251,N_35798,N_35079);
nand U36252 (N_36252,N_35935,N_35703);
nor U36253 (N_36253,N_35597,N_35050);
xnor U36254 (N_36254,N_35443,N_35863);
and U36255 (N_36255,N_35762,N_35023);
or U36256 (N_36256,N_35389,N_35757);
or U36257 (N_36257,N_35093,N_35858);
or U36258 (N_36258,N_35499,N_35637);
or U36259 (N_36259,N_35442,N_35635);
and U36260 (N_36260,N_35242,N_35705);
xor U36261 (N_36261,N_35110,N_35914);
or U36262 (N_36262,N_35377,N_35257);
and U36263 (N_36263,N_35702,N_35553);
nand U36264 (N_36264,N_35680,N_35810);
nand U36265 (N_36265,N_35789,N_35572);
and U36266 (N_36266,N_35800,N_35095);
or U36267 (N_36267,N_35183,N_35506);
and U36268 (N_36268,N_35352,N_35105);
nor U36269 (N_36269,N_35783,N_35339);
xnor U36270 (N_36270,N_35446,N_35589);
xnor U36271 (N_36271,N_35372,N_35514);
or U36272 (N_36272,N_35731,N_35433);
xnor U36273 (N_36273,N_35201,N_35615);
nor U36274 (N_36274,N_35925,N_35859);
or U36275 (N_36275,N_35973,N_35871);
xnor U36276 (N_36276,N_35078,N_35420);
nand U36277 (N_36277,N_35855,N_35835);
and U36278 (N_36278,N_35649,N_35736);
or U36279 (N_36279,N_35689,N_35943);
xnor U36280 (N_36280,N_35684,N_35421);
xor U36281 (N_36281,N_35194,N_35486);
or U36282 (N_36282,N_35579,N_35205);
nand U36283 (N_36283,N_35460,N_35168);
or U36284 (N_36284,N_35272,N_35586);
and U36285 (N_36285,N_35968,N_35872);
or U36286 (N_36286,N_35604,N_35687);
nor U36287 (N_36287,N_35245,N_35804);
xor U36288 (N_36288,N_35701,N_35624);
xnor U36289 (N_36289,N_35941,N_35231);
or U36290 (N_36290,N_35716,N_35822);
and U36291 (N_36291,N_35378,N_35217);
and U36292 (N_36292,N_35357,N_35814);
or U36293 (N_36293,N_35764,N_35876);
and U36294 (N_36294,N_35326,N_35392);
or U36295 (N_36295,N_35997,N_35921);
xor U36296 (N_36296,N_35775,N_35018);
xor U36297 (N_36297,N_35483,N_35365);
or U36298 (N_36298,N_35522,N_35894);
and U36299 (N_36299,N_35371,N_35883);
nand U36300 (N_36300,N_35962,N_35278);
xor U36301 (N_36301,N_35895,N_35241);
nand U36302 (N_36302,N_35103,N_35343);
xor U36303 (N_36303,N_35200,N_35243);
nor U36304 (N_36304,N_35975,N_35037);
or U36305 (N_36305,N_35239,N_35539);
nor U36306 (N_36306,N_35212,N_35889);
nand U36307 (N_36307,N_35793,N_35383);
and U36308 (N_36308,N_35544,N_35484);
nand U36309 (N_36309,N_35423,N_35070);
nand U36310 (N_36310,N_35022,N_35400);
or U36311 (N_36311,N_35791,N_35742);
xor U36312 (N_36312,N_35627,N_35395);
xnor U36313 (N_36313,N_35445,N_35729);
xor U36314 (N_36314,N_35393,N_35479);
or U36315 (N_36315,N_35998,N_35342);
nor U36316 (N_36316,N_35751,N_35208);
nor U36317 (N_36317,N_35305,N_35567);
xnor U36318 (N_36318,N_35082,N_35236);
xnor U36319 (N_36319,N_35838,N_35175);
nand U36320 (N_36320,N_35309,N_35566);
and U36321 (N_36321,N_35628,N_35490);
nand U36322 (N_36322,N_35379,N_35422);
or U36323 (N_36323,N_35598,N_35675);
nand U36324 (N_36324,N_35813,N_35630);
xor U36325 (N_36325,N_35581,N_35778);
or U36326 (N_36326,N_35189,N_35096);
nand U36327 (N_36327,N_35681,N_35546);
and U36328 (N_36328,N_35639,N_35358);
nor U36329 (N_36329,N_35163,N_35192);
nor U36330 (N_36330,N_35142,N_35543);
or U36331 (N_36331,N_35708,N_35003);
nand U36332 (N_36332,N_35228,N_35857);
or U36333 (N_36333,N_35165,N_35916);
and U36334 (N_36334,N_35081,N_35451);
and U36335 (N_36335,N_35481,N_35010);
xor U36336 (N_36336,N_35154,N_35350);
nor U36337 (N_36337,N_35133,N_35556);
xnor U36338 (N_36338,N_35431,N_35060);
nor U36339 (N_36339,N_35909,N_35603);
nor U36340 (N_36340,N_35564,N_35492);
nand U36341 (N_36341,N_35888,N_35602);
nor U36342 (N_36342,N_35511,N_35229);
and U36343 (N_36343,N_35934,N_35470);
xor U36344 (N_36344,N_35001,N_35512);
xnor U36345 (N_36345,N_35185,N_35540);
nor U36346 (N_36346,N_35299,N_35930);
and U36347 (N_36347,N_35985,N_35363);
nand U36348 (N_36348,N_35258,N_35678);
and U36349 (N_36349,N_35348,N_35831);
or U36350 (N_36350,N_35907,N_35306);
nor U36351 (N_36351,N_35462,N_35279);
or U36352 (N_36352,N_35488,N_35472);
or U36353 (N_36353,N_35549,N_35927);
nor U36354 (N_36354,N_35668,N_35301);
nand U36355 (N_36355,N_35016,N_35704);
nor U36356 (N_36356,N_35160,N_35583);
nor U36357 (N_36357,N_35972,N_35140);
and U36358 (N_36358,N_35276,N_35253);
nor U36359 (N_36359,N_35834,N_35323);
and U36360 (N_36360,N_35868,N_35693);
xor U36361 (N_36361,N_35444,N_35746);
nand U36362 (N_36362,N_35046,N_35981);
nor U36363 (N_36363,N_35753,N_35355);
nor U36364 (N_36364,N_35273,N_35819);
xnor U36365 (N_36365,N_35971,N_35254);
nor U36366 (N_36366,N_35038,N_35109);
xor U36367 (N_36367,N_35114,N_35999);
or U36368 (N_36368,N_35609,N_35088);
nand U36369 (N_36369,N_35706,N_35643);
xor U36370 (N_36370,N_35594,N_35531);
and U36371 (N_36371,N_35761,N_35824);
or U36372 (N_36372,N_35854,N_35809);
and U36373 (N_36373,N_35785,N_35264);
nor U36374 (N_36374,N_35266,N_35468);
and U36375 (N_36375,N_35654,N_35187);
xnor U36376 (N_36376,N_35749,N_35180);
or U36377 (N_36377,N_35482,N_35503);
or U36378 (N_36378,N_35554,N_35755);
or U36379 (N_36379,N_35601,N_35285);
and U36380 (N_36380,N_35897,N_35268);
or U36381 (N_36381,N_35177,N_35222);
nand U36382 (N_36382,N_35585,N_35805);
nand U36383 (N_36383,N_35149,N_35184);
or U36384 (N_36384,N_35480,N_35308);
nor U36385 (N_36385,N_35310,N_35796);
or U36386 (N_36386,N_35900,N_35610);
or U36387 (N_36387,N_35645,N_35107);
and U36388 (N_36388,N_35458,N_35776);
and U36389 (N_36389,N_35625,N_35319);
or U36390 (N_36390,N_35406,N_35436);
nor U36391 (N_36391,N_35054,N_35024);
xor U36392 (N_36392,N_35845,N_35534);
xor U36393 (N_36393,N_35368,N_35271);
and U36394 (N_36394,N_35246,N_35359);
or U36395 (N_36395,N_35216,N_35608);
and U36396 (N_36396,N_35555,N_35957);
and U36397 (N_36397,N_35519,N_35526);
and U36398 (N_36398,N_35634,N_35686);
and U36399 (N_36399,N_35002,N_35080);
and U36400 (N_36400,N_35447,N_35198);
and U36401 (N_36401,N_35227,N_35915);
nor U36402 (N_36402,N_35112,N_35148);
xnor U36403 (N_36403,N_35724,N_35403);
or U36404 (N_36404,N_35367,N_35827);
xnor U36405 (N_36405,N_35014,N_35820);
nor U36406 (N_36406,N_35017,N_35559);
or U36407 (N_36407,N_35459,N_35551);
nand U36408 (N_36408,N_35230,N_35068);
xor U36409 (N_36409,N_35516,N_35951);
xor U36410 (N_36410,N_35723,N_35588);
or U36411 (N_36411,N_35734,N_35255);
and U36412 (N_36412,N_35712,N_35410);
or U36413 (N_36413,N_35176,N_35428);
xnor U36414 (N_36414,N_35692,N_35015);
and U36415 (N_36415,N_35691,N_35092);
nor U36416 (N_36416,N_35463,N_35401);
and U36417 (N_36417,N_35417,N_35886);
xor U36418 (N_36418,N_35297,N_35641);
xor U36419 (N_36419,N_35803,N_35344);
or U36420 (N_36420,N_35781,N_35335);
and U36421 (N_36421,N_35673,N_35432);
and U36422 (N_36422,N_35071,N_35296);
nand U36423 (N_36423,N_35795,N_35638);
xnor U36424 (N_36424,N_35867,N_35984);
or U36425 (N_36425,N_35340,N_35537);
nor U36426 (N_36426,N_35047,N_35146);
xnor U36427 (N_36427,N_35837,N_35121);
or U36428 (N_36428,N_35905,N_35898);
nor U36429 (N_36429,N_35966,N_35156);
nand U36430 (N_36430,N_35102,N_35618);
xor U36431 (N_36431,N_35351,N_35920);
nor U36432 (N_36432,N_35220,N_35979);
and U36433 (N_36433,N_35008,N_35256);
and U36434 (N_36434,N_35147,N_35331);
and U36435 (N_36435,N_35111,N_35665);
nor U36436 (N_36436,N_35607,N_35982);
nor U36437 (N_36437,N_35126,N_35172);
nand U36438 (N_36438,N_35818,N_35694);
nand U36439 (N_36439,N_35765,N_35792);
or U36440 (N_36440,N_35467,N_35977);
nand U36441 (N_36441,N_35452,N_35561);
or U36442 (N_36442,N_35772,N_35937);
nand U36443 (N_36443,N_35605,N_35416);
nor U36444 (N_36444,N_35509,N_35169);
nand U36445 (N_36445,N_35748,N_35733);
or U36446 (N_36446,N_35113,N_35077);
and U36447 (N_36447,N_35621,N_35124);
or U36448 (N_36448,N_35667,N_35816);
nor U36449 (N_36449,N_35051,N_35036);
and U36450 (N_36450,N_35504,N_35846);
or U36451 (N_36451,N_35782,N_35777);
xnor U36452 (N_36452,N_35040,N_35011);
or U36453 (N_36453,N_35787,N_35414);
nor U36454 (N_36454,N_35744,N_35730);
nor U36455 (N_36455,N_35269,N_35260);
or U36456 (N_36456,N_35455,N_35958);
nor U36457 (N_36457,N_35396,N_35636);
or U36458 (N_36458,N_35592,N_35861);
nand U36459 (N_36459,N_35322,N_35487);
nand U36460 (N_36460,N_35964,N_35072);
nor U36461 (N_36461,N_35438,N_35923);
or U36462 (N_36462,N_35632,N_35878);
and U36463 (N_36463,N_35353,N_35946);
nand U36464 (N_36464,N_35758,N_35012);
or U36465 (N_36465,N_35195,N_35799);
nor U36466 (N_36466,N_35100,N_35426);
nand U36467 (N_36467,N_35874,N_35049);
nand U36468 (N_36468,N_35547,N_35275);
or U36469 (N_36469,N_35527,N_35910);
and U36470 (N_36470,N_35122,N_35304);
or U36471 (N_36471,N_35974,N_35429);
and U36472 (N_36472,N_35976,N_35784);
and U36473 (N_36473,N_35108,N_35518);
or U36474 (N_36474,N_35674,N_35893);
or U36475 (N_36475,N_35405,N_35887);
nor U36476 (N_36476,N_35034,N_35718);
nor U36477 (N_36477,N_35994,N_35695);
and U36478 (N_36478,N_35473,N_35218);
nand U36479 (N_36479,N_35885,N_35461);
and U36480 (N_36480,N_35917,N_35489);
and U36481 (N_36481,N_35595,N_35980);
nor U36482 (N_36482,N_35743,N_35978);
or U36483 (N_36483,N_35244,N_35491);
nand U36484 (N_36484,N_35007,N_35106);
xor U36485 (N_36485,N_35261,N_35065);
nand U36486 (N_36486,N_35388,N_35763);
nand U36487 (N_36487,N_35009,N_35542);
xnor U36488 (N_36488,N_35129,N_35381);
nor U36489 (N_36489,N_35873,N_35324);
xnor U36490 (N_36490,N_35802,N_35311);
or U36491 (N_36491,N_35580,N_35931);
xnor U36492 (N_36492,N_35374,N_35197);
nand U36493 (N_36493,N_35120,N_35525);
nor U36494 (N_36494,N_35655,N_35360);
and U36495 (N_36495,N_35199,N_35157);
xor U36496 (N_36496,N_35593,N_35233);
and U36497 (N_36497,N_35727,N_35474);
nand U36498 (N_36498,N_35370,N_35469);
and U36499 (N_36499,N_35341,N_35171);
nor U36500 (N_36500,N_35086,N_35910);
or U36501 (N_36501,N_35701,N_35273);
nand U36502 (N_36502,N_35217,N_35698);
nor U36503 (N_36503,N_35352,N_35531);
and U36504 (N_36504,N_35176,N_35197);
or U36505 (N_36505,N_35551,N_35141);
xnor U36506 (N_36506,N_35745,N_35969);
or U36507 (N_36507,N_35138,N_35178);
nand U36508 (N_36508,N_35995,N_35620);
or U36509 (N_36509,N_35664,N_35416);
nand U36510 (N_36510,N_35291,N_35426);
and U36511 (N_36511,N_35503,N_35062);
and U36512 (N_36512,N_35943,N_35076);
nor U36513 (N_36513,N_35290,N_35063);
or U36514 (N_36514,N_35010,N_35915);
and U36515 (N_36515,N_35756,N_35587);
and U36516 (N_36516,N_35595,N_35897);
and U36517 (N_36517,N_35508,N_35467);
nand U36518 (N_36518,N_35717,N_35951);
nor U36519 (N_36519,N_35873,N_35291);
nand U36520 (N_36520,N_35846,N_35480);
xor U36521 (N_36521,N_35601,N_35497);
nor U36522 (N_36522,N_35857,N_35760);
or U36523 (N_36523,N_35956,N_35343);
or U36524 (N_36524,N_35709,N_35115);
or U36525 (N_36525,N_35623,N_35587);
nand U36526 (N_36526,N_35162,N_35134);
xnor U36527 (N_36527,N_35282,N_35777);
nor U36528 (N_36528,N_35864,N_35696);
nand U36529 (N_36529,N_35709,N_35737);
and U36530 (N_36530,N_35179,N_35249);
or U36531 (N_36531,N_35185,N_35755);
nand U36532 (N_36532,N_35897,N_35654);
xnor U36533 (N_36533,N_35796,N_35726);
nand U36534 (N_36534,N_35403,N_35051);
nor U36535 (N_36535,N_35536,N_35776);
and U36536 (N_36536,N_35559,N_35997);
and U36537 (N_36537,N_35520,N_35072);
nand U36538 (N_36538,N_35321,N_35183);
or U36539 (N_36539,N_35252,N_35671);
or U36540 (N_36540,N_35058,N_35441);
and U36541 (N_36541,N_35534,N_35817);
nor U36542 (N_36542,N_35148,N_35889);
nand U36543 (N_36543,N_35745,N_35644);
xnor U36544 (N_36544,N_35693,N_35452);
nor U36545 (N_36545,N_35829,N_35784);
or U36546 (N_36546,N_35033,N_35546);
or U36547 (N_36547,N_35924,N_35380);
or U36548 (N_36548,N_35892,N_35210);
nor U36549 (N_36549,N_35278,N_35364);
and U36550 (N_36550,N_35342,N_35114);
and U36551 (N_36551,N_35427,N_35675);
and U36552 (N_36552,N_35373,N_35782);
or U36553 (N_36553,N_35610,N_35303);
and U36554 (N_36554,N_35503,N_35173);
nand U36555 (N_36555,N_35237,N_35265);
nor U36556 (N_36556,N_35725,N_35611);
xor U36557 (N_36557,N_35678,N_35713);
nand U36558 (N_36558,N_35409,N_35466);
and U36559 (N_36559,N_35833,N_35951);
and U36560 (N_36560,N_35322,N_35085);
and U36561 (N_36561,N_35907,N_35096);
and U36562 (N_36562,N_35108,N_35898);
xnor U36563 (N_36563,N_35015,N_35735);
nor U36564 (N_36564,N_35141,N_35662);
and U36565 (N_36565,N_35703,N_35286);
and U36566 (N_36566,N_35642,N_35187);
xnor U36567 (N_36567,N_35498,N_35851);
and U36568 (N_36568,N_35452,N_35956);
or U36569 (N_36569,N_35072,N_35664);
nor U36570 (N_36570,N_35809,N_35419);
nor U36571 (N_36571,N_35966,N_35560);
and U36572 (N_36572,N_35669,N_35965);
nand U36573 (N_36573,N_35780,N_35221);
nand U36574 (N_36574,N_35187,N_35338);
and U36575 (N_36575,N_35273,N_35372);
nand U36576 (N_36576,N_35265,N_35543);
or U36577 (N_36577,N_35441,N_35167);
nor U36578 (N_36578,N_35077,N_35997);
or U36579 (N_36579,N_35589,N_35959);
or U36580 (N_36580,N_35100,N_35593);
nand U36581 (N_36581,N_35538,N_35445);
nor U36582 (N_36582,N_35125,N_35277);
or U36583 (N_36583,N_35487,N_35219);
and U36584 (N_36584,N_35262,N_35131);
xnor U36585 (N_36585,N_35728,N_35892);
xnor U36586 (N_36586,N_35469,N_35660);
and U36587 (N_36587,N_35612,N_35430);
and U36588 (N_36588,N_35450,N_35366);
nand U36589 (N_36589,N_35781,N_35945);
or U36590 (N_36590,N_35007,N_35072);
or U36591 (N_36591,N_35259,N_35654);
and U36592 (N_36592,N_35728,N_35367);
and U36593 (N_36593,N_35247,N_35630);
nor U36594 (N_36594,N_35441,N_35854);
or U36595 (N_36595,N_35037,N_35459);
nor U36596 (N_36596,N_35951,N_35613);
and U36597 (N_36597,N_35960,N_35028);
nor U36598 (N_36598,N_35338,N_35214);
nor U36599 (N_36599,N_35729,N_35309);
or U36600 (N_36600,N_35275,N_35249);
nand U36601 (N_36601,N_35400,N_35638);
or U36602 (N_36602,N_35947,N_35754);
nor U36603 (N_36603,N_35495,N_35362);
nand U36604 (N_36604,N_35185,N_35437);
nand U36605 (N_36605,N_35114,N_35883);
and U36606 (N_36606,N_35034,N_35430);
or U36607 (N_36607,N_35512,N_35838);
nand U36608 (N_36608,N_35503,N_35919);
xor U36609 (N_36609,N_35145,N_35624);
and U36610 (N_36610,N_35705,N_35715);
xnor U36611 (N_36611,N_35718,N_35100);
or U36612 (N_36612,N_35834,N_35824);
or U36613 (N_36613,N_35738,N_35065);
or U36614 (N_36614,N_35817,N_35714);
nor U36615 (N_36615,N_35948,N_35604);
nand U36616 (N_36616,N_35194,N_35440);
xor U36617 (N_36617,N_35982,N_35585);
xor U36618 (N_36618,N_35491,N_35778);
xnor U36619 (N_36619,N_35410,N_35044);
xnor U36620 (N_36620,N_35847,N_35782);
nor U36621 (N_36621,N_35434,N_35328);
nor U36622 (N_36622,N_35758,N_35260);
nor U36623 (N_36623,N_35345,N_35491);
nand U36624 (N_36624,N_35229,N_35086);
nor U36625 (N_36625,N_35306,N_35175);
nor U36626 (N_36626,N_35768,N_35945);
nor U36627 (N_36627,N_35637,N_35800);
nor U36628 (N_36628,N_35212,N_35947);
nor U36629 (N_36629,N_35852,N_35247);
nand U36630 (N_36630,N_35278,N_35199);
or U36631 (N_36631,N_35254,N_35801);
nand U36632 (N_36632,N_35776,N_35703);
nand U36633 (N_36633,N_35088,N_35128);
or U36634 (N_36634,N_35405,N_35085);
nand U36635 (N_36635,N_35673,N_35040);
and U36636 (N_36636,N_35403,N_35104);
xnor U36637 (N_36637,N_35992,N_35990);
nor U36638 (N_36638,N_35404,N_35480);
xnor U36639 (N_36639,N_35319,N_35156);
and U36640 (N_36640,N_35915,N_35016);
xnor U36641 (N_36641,N_35762,N_35647);
or U36642 (N_36642,N_35903,N_35979);
or U36643 (N_36643,N_35684,N_35795);
nand U36644 (N_36644,N_35235,N_35987);
xor U36645 (N_36645,N_35488,N_35280);
and U36646 (N_36646,N_35230,N_35095);
or U36647 (N_36647,N_35762,N_35939);
or U36648 (N_36648,N_35728,N_35786);
nor U36649 (N_36649,N_35264,N_35659);
or U36650 (N_36650,N_35727,N_35048);
or U36651 (N_36651,N_35319,N_35631);
nand U36652 (N_36652,N_35825,N_35409);
or U36653 (N_36653,N_35388,N_35968);
nor U36654 (N_36654,N_35212,N_35140);
nand U36655 (N_36655,N_35268,N_35006);
nand U36656 (N_36656,N_35445,N_35131);
nand U36657 (N_36657,N_35191,N_35719);
nand U36658 (N_36658,N_35081,N_35065);
xnor U36659 (N_36659,N_35554,N_35480);
or U36660 (N_36660,N_35154,N_35584);
nand U36661 (N_36661,N_35543,N_35042);
nand U36662 (N_36662,N_35904,N_35100);
and U36663 (N_36663,N_35071,N_35776);
and U36664 (N_36664,N_35807,N_35235);
and U36665 (N_36665,N_35296,N_35190);
nor U36666 (N_36666,N_35903,N_35605);
xor U36667 (N_36667,N_35119,N_35407);
nor U36668 (N_36668,N_35408,N_35433);
xnor U36669 (N_36669,N_35491,N_35713);
nand U36670 (N_36670,N_35861,N_35372);
xnor U36671 (N_36671,N_35808,N_35233);
or U36672 (N_36672,N_35997,N_35530);
nor U36673 (N_36673,N_35274,N_35912);
xor U36674 (N_36674,N_35125,N_35458);
or U36675 (N_36675,N_35718,N_35846);
and U36676 (N_36676,N_35665,N_35590);
xor U36677 (N_36677,N_35752,N_35857);
nand U36678 (N_36678,N_35803,N_35430);
and U36679 (N_36679,N_35742,N_35243);
and U36680 (N_36680,N_35435,N_35057);
and U36681 (N_36681,N_35634,N_35418);
xor U36682 (N_36682,N_35387,N_35759);
nor U36683 (N_36683,N_35787,N_35638);
and U36684 (N_36684,N_35717,N_35339);
nand U36685 (N_36685,N_35650,N_35587);
and U36686 (N_36686,N_35101,N_35850);
nand U36687 (N_36687,N_35399,N_35756);
and U36688 (N_36688,N_35941,N_35535);
xnor U36689 (N_36689,N_35702,N_35181);
and U36690 (N_36690,N_35647,N_35804);
xnor U36691 (N_36691,N_35146,N_35160);
and U36692 (N_36692,N_35228,N_35968);
xnor U36693 (N_36693,N_35604,N_35964);
nor U36694 (N_36694,N_35332,N_35676);
or U36695 (N_36695,N_35586,N_35560);
and U36696 (N_36696,N_35188,N_35044);
or U36697 (N_36697,N_35872,N_35135);
and U36698 (N_36698,N_35579,N_35713);
nand U36699 (N_36699,N_35828,N_35552);
xnor U36700 (N_36700,N_35952,N_35706);
or U36701 (N_36701,N_35722,N_35111);
and U36702 (N_36702,N_35041,N_35410);
nand U36703 (N_36703,N_35680,N_35831);
nand U36704 (N_36704,N_35745,N_35573);
or U36705 (N_36705,N_35665,N_35504);
and U36706 (N_36706,N_35417,N_35814);
nor U36707 (N_36707,N_35070,N_35794);
nor U36708 (N_36708,N_35390,N_35537);
or U36709 (N_36709,N_35477,N_35273);
xnor U36710 (N_36710,N_35471,N_35231);
xor U36711 (N_36711,N_35336,N_35015);
and U36712 (N_36712,N_35597,N_35905);
or U36713 (N_36713,N_35086,N_35155);
and U36714 (N_36714,N_35676,N_35742);
nand U36715 (N_36715,N_35689,N_35348);
nor U36716 (N_36716,N_35641,N_35938);
or U36717 (N_36717,N_35066,N_35930);
or U36718 (N_36718,N_35996,N_35748);
nor U36719 (N_36719,N_35240,N_35649);
xnor U36720 (N_36720,N_35669,N_35355);
xnor U36721 (N_36721,N_35389,N_35580);
nor U36722 (N_36722,N_35649,N_35333);
or U36723 (N_36723,N_35235,N_35753);
and U36724 (N_36724,N_35808,N_35694);
xor U36725 (N_36725,N_35457,N_35111);
and U36726 (N_36726,N_35611,N_35428);
or U36727 (N_36727,N_35172,N_35280);
nor U36728 (N_36728,N_35301,N_35895);
xor U36729 (N_36729,N_35568,N_35900);
nand U36730 (N_36730,N_35530,N_35156);
and U36731 (N_36731,N_35271,N_35863);
xnor U36732 (N_36732,N_35000,N_35854);
xnor U36733 (N_36733,N_35872,N_35266);
xnor U36734 (N_36734,N_35116,N_35000);
nor U36735 (N_36735,N_35556,N_35124);
and U36736 (N_36736,N_35019,N_35720);
or U36737 (N_36737,N_35525,N_35502);
and U36738 (N_36738,N_35372,N_35561);
and U36739 (N_36739,N_35997,N_35796);
and U36740 (N_36740,N_35260,N_35370);
or U36741 (N_36741,N_35475,N_35184);
xnor U36742 (N_36742,N_35481,N_35656);
nand U36743 (N_36743,N_35285,N_35528);
or U36744 (N_36744,N_35807,N_35507);
xor U36745 (N_36745,N_35044,N_35085);
nor U36746 (N_36746,N_35048,N_35185);
or U36747 (N_36747,N_35042,N_35838);
nor U36748 (N_36748,N_35771,N_35897);
nand U36749 (N_36749,N_35432,N_35656);
and U36750 (N_36750,N_35343,N_35989);
nand U36751 (N_36751,N_35741,N_35769);
or U36752 (N_36752,N_35720,N_35324);
and U36753 (N_36753,N_35908,N_35449);
nand U36754 (N_36754,N_35061,N_35114);
nor U36755 (N_36755,N_35287,N_35698);
nor U36756 (N_36756,N_35439,N_35382);
nor U36757 (N_36757,N_35388,N_35488);
nor U36758 (N_36758,N_35529,N_35476);
xnor U36759 (N_36759,N_35821,N_35585);
or U36760 (N_36760,N_35640,N_35555);
xnor U36761 (N_36761,N_35745,N_35586);
and U36762 (N_36762,N_35981,N_35914);
nor U36763 (N_36763,N_35138,N_35036);
nor U36764 (N_36764,N_35435,N_35275);
xor U36765 (N_36765,N_35795,N_35522);
nor U36766 (N_36766,N_35883,N_35304);
or U36767 (N_36767,N_35866,N_35102);
nand U36768 (N_36768,N_35297,N_35506);
nor U36769 (N_36769,N_35231,N_35671);
nor U36770 (N_36770,N_35711,N_35480);
and U36771 (N_36771,N_35745,N_35172);
or U36772 (N_36772,N_35610,N_35865);
and U36773 (N_36773,N_35112,N_35660);
and U36774 (N_36774,N_35458,N_35419);
xnor U36775 (N_36775,N_35852,N_35215);
xnor U36776 (N_36776,N_35610,N_35409);
nand U36777 (N_36777,N_35051,N_35598);
and U36778 (N_36778,N_35799,N_35986);
and U36779 (N_36779,N_35988,N_35717);
nand U36780 (N_36780,N_35926,N_35455);
nand U36781 (N_36781,N_35540,N_35189);
nor U36782 (N_36782,N_35677,N_35385);
or U36783 (N_36783,N_35564,N_35092);
and U36784 (N_36784,N_35383,N_35398);
xor U36785 (N_36785,N_35742,N_35962);
nand U36786 (N_36786,N_35299,N_35072);
or U36787 (N_36787,N_35235,N_35171);
xor U36788 (N_36788,N_35847,N_35987);
nor U36789 (N_36789,N_35316,N_35781);
nor U36790 (N_36790,N_35606,N_35079);
nand U36791 (N_36791,N_35448,N_35215);
or U36792 (N_36792,N_35250,N_35057);
nand U36793 (N_36793,N_35956,N_35382);
nand U36794 (N_36794,N_35860,N_35350);
xor U36795 (N_36795,N_35297,N_35201);
or U36796 (N_36796,N_35574,N_35722);
nor U36797 (N_36797,N_35419,N_35057);
or U36798 (N_36798,N_35881,N_35571);
and U36799 (N_36799,N_35417,N_35694);
nand U36800 (N_36800,N_35367,N_35338);
xnor U36801 (N_36801,N_35588,N_35894);
nand U36802 (N_36802,N_35591,N_35183);
or U36803 (N_36803,N_35868,N_35804);
and U36804 (N_36804,N_35160,N_35532);
nor U36805 (N_36805,N_35367,N_35736);
nand U36806 (N_36806,N_35858,N_35155);
and U36807 (N_36807,N_35665,N_35443);
xor U36808 (N_36808,N_35989,N_35357);
xnor U36809 (N_36809,N_35181,N_35024);
nand U36810 (N_36810,N_35605,N_35485);
xnor U36811 (N_36811,N_35166,N_35390);
nand U36812 (N_36812,N_35156,N_35682);
nor U36813 (N_36813,N_35817,N_35606);
nand U36814 (N_36814,N_35569,N_35261);
or U36815 (N_36815,N_35678,N_35965);
or U36816 (N_36816,N_35009,N_35778);
and U36817 (N_36817,N_35587,N_35199);
and U36818 (N_36818,N_35158,N_35836);
nor U36819 (N_36819,N_35416,N_35499);
or U36820 (N_36820,N_35590,N_35271);
or U36821 (N_36821,N_35620,N_35930);
nand U36822 (N_36822,N_35979,N_35032);
xor U36823 (N_36823,N_35471,N_35438);
nor U36824 (N_36824,N_35294,N_35771);
nor U36825 (N_36825,N_35753,N_35063);
or U36826 (N_36826,N_35768,N_35414);
nor U36827 (N_36827,N_35608,N_35178);
and U36828 (N_36828,N_35203,N_35382);
nor U36829 (N_36829,N_35334,N_35937);
xor U36830 (N_36830,N_35570,N_35449);
and U36831 (N_36831,N_35962,N_35386);
nand U36832 (N_36832,N_35807,N_35656);
nand U36833 (N_36833,N_35357,N_35552);
and U36834 (N_36834,N_35299,N_35679);
or U36835 (N_36835,N_35468,N_35708);
xor U36836 (N_36836,N_35062,N_35668);
nand U36837 (N_36837,N_35068,N_35588);
xor U36838 (N_36838,N_35496,N_35168);
xnor U36839 (N_36839,N_35490,N_35794);
and U36840 (N_36840,N_35457,N_35199);
nor U36841 (N_36841,N_35659,N_35545);
nor U36842 (N_36842,N_35384,N_35822);
xnor U36843 (N_36843,N_35800,N_35116);
and U36844 (N_36844,N_35732,N_35701);
nor U36845 (N_36845,N_35584,N_35918);
or U36846 (N_36846,N_35406,N_35786);
nor U36847 (N_36847,N_35218,N_35466);
and U36848 (N_36848,N_35031,N_35687);
and U36849 (N_36849,N_35411,N_35858);
and U36850 (N_36850,N_35255,N_35991);
or U36851 (N_36851,N_35657,N_35245);
nor U36852 (N_36852,N_35166,N_35519);
or U36853 (N_36853,N_35073,N_35306);
nor U36854 (N_36854,N_35498,N_35166);
or U36855 (N_36855,N_35163,N_35793);
and U36856 (N_36856,N_35123,N_35927);
nor U36857 (N_36857,N_35933,N_35693);
xnor U36858 (N_36858,N_35221,N_35585);
or U36859 (N_36859,N_35834,N_35373);
or U36860 (N_36860,N_35488,N_35094);
nor U36861 (N_36861,N_35656,N_35668);
xor U36862 (N_36862,N_35884,N_35104);
xor U36863 (N_36863,N_35261,N_35268);
xnor U36864 (N_36864,N_35930,N_35140);
nor U36865 (N_36865,N_35757,N_35748);
nand U36866 (N_36866,N_35623,N_35328);
and U36867 (N_36867,N_35978,N_35878);
nor U36868 (N_36868,N_35017,N_35943);
or U36869 (N_36869,N_35261,N_35455);
nor U36870 (N_36870,N_35096,N_35520);
and U36871 (N_36871,N_35060,N_35727);
nand U36872 (N_36872,N_35107,N_35901);
nand U36873 (N_36873,N_35527,N_35729);
or U36874 (N_36874,N_35172,N_35023);
xor U36875 (N_36875,N_35007,N_35397);
and U36876 (N_36876,N_35863,N_35027);
and U36877 (N_36877,N_35101,N_35972);
nor U36878 (N_36878,N_35076,N_35276);
or U36879 (N_36879,N_35339,N_35221);
and U36880 (N_36880,N_35597,N_35739);
nand U36881 (N_36881,N_35360,N_35700);
nor U36882 (N_36882,N_35432,N_35268);
nand U36883 (N_36883,N_35526,N_35821);
nand U36884 (N_36884,N_35553,N_35208);
nor U36885 (N_36885,N_35689,N_35454);
xnor U36886 (N_36886,N_35513,N_35658);
xor U36887 (N_36887,N_35140,N_35237);
nand U36888 (N_36888,N_35794,N_35304);
nor U36889 (N_36889,N_35958,N_35604);
nand U36890 (N_36890,N_35889,N_35630);
and U36891 (N_36891,N_35853,N_35549);
and U36892 (N_36892,N_35646,N_35680);
or U36893 (N_36893,N_35756,N_35044);
nor U36894 (N_36894,N_35083,N_35193);
nor U36895 (N_36895,N_35966,N_35200);
nand U36896 (N_36896,N_35750,N_35941);
xor U36897 (N_36897,N_35754,N_35324);
nand U36898 (N_36898,N_35161,N_35491);
or U36899 (N_36899,N_35861,N_35587);
or U36900 (N_36900,N_35379,N_35488);
xnor U36901 (N_36901,N_35416,N_35762);
or U36902 (N_36902,N_35852,N_35878);
nor U36903 (N_36903,N_35754,N_35566);
or U36904 (N_36904,N_35280,N_35370);
or U36905 (N_36905,N_35648,N_35114);
and U36906 (N_36906,N_35965,N_35485);
nor U36907 (N_36907,N_35006,N_35970);
and U36908 (N_36908,N_35095,N_35495);
and U36909 (N_36909,N_35466,N_35730);
and U36910 (N_36910,N_35257,N_35621);
and U36911 (N_36911,N_35020,N_35196);
xor U36912 (N_36912,N_35840,N_35781);
or U36913 (N_36913,N_35442,N_35759);
nand U36914 (N_36914,N_35055,N_35239);
and U36915 (N_36915,N_35828,N_35754);
nor U36916 (N_36916,N_35922,N_35717);
and U36917 (N_36917,N_35917,N_35760);
and U36918 (N_36918,N_35443,N_35357);
nand U36919 (N_36919,N_35180,N_35364);
nand U36920 (N_36920,N_35531,N_35553);
and U36921 (N_36921,N_35623,N_35111);
xor U36922 (N_36922,N_35883,N_35687);
nor U36923 (N_36923,N_35871,N_35493);
xor U36924 (N_36924,N_35461,N_35669);
or U36925 (N_36925,N_35101,N_35318);
nor U36926 (N_36926,N_35868,N_35469);
nor U36927 (N_36927,N_35569,N_35628);
nand U36928 (N_36928,N_35544,N_35203);
xnor U36929 (N_36929,N_35493,N_35295);
and U36930 (N_36930,N_35101,N_35168);
xnor U36931 (N_36931,N_35675,N_35733);
nor U36932 (N_36932,N_35839,N_35956);
nand U36933 (N_36933,N_35471,N_35026);
and U36934 (N_36934,N_35976,N_35756);
xor U36935 (N_36935,N_35353,N_35165);
nand U36936 (N_36936,N_35926,N_35487);
and U36937 (N_36937,N_35862,N_35075);
nor U36938 (N_36938,N_35213,N_35185);
xnor U36939 (N_36939,N_35640,N_35414);
and U36940 (N_36940,N_35868,N_35658);
nand U36941 (N_36941,N_35261,N_35880);
or U36942 (N_36942,N_35415,N_35495);
or U36943 (N_36943,N_35009,N_35888);
and U36944 (N_36944,N_35017,N_35204);
xor U36945 (N_36945,N_35561,N_35411);
and U36946 (N_36946,N_35692,N_35972);
nor U36947 (N_36947,N_35353,N_35838);
xnor U36948 (N_36948,N_35938,N_35813);
or U36949 (N_36949,N_35335,N_35271);
and U36950 (N_36950,N_35342,N_35426);
or U36951 (N_36951,N_35828,N_35006);
and U36952 (N_36952,N_35783,N_35408);
nor U36953 (N_36953,N_35102,N_35982);
and U36954 (N_36954,N_35560,N_35899);
nand U36955 (N_36955,N_35706,N_35442);
xor U36956 (N_36956,N_35004,N_35834);
nand U36957 (N_36957,N_35036,N_35659);
or U36958 (N_36958,N_35020,N_35891);
and U36959 (N_36959,N_35961,N_35810);
xor U36960 (N_36960,N_35416,N_35742);
and U36961 (N_36961,N_35580,N_35507);
xnor U36962 (N_36962,N_35860,N_35579);
and U36963 (N_36963,N_35010,N_35151);
xnor U36964 (N_36964,N_35167,N_35876);
and U36965 (N_36965,N_35473,N_35977);
nand U36966 (N_36966,N_35842,N_35975);
or U36967 (N_36967,N_35493,N_35161);
nor U36968 (N_36968,N_35249,N_35485);
and U36969 (N_36969,N_35599,N_35112);
and U36970 (N_36970,N_35724,N_35043);
and U36971 (N_36971,N_35169,N_35342);
and U36972 (N_36972,N_35189,N_35623);
nor U36973 (N_36973,N_35322,N_35730);
xor U36974 (N_36974,N_35688,N_35796);
nor U36975 (N_36975,N_35184,N_35510);
and U36976 (N_36976,N_35312,N_35145);
or U36977 (N_36977,N_35867,N_35142);
xnor U36978 (N_36978,N_35250,N_35983);
and U36979 (N_36979,N_35297,N_35011);
nand U36980 (N_36980,N_35767,N_35056);
nand U36981 (N_36981,N_35615,N_35459);
nor U36982 (N_36982,N_35099,N_35892);
nand U36983 (N_36983,N_35424,N_35702);
nand U36984 (N_36984,N_35139,N_35969);
nor U36985 (N_36985,N_35677,N_35416);
xnor U36986 (N_36986,N_35601,N_35509);
xor U36987 (N_36987,N_35829,N_35795);
nor U36988 (N_36988,N_35731,N_35790);
and U36989 (N_36989,N_35303,N_35949);
and U36990 (N_36990,N_35295,N_35086);
xnor U36991 (N_36991,N_35571,N_35165);
and U36992 (N_36992,N_35176,N_35800);
nand U36993 (N_36993,N_35995,N_35524);
nor U36994 (N_36994,N_35940,N_35748);
or U36995 (N_36995,N_35265,N_35736);
nor U36996 (N_36996,N_35457,N_35312);
and U36997 (N_36997,N_35610,N_35911);
nand U36998 (N_36998,N_35917,N_35607);
nor U36999 (N_36999,N_35700,N_35230);
nor U37000 (N_37000,N_36090,N_36063);
nor U37001 (N_37001,N_36212,N_36539);
and U37002 (N_37002,N_36080,N_36532);
xnor U37003 (N_37003,N_36109,N_36643);
or U37004 (N_37004,N_36546,N_36297);
nor U37005 (N_37005,N_36217,N_36913);
nand U37006 (N_37006,N_36085,N_36267);
or U37007 (N_37007,N_36824,N_36461);
nand U37008 (N_37008,N_36438,N_36499);
or U37009 (N_37009,N_36186,N_36823);
nand U37010 (N_37010,N_36455,N_36638);
nand U37011 (N_37011,N_36042,N_36929);
nor U37012 (N_37012,N_36954,N_36431);
nor U37013 (N_37013,N_36460,N_36489);
nand U37014 (N_37014,N_36124,N_36915);
nand U37015 (N_37015,N_36066,N_36030);
nor U37016 (N_37016,N_36322,N_36477);
or U37017 (N_37017,N_36992,N_36382);
nor U37018 (N_37018,N_36896,N_36414);
nand U37019 (N_37019,N_36263,N_36513);
nand U37020 (N_37020,N_36337,N_36588);
nand U37021 (N_37021,N_36181,N_36418);
nand U37022 (N_37022,N_36260,N_36250);
or U37023 (N_37023,N_36770,N_36701);
xnor U37024 (N_37024,N_36449,N_36122);
or U37025 (N_37025,N_36453,N_36016);
or U37026 (N_37026,N_36517,N_36820);
nor U37027 (N_37027,N_36490,N_36482);
xnor U37028 (N_37028,N_36028,N_36926);
nor U37029 (N_37029,N_36619,N_36190);
nand U37030 (N_37030,N_36525,N_36007);
and U37031 (N_37031,N_36290,N_36386);
and U37032 (N_37032,N_36423,N_36467);
xnor U37033 (N_37033,N_36991,N_36253);
or U37034 (N_37034,N_36395,N_36686);
nand U37035 (N_37035,N_36091,N_36218);
xnor U37036 (N_37036,N_36202,N_36331);
or U37037 (N_37037,N_36728,N_36964);
and U37038 (N_37038,N_36027,N_36226);
and U37039 (N_37039,N_36623,N_36147);
xnor U37040 (N_37040,N_36236,N_36861);
and U37041 (N_37041,N_36156,N_36501);
nand U37042 (N_37042,N_36578,N_36123);
nand U37043 (N_37043,N_36401,N_36357);
and U37044 (N_37044,N_36478,N_36606);
nand U37045 (N_37045,N_36246,N_36448);
nand U37046 (N_37046,N_36220,N_36555);
nand U37047 (N_37047,N_36474,N_36161);
xnor U37048 (N_37048,N_36613,N_36818);
and U37049 (N_37049,N_36249,N_36120);
xnor U37050 (N_37050,N_36082,N_36367);
or U37051 (N_37051,N_36551,N_36494);
nor U37052 (N_37052,N_36328,N_36305);
or U37053 (N_37053,N_36536,N_36222);
xor U37054 (N_37054,N_36316,N_36971);
xor U37055 (N_37055,N_36115,N_36271);
nor U37056 (N_37056,N_36177,N_36458);
xor U37057 (N_37057,N_36409,N_36862);
nor U37058 (N_37058,N_36544,N_36822);
nand U37059 (N_37059,N_36607,N_36303);
xnor U37060 (N_37060,N_36003,N_36352);
nor U37061 (N_37061,N_36302,N_36348);
nor U37062 (N_37062,N_36265,N_36918);
nand U37063 (N_37063,N_36724,N_36998);
xor U37064 (N_37064,N_36668,N_36570);
and U37065 (N_37065,N_36432,N_36070);
or U37066 (N_37066,N_36615,N_36947);
nor U37067 (N_37067,N_36841,N_36855);
xor U37068 (N_37068,N_36796,N_36493);
and U37069 (N_37069,N_36074,N_36987);
and U37070 (N_37070,N_36366,N_36900);
or U37071 (N_37071,N_36663,N_36596);
or U37072 (N_37072,N_36436,N_36447);
nand U37073 (N_37073,N_36858,N_36782);
and U37074 (N_37074,N_36426,N_36173);
xor U37075 (N_37075,N_36330,N_36692);
or U37076 (N_37076,N_36683,N_36377);
or U37077 (N_37077,N_36069,N_36373);
nand U37078 (N_37078,N_36046,N_36283);
and U37079 (N_37079,N_36771,N_36153);
xnor U37080 (N_37080,N_36295,N_36909);
and U37081 (N_37081,N_36644,N_36952);
xnor U37082 (N_37082,N_36150,N_36761);
and U37083 (N_37083,N_36864,N_36139);
xnor U37084 (N_37084,N_36107,N_36905);
or U37085 (N_37085,N_36203,N_36565);
nand U37086 (N_37086,N_36895,N_36384);
xnor U37087 (N_37087,N_36088,N_36700);
xor U37088 (N_37088,N_36463,N_36924);
xnor U37089 (N_37089,N_36158,N_36691);
or U37090 (N_37090,N_36289,N_36550);
xnor U37091 (N_37091,N_36865,N_36104);
nand U37092 (N_37092,N_36257,N_36885);
nor U37093 (N_37093,N_36970,N_36747);
and U37094 (N_37094,N_36183,N_36325);
nand U37095 (N_37095,N_36799,N_36151);
nand U37096 (N_37096,N_36312,N_36777);
nor U37097 (N_37097,N_36041,N_36456);
xnor U37098 (N_37098,N_36067,N_36335);
and U37099 (N_37099,N_36197,N_36149);
and U37100 (N_37100,N_36060,N_36038);
xnor U37101 (N_37101,N_36043,N_36506);
nor U37102 (N_37102,N_36802,N_36018);
or U37103 (N_37103,N_36631,N_36745);
xnor U37104 (N_37104,N_36825,N_36937);
or U37105 (N_37105,N_36755,N_36008);
xnor U37106 (N_37106,N_36317,N_36087);
nor U37107 (N_37107,N_36098,N_36645);
and U37108 (N_37108,N_36052,N_36979);
nand U37109 (N_37109,N_36670,N_36966);
nor U37110 (N_37110,N_36882,N_36783);
xor U37111 (N_37111,N_36627,N_36089);
xnor U37112 (N_37112,N_36336,N_36727);
nand U37113 (N_37113,N_36793,N_36968);
and U37114 (N_37114,N_36451,N_36342);
and U37115 (N_37115,N_36651,N_36450);
xor U37116 (N_37116,N_36393,N_36636);
and U37117 (N_37117,N_36339,N_36024);
xnor U37118 (N_37118,N_36713,N_36108);
nand U37119 (N_37119,N_36372,N_36790);
and U37120 (N_37120,N_36049,N_36326);
nor U37121 (N_37121,N_36208,N_36320);
nor U37122 (N_37122,N_36816,N_36817);
and U37123 (N_37123,N_36381,N_36928);
nor U37124 (N_37124,N_36398,N_36084);
xor U37125 (N_37125,N_36571,N_36764);
nor U37126 (N_37126,N_36752,N_36813);
or U37127 (N_37127,N_36657,N_36040);
and U37128 (N_37128,N_36511,N_36914);
and U37129 (N_37129,N_36065,N_36428);
and U37130 (N_37130,N_36152,N_36094);
or U37131 (N_37131,N_36845,N_36219);
nand U37132 (N_37132,N_36308,N_36883);
or U37133 (N_37133,N_36726,N_36575);
nor U37134 (N_37134,N_36130,N_36803);
and U37135 (N_37135,N_36666,N_36963);
and U37136 (N_37136,N_36829,N_36284);
and U37137 (N_37137,N_36200,N_36170);
or U37138 (N_37138,N_36189,N_36270);
or U37139 (N_37139,N_36961,N_36637);
and U37140 (N_37140,N_36288,N_36689);
or U37141 (N_37141,N_36681,N_36597);
nand U37142 (N_37142,N_36852,N_36949);
or U37143 (N_37143,N_36719,N_36664);
and U37144 (N_37144,N_36344,N_36660);
nor U37145 (N_37145,N_36695,N_36945);
xnor U37146 (N_37146,N_36345,N_36138);
or U37147 (N_37147,N_36406,N_36894);
xnor U37148 (N_37148,N_36475,N_36736);
or U37149 (N_37149,N_36598,N_36658);
xor U37150 (N_37150,N_36955,N_36983);
and U37151 (N_37151,N_36213,N_36936);
nand U37152 (N_37152,N_36001,N_36471);
and U37153 (N_37153,N_36440,N_36380);
nand U37154 (N_37154,N_36699,N_36577);
nor U37155 (N_37155,N_36560,N_36402);
xnor U37156 (N_37156,N_36648,N_36647);
xnor U37157 (N_37157,N_36687,N_36445);
or U37158 (N_37158,N_36140,N_36806);
or U37159 (N_37159,N_36311,N_36053);
or U37160 (N_37160,N_36113,N_36653);
nor U37161 (N_37161,N_36103,N_36733);
nand U37162 (N_37162,N_36282,N_36388);
nand U37163 (N_37163,N_36775,N_36723);
nor U37164 (N_37164,N_36935,N_36280);
and U37165 (N_37165,N_36300,N_36285);
or U37166 (N_37166,N_36237,N_36839);
nor U37167 (N_37167,N_36235,N_36781);
or U37168 (N_37168,N_36143,N_36856);
nor U37169 (N_37169,N_36674,N_36809);
nor U37170 (N_37170,N_36141,N_36356);
and U37171 (N_37171,N_36911,N_36828);
or U37172 (N_37172,N_36661,N_36669);
nand U37173 (N_37173,N_36843,N_36223);
or U37174 (N_37174,N_36500,N_36950);
and U37175 (N_37175,N_36628,N_36368);
nand U37176 (N_37176,N_36621,N_36299);
and U37177 (N_37177,N_36616,N_36880);
nand U37178 (N_37178,N_36403,N_36465);
nor U37179 (N_37179,N_36227,N_36920);
nand U37180 (N_37180,N_36160,N_36278);
or U37181 (N_37181,N_36005,N_36452);
or U37182 (N_37182,N_36370,N_36605);
and U37183 (N_37183,N_36840,N_36045);
nor U37184 (N_37184,N_36239,N_36096);
xor U37185 (N_37185,N_36266,N_36364);
nor U37186 (N_37186,N_36910,N_36556);
nand U37187 (N_37187,N_36705,N_36769);
and U37188 (N_37188,N_36762,N_36583);
nand U37189 (N_37189,N_36917,N_36753);
or U37190 (N_37190,N_36626,N_36412);
and U37191 (N_37191,N_36587,N_36276);
nor U37192 (N_37192,N_36291,N_36850);
or U37193 (N_37193,N_36433,N_36415);
and U37194 (N_37194,N_36590,N_36343);
xor U37195 (N_37195,N_36847,N_36547);
and U37196 (N_37196,N_36015,N_36182);
or U37197 (N_37197,N_36430,N_36092);
nor U37198 (N_37198,N_36720,N_36977);
xor U37199 (N_37199,N_36132,N_36044);
nor U37200 (N_37200,N_36688,N_36327);
nor U37201 (N_37201,N_36792,N_36863);
nand U37202 (N_37202,N_36240,N_36941);
nand U37203 (N_37203,N_36351,N_36420);
nand U37204 (N_37204,N_36021,N_36989);
xor U37205 (N_37205,N_36545,N_36309);
or U37206 (N_37206,N_36932,N_36960);
xnor U37207 (N_37207,N_36017,N_36011);
and U37208 (N_37208,N_36298,N_36938);
and U37209 (N_37209,N_36599,N_36013);
or U37210 (N_37210,N_36927,N_36527);
nand U37211 (N_37211,N_36757,N_36396);
nand U37212 (N_37212,N_36110,N_36617);
or U37213 (N_37213,N_36574,N_36842);
nor U37214 (N_37214,N_36441,N_36698);
xor U37215 (N_37215,N_36526,N_36780);
nor U37216 (N_37216,N_36710,N_36215);
nor U37217 (N_37217,N_36665,N_36939);
xor U37218 (N_37218,N_36488,N_36640);
xnor U37219 (N_37219,N_36304,N_36602);
xor U37220 (N_37220,N_36329,N_36662);
and U37221 (N_37221,N_36749,N_36164);
or U37222 (N_37222,N_36552,N_36774);
or U37223 (N_37223,N_36064,N_36247);
xnor U37224 (N_37224,N_36006,N_36930);
nor U37225 (N_37225,N_36262,N_36951);
xnor U37226 (N_37226,N_36756,N_36778);
or U37227 (N_37227,N_36633,N_36287);
or U37228 (N_37228,N_36025,N_36333);
nand U37229 (N_37229,N_36767,N_36819);
and U37230 (N_37230,N_36677,N_36101);
nor U37231 (N_37231,N_36534,N_36870);
or U37232 (N_37232,N_36540,N_36982);
nor U37233 (N_37233,N_36646,N_36608);
and U37234 (N_37234,N_36010,N_36221);
xnor U37235 (N_37235,N_36472,N_36034);
xnor U37236 (N_37236,N_36561,N_36542);
or U37237 (N_37237,N_36721,N_36154);
nor U37238 (N_37238,N_36776,N_36634);
nand U37239 (N_37239,N_36077,N_36437);
nor U37240 (N_37240,N_36039,N_36717);
xnor U37241 (N_37241,N_36514,N_36324);
nand U37242 (N_37242,N_36427,N_36632);
and U37243 (N_37243,N_36789,N_36272);
nor U37244 (N_37244,N_36521,N_36051);
nor U37245 (N_37245,N_36697,N_36166);
and U37246 (N_37246,N_36136,N_36269);
and U37247 (N_37247,N_36023,N_36273);
xnor U37248 (N_37248,N_36496,N_36256);
or U37249 (N_37249,N_36424,N_36296);
xor U37250 (N_37250,N_36376,N_36944);
and U37251 (N_37251,N_36603,N_36157);
nor U37252 (N_37252,N_36854,N_36392);
xnor U37253 (N_37253,N_36682,N_36965);
nor U37254 (N_37254,N_36833,N_36076);
nor U37255 (N_37255,N_36563,N_36421);
or U37256 (N_37256,N_36711,N_36838);
xnor U37257 (N_37257,N_36245,N_36904);
xor U37258 (N_37258,N_36252,N_36061);
or U37259 (N_37259,N_36358,N_36919);
or U37260 (N_37260,N_36314,N_36898);
nor U37261 (N_37261,N_36740,N_36174);
nand U37262 (N_37262,N_36146,N_36468);
nor U37263 (N_37263,N_36429,N_36586);
xor U37264 (N_37264,N_36071,N_36884);
nand U37265 (N_37265,N_36012,N_36612);
nor U37266 (N_37266,N_36207,N_36879);
xor U37267 (N_37267,N_36836,N_36693);
nand U37268 (N_37268,N_36837,N_36168);
nand U37269 (N_37269,N_36476,N_36385);
or U37270 (N_37270,N_36102,N_36844);
or U37271 (N_37271,N_36625,N_36785);
and U37272 (N_37272,N_36261,N_36002);
xnor U37273 (N_37273,N_36172,N_36375);
nor U37274 (N_37274,N_36933,N_36251);
xor U37275 (N_37275,N_36095,N_36125);
or U37276 (N_37276,N_36338,N_36593);
nor U37277 (N_37277,N_36155,N_36830);
xor U37278 (N_37278,N_36121,N_36528);
nand U37279 (N_37279,N_36957,N_36347);
nor U37280 (N_37280,N_36872,N_36078);
nor U37281 (N_37281,N_36228,N_36811);
nand U37282 (N_37282,N_36417,N_36443);
xor U37283 (N_37283,N_36874,N_36614);
nand U37284 (N_37284,N_36033,N_36642);
nand U37285 (N_37285,N_36871,N_36425);
nor U37286 (N_37286,N_36600,N_36656);
nand U37287 (N_37287,N_36029,N_36622);
xor U37288 (N_37288,N_36159,N_36654);
nand U37289 (N_37289,N_36307,N_36188);
xnor U37290 (N_37290,N_36916,N_36784);
and U37291 (N_37291,N_36579,N_36162);
and U37292 (N_37292,N_36473,N_36718);
nor U37293 (N_37293,N_36259,N_36592);
nor U37294 (N_37294,N_36797,N_36881);
nor U37295 (N_37295,N_36869,N_36175);
or U37296 (N_37296,N_36196,N_36243);
or U37297 (N_37297,N_36313,N_36184);
or U37298 (N_37298,N_36649,N_36503);
xnor U37299 (N_37299,N_36541,N_36671);
and U37300 (N_37300,N_36958,N_36310);
nor U37301 (N_37301,N_36652,N_36859);
nor U37302 (N_37302,N_36585,N_36846);
nor U37303 (N_37303,N_36899,N_36504);
nand U37304 (N_37304,N_36004,N_36897);
nand U37305 (N_37305,N_36976,N_36334);
nor U37306 (N_37306,N_36079,N_36630);
nand U37307 (N_37307,N_36306,N_36281);
and U37308 (N_37308,N_36073,N_36609);
xnor U37309 (N_37309,N_36734,N_36210);
nand U37310 (N_37310,N_36036,N_36773);
and U37311 (N_37311,N_36187,N_36454);
nand U37312 (N_37312,N_36179,N_36748);
xor U37313 (N_37313,N_36572,N_36974);
xor U37314 (N_37314,N_36568,N_36730);
or U37315 (N_37315,N_36584,N_36980);
nand U37316 (N_37316,N_36582,N_36535);
nor U37317 (N_37317,N_36759,N_36529);
xor U37318 (N_37318,N_36554,N_36349);
nor U37319 (N_37319,N_36516,N_36072);
xor U37320 (N_37320,N_36047,N_36754);
and U37321 (N_37321,N_36994,N_36301);
nor U37322 (N_37322,N_36274,N_36134);
xor U37323 (N_37323,N_36408,N_36026);
and U37324 (N_37324,N_36419,N_36901);
nand U37325 (N_37325,N_36907,N_36435);
nor U37326 (N_37326,N_36031,N_36779);
nand U37327 (N_37327,N_36531,N_36741);
xor U37328 (N_37328,N_36673,N_36515);
and U37329 (N_37329,N_36931,N_36389);
nand U37330 (N_37330,N_36831,N_36332);
and U37331 (N_37331,N_36925,N_36050);
nand U37332 (N_37332,N_36997,N_36746);
and U37333 (N_37333,N_36804,N_36549);
or U37334 (N_37334,N_36795,N_36486);
or U37335 (N_37335,N_36163,N_36834);
and U37336 (N_37336,N_36000,N_36601);
xnor U37337 (N_37337,N_36875,N_36610);
or U37338 (N_37338,N_36808,N_36321);
nand U37339 (N_37339,N_36341,N_36100);
nand U37340 (N_37340,N_36712,N_36204);
and U37341 (N_37341,N_36851,N_36685);
nand U37342 (N_37342,N_36127,N_36969);
nor U37343 (N_37343,N_36469,N_36890);
and U37344 (N_37344,N_36975,N_36946);
nand U37345 (N_37345,N_36943,N_36464);
nor U37346 (N_37346,N_36180,N_36562);
or U37347 (N_37347,N_36760,N_36812);
and U37348 (N_37348,N_36893,N_36201);
xnor U37349 (N_37349,N_36707,N_36242);
nor U37350 (N_37350,N_36275,N_36888);
xnor U37351 (N_37351,N_36319,N_36457);
or U37352 (N_37352,N_36399,N_36675);
and U37353 (N_37353,N_36144,N_36264);
nor U37354 (N_37354,N_36559,N_36097);
nor U37355 (N_37355,N_36397,N_36354);
and U37356 (N_37356,N_36020,N_36735);
and U37357 (N_37357,N_36714,N_36581);
or U37358 (N_37358,N_36611,N_36510);
xnor U37359 (N_37359,N_36199,N_36485);
nand U37360 (N_37360,N_36566,N_36106);
and U37361 (N_37361,N_36986,N_36737);
or U37362 (N_37362,N_36075,N_36860);
or U37363 (N_37363,N_36194,N_36903);
and U37364 (N_37364,N_36378,N_36410);
xnor U37365 (N_37365,N_36873,N_36206);
or U37366 (N_37366,N_36277,N_36953);
or U37367 (N_37367,N_36362,N_36524);
xnor U37368 (N_37368,N_36487,N_36238);
or U37369 (N_37369,N_36672,N_36119);
nor U37370 (N_37370,N_36548,N_36543);
nor U37371 (N_37371,N_36791,N_36400);
nor U37372 (N_37372,N_36922,N_36887);
or U37373 (N_37373,N_36404,N_36086);
nand U37374 (N_37374,N_36772,N_36763);
nand U37375 (N_37375,N_36832,N_36744);
nand U37376 (N_37376,N_36371,N_36878);
nand U37377 (N_37377,N_36178,N_36620);
xnor U37378 (N_37378,N_36191,N_36148);
nand U37379 (N_37379,N_36973,N_36618);
nand U37380 (N_37380,N_36462,N_36886);
and U37381 (N_37381,N_36035,N_36491);
nand U37382 (N_37382,N_36497,N_36444);
or U37383 (N_37383,N_36083,N_36232);
nand U37384 (N_37384,N_36810,N_36948);
xor U37385 (N_37385,N_36137,N_36248);
nor U37386 (N_37386,N_36522,N_36117);
and U37387 (N_37387,N_36323,N_36126);
and U37388 (N_37388,N_36750,N_36231);
nand U37389 (N_37389,N_36629,N_36416);
nand U37390 (N_37390,N_36690,N_36996);
nand U37391 (N_37391,N_36470,N_36765);
and U37392 (N_37392,N_36679,N_36258);
xor U37393 (N_37393,N_36224,N_36165);
xor U37394 (N_37394,N_36116,N_36787);
nand U37395 (N_37395,N_36567,N_36678);
nor U37396 (N_37396,N_36214,N_36519);
nand U37397 (N_37397,N_36365,N_36537);
nand U37398 (N_37398,N_36434,N_36093);
and U37399 (N_37399,N_36422,N_36889);
nor U37400 (N_37400,N_36286,N_36959);
nor U37401 (N_37401,N_36255,N_36484);
and U37402 (N_37402,N_36580,N_36739);
nand U37403 (N_37403,N_36659,N_36999);
xor U37404 (N_37404,N_36105,N_36411);
and U37405 (N_37405,N_36355,N_36131);
xnor U37406 (N_37406,N_36059,N_36868);
or U37407 (N_37407,N_36145,N_36650);
and U37408 (N_37408,N_36553,N_36192);
nor U37409 (N_37409,N_36967,N_36849);
nor U37410 (N_37410,N_36479,N_36315);
xor U37411 (N_37411,N_36507,N_36171);
nand U37412 (N_37412,N_36268,N_36538);
or U37413 (N_37413,N_36230,N_36369);
nand U37414 (N_37414,N_36934,N_36706);
and U37415 (N_37415,N_36244,N_36211);
xnor U37416 (N_37416,N_36942,N_36908);
and U37417 (N_37417,N_36294,N_36480);
xor U37418 (N_37418,N_36694,N_36805);
xor U37419 (N_37419,N_36512,N_36557);
and U37420 (N_37420,N_36019,N_36835);
or U37421 (N_37421,N_36738,N_36198);
nor U37422 (N_37422,N_36481,N_36359);
or U37423 (N_37423,N_36940,N_36995);
nor U37424 (N_37424,N_36234,N_36923);
nand U37425 (N_37425,N_36702,N_36466);
or U37426 (N_37426,N_36054,N_36340);
nor U37427 (N_37427,N_36877,N_36483);
and U37428 (N_37428,N_36099,N_36984);
or U37429 (N_37429,N_36722,N_36169);
or U37430 (N_37430,N_36185,N_36379);
or U37431 (N_37431,N_36225,N_36533);
nor U37432 (N_37432,N_36815,N_36193);
nor U37433 (N_37433,N_36062,N_36798);
nor U37434 (N_37434,N_36857,N_36676);
nor U37435 (N_37435,N_36680,N_36696);
nand U37436 (N_37436,N_36209,N_36639);
or U37437 (N_37437,N_36055,N_36014);
nor U37438 (N_37438,N_36081,N_36135);
or U37439 (N_37439,N_36635,N_36725);
and U37440 (N_37440,N_36786,N_36508);
xor U37441 (N_37441,N_36442,N_36361);
or U37442 (N_37442,N_36751,N_36892);
nand U37443 (N_37443,N_36254,N_36704);
nand U37444 (N_37444,N_36867,N_36413);
or U37445 (N_37445,N_36057,N_36518);
xor U37446 (N_37446,N_36363,N_36807);
and U37447 (N_37447,N_36800,N_36794);
nor U37448 (N_37448,N_36118,N_36111);
nand U37449 (N_37449,N_36293,N_36569);
nand U37450 (N_37450,N_36374,N_36048);
or U37451 (N_37451,N_36233,N_36827);
xnor U37452 (N_37452,N_36205,N_36848);
or U37453 (N_37453,N_36394,N_36716);
nor U37454 (N_37454,N_36128,N_36390);
and U37455 (N_37455,N_36576,N_36439);
or U37456 (N_37456,N_36821,N_36530);
or U37457 (N_37457,N_36826,N_36558);
nand U37458 (N_37458,N_36353,N_36405);
or U37459 (N_37459,N_36766,N_36505);
and U37460 (N_37460,N_36921,N_36129);
and U37461 (N_37461,N_36523,N_36906);
xnor U37462 (N_37462,N_36167,N_36520);
nand U37463 (N_37463,N_36801,N_36891);
nor U37464 (N_37464,N_36407,N_36279);
nor U37465 (N_37465,N_36956,N_36009);
nand U37466 (N_37466,N_36972,N_36037);
nor U37467 (N_37467,N_36350,N_36981);
or U37468 (N_37468,N_36708,N_36731);
or U37469 (N_37469,N_36758,N_36391);
and U37470 (N_37470,N_36564,N_36495);
and U37471 (N_37471,N_36068,N_36216);
and U37472 (N_37472,N_36022,N_36641);
nor U37473 (N_37473,N_36993,N_36176);
and U37474 (N_37474,N_36814,N_36058);
and U37475 (N_37475,N_36742,N_36318);
or U37476 (N_37476,N_36684,N_36667);
nor U37477 (N_37477,N_36743,N_36978);
nor U37478 (N_37478,N_36229,N_36133);
xnor U37479 (N_37479,N_36732,N_36502);
or U37480 (N_37480,N_36990,N_36715);
nand U37481 (N_37481,N_36387,N_36985);
nor U37482 (N_37482,N_36112,N_36292);
nand U37483 (N_37483,N_36788,N_36498);
nor U37484 (N_37484,N_36595,N_36589);
xor U37485 (N_37485,N_36902,N_36591);
xor U37486 (N_37486,N_36383,N_36346);
and U37487 (N_37487,N_36853,N_36866);
nand U37488 (N_37488,N_36604,N_36729);
or U37489 (N_37489,N_36768,N_36962);
xnor U37490 (N_37490,N_36241,N_36114);
and U37491 (N_37491,N_36195,N_36703);
or U37492 (N_37492,N_36446,N_36056);
nor U37493 (N_37493,N_36509,N_36709);
xnor U37494 (N_37494,N_36492,N_36032);
nand U37495 (N_37495,N_36573,N_36988);
nor U37496 (N_37496,N_36876,N_36594);
or U37497 (N_37497,N_36142,N_36655);
xor U37498 (N_37498,N_36912,N_36459);
and U37499 (N_37499,N_36360,N_36624);
or U37500 (N_37500,N_36856,N_36031);
or U37501 (N_37501,N_36302,N_36058);
nand U37502 (N_37502,N_36824,N_36021);
nor U37503 (N_37503,N_36070,N_36170);
nor U37504 (N_37504,N_36913,N_36479);
or U37505 (N_37505,N_36597,N_36002);
nor U37506 (N_37506,N_36388,N_36220);
or U37507 (N_37507,N_36230,N_36070);
or U37508 (N_37508,N_36911,N_36807);
nand U37509 (N_37509,N_36676,N_36590);
or U37510 (N_37510,N_36360,N_36676);
and U37511 (N_37511,N_36954,N_36387);
or U37512 (N_37512,N_36353,N_36842);
nor U37513 (N_37513,N_36603,N_36007);
xnor U37514 (N_37514,N_36998,N_36825);
xnor U37515 (N_37515,N_36016,N_36928);
nor U37516 (N_37516,N_36309,N_36387);
nand U37517 (N_37517,N_36724,N_36879);
nor U37518 (N_37518,N_36615,N_36013);
nor U37519 (N_37519,N_36692,N_36403);
or U37520 (N_37520,N_36717,N_36307);
nand U37521 (N_37521,N_36860,N_36088);
and U37522 (N_37522,N_36650,N_36412);
or U37523 (N_37523,N_36946,N_36805);
xor U37524 (N_37524,N_36146,N_36603);
or U37525 (N_37525,N_36692,N_36546);
nand U37526 (N_37526,N_36747,N_36272);
or U37527 (N_37527,N_36583,N_36816);
nor U37528 (N_37528,N_36480,N_36080);
xnor U37529 (N_37529,N_36921,N_36627);
nor U37530 (N_37530,N_36249,N_36168);
or U37531 (N_37531,N_36259,N_36752);
nor U37532 (N_37532,N_36870,N_36233);
nand U37533 (N_37533,N_36054,N_36989);
and U37534 (N_37534,N_36759,N_36073);
and U37535 (N_37535,N_36132,N_36885);
nor U37536 (N_37536,N_36520,N_36375);
and U37537 (N_37537,N_36703,N_36322);
nand U37538 (N_37538,N_36044,N_36281);
or U37539 (N_37539,N_36489,N_36609);
or U37540 (N_37540,N_36707,N_36710);
nand U37541 (N_37541,N_36190,N_36155);
xor U37542 (N_37542,N_36485,N_36333);
xor U37543 (N_37543,N_36716,N_36111);
nor U37544 (N_37544,N_36359,N_36665);
and U37545 (N_37545,N_36141,N_36146);
and U37546 (N_37546,N_36182,N_36203);
xor U37547 (N_37547,N_36230,N_36728);
and U37548 (N_37548,N_36380,N_36024);
nor U37549 (N_37549,N_36708,N_36278);
xnor U37550 (N_37550,N_36141,N_36769);
or U37551 (N_37551,N_36862,N_36109);
or U37552 (N_37552,N_36057,N_36302);
nor U37553 (N_37553,N_36810,N_36946);
xnor U37554 (N_37554,N_36391,N_36538);
or U37555 (N_37555,N_36700,N_36687);
nor U37556 (N_37556,N_36119,N_36716);
or U37557 (N_37557,N_36157,N_36760);
nor U37558 (N_37558,N_36644,N_36222);
xor U37559 (N_37559,N_36822,N_36050);
or U37560 (N_37560,N_36824,N_36380);
nand U37561 (N_37561,N_36627,N_36874);
or U37562 (N_37562,N_36497,N_36245);
xor U37563 (N_37563,N_36864,N_36576);
nor U37564 (N_37564,N_36752,N_36960);
nand U37565 (N_37565,N_36941,N_36654);
or U37566 (N_37566,N_36816,N_36096);
nand U37567 (N_37567,N_36652,N_36114);
or U37568 (N_37568,N_36102,N_36799);
nor U37569 (N_37569,N_36048,N_36663);
nand U37570 (N_37570,N_36490,N_36910);
nand U37571 (N_37571,N_36096,N_36727);
nor U37572 (N_37572,N_36001,N_36125);
xnor U37573 (N_37573,N_36145,N_36676);
and U37574 (N_37574,N_36689,N_36641);
nor U37575 (N_37575,N_36542,N_36609);
nand U37576 (N_37576,N_36543,N_36896);
nor U37577 (N_37577,N_36948,N_36983);
nand U37578 (N_37578,N_36044,N_36673);
or U37579 (N_37579,N_36321,N_36701);
nand U37580 (N_37580,N_36219,N_36973);
and U37581 (N_37581,N_36048,N_36806);
and U37582 (N_37582,N_36704,N_36998);
and U37583 (N_37583,N_36754,N_36787);
nor U37584 (N_37584,N_36216,N_36562);
and U37585 (N_37585,N_36877,N_36691);
and U37586 (N_37586,N_36808,N_36386);
nor U37587 (N_37587,N_36198,N_36571);
or U37588 (N_37588,N_36636,N_36607);
and U37589 (N_37589,N_36059,N_36745);
xor U37590 (N_37590,N_36108,N_36063);
nor U37591 (N_37591,N_36902,N_36581);
nor U37592 (N_37592,N_36363,N_36332);
and U37593 (N_37593,N_36999,N_36457);
nand U37594 (N_37594,N_36294,N_36845);
and U37595 (N_37595,N_36437,N_36040);
nor U37596 (N_37596,N_36810,N_36083);
nand U37597 (N_37597,N_36419,N_36048);
nor U37598 (N_37598,N_36197,N_36824);
xnor U37599 (N_37599,N_36781,N_36008);
and U37600 (N_37600,N_36684,N_36677);
and U37601 (N_37601,N_36728,N_36482);
or U37602 (N_37602,N_36513,N_36237);
or U37603 (N_37603,N_36965,N_36061);
xnor U37604 (N_37604,N_36022,N_36096);
xor U37605 (N_37605,N_36452,N_36415);
and U37606 (N_37606,N_36876,N_36862);
or U37607 (N_37607,N_36629,N_36443);
xor U37608 (N_37608,N_36122,N_36630);
and U37609 (N_37609,N_36632,N_36245);
xnor U37610 (N_37610,N_36288,N_36179);
nor U37611 (N_37611,N_36957,N_36115);
nor U37612 (N_37612,N_36475,N_36530);
nand U37613 (N_37613,N_36308,N_36425);
and U37614 (N_37614,N_36026,N_36561);
nor U37615 (N_37615,N_36326,N_36413);
xnor U37616 (N_37616,N_36564,N_36100);
nand U37617 (N_37617,N_36115,N_36692);
and U37618 (N_37618,N_36149,N_36252);
nor U37619 (N_37619,N_36219,N_36794);
xnor U37620 (N_37620,N_36900,N_36721);
nor U37621 (N_37621,N_36743,N_36334);
nor U37622 (N_37622,N_36603,N_36386);
nand U37623 (N_37623,N_36255,N_36293);
nand U37624 (N_37624,N_36242,N_36189);
nor U37625 (N_37625,N_36288,N_36040);
nor U37626 (N_37626,N_36747,N_36421);
xnor U37627 (N_37627,N_36566,N_36972);
nand U37628 (N_37628,N_36388,N_36765);
nor U37629 (N_37629,N_36886,N_36240);
and U37630 (N_37630,N_36094,N_36823);
xnor U37631 (N_37631,N_36160,N_36075);
nand U37632 (N_37632,N_36934,N_36571);
xnor U37633 (N_37633,N_36014,N_36464);
nor U37634 (N_37634,N_36948,N_36601);
nand U37635 (N_37635,N_36192,N_36289);
or U37636 (N_37636,N_36676,N_36764);
xor U37637 (N_37637,N_36745,N_36585);
or U37638 (N_37638,N_36667,N_36783);
or U37639 (N_37639,N_36962,N_36781);
or U37640 (N_37640,N_36811,N_36340);
and U37641 (N_37641,N_36154,N_36882);
or U37642 (N_37642,N_36923,N_36278);
nand U37643 (N_37643,N_36834,N_36990);
or U37644 (N_37644,N_36048,N_36946);
nand U37645 (N_37645,N_36874,N_36699);
nor U37646 (N_37646,N_36667,N_36043);
nor U37647 (N_37647,N_36829,N_36735);
nand U37648 (N_37648,N_36926,N_36343);
nand U37649 (N_37649,N_36843,N_36890);
xor U37650 (N_37650,N_36348,N_36531);
nor U37651 (N_37651,N_36150,N_36185);
and U37652 (N_37652,N_36039,N_36595);
or U37653 (N_37653,N_36499,N_36039);
nor U37654 (N_37654,N_36888,N_36663);
xnor U37655 (N_37655,N_36555,N_36465);
nor U37656 (N_37656,N_36767,N_36261);
xnor U37657 (N_37657,N_36951,N_36641);
or U37658 (N_37658,N_36603,N_36013);
nor U37659 (N_37659,N_36766,N_36144);
nor U37660 (N_37660,N_36513,N_36680);
nor U37661 (N_37661,N_36263,N_36742);
xnor U37662 (N_37662,N_36472,N_36803);
and U37663 (N_37663,N_36066,N_36606);
and U37664 (N_37664,N_36294,N_36086);
nand U37665 (N_37665,N_36866,N_36924);
nor U37666 (N_37666,N_36156,N_36438);
xor U37667 (N_37667,N_36534,N_36176);
xnor U37668 (N_37668,N_36752,N_36123);
nor U37669 (N_37669,N_36301,N_36628);
xor U37670 (N_37670,N_36355,N_36493);
xnor U37671 (N_37671,N_36980,N_36930);
and U37672 (N_37672,N_36290,N_36200);
and U37673 (N_37673,N_36631,N_36681);
nor U37674 (N_37674,N_36029,N_36344);
or U37675 (N_37675,N_36674,N_36961);
xor U37676 (N_37676,N_36419,N_36806);
and U37677 (N_37677,N_36348,N_36175);
xor U37678 (N_37678,N_36119,N_36833);
xnor U37679 (N_37679,N_36537,N_36147);
or U37680 (N_37680,N_36650,N_36240);
nand U37681 (N_37681,N_36619,N_36623);
or U37682 (N_37682,N_36203,N_36088);
or U37683 (N_37683,N_36907,N_36585);
xnor U37684 (N_37684,N_36171,N_36660);
or U37685 (N_37685,N_36510,N_36166);
nor U37686 (N_37686,N_36686,N_36301);
and U37687 (N_37687,N_36108,N_36653);
or U37688 (N_37688,N_36172,N_36077);
and U37689 (N_37689,N_36907,N_36670);
and U37690 (N_37690,N_36060,N_36534);
xnor U37691 (N_37691,N_36445,N_36859);
or U37692 (N_37692,N_36391,N_36676);
or U37693 (N_37693,N_36681,N_36546);
and U37694 (N_37694,N_36329,N_36486);
xor U37695 (N_37695,N_36423,N_36429);
and U37696 (N_37696,N_36132,N_36696);
nor U37697 (N_37697,N_36745,N_36269);
or U37698 (N_37698,N_36978,N_36767);
nand U37699 (N_37699,N_36049,N_36781);
or U37700 (N_37700,N_36071,N_36093);
xnor U37701 (N_37701,N_36857,N_36023);
nor U37702 (N_37702,N_36833,N_36802);
and U37703 (N_37703,N_36096,N_36142);
or U37704 (N_37704,N_36551,N_36602);
xor U37705 (N_37705,N_36724,N_36183);
nor U37706 (N_37706,N_36831,N_36023);
nand U37707 (N_37707,N_36370,N_36716);
nor U37708 (N_37708,N_36377,N_36838);
and U37709 (N_37709,N_36265,N_36032);
xnor U37710 (N_37710,N_36838,N_36494);
and U37711 (N_37711,N_36334,N_36782);
nand U37712 (N_37712,N_36657,N_36171);
nor U37713 (N_37713,N_36694,N_36142);
or U37714 (N_37714,N_36543,N_36070);
or U37715 (N_37715,N_36504,N_36033);
and U37716 (N_37716,N_36148,N_36710);
xnor U37717 (N_37717,N_36740,N_36617);
nor U37718 (N_37718,N_36684,N_36048);
and U37719 (N_37719,N_36117,N_36112);
nor U37720 (N_37720,N_36532,N_36530);
xor U37721 (N_37721,N_36926,N_36005);
xnor U37722 (N_37722,N_36510,N_36111);
nand U37723 (N_37723,N_36566,N_36830);
or U37724 (N_37724,N_36679,N_36703);
or U37725 (N_37725,N_36943,N_36300);
nor U37726 (N_37726,N_36662,N_36202);
and U37727 (N_37727,N_36585,N_36544);
nor U37728 (N_37728,N_36814,N_36844);
nand U37729 (N_37729,N_36291,N_36615);
nand U37730 (N_37730,N_36869,N_36212);
xor U37731 (N_37731,N_36837,N_36041);
xor U37732 (N_37732,N_36881,N_36028);
or U37733 (N_37733,N_36885,N_36988);
nor U37734 (N_37734,N_36495,N_36527);
nand U37735 (N_37735,N_36576,N_36454);
xnor U37736 (N_37736,N_36278,N_36075);
xor U37737 (N_37737,N_36118,N_36426);
or U37738 (N_37738,N_36046,N_36735);
and U37739 (N_37739,N_36368,N_36117);
and U37740 (N_37740,N_36285,N_36870);
or U37741 (N_37741,N_36232,N_36905);
nand U37742 (N_37742,N_36329,N_36285);
nor U37743 (N_37743,N_36509,N_36653);
nand U37744 (N_37744,N_36336,N_36841);
and U37745 (N_37745,N_36467,N_36925);
xor U37746 (N_37746,N_36782,N_36615);
and U37747 (N_37747,N_36604,N_36514);
nand U37748 (N_37748,N_36892,N_36163);
nor U37749 (N_37749,N_36647,N_36514);
or U37750 (N_37750,N_36040,N_36543);
xor U37751 (N_37751,N_36985,N_36243);
xnor U37752 (N_37752,N_36146,N_36109);
xnor U37753 (N_37753,N_36918,N_36052);
xnor U37754 (N_37754,N_36671,N_36783);
xor U37755 (N_37755,N_36120,N_36363);
nand U37756 (N_37756,N_36105,N_36377);
and U37757 (N_37757,N_36975,N_36123);
xnor U37758 (N_37758,N_36146,N_36259);
nand U37759 (N_37759,N_36677,N_36757);
nor U37760 (N_37760,N_36459,N_36168);
or U37761 (N_37761,N_36383,N_36434);
nand U37762 (N_37762,N_36491,N_36993);
nand U37763 (N_37763,N_36506,N_36203);
or U37764 (N_37764,N_36773,N_36211);
nor U37765 (N_37765,N_36333,N_36691);
nand U37766 (N_37766,N_36916,N_36716);
or U37767 (N_37767,N_36950,N_36238);
or U37768 (N_37768,N_36991,N_36435);
nor U37769 (N_37769,N_36670,N_36249);
nand U37770 (N_37770,N_36070,N_36585);
and U37771 (N_37771,N_36655,N_36614);
and U37772 (N_37772,N_36303,N_36772);
or U37773 (N_37773,N_36526,N_36051);
or U37774 (N_37774,N_36967,N_36534);
nor U37775 (N_37775,N_36462,N_36669);
xnor U37776 (N_37776,N_36344,N_36702);
or U37777 (N_37777,N_36681,N_36730);
nor U37778 (N_37778,N_36508,N_36379);
xnor U37779 (N_37779,N_36021,N_36622);
xnor U37780 (N_37780,N_36141,N_36478);
and U37781 (N_37781,N_36850,N_36885);
nand U37782 (N_37782,N_36801,N_36450);
or U37783 (N_37783,N_36776,N_36574);
and U37784 (N_37784,N_36932,N_36795);
xor U37785 (N_37785,N_36697,N_36599);
nand U37786 (N_37786,N_36765,N_36274);
or U37787 (N_37787,N_36654,N_36734);
and U37788 (N_37788,N_36924,N_36440);
and U37789 (N_37789,N_36090,N_36382);
or U37790 (N_37790,N_36968,N_36940);
or U37791 (N_37791,N_36044,N_36454);
and U37792 (N_37792,N_36236,N_36545);
xor U37793 (N_37793,N_36366,N_36443);
nor U37794 (N_37794,N_36060,N_36017);
xor U37795 (N_37795,N_36995,N_36111);
nand U37796 (N_37796,N_36154,N_36008);
or U37797 (N_37797,N_36317,N_36403);
nand U37798 (N_37798,N_36557,N_36678);
nor U37799 (N_37799,N_36817,N_36396);
or U37800 (N_37800,N_36815,N_36653);
nor U37801 (N_37801,N_36256,N_36028);
and U37802 (N_37802,N_36056,N_36212);
nor U37803 (N_37803,N_36982,N_36326);
xor U37804 (N_37804,N_36571,N_36606);
and U37805 (N_37805,N_36831,N_36746);
nor U37806 (N_37806,N_36305,N_36185);
or U37807 (N_37807,N_36536,N_36879);
nand U37808 (N_37808,N_36709,N_36688);
or U37809 (N_37809,N_36545,N_36405);
nand U37810 (N_37810,N_36662,N_36480);
xnor U37811 (N_37811,N_36781,N_36816);
and U37812 (N_37812,N_36872,N_36932);
nand U37813 (N_37813,N_36377,N_36645);
xor U37814 (N_37814,N_36097,N_36317);
xor U37815 (N_37815,N_36890,N_36498);
xor U37816 (N_37816,N_36110,N_36385);
or U37817 (N_37817,N_36810,N_36819);
nand U37818 (N_37818,N_36284,N_36610);
or U37819 (N_37819,N_36685,N_36979);
and U37820 (N_37820,N_36508,N_36565);
nand U37821 (N_37821,N_36287,N_36147);
or U37822 (N_37822,N_36388,N_36277);
or U37823 (N_37823,N_36900,N_36862);
nand U37824 (N_37824,N_36548,N_36564);
and U37825 (N_37825,N_36899,N_36301);
nor U37826 (N_37826,N_36430,N_36583);
nor U37827 (N_37827,N_36418,N_36096);
nand U37828 (N_37828,N_36491,N_36666);
and U37829 (N_37829,N_36405,N_36883);
nor U37830 (N_37830,N_36383,N_36007);
or U37831 (N_37831,N_36785,N_36309);
xor U37832 (N_37832,N_36973,N_36445);
xnor U37833 (N_37833,N_36208,N_36731);
xor U37834 (N_37834,N_36649,N_36036);
and U37835 (N_37835,N_36789,N_36268);
and U37836 (N_37836,N_36008,N_36513);
or U37837 (N_37837,N_36872,N_36255);
nand U37838 (N_37838,N_36042,N_36354);
nand U37839 (N_37839,N_36176,N_36745);
or U37840 (N_37840,N_36187,N_36908);
and U37841 (N_37841,N_36729,N_36115);
xnor U37842 (N_37842,N_36652,N_36032);
nand U37843 (N_37843,N_36773,N_36858);
nand U37844 (N_37844,N_36004,N_36272);
or U37845 (N_37845,N_36630,N_36533);
xor U37846 (N_37846,N_36261,N_36474);
nor U37847 (N_37847,N_36581,N_36530);
nor U37848 (N_37848,N_36030,N_36347);
or U37849 (N_37849,N_36659,N_36015);
xnor U37850 (N_37850,N_36224,N_36909);
xnor U37851 (N_37851,N_36584,N_36019);
or U37852 (N_37852,N_36510,N_36008);
and U37853 (N_37853,N_36315,N_36330);
nand U37854 (N_37854,N_36461,N_36923);
and U37855 (N_37855,N_36812,N_36595);
or U37856 (N_37856,N_36180,N_36817);
nand U37857 (N_37857,N_36477,N_36741);
nor U37858 (N_37858,N_36598,N_36125);
nand U37859 (N_37859,N_36803,N_36397);
or U37860 (N_37860,N_36952,N_36757);
xor U37861 (N_37861,N_36898,N_36135);
nor U37862 (N_37862,N_36560,N_36859);
nor U37863 (N_37863,N_36518,N_36245);
nor U37864 (N_37864,N_36723,N_36471);
or U37865 (N_37865,N_36624,N_36371);
xor U37866 (N_37866,N_36809,N_36442);
or U37867 (N_37867,N_36126,N_36521);
xnor U37868 (N_37868,N_36215,N_36167);
and U37869 (N_37869,N_36748,N_36286);
nor U37870 (N_37870,N_36401,N_36113);
xnor U37871 (N_37871,N_36302,N_36895);
nor U37872 (N_37872,N_36210,N_36687);
and U37873 (N_37873,N_36722,N_36756);
and U37874 (N_37874,N_36716,N_36859);
or U37875 (N_37875,N_36390,N_36833);
or U37876 (N_37876,N_36758,N_36581);
or U37877 (N_37877,N_36606,N_36912);
nor U37878 (N_37878,N_36406,N_36276);
or U37879 (N_37879,N_36743,N_36511);
or U37880 (N_37880,N_36154,N_36661);
nand U37881 (N_37881,N_36724,N_36918);
nor U37882 (N_37882,N_36829,N_36540);
nor U37883 (N_37883,N_36137,N_36613);
nand U37884 (N_37884,N_36891,N_36666);
and U37885 (N_37885,N_36491,N_36331);
nand U37886 (N_37886,N_36321,N_36081);
xnor U37887 (N_37887,N_36915,N_36261);
nor U37888 (N_37888,N_36366,N_36232);
nor U37889 (N_37889,N_36226,N_36774);
and U37890 (N_37890,N_36576,N_36360);
nor U37891 (N_37891,N_36196,N_36673);
nand U37892 (N_37892,N_36168,N_36343);
and U37893 (N_37893,N_36671,N_36124);
xor U37894 (N_37894,N_36148,N_36722);
and U37895 (N_37895,N_36233,N_36293);
xor U37896 (N_37896,N_36486,N_36721);
nand U37897 (N_37897,N_36203,N_36431);
or U37898 (N_37898,N_36393,N_36341);
nor U37899 (N_37899,N_36210,N_36464);
xor U37900 (N_37900,N_36402,N_36868);
nor U37901 (N_37901,N_36898,N_36981);
xor U37902 (N_37902,N_36464,N_36892);
or U37903 (N_37903,N_36711,N_36759);
and U37904 (N_37904,N_36110,N_36634);
xnor U37905 (N_37905,N_36490,N_36047);
or U37906 (N_37906,N_36162,N_36938);
and U37907 (N_37907,N_36162,N_36197);
or U37908 (N_37908,N_36727,N_36689);
nor U37909 (N_37909,N_36548,N_36896);
nand U37910 (N_37910,N_36581,N_36518);
nor U37911 (N_37911,N_36458,N_36664);
or U37912 (N_37912,N_36626,N_36877);
nor U37913 (N_37913,N_36753,N_36610);
nand U37914 (N_37914,N_36410,N_36934);
xnor U37915 (N_37915,N_36238,N_36101);
nor U37916 (N_37916,N_36807,N_36582);
or U37917 (N_37917,N_36292,N_36919);
xnor U37918 (N_37918,N_36916,N_36865);
or U37919 (N_37919,N_36921,N_36654);
and U37920 (N_37920,N_36766,N_36213);
nand U37921 (N_37921,N_36122,N_36337);
nor U37922 (N_37922,N_36882,N_36147);
and U37923 (N_37923,N_36755,N_36577);
nor U37924 (N_37924,N_36468,N_36056);
and U37925 (N_37925,N_36574,N_36853);
or U37926 (N_37926,N_36106,N_36290);
nand U37927 (N_37927,N_36782,N_36458);
xnor U37928 (N_37928,N_36250,N_36678);
or U37929 (N_37929,N_36892,N_36221);
nand U37930 (N_37930,N_36848,N_36413);
xnor U37931 (N_37931,N_36769,N_36380);
xnor U37932 (N_37932,N_36233,N_36323);
nor U37933 (N_37933,N_36213,N_36168);
nor U37934 (N_37934,N_36426,N_36772);
or U37935 (N_37935,N_36375,N_36374);
or U37936 (N_37936,N_36830,N_36347);
or U37937 (N_37937,N_36012,N_36730);
and U37938 (N_37938,N_36748,N_36016);
xnor U37939 (N_37939,N_36355,N_36707);
nand U37940 (N_37940,N_36706,N_36025);
nand U37941 (N_37941,N_36467,N_36239);
and U37942 (N_37942,N_36413,N_36725);
xnor U37943 (N_37943,N_36367,N_36693);
and U37944 (N_37944,N_36465,N_36341);
nor U37945 (N_37945,N_36375,N_36280);
nor U37946 (N_37946,N_36465,N_36280);
nor U37947 (N_37947,N_36367,N_36002);
and U37948 (N_37948,N_36225,N_36532);
and U37949 (N_37949,N_36829,N_36661);
nand U37950 (N_37950,N_36898,N_36498);
nor U37951 (N_37951,N_36612,N_36764);
xnor U37952 (N_37952,N_36228,N_36551);
and U37953 (N_37953,N_36770,N_36388);
and U37954 (N_37954,N_36558,N_36255);
and U37955 (N_37955,N_36223,N_36507);
nor U37956 (N_37956,N_36047,N_36383);
and U37957 (N_37957,N_36412,N_36078);
or U37958 (N_37958,N_36592,N_36726);
and U37959 (N_37959,N_36783,N_36504);
and U37960 (N_37960,N_36198,N_36826);
and U37961 (N_37961,N_36922,N_36747);
and U37962 (N_37962,N_36241,N_36204);
xnor U37963 (N_37963,N_36777,N_36787);
nand U37964 (N_37964,N_36830,N_36179);
or U37965 (N_37965,N_36164,N_36206);
xor U37966 (N_37966,N_36355,N_36874);
or U37967 (N_37967,N_36268,N_36114);
or U37968 (N_37968,N_36094,N_36735);
nor U37969 (N_37969,N_36889,N_36330);
and U37970 (N_37970,N_36844,N_36229);
and U37971 (N_37971,N_36378,N_36385);
and U37972 (N_37972,N_36715,N_36910);
nor U37973 (N_37973,N_36685,N_36295);
xnor U37974 (N_37974,N_36733,N_36626);
and U37975 (N_37975,N_36269,N_36599);
or U37976 (N_37976,N_36874,N_36991);
nor U37977 (N_37977,N_36647,N_36907);
and U37978 (N_37978,N_36203,N_36702);
and U37979 (N_37979,N_36563,N_36756);
nand U37980 (N_37980,N_36059,N_36596);
xnor U37981 (N_37981,N_36471,N_36383);
nor U37982 (N_37982,N_36649,N_36123);
or U37983 (N_37983,N_36526,N_36778);
xnor U37984 (N_37984,N_36686,N_36937);
or U37985 (N_37985,N_36174,N_36507);
nand U37986 (N_37986,N_36049,N_36391);
nor U37987 (N_37987,N_36600,N_36215);
nand U37988 (N_37988,N_36526,N_36575);
and U37989 (N_37989,N_36180,N_36292);
nand U37990 (N_37990,N_36976,N_36175);
nor U37991 (N_37991,N_36363,N_36673);
xor U37992 (N_37992,N_36995,N_36038);
or U37993 (N_37993,N_36853,N_36972);
xor U37994 (N_37994,N_36276,N_36346);
and U37995 (N_37995,N_36790,N_36519);
or U37996 (N_37996,N_36100,N_36360);
and U37997 (N_37997,N_36794,N_36340);
nor U37998 (N_37998,N_36041,N_36413);
nand U37999 (N_37999,N_36139,N_36112);
or U38000 (N_38000,N_37495,N_37104);
nor U38001 (N_38001,N_37463,N_37434);
and U38002 (N_38002,N_37953,N_37524);
nor U38003 (N_38003,N_37343,N_37082);
xor U38004 (N_38004,N_37115,N_37590);
or U38005 (N_38005,N_37186,N_37476);
or U38006 (N_38006,N_37538,N_37973);
xor U38007 (N_38007,N_37628,N_37257);
and U38008 (N_38008,N_37983,N_37125);
nor U38009 (N_38009,N_37854,N_37484);
xnor U38010 (N_38010,N_37736,N_37711);
nor U38011 (N_38011,N_37169,N_37444);
xor U38012 (N_38012,N_37056,N_37540);
xnor U38013 (N_38013,N_37893,N_37837);
nor U38014 (N_38014,N_37282,N_37647);
nand U38015 (N_38015,N_37043,N_37634);
nor U38016 (N_38016,N_37829,N_37998);
xor U38017 (N_38017,N_37521,N_37702);
nor U38018 (N_38018,N_37431,N_37354);
nand U38019 (N_38019,N_37695,N_37742);
xor U38020 (N_38020,N_37892,N_37818);
or U38021 (N_38021,N_37767,N_37297);
or U38022 (N_38022,N_37166,N_37122);
nand U38023 (N_38023,N_37038,N_37578);
and U38024 (N_38024,N_37300,N_37630);
and U38025 (N_38025,N_37821,N_37008);
xor U38026 (N_38026,N_37205,N_37280);
and U38027 (N_38027,N_37743,N_37157);
or U38028 (N_38028,N_37775,N_37027);
xnor U38029 (N_38029,N_37888,N_37853);
xnor U38030 (N_38030,N_37366,N_37926);
and U38031 (N_38031,N_37648,N_37600);
nor U38032 (N_38032,N_37774,N_37065);
or U38033 (N_38033,N_37571,N_37371);
nor U38034 (N_38034,N_37701,N_37867);
or U38035 (N_38035,N_37505,N_37135);
nor U38036 (N_38036,N_37248,N_37241);
or U38037 (N_38037,N_37962,N_37093);
nand U38038 (N_38038,N_37996,N_37734);
nor U38039 (N_38039,N_37076,N_37078);
nand U38040 (N_38040,N_37069,N_37652);
nand U38041 (N_38041,N_37058,N_37003);
or U38042 (N_38042,N_37650,N_37506);
or U38043 (N_38043,N_37461,N_37771);
nor U38044 (N_38044,N_37547,N_37335);
nand U38045 (N_38045,N_37117,N_37311);
nand U38046 (N_38046,N_37869,N_37703);
nand U38047 (N_38047,N_37095,N_37288);
xnor U38048 (N_38048,N_37527,N_37929);
or U38049 (N_38049,N_37567,N_37331);
nor U38050 (N_38050,N_37856,N_37174);
and U38051 (N_38051,N_37201,N_37026);
or U38052 (N_38052,N_37320,N_37988);
and U38053 (N_38053,N_37964,N_37100);
and U38054 (N_38054,N_37295,N_37671);
nor U38055 (N_38055,N_37637,N_37274);
xor U38056 (N_38056,N_37194,N_37290);
xor U38057 (N_38057,N_37001,N_37945);
nor U38058 (N_38058,N_37429,N_37594);
and U38059 (N_38059,N_37522,N_37633);
nand U38060 (N_38060,N_37750,N_37807);
nand U38061 (N_38061,N_37979,N_37266);
or U38062 (N_38062,N_37519,N_37490);
or U38063 (N_38063,N_37155,N_37681);
and U38064 (N_38064,N_37817,N_37941);
nor U38065 (N_38065,N_37086,N_37209);
and U38066 (N_38066,N_37968,N_37468);
and U38067 (N_38067,N_37672,N_37876);
or U38068 (N_38068,N_37179,N_37757);
or U38069 (N_38069,N_37258,N_37810);
or U38070 (N_38070,N_37931,N_37077);
or U38071 (N_38071,N_37609,N_37044);
xnor U38072 (N_38072,N_37970,N_37760);
xor U38073 (N_38073,N_37314,N_37351);
xor U38074 (N_38074,N_37377,N_37855);
xor U38075 (N_38075,N_37756,N_37606);
or U38076 (N_38076,N_37824,N_37062);
nor U38077 (N_38077,N_37942,N_37251);
nand U38078 (N_38078,N_37339,N_37987);
nand U38079 (N_38079,N_37134,N_37891);
and U38080 (N_38080,N_37799,N_37961);
nor U38081 (N_38081,N_37577,N_37801);
xor U38082 (N_38082,N_37641,N_37114);
and U38083 (N_38083,N_37148,N_37747);
nor U38084 (N_38084,N_37032,N_37212);
or U38085 (N_38085,N_37328,N_37791);
and U38086 (N_38086,N_37697,N_37886);
nor U38087 (N_38087,N_37758,N_37414);
or U38088 (N_38088,N_37805,N_37327);
nand U38089 (N_38089,N_37809,N_37140);
and U38090 (N_38090,N_37399,N_37683);
or U38091 (N_38091,N_37502,N_37604);
nor U38092 (N_38092,N_37727,N_37948);
and U38093 (N_38093,N_37132,N_37237);
or U38094 (N_38094,N_37828,N_37441);
nand U38095 (N_38095,N_37080,N_37124);
xor U38096 (N_38096,N_37560,N_37548);
nand U38097 (N_38097,N_37191,N_37501);
nor U38098 (N_38098,N_37835,N_37638);
and U38099 (N_38099,N_37066,N_37773);
nor U38100 (N_38100,N_37706,N_37993);
and U38101 (N_38101,N_37507,N_37665);
nor U38102 (N_38102,N_37470,N_37811);
and U38103 (N_38103,N_37384,N_37875);
nand U38104 (N_38104,N_37025,N_37557);
xnor U38105 (N_38105,N_37798,N_37240);
nand U38106 (N_38106,N_37880,N_37160);
and U38107 (N_38107,N_37704,N_37222);
and U38108 (N_38108,N_37218,N_37050);
xor U38109 (N_38109,N_37733,N_37698);
nor U38110 (N_38110,N_37089,N_37190);
nor U38111 (N_38111,N_37659,N_37518);
or U38112 (N_38112,N_37284,N_37784);
and U38113 (N_38113,N_37656,N_37735);
or U38114 (N_38114,N_37489,N_37040);
nor U38115 (N_38115,N_37778,N_37270);
and U38116 (N_38116,N_37388,N_37060);
xnor U38117 (N_38117,N_37595,N_37553);
and U38118 (N_38118,N_37075,N_37419);
nor U38119 (N_38119,N_37843,N_37966);
nor U38120 (N_38120,N_37304,N_37716);
xor U38121 (N_38121,N_37833,N_37305);
xnor U38122 (N_38122,N_37903,N_37618);
xor U38123 (N_38123,N_37477,N_37667);
or U38124 (N_38124,N_37849,N_37107);
and U38125 (N_38125,N_37021,N_37316);
nand U38126 (N_38126,N_37513,N_37611);
and U38127 (N_38127,N_37857,N_37797);
nand U38128 (N_38128,N_37686,N_37421);
nor U38129 (N_38129,N_37183,N_37907);
or U38130 (N_38130,N_37460,N_37459);
xnor U38131 (N_38131,N_37199,N_37841);
and U38132 (N_38132,N_37550,N_37275);
nor U38133 (N_38133,N_37063,N_37203);
nor U38134 (N_38134,N_37916,N_37786);
xnor U38135 (N_38135,N_37789,N_37874);
and U38136 (N_38136,N_37464,N_37079);
xnor U38137 (N_38137,N_37769,N_37616);
nor U38138 (N_38138,N_37908,N_37448);
xnor U38139 (N_38139,N_37188,N_37914);
xnor U38140 (N_38140,N_37635,N_37109);
xor U38141 (N_38141,N_37765,N_37016);
nor U38142 (N_38142,N_37860,N_37227);
and U38143 (N_38143,N_37906,N_37899);
and U38144 (N_38144,N_37951,N_37674);
and U38145 (N_38145,N_37192,N_37121);
nor U38146 (N_38146,N_37369,N_37536);
nand U38147 (N_38147,N_37555,N_37272);
and U38148 (N_38148,N_37197,N_37673);
and U38149 (N_38149,N_37720,N_37868);
nor U38150 (N_38150,N_37059,N_37465);
xnor U38151 (N_38151,N_37048,N_37509);
nand U38152 (N_38152,N_37376,N_37110);
nand U38153 (N_38153,N_37726,N_37932);
and U38154 (N_38154,N_37622,N_37176);
nand U38155 (N_38155,N_37103,N_37232);
nor U38156 (N_38156,N_37885,N_37137);
and U38157 (N_38157,N_37276,N_37820);
nand U38158 (N_38158,N_37046,N_37310);
nand U38159 (N_38159,N_37710,N_37812);
or U38160 (N_38160,N_37426,N_37644);
xor U38161 (N_38161,N_37952,N_37020);
xor U38162 (N_38162,N_37009,N_37229);
nand U38163 (N_38163,N_37440,N_37823);
xor U38164 (N_38164,N_37034,N_37549);
nor U38165 (N_38165,N_37416,N_37233);
and U38166 (N_38166,N_37491,N_37091);
xnor U38167 (N_38167,N_37261,N_37442);
xor U38168 (N_38168,N_37541,N_37787);
or U38169 (N_38169,N_37989,N_37839);
nor U38170 (N_38170,N_37279,N_37204);
or U38171 (N_38171,N_37792,N_37569);
nand U38172 (N_38172,N_37564,N_37333);
nand U38173 (N_38173,N_37515,N_37688);
xnor U38174 (N_38174,N_37360,N_37613);
nand U38175 (N_38175,N_37684,N_37363);
xnor U38176 (N_38176,N_37106,N_37017);
nand U38177 (N_38177,N_37680,N_37958);
nor U38178 (N_38178,N_37643,N_37943);
or U38179 (N_38179,N_37269,N_37146);
and U38180 (N_38180,N_37921,N_37764);
xnor U38181 (N_38181,N_37127,N_37572);
xnor U38182 (N_38182,N_37693,N_37937);
and U38183 (N_38183,N_37249,N_37709);
nand U38184 (N_38184,N_37991,N_37894);
or U38185 (N_38185,N_37877,N_37895);
or U38186 (N_38186,N_37011,N_37031);
xnor U38187 (N_38187,N_37037,N_37239);
nand U38188 (N_38188,N_37386,N_37424);
xor U38189 (N_38189,N_37189,N_37412);
xor U38190 (N_38190,N_37859,N_37910);
nand U38191 (N_38191,N_37356,N_37761);
and U38192 (N_38192,N_37878,N_37030);
nand U38193 (N_38193,N_37568,N_37654);
xor U38194 (N_38194,N_37221,N_37623);
or U38195 (N_38195,N_37847,N_37319);
and U38196 (N_38196,N_37940,N_37512);
nand U38197 (N_38197,N_37340,N_37514);
nand U38198 (N_38198,N_37479,N_37969);
and U38199 (N_38199,N_37587,N_37170);
nand U38200 (N_38200,N_37579,N_37342);
and U38201 (N_38201,N_37938,N_37640);
or U38202 (N_38202,N_37023,N_37788);
nor U38203 (N_38203,N_37934,N_37108);
and U38204 (N_38204,N_37884,N_37840);
nor U38205 (N_38205,N_37748,N_37281);
xor U38206 (N_38206,N_37158,N_37803);
and U38207 (N_38207,N_37528,N_37483);
or U38208 (N_38208,N_37088,N_37129);
nor U38209 (N_38209,N_37959,N_37777);
nor U38210 (N_38210,N_37289,N_37375);
or U38211 (N_38211,N_37175,N_37359);
xor U38212 (N_38212,N_37168,N_37225);
and U38213 (N_38213,N_37430,N_37971);
nand U38214 (N_38214,N_37374,N_37024);
nor U38215 (N_38215,N_37466,N_37350);
nor U38216 (N_38216,N_37474,N_37585);
and U38217 (N_38217,N_37919,N_37586);
nand U38218 (N_38218,N_37144,N_37796);
nand U38219 (N_38219,N_37014,N_37167);
xor U38220 (N_38220,N_37309,N_37171);
nor U38221 (N_38221,N_37762,N_37415);
nor U38222 (N_38222,N_37262,N_37051);
or U38223 (N_38223,N_37398,N_37631);
xor U38224 (N_38224,N_37226,N_37214);
or U38225 (N_38225,N_37012,N_37722);
nor U38226 (N_38226,N_37111,N_37508);
or U38227 (N_38227,N_37882,N_37230);
and U38228 (N_38228,N_37180,N_37213);
nand U38229 (N_38229,N_37678,N_37890);
xnor U38230 (N_38230,N_37329,N_37341);
nor U38231 (N_38231,N_37531,N_37596);
or U38232 (N_38232,N_37403,N_37898);
and U38233 (N_38233,N_37482,N_37871);
nor U38234 (N_38234,N_37956,N_37944);
and U38235 (N_38235,N_37345,N_37763);
and U38236 (N_38236,N_37177,N_37128);
nand U38237 (N_38237,N_37662,N_37361);
nand U38238 (N_38238,N_37151,N_37348);
and U38239 (N_38239,N_37902,N_37713);
or U38240 (N_38240,N_37692,N_37670);
nand U38241 (N_38241,N_37954,N_37162);
nand U38242 (N_38242,N_37285,N_37957);
nand U38243 (N_38243,N_37315,N_37219);
nor U38244 (N_38244,N_37112,N_37367);
nand U38245 (N_38245,N_37783,N_37928);
and U38246 (N_38246,N_37487,N_37301);
xor U38247 (N_38247,N_37780,N_37696);
or U38248 (N_38248,N_37385,N_37287);
nor U38249 (N_38249,N_37486,N_37831);
nand U38250 (N_38250,N_37981,N_37980);
xnor U38251 (N_38251,N_37534,N_37738);
xnor U38252 (N_38252,N_37368,N_37049);
or U38253 (N_38253,N_37246,N_37752);
nand U38254 (N_38254,N_37588,N_37566);
nand U38255 (N_38255,N_37717,N_37516);
nand U38256 (N_38256,N_37299,N_37992);
and U38257 (N_38257,N_37323,N_37744);
nor U38258 (N_38258,N_37675,N_37277);
and U38259 (N_38259,N_37563,N_37617);
nor U38260 (N_38260,N_37267,N_37126);
xor U38261 (N_38261,N_37923,N_37715);
xnor U38262 (N_38262,N_37410,N_37498);
xor U38263 (N_38263,N_37172,N_37754);
and U38264 (N_38264,N_37325,N_37689);
xor U38265 (N_38265,N_37963,N_37532);
nor U38266 (N_38266,N_37317,N_37094);
nor U38267 (N_38267,N_37994,N_37409);
and U38268 (N_38268,N_37061,N_37161);
nor U38269 (N_38269,N_37592,N_37520);
or U38270 (N_38270,N_37887,N_37946);
nor U38271 (N_38271,N_37150,N_37456);
and U38272 (N_38272,N_37781,N_37278);
nor U38273 (N_38273,N_37790,N_37620);
xor U38274 (N_38274,N_37364,N_37755);
xnor U38275 (N_38275,N_37863,N_37447);
nor U38276 (N_38276,N_37446,N_37098);
or U38277 (N_38277,N_37917,N_37939);
xnor U38278 (N_38278,N_37215,N_37608);
nand U38279 (N_38279,N_37185,N_37985);
or U38280 (N_38280,N_37815,N_37362);
xnor U38281 (N_38281,N_37253,N_37308);
and U38282 (N_38282,N_37729,N_37925);
nor U38283 (N_38283,N_37220,N_37804);
xor U38284 (N_38284,N_37256,N_37208);
or U38285 (N_38285,N_37254,N_37453);
and U38286 (N_38286,N_37615,N_37223);
nor U38287 (N_38287,N_37268,N_37451);
and U38288 (N_38288,N_37480,N_37806);
nand U38289 (N_38289,N_37632,N_37605);
and U38290 (N_38290,N_37224,N_37390);
xnor U38291 (N_38291,N_37712,N_37200);
nor U38292 (N_38292,N_37420,N_37196);
xor U38293 (N_38293,N_37164,N_37723);
and U38294 (N_38294,N_37601,N_37552);
nand U38295 (N_38295,N_37437,N_37813);
and U38296 (N_38296,N_37039,N_37475);
xor U38297 (N_38297,N_37153,N_37533);
xor U38298 (N_38298,N_37574,N_37033);
nor U38299 (N_38299,N_37271,N_37131);
or U38300 (N_38300,N_37666,N_37646);
nor U38301 (N_38301,N_37101,N_37006);
nor U38302 (N_38302,N_37873,N_37092);
nor U38303 (N_38303,N_37458,N_37610);
or U38304 (N_38304,N_37858,N_37298);
and U38305 (N_38305,N_37142,N_37090);
nand U38306 (N_38306,N_37234,N_37235);
or U38307 (N_38307,N_37685,N_37379);
xor U38308 (N_38308,N_37583,N_37013);
nor U38309 (N_38309,N_37318,N_37313);
or U38310 (N_38310,N_37496,N_37064);
or U38311 (N_38311,N_37243,N_37344);
and U38312 (N_38312,N_37332,N_37005);
nor U38313 (N_38313,N_37478,N_37402);
and U38314 (N_38314,N_37669,N_37147);
or U38315 (N_38315,N_37417,N_37753);
and U38316 (N_38316,N_37370,N_37373);
and U38317 (N_38317,N_37488,N_37770);
and U38318 (N_38318,N_37772,N_37238);
xnor U38319 (N_38319,N_37614,N_37639);
or U38320 (N_38320,N_37494,N_37492);
and U38321 (N_38321,N_37544,N_37655);
and U38322 (N_38322,N_37292,N_37141);
and U38323 (N_38323,N_37768,N_37740);
xnor U38324 (N_38324,N_37349,N_37607);
xnor U38325 (N_38325,N_37982,N_37822);
and U38326 (N_38326,N_37250,N_37975);
or U38327 (N_38327,N_37156,N_37473);
nand U38328 (N_38328,N_37986,N_37010);
nor U38329 (N_38329,N_37102,N_37896);
xor U38330 (N_38330,N_37467,N_37739);
xnor U38331 (N_38331,N_37418,N_37759);
nor U38332 (N_38332,N_37751,N_37326);
nor U38333 (N_38333,N_37582,N_37904);
and U38334 (N_38334,N_37559,N_37015);
nor U38335 (N_38335,N_37439,N_37452);
and U38336 (N_38336,N_37499,N_37936);
nand U38337 (N_38337,N_37556,N_37182);
and U38338 (N_38338,N_37997,N_37035);
nor U38339 (N_38339,N_37422,N_37438);
nor U38340 (N_38340,N_37428,N_37526);
xor U38341 (N_38341,N_37842,N_37336);
and U38342 (N_38342,N_37372,N_37537);
or U38343 (N_38343,N_37028,N_37057);
nand U38344 (N_38344,N_37265,N_37661);
and U38345 (N_38345,N_37500,N_37252);
nor U38346 (N_38346,N_37865,N_37105);
nand U38347 (N_38347,N_37776,N_37511);
nand U38348 (N_38348,N_37668,N_37730);
xnor U38349 (N_38349,N_37658,N_37724);
xnor U38350 (N_38350,N_37136,N_37636);
nand U38351 (N_38351,N_37307,N_37503);
nand U38352 (N_38352,N_37004,N_37321);
xor U38353 (N_38353,N_37469,N_37990);
nand U38354 (N_38354,N_37068,N_37383);
and U38355 (N_38355,N_37927,N_37691);
nand U38356 (N_38356,N_37741,N_37955);
or U38357 (N_38357,N_37255,N_37879);
xnor U38358 (N_38358,N_37389,N_37913);
nor U38359 (N_38359,N_37423,N_37029);
nand U38360 (N_38360,N_37445,N_37497);
xnor U38361 (N_38361,N_37581,N_37664);
and U38362 (N_38362,N_37481,N_37154);
or U38363 (N_38363,N_37337,N_37974);
or U38364 (N_38364,N_37626,N_37380);
nor U38365 (N_38365,N_37401,N_37651);
and U38366 (N_38366,N_37085,N_37901);
nor U38367 (N_38367,N_37334,N_37603);
and U38368 (N_38368,N_37054,N_37976);
nand U38369 (N_38369,N_37306,N_37260);
nand U38370 (N_38370,N_37705,N_37999);
xor U38371 (N_38371,N_37145,N_37832);
or U38372 (N_38372,N_37679,N_37097);
nand U38373 (N_38373,N_37291,N_37960);
xor U38374 (N_38374,N_37216,N_37041);
nand U38375 (N_38375,N_37217,N_37800);
and U38376 (N_38376,N_37573,N_37677);
nand U38377 (N_38377,N_37909,N_37303);
xnor U38378 (N_38378,N_37852,N_37794);
and U38379 (N_38379,N_37766,N_37714);
xnor U38380 (N_38380,N_37845,N_37074);
nor U38381 (N_38381,N_37036,N_37396);
or U38382 (N_38382,N_37391,N_37346);
and U38383 (N_38383,N_37627,N_37814);
xor U38384 (N_38384,N_37259,N_37352);
nor U38385 (N_38385,N_37053,N_37357);
nand U38386 (N_38386,N_37707,N_37785);
and U38387 (N_38387,N_37198,N_37202);
and U38388 (N_38388,N_37413,N_37493);
nor U38389 (N_38389,N_37864,N_37393);
nand U38390 (N_38390,N_37067,N_37836);
or U38391 (N_38391,N_37378,N_37721);
nand U38392 (N_38392,N_37745,N_37206);
xor U38393 (N_38393,N_37118,N_37330);
xnor U38394 (N_38394,N_37851,N_37324);
nand U38395 (N_38395,N_37687,N_37457);
xnor U38396 (N_38396,N_37296,N_37073);
or U38397 (N_38397,N_37599,N_37558);
and U38398 (N_38398,N_37850,N_37455);
and U38399 (N_38399,N_37924,N_37407);
nand U38400 (N_38400,N_37642,N_37535);
or U38401 (N_38401,N_37302,N_37247);
nor U38402 (N_38402,N_37381,N_37264);
nor U38403 (N_38403,N_37338,N_37143);
nand U38404 (N_38404,N_37485,N_37159);
nand U38405 (N_38405,N_37542,N_37228);
xor U38406 (N_38406,N_37123,N_37793);
xor U38407 (N_38407,N_37621,N_37816);
nand U38408 (N_38408,N_37149,N_37554);
or U38409 (N_38409,N_37187,N_37072);
and U38410 (N_38410,N_37897,N_37052);
xnor U38411 (N_38411,N_37718,N_37645);
nor U38412 (N_38412,N_37565,N_37139);
or U38413 (N_38413,N_37242,N_37207);
or U38414 (N_38414,N_37195,N_37593);
nand U38415 (N_38415,N_37930,N_37427);
or U38416 (N_38416,N_37737,N_37676);
xnor U38417 (N_38417,N_37872,N_37462);
nor U38418 (N_38418,N_37995,N_37694);
xnor U38419 (N_38419,N_37912,N_37570);
and U38420 (N_38420,N_37649,N_37096);
nand U38421 (N_38421,N_37819,N_37070);
nor U38422 (N_38422,N_37984,N_37663);
nand U38423 (N_38423,N_37152,N_37408);
nor U38424 (N_38424,N_37165,N_37844);
nand U38425 (N_38425,N_37083,N_37263);
nor U38426 (N_38426,N_37825,N_37504);
and U38427 (N_38427,N_37947,N_37862);
nor U38428 (N_38428,N_37099,N_37530);
and U38429 (N_38429,N_37965,N_37353);
xor U38430 (N_38430,N_37400,N_37425);
nor U38431 (N_38431,N_37113,N_37950);
nand U38432 (N_38432,N_37087,N_37436);
or U38433 (N_38433,N_37795,N_37861);
xnor U38434 (N_38434,N_37978,N_37236);
and U38435 (N_38435,N_37231,N_37523);
xor U38436 (N_38436,N_37597,N_37081);
nor U38437 (N_38437,N_37883,N_37905);
xor U38438 (N_38438,N_37355,N_37731);
nand U38439 (N_38439,N_37808,N_37517);
nand U38440 (N_38440,N_37625,N_37245);
nor U38441 (N_38441,N_37286,N_37294);
and U38442 (N_38442,N_37866,N_37432);
and U38443 (N_38443,N_37071,N_37055);
xor U38444 (N_38444,N_37181,N_37629);
xor U38445 (N_38445,N_37347,N_37591);
nand U38446 (N_38446,N_37018,N_37967);
and U38447 (N_38447,N_37690,N_37312);
xor U38448 (N_38448,N_37454,N_37163);
xnor U38449 (N_38449,N_37404,N_37543);
or U38450 (N_38450,N_37283,N_37395);
or U38451 (N_38451,N_37700,N_37682);
nor U38452 (N_38452,N_37915,N_37660);
xor U38453 (N_38453,N_37719,N_37826);
nand U38454 (N_38454,N_37472,N_37173);
nand U38455 (N_38455,N_37619,N_37116);
xnor U38456 (N_38456,N_37598,N_37551);
or U38457 (N_38457,N_37133,N_37575);
xor U38458 (N_38458,N_37657,N_37387);
nand U38459 (N_38459,N_37562,N_37580);
xor U38460 (N_38460,N_37708,N_37602);
nand U38461 (N_38461,N_37920,N_37529);
xnor U38462 (N_38462,N_37244,N_37830);
nand U38463 (N_38463,N_37002,N_37870);
nor U38464 (N_38464,N_37435,N_37918);
and U38465 (N_38465,N_37119,N_37802);
xnor U38466 (N_38466,N_37977,N_37834);
xor U38467 (N_38467,N_37911,N_37848);
and U38468 (N_38468,N_37972,N_37405);
nand U38469 (N_38469,N_37546,N_37193);
nand U38470 (N_38470,N_37047,N_37443);
xor U38471 (N_38471,N_37732,N_37433);
nand U38472 (N_38472,N_37138,N_37782);
or U38473 (N_38473,N_37881,N_37900);
nand U38474 (N_38474,N_37545,N_37392);
nor U38475 (N_38475,N_37728,N_37725);
nor U38476 (N_38476,N_37406,N_37846);
and U38477 (N_38477,N_37949,N_37293);
xor U38478 (N_38478,N_37210,N_37365);
and U38479 (N_38479,N_37749,N_37576);
xor U38480 (N_38480,N_37019,N_37699);
nand U38481 (N_38481,N_37394,N_37022);
nand U38482 (N_38482,N_37007,N_37397);
nand U38483 (N_38483,N_37449,N_37184);
nand U38484 (N_38484,N_37612,N_37130);
nand U38485 (N_38485,N_37838,N_37624);
and U38486 (N_38486,N_37746,N_37889);
and U38487 (N_38487,N_37000,N_37084);
or U38488 (N_38488,N_37358,N_37045);
nor U38489 (N_38489,N_37653,N_37539);
xor U38490 (N_38490,N_37561,N_37933);
xor U38491 (N_38491,N_37922,N_37471);
xor U38492 (N_38492,N_37211,N_37510);
xor U38493 (N_38493,N_37450,N_37322);
and U38494 (N_38494,N_37827,N_37779);
and U38495 (N_38495,N_37584,N_37273);
nor U38496 (N_38496,N_37120,N_37042);
nand U38497 (N_38497,N_37178,N_37935);
nor U38498 (N_38498,N_37382,N_37411);
nor U38499 (N_38499,N_37589,N_37525);
nand U38500 (N_38500,N_37888,N_37587);
nand U38501 (N_38501,N_37199,N_37922);
nor U38502 (N_38502,N_37191,N_37100);
and U38503 (N_38503,N_37412,N_37536);
or U38504 (N_38504,N_37108,N_37419);
and U38505 (N_38505,N_37708,N_37576);
or U38506 (N_38506,N_37048,N_37798);
and U38507 (N_38507,N_37446,N_37865);
xnor U38508 (N_38508,N_37862,N_37533);
nand U38509 (N_38509,N_37708,N_37574);
nand U38510 (N_38510,N_37157,N_37718);
nand U38511 (N_38511,N_37714,N_37460);
and U38512 (N_38512,N_37972,N_37722);
nand U38513 (N_38513,N_37664,N_37485);
nor U38514 (N_38514,N_37699,N_37835);
nor U38515 (N_38515,N_37184,N_37540);
nor U38516 (N_38516,N_37496,N_37836);
and U38517 (N_38517,N_37561,N_37501);
and U38518 (N_38518,N_37639,N_37035);
and U38519 (N_38519,N_37087,N_37149);
and U38520 (N_38520,N_37134,N_37632);
xor U38521 (N_38521,N_37757,N_37719);
nand U38522 (N_38522,N_37261,N_37970);
and U38523 (N_38523,N_37039,N_37579);
nand U38524 (N_38524,N_37131,N_37507);
xnor U38525 (N_38525,N_37702,N_37302);
nor U38526 (N_38526,N_37612,N_37669);
nor U38527 (N_38527,N_37870,N_37126);
nor U38528 (N_38528,N_37055,N_37623);
nor U38529 (N_38529,N_37363,N_37231);
xnor U38530 (N_38530,N_37934,N_37601);
nor U38531 (N_38531,N_37990,N_37750);
nor U38532 (N_38532,N_37395,N_37972);
or U38533 (N_38533,N_37426,N_37813);
and U38534 (N_38534,N_37246,N_37748);
xor U38535 (N_38535,N_37768,N_37794);
nor U38536 (N_38536,N_37076,N_37880);
nor U38537 (N_38537,N_37568,N_37859);
and U38538 (N_38538,N_37867,N_37647);
xnor U38539 (N_38539,N_37744,N_37535);
nand U38540 (N_38540,N_37377,N_37210);
nor U38541 (N_38541,N_37280,N_37842);
xnor U38542 (N_38542,N_37113,N_37968);
and U38543 (N_38543,N_37603,N_37282);
nand U38544 (N_38544,N_37137,N_37593);
or U38545 (N_38545,N_37767,N_37084);
xnor U38546 (N_38546,N_37293,N_37157);
and U38547 (N_38547,N_37435,N_37980);
nand U38548 (N_38548,N_37601,N_37171);
and U38549 (N_38549,N_37976,N_37144);
nor U38550 (N_38550,N_37935,N_37363);
nor U38551 (N_38551,N_37255,N_37283);
xor U38552 (N_38552,N_37296,N_37316);
and U38553 (N_38553,N_37514,N_37695);
xor U38554 (N_38554,N_37108,N_37113);
xor U38555 (N_38555,N_37406,N_37788);
nor U38556 (N_38556,N_37982,N_37284);
nand U38557 (N_38557,N_37046,N_37123);
xor U38558 (N_38558,N_37134,N_37915);
and U38559 (N_38559,N_37423,N_37478);
nor U38560 (N_38560,N_37190,N_37260);
nand U38561 (N_38561,N_37815,N_37175);
nor U38562 (N_38562,N_37724,N_37628);
nor U38563 (N_38563,N_37487,N_37422);
or U38564 (N_38564,N_37509,N_37638);
xnor U38565 (N_38565,N_37680,N_37702);
xnor U38566 (N_38566,N_37924,N_37647);
and U38567 (N_38567,N_37652,N_37909);
xor U38568 (N_38568,N_37421,N_37953);
nand U38569 (N_38569,N_37739,N_37990);
or U38570 (N_38570,N_37081,N_37073);
nand U38571 (N_38571,N_37161,N_37029);
xor U38572 (N_38572,N_37324,N_37790);
nor U38573 (N_38573,N_37472,N_37859);
xnor U38574 (N_38574,N_37532,N_37985);
or U38575 (N_38575,N_37946,N_37496);
and U38576 (N_38576,N_37497,N_37087);
xor U38577 (N_38577,N_37710,N_37862);
or U38578 (N_38578,N_37197,N_37597);
xnor U38579 (N_38579,N_37410,N_37100);
nand U38580 (N_38580,N_37205,N_37513);
xnor U38581 (N_38581,N_37566,N_37754);
nand U38582 (N_38582,N_37031,N_37770);
nor U38583 (N_38583,N_37987,N_37985);
xnor U38584 (N_38584,N_37306,N_37171);
and U38585 (N_38585,N_37277,N_37093);
and U38586 (N_38586,N_37675,N_37136);
xor U38587 (N_38587,N_37671,N_37693);
nand U38588 (N_38588,N_37973,N_37052);
nor U38589 (N_38589,N_37283,N_37305);
nand U38590 (N_38590,N_37707,N_37253);
or U38591 (N_38591,N_37214,N_37229);
nand U38592 (N_38592,N_37606,N_37711);
nor U38593 (N_38593,N_37608,N_37338);
xor U38594 (N_38594,N_37434,N_37376);
nor U38595 (N_38595,N_37953,N_37121);
xnor U38596 (N_38596,N_37125,N_37654);
or U38597 (N_38597,N_37878,N_37520);
or U38598 (N_38598,N_37362,N_37822);
or U38599 (N_38599,N_37218,N_37610);
xor U38600 (N_38600,N_37762,N_37840);
xor U38601 (N_38601,N_37194,N_37996);
nor U38602 (N_38602,N_37129,N_37584);
nand U38603 (N_38603,N_37791,N_37560);
nand U38604 (N_38604,N_37818,N_37050);
or U38605 (N_38605,N_37984,N_37003);
or U38606 (N_38606,N_37785,N_37701);
nor U38607 (N_38607,N_37693,N_37769);
nor U38608 (N_38608,N_37893,N_37724);
xor U38609 (N_38609,N_37422,N_37102);
nor U38610 (N_38610,N_37717,N_37391);
nand U38611 (N_38611,N_37538,N_37599);
xnor U38612 (N_38612,N_37529,N_37383);
xor U38613 (N_38613,N_37349,N_37986);
or U38614 (N_38614,N_37850,N_37606);
and U38615 (N_38615,N_37275,N_37149);
xnor U38616 (N_38616,N_37736,N_37404);
nand U38617 (N_38617,N_37963,N_37698);
and U38618 (N_38618,N_37061,N_37792);
nand U38619 (N_38619,N_37005,N_37050);
nand U38620 (N_38620,N_37915,N_37796);
nor U38621 (N_38621,N_37233,N_37176);
or U38622 (N_38622,N_37746,N_37455);
nor U38623 (N_38623,N_37402,N_37045);
nor U38624 (N_38624,N_37425,N_37271);
and U38625 (N_38625,N_37111,N_37569);
or U38626 (N_38626,N_37698,N_37824);
nor U38627 (N_38627,N_37339,N_37050);
xor U38628 (N_38628,N_37737,N_37457);
or U38629 (N_38629,N_37640,N_37119);
nand U38630 (N_38630,N_37984,N_37956);
or U38631 (N_38631,N_37122,N_37727);
nand U38632 (N_38632,N_37144,N_37233);
and U38633 (N_38633,N_37348,N_37830);
xor U38634 (N_38634,N_37554,N_37689);
and U38635 (N_38635,N_37407,N_37829);
nor U38636 (N_38636,N_37367,N_37140);
xor U38637 (N_38637,N_37665,N_37383);
or U38638 (N_38638,N_37390,N_37534);
xor U38639 (N_38639,N_37416,N_37504);
xnor U38640 (N_38640,N_37034,N_37083);
nand U38641 (N_38641,N_37269,N_37740);
nand U38642 (N_38642,N_37723,N_37537);
xnor U38643 (N_38643,N_37260,N_37452);
nand U38644 (N_38644,N_37763,N_37084);
or U38645 (N_38645,N_37029,N_37020);
or U38646 (N_38646,N_37163,N_37254);
or U38647 (N_38647,N_37707,N_37971);
and U38648 (N_38648,N_37127,N_37032);
or U38649 (N_38649,N_37650,N_37723);
or U38650 (N_38650,N_37570,N_37596);
and U38651 (N_38651,N_37759,N_37826);
nor U38652 (N_38652,N_37665,N_37547);
nor U38653 (N_38653,N_37570,N_37948);
xnor U38654 (N_38654,N_37720,N_37554);
xor U38655 (N_38655,N_37423,N_37905);
nor U38656 (N_38656,N_37684,N_37024);
xor U38657 (N_38657,N_37679,N_37089);
xor U38658 (N_38658,N_37627,N_37576);
nor U38659 (N_38659,N_37531,N_37170);
nor U38660 (N_38660,N_37189,N_37449);
or U38661 (N_38661,N_37469,N_37485);
nand U38662 (N_38662,N_37904,N_37900);
and U38663 (N_38663,N_37452,N_37806);
nand U38664 (N_38664,N_37746,N_37901);
nor U38665 (N_38665,N_37609,N_37034);
nand U38666 (N_38666,N_37120,N_37936);
and U38667 (N_38667,N_37744,N_37950);
or U38668 (N_38668,N_37490,N_37105);
nand U38669 (N_38669,N_37092,N_37870);
xnor U38670 (N_38670,N_37725,N_37199);
xor U38671 (N_38671,N_37032,N_37439);
xnor U38672 (N_38672,N_37828,N_37115);
nand U38673 (N_38673,N_37529,N_37151);
or U38674 (N_38674,N_37701,N_37439);
nand U38675 (N_38675,N_37889,N_37552);
or U38676 (N_38676,N_37253,N_37714);
or U38677 (N_38677,N_37142,N_37566);
xnor U38678 (N_38678,N_37149,N_37560);
and U38679 (N_38679,N_37687,N_37679);
nor U38680 (N_38680,N_37830,N_37312);
and U38681 (N_38681,N_37570,N_37719);
nor U38682 (N_38682,N_37638,N_37483);
nor U38683 (N_38683,N_37698,N_37851);
xnor U38684 (N_38684,N_37012,N_37076);
or U38685 (N_38685,N_37385,N_37930);
xor U38686 (N_38686,N_37441,N_37990);
xnor U38687 (N_38687,N_37075,N_37743);
and U38688 (N_38688,N_37618,N_37142);
or U38689 (N_38689,N_37450,N_37287);
xor U38690 (N_38690,N_37551,N_37050);
and U38691 (N_38691,N_37184,N_37458);
nand U38692 (N_38692,N_37790,N_37049);
and U38693 (N_38693,N_37448,N_37005);
and U38694 (N_38694,N_37710,N_37228);
or U38695 (N_38695,N_37198,N_37500);
nand U38696 (N_38696,N_37681,N_37950);
xnor U38697 (N_38697,N_37435,N_37953);
nand U38698 (N_38698,N_37633,N_37517);
or U38699 (N_38699,N_37774,N_37941);
and U38700 (N_38700,N_37658,N_37756);
nand U38701 (N_38701,N_37765,N_37349);
nor U38702 (N_38702,N_37782,N_37612);
nand U38703 (N_38703,N_37284,N_37017);
or U38704 (N_38704,N_37686,N_37445);
nand U38705 (N_38705,N_37394,N_37348);
nor U38706 (N_38706,N_37519,N_37995);
nand U38707 (N_38707,N_37798,N_37843);
and U38708 (N_38708,N_37579,N_37818);
xor U38709 (N_38709,N_37149,N_37960);
xor U38710 (N_38710,N_37784,N_37235);
or U38711 (N_38711,N_37908,N_37403);
nor U38712 (N_38712,N_37550,N_37293);
nand U38713 (N_38713,N_37505,N_37079);
nor U38714 (N_38714,N_37791,N_37568);
or U38715 (N_38715,N_37511,N_37375);
nand U38716 (N_38716,N_37826,N_37754);
nor U38717 (N_38717,N_37002,N_37645);
nand U38718 (N_38718,N_37061,N_37408);
nor U38719 (N_38719,N_37993,N_37513);
nor U38720 (N_38720,N_37067,N_37944);
or U38721 (N_38721,N_37440,N_37867);
and U38722 (N_38722,N_37894,N_37036);
xnor U38723 (N_38723,N_37628,N_37871);
xor U38724 (N_38724,N_37285,N_37970);
xnor U38725 (N_38725,N_37970,N_37634);
and U38726 (N_38726,N_37073,N_37349);
xor U38727 (N_38727,N_37767,N_37485);
xor U38728 (N_38728,N_37216,N_37401);
nand U38729 (N_38729,N_37211,N_37927);
and U38730 (N_38730,N_37700,N_37699);
nand U38731 (N_38731,N_37796,N_37585);
and U38732 (N_38732,N_37442,N_37811);
xnor U38733 (N_38733,N_37228,N_37902);
or U38734 (N_38734,N_37213,N_37210);
nand U38735 (N_38735,N_37900,N_37739);
or U38736 (N_38736,N_37539,N_37832);
or U38737 (N_38737,N_37250,N_37598);
xor U38738 (N_38738,N_37534,N_37882);
or U38739 (N_38739,N_37077,N_37246);
xor U38740 (N_38740,N_37693,N_37217);
nor U38741 (N_38741,N_37084,N_37552);
xor U38742 (N_38742,N_37113,N_37461);
or U38743 (N_38743,N_37918,N_37500);
or U38744 (N_38744,N_37980,N_37921);
or U38745 (N_38745,N_37229,N_37949);
nor U38746 (N_38746,N_37512,N_37882);
and U38747 (N_38747,N_37179,N_37775);
and U38748 (N_38748,N_37682,N_37275);
and U38749 (N_38749,N_37614,N_37552);
nor U38750 (N_38750,N_37955,N_37353);
nand U38751 (N_38751,N_37652,N_37756);
or U38752 (N_38752,N_37689,N_37322);
or U38753 (N_38753,N_37241,N_37428);
and U38754 (N_38754,N_37136,N_37268);
xor U38755 (N_38755,N_37676,N_37144);
xor U38756 (N_38756,N_37183,N_37531);
nor U38757 (N_38757,N_37131,N_37035);
nor U38758 (N_38758,N_37938,N_37765);
or U38759 (N_38759,N_37925,N_37071);
nor U38760 (N_38760,N_37009,N_37496);
xor U38761 (N_38761,N_37927,N_37093);
or U38762 (N_38762,N_37943,N_37213);
nor U38763 (N_38763,N_37897,N_37833);
and U38764 (N_38764,N_37450,N_37412);
nor U38765 (N_38765,N_37063,N_37247);
and U38766 (N_38766,N_37496,N_37796);
nor U38767 (N_38767,N_37075,N_37323);
nand U38768 (N_38768,N_37851,N_37898);
xor U38769 (N_38769,N_37357,N_37305);
nand U38770 (N_38770,N_37794,N_37641);
nand U38771 (N_38771,N_37343,N_37809);
nor U38772 (N_38772,N_37558,N_37456);
and U38773 (N_38773,N_37195,N_37728);
or U38774 (N_38774,N_37489,N_37978);
nand U38775 (N_38775,N_37244,N_37577);
or U38776 (N_38776,N_37473,N_37484);
nor U38777 (N_38777,N_37188,N_37696);
nor U38778 (N_38778,N_37460,N_37803);
xnor U38779 (N_38779,N_37817,N_37847);
and U38780 (N_38780,N_37568,N_37854);
or U38781 (N_38781,N_37807,N_37595);
nand U38782 (N_38782,N_37132,N_37752);
or U38783 (N_38783,N_37547,N_37284);
or U38784 (N_38784,N_37852,N_37103);
or U38785 (N_38785,N_37564,N_37627);
and U38786 (N_38786,N_37520,N_37510);
nor U38787 (N_38787,N_37086,N_37220);
nor U38788 (N_38788,N_37243,N_37551);
nor U38789 (N_38789,N_37265,N_37392);
nor U38790 (N_38790,N_37243,N_37619);
nand U38791 (N_38791,N_37563,N_37933);
or U38792 (N_38792,N_37255,N_37396);
nand U38793 (N_38793,N_37494,N_37478);
xnor U38794 (N_38794,N_37663,N_37221);
nand U38795 (N_38795,N_37431,N_37629);
or U38796 (N_38796,N_37393,N_37581);
and U38797 (N_38797,N_37395,N_37917);
nor U38798 (N_38798,N_37641,N_37543);
nor U38799 (N_38799,N_37452,N_37082);
and U38800 (N_38800,N_37587,N_37333);
and U38801 (N_38801,N_37557,N_37510);
and U38802 (N_38802,N_37377,N_37378);
nand U38803 (N_38803,N_37940,N_37458);
or U38804 (N_38804,N_37536,N_37549);
and U38805 (N_38805,N_37843,N_37284);
or U38806 (N_38806,N_37876,N_37977);
and U38807 (N_38807,N_37852,N_37861);
nor U38808 (N_38808,N_37280,N_37485);
nand U38809 (N_38809,N_37106,N_37286);
or U38810 (N_38810,N_37289,N_37242);
nor U38811 (N_38811,N_37093,N_37611);
or U38812 (N_38812,N_37916,N_37249);
xnor U38813 (N_38813,N_37179,N_37140);
nand U38814 (N_38814,N_37890,N_37595);
nand U38815 (N_38815,N_37253,N_37898);
nand U38816 (N_38816,N_37520,N_37560);
or U38817 (N_38817,N_37228,N_37766);
or U38818 (N_38818,N_37564,N_37515);
nor U38819 (N_38819,N_37107,N_37388);
xnor U38820 (N_38820,N_37594,N_37347);
xor U38821 (N_38821,N_37511,N_37226);
and U38822 (N_38822,N_37101,N_37168);
xnor U38823 (N_38823,N_37656,N_37027);
or U38824 (N_38824,N_37520,N_37684);
and U38825 (N_38825,N_37475,N_37473);
nand U38826 (N_38826,N_37251,N_37990);
nor U38827 (N_38827,N_37730,N_37521);
and U38828 (N_38828,N_37668,N_37086);
and U38829 (N_38829,N_37265,N_37171);
nor U38830 (N_38830,N_37106,N_37207);
nor U38831 (N_38831,N_37140,N_37277);
nor U38832 (N_38832,N_37471,N_37397);
nand U38833 (N_38833,N_37981,N_37248);
and U38834 (N_38834,N_37368,N_37295);
xnor U38835 (N_38835,N_37552,N_37541);
and U38836 (N_38836,N_37791,N_37130);
xor U38837 (N_38837,N_37038,N_37948);
xnor U38838 (N_38838,N_37980,N_37730);
nand U38839 (N_38839,N_37592,N_37502);
or U38840 (N_38840,N_37664,N_37757);
nor U38841 (N_38841,N_37471,N_37432);
nor U38842 (N_38842,N_37266,N_37487);
and U38843 (N_38843,N_37794,N_37396);
or U38844 (N_38844,N_37604,N_37204);
xor U38845 (N_38845,N_37131,N_37296);
xor U38846 (N_38846,N_37945,N_37058);
nor U38847 (N_38847,N_37557,N_37632);
and U38848 (N_38848,N_37460,N_37978);
and U38849 (N_38849,N_37934,N_37212);
nor U38850 (N_38850,N_37299,N_37855);
nand U38851 (N_38851,N_37537,N_37789);
and U38852 (N_38852,N_37262,N_37384);
nor U38853 (N_38853,N_37605,N_37053);
nor U38854 (N_38854,N_37685,N_37914);
and U38855 (N_38855,N_37908,N_37606);
nor U38856 (N_38856,N_37755,N_37771);
and U38857 (N_38857,N_37288,N_37030);
xnor U38858 (N_38858,N_37846,N_37229);
nand U38859 (N_38859,N_37678,N_37422);
or U38860 (N_38860,N_37072,N_37985);
nor U38861 (N_38861,N_37096,N_37645);
xor U38862 (N_38862,N_37322,N_37015);
nor U38863 (N_38863,N_37042,N_37556);
nand U38864 (N_38864,N_37195,N_37604);
nor U38865 (N_38865,N_37927,N_37019);
and U38866 (N_38866,N_37048,N_37431);
and U38867 (N_38867,N_37743,N_37499);
or U38868 (N_38868,N_37528,N_37986);
and U38869 (N_38869,N_37708,N_37084);
nand U38870 (N_38870,N_37848,N_37166);
nand U38871 (N_38871,N_37820,N_37926);
xnor U38872 (N_38872,N_37661,N_37654);
xor U38873 (N_38873,N_37655,N_37921);
xnor U38874 (N_38874,N_37402,N_37454);
or U38875 (N_38875,N_37280,N_37239);
or U38876 (N_38876,N_37830,N_37089);
or U38877 (N_38877,N_37166,N_37463);
xor U38878 (N_38878,N_37836,N_37476);
nor U38879 (N_38879,N_37164,N_37632);
and U38880 (N_38880,N_37239,N_37873);
nor U38881 (N_38881,N_37077,N_37819);
nor U38882 (N_38882,N_37844,N_37628);
xnor U38883 (N_38883,N_37279,N_37269);
xor U38884 (N_38884,N_37099,N_37717);
xnor U38885 (N_38885,N_37138,N_37738);
nand U38886 (N_38886,N_37313,N_37194);
nor U38887 (N_38887,N_37969,N_37472);
nor U38888 (N_38888,N_37527,N_37932);
nor U38889 (N_38889,N_37281,N_37713);
nor U38890 (N_38890,N_37115,N_37336);
xor U38891 (N_38891,N_37111,N_37178);
or U38892 (N_38892,N_37609,N_37340);
and U38893 (N_38893,N_37443,N_37052);
and U38894 (N_38894,N_37184,N_37074);
nor U38895 (N_38895,N_37344,N_37829);
nor U38896 (N_38896,N_37092,N_37849);
nand U38897 (N_38897,N_37827,N_37286);
and U38898 (N_38898,N_37627,N_37504);
and U38899 (N_38899,N_37456,N_37292);
xor U38900 (N_38900,N_37953,N_37394);
and U38901 (N_38901,N_37652,N_37666);
nor U38902 (N_38902,N_37027,N_37142);
or U38903 (N_38903,N_37934,N_37545);
nand U38904 (N_38904,N_37753,N_37497);
and U38905 (N_38905,N_37572,N_37891);
nand U38906 (N_38906,N_37906,N_37380);
xnor U38907 (N_38907,N_37825,N_37191);
and U38908 (N_38908,N_37210,N_37181);
nor U38909 (N_38909,N_37053,N_37320);
nor U38910 (N_38910,N_37565,N_37267);
xnor U38911 (N_38911,N_37954,N_37690);
or U38912 (N_38912,N_37194,N_37023);
xor U38913 (N_38913,N_37317,N_37492);
and U38914 (N_38914,N_37758,N_37850);
xor U38915 (N_38915,N_37754,N_37852);
or U38916 (N_38916,N_37851,N_37789);
or U38917 (N_38917,N_37990,N_37406);
nand U38918 (N_38918,N_37431,N_37006);
nor U38919 (N_38919,N_37574,N_37749);
nor U38920 (N_38920,N_37076,N_37228);
nand U38921 (N_38921,N_37520,N_37069);
and U38922 (N_38922,N_37839,N_37999);
xnor U38923 (N_38923,N_37522,N_37259);
nand U38924 (N_38924,N_37040,N_37669);
and U38925 (N_38925,N_37416,N_37677);
and U38926 (N_38926,N_37612,N_37215);
xnor U38927 (N_38927,N_37885,N_37261);
xnor U38928 (N_38928,N_37099,N_37180);
nand U38929 (N_38929,N_37468,N_37540);
xnor U38930 (N_38930,N_37375,N_37791);
xnor U38931 (N_38931,N_37247,N_37679);
nor U38932 (N_38932,N_37035,N_37096);
xor U38933 (N_38933,N_37072,N_37977);
xor U38934 (N_38934,N_37020,N_37247);
and U38935 (N_38935,N_37420,N_37783);
or U38936 (N_38936,N_37444,N_37071);
xnor U38937 (N_38937,N_37155,N_37044);
or U38938 (N_38938,N_37518,N_37371);
xnor U38939 (N_38939,N_37567,N_37644);
xnor U38940 (N_38940,N_37209,N_37269);
nand U38941 (N_38941,N_37916,N_37920);
nor U38942 (N_38942,N_37910,N_37778);
xor U38943 (N_38943,N_37802,N_37126);
xor U38944 (N_38944,N_37236,N_37122);
and U38945 (N_38945,N_37449,N_37267);
or U38946 (N_38946,N_37476,N_37474);
or U38947 (N_38947,N_37584,N_37014);
and U38948 (N_38948,N_37706,N_37694);
nor U38949 (N_38949,N_37319,N_37489);
or U38950 (N_38950,N_37997,N_37430);
and U38951 (N_38951,N_37780,N_37945);
nor U38952 (N_38952,N_37107,N_37085);
nand U38953 (N_38953,N_37112,N_37182);
nor U38954 (N_38954,N_37315,N_37193);
nor U38955 (N_38955,N_37378,N_37922);
xor U38956 (N_38956,N_37310,N_37143);
nand U38957 (N_38957,N_37857,N_37922);
nor U38958 (N_38958,N_37387,N_37627);
xor U38959 (N_38959,N_37199,N_37162);
and U38960 (N_38960,N_37818,N_37986);
and U38961 (N_38961,N_37520,N_37506);
nand U38962 (N_38962,N_37422,N_37483);
nand U38963 (N_38963,N_37186,N_37173);
and U38964 (N_38964,N_37064,N_37612);
and U38965 (N_38965,N_37227,N_37412);
and U38966 (N_38966,N_37738,N_37970);
xor U38967 (N_38967,N_37155,N_37371);
and U38968 (N_38968,N_37277,N_37453);
nand U38969 (N_38969,N_37627,N_37738);
xnor U38970 (N_38970,N_37670,N_37536);
nand U38971 (N_38971,N_37908,N_37248);
xor U38972 (N_38972,N_37695,N_37128);
nor U38973 (N_38973,N_37178,N_37755);
or U38974 (N_38974,N_37482,N_37810);
nor U38975 (N_38975,N_37408,N_37905);
nor U38976 (N_38976,N_37612,N_37027);
or U38977 (N_38977,N_37416,N_37115);
nand U38978 (N_38978,N_37139,N_37014);
nor U38979 (N_38979,N_37385,N_37836);
and U38980 (N_38980,N_37591,N_37498);
and U38981 (N_38981,N_37718,N_37858);
nor U38982 (N_38982,N_37608,N_37385);
and U38983 (N_38983,N_37485,N_37846);
xnor U38984 (N_38984,N_37981,N_37154);
or U38985 (N_38985,N_37871,N_37052);
or U38986 (N_38986,N_37942,N_37579);
nor U38987 (N_38987,N_37975,N_37093);
and U38988 (N_38988,N_37322,N_37036);
and U38989 (N_38989,N_37526,N_37577);
xnor U38990 (N_38990,N_37233,N_37951);
nand U38991 (N_38991,N_37732,N_37316);
and U38992 (N_38992,N_37988,N_37805);
xnor U38993 (N_38993,N_37439,N_37913);
or U38994 (N_38994,N_37635,N_37466);
or U38995 (N_38995,N_37373,N_37254);
and U38996 (N_38996,N_37182,N_37916);
xor U38997 (N_38997,N_37329,N_37902);
and U38998 (N_38998,N_37795,N_37676);
nand U38999 (N_38999,N_37264,N_37984);
nor U39000 (N_39000,N_38857,N_38284);
xor U39001 (N_39001,N_38256,N_38506);
and U39002 (N_39002,N_38898,N_38448);
or U39003 (N_39003,N_38627,N_38524);
or U39004 (N_39004,N_38858,N_38850);
nor U39005 (N_39005,N_38690,N_38433);
nor U39006 (N_39006,N_38855,N_38501);
nor U39007 (N_39007,N_38413,N_38702);
xnor U39008 (N_39008,N_38882,N_38359);
and U39009 (N_39009,N_38689,N_38464);
xnor U39010 (N_39010,N_38562,N_38207);
xor U39011 (N_39011,N_38128,N_38036);
or U39012 (N_39012,N_38814,N_38537);
nand U39013 (N_39013,N_38726,N_38912);
nand U39014 (N_39014,N_38680,N_38720);
nor U39015 (N_39015,N_38539,N_38233);
or U39016 (N_39016,N_38015,N_38333);
and U39017 (N_39017,N_38989,N_38826);
xor U39018 (N_39018,N_38823,N_38107);
nand U39019 (N_39019,N_38495,N_38148);
and U39020 (N_39020,N_38301,N_38065);
nand U39021 (N_39021,N_38336,N_38727);
xnor U39022 (N_39022,N_38124,N_38693);
xor U39023 (N_39023,N_38743,N_38371);
xnor U39024 (N_39024,N_38719,N_38566);
nand U39025 (N_39025,N_38410,N_38567);
and U39026 (N_39026,N_38018,N_38615);
nor U39027 (N_39027,N_38304,N_38637);
nor U39028 (N_39028,N_38430,N_38951);
or U39029 (N_39029,N_38210,N_38815);
xnor U39030 (N_39030,N_38253,N_38290);
xnor U39031 (N_39031,N_38466,N_38728);
xnor U39032 (N_39032,N_38902,N_38579);
nand U39033 (N_39033,N_38157,N_38473);
or U39034 (N_39034,N_38922,N_38964);
nand U39035 (N_39035,N_38249,N_38168);
nand U39036 (N_39036,N_38777,N_38972);
and U39037 (N_39037,N_38252,N_38362);
nand U39038 (N_39038,N_38664,N_38663);
nor U39039 (N_39039,N_38507,N_38668);
nor U39040 (N_39040,N_38365,N_38205);
nand U39041 (N_39041,N_38748,N_38717);
nor U39042 (N_39042,N_38041,N_38971);
nor U39043 (N_39043,N_38025,N_38799);
xnor U39044 (N_39044,N_38986,N_38551);
or U39045 (N_39045,N_38062,N_38797);
nand U39046 (N_39046,N_38741,N_38950);
nor U39047 (N_39047,N_38051,N_38153);
nand U39048 (N_39048,N_38774,N_38840);
and U39049 (N_39049,N_38395,N_38776);
nand U39050 (N_39050,N_38809,N_38924);
xnor U39051 (N_39051,N_38530,N_38127);
and U39052 (N_39052,N_38186,N_38274);
nor U39053 (N_39053,N_38242,N_38837);
and U39054 (N_39054,N_38665,N_38595);
and U39055 (N_39055,N_38251,N_38461);
xnor U39056 (N_39056,N_38164,N_38259);
nor U39057 (N_39057,N_38778,N_38600);
or U39058 (N_39058,N_38597,N_38588);
nor U39059 (N_39059,N_38869,N_38784);
xor U39060 (N_39060,N_38052,N_38240);
xor U39061 (N_39061,N_38174,N_38508);
nor U39062 (N_39062,N_38347,N_38111);
and U39063 (N_39063,N_38411,N_38047);
and U39064 (N_39064,N_38773,N_38278);
or U39065 (N_39065,N_38158,N_38675);
and U39066 (N_39066,N_38305,N_38628);
nor U39067 (N_39067,N_38403,N_38428);
xor U39068 (N_39068,N_38571,N_38548);
or U39069 (N_39069,N_38187,N_38752);
xnor U39070 (N_39070,N_38300,N_38463);
xor U39071 (N_39071,N_38522,N_38106);
nor U39072 (N_39072,N_38173,N_38180);
or U39073 (N_39073,N_38594,N_38800);
nand U39074 (N_39074,N_38004,N_38948);
xnor U39075 (N_39075,N_38575,N_38745);
xnor U39076 (N_39076,N_38344,N_38839);
nor U39077 (N_39077,N_38272,N_38149);
nor U39078 (N_39078,N_38311,N_38360);
and U39079 (N_39079,N_38293,N_38490);
and U39080 (N_39080,N_38959,N_38346);
nand U39081 (N_39081,N_38331,N_38974);
and U39082 (N_39082,N_38555,N_38457);
nand U39083 (N_39083,N_38434,N_38616);
and U39084 (N_39084,N_38150,N_38324);
xnor U39085 (N_39085,N_38481,N_38831);
or U39086 (N_39086,N_38611,N_38043);
nand U39087 (N_39087,N_38833,N_38913);
nor U39088 (N_39088,N_38527,N_38125);
xnor U39089 (N_39089,N_38298,N_38984);
and U39090 (N_39090,N_38236,N_38269);
nor U39091 (N_39091,N_38423,N_38746);
and U39092 (N_39092,N_38289,N_38165);
or U39093 (N_39093,N_38028,N_38443);
and U39094 (N_39094,N_38783,N_38294);
nor U39095 (N_39095,N_38729,N_38722);
or U39096 (N_39096,N_38063,N_38266);
nand U39097 (N_39097,N_38904,N_38055);
or U39098 (N_39098,N_38110,N_38868);
and U39099 (N_39099,N_38910,N_38667);
xnor U39100 (N_39100,N_38970,N_38985);
and U39101 (N_39101,N_38183,N_38112);
nor U39102 (N_39102,N_38909,N_38963);
and U39103 (N_39103,N_38515,N_38458);
nor U39104 (N_39104,N_38193,N_38644);
and U39105 (N_39105,N_38129,N_38085);
xnor U39106 (N_39106,N_38140,N_38343);
or U39107 (N_39107,N_38923,N_38864);
nand U39108 (N_39108,N_38711,N_38008);
xor U39109 (N_39109,N_38400,N_38966);
xnor U39110 (N_39110,N_38138,N_38132);
xnor U39111 (N_39111,N_38633,N_38231);
xor U39112 (N_39112,N_38647,N_38947);
nand U39113 (N_39113,N_38345,N_38209);
nand U39114 (N_39114,N_38027,N_38459);
or U39115 (N_39115,N_38396,N_38279);
nand U39116 (N_39116,N_38061,N_38334);
nor U39117 (N_39117,N_38834,N_38813);
nand U39118 (N_39118,N_38368,N_38906);
nand U39119 (N_39119,N_38011,N_38544);
and U39120 (N_39120,N_38988,N_38682);
or U39121 (N_39121,N_38021,N_38218);
or U39122 (N_39122,N_38216,N_38763);
nand U39123 (N_39123,N_38980,N_38885);
xor U39124 (N_39124,N_38176,N_38213);
nand U39125 (N_39125,N_38642,N_38603);
and U39126 (N_39126,N_38029,N_38019);
xnor U39127 (N_39127,N_38066,N_38824);
and U39128 (N_39128,N_38918,N_38446);
xor U39129 (N_39129,N_38387,N_38751);
nor U39130 (N_39130,N_38325,N_38709);
nand U39131 (N_39131,N_38679,N_38104);
nand U39132 (N_39132,N_38366,N_38756);
and U39133 (N_39133,N_38979,N_38535);
xnor U39134 (N_39134,N_38856,N_38944);
xor U39135 (N_39135,N_38648,N_38811);
or U39136 (N_39136,N_38312,N_38761);
nor U39137 (N_39137,N_38131,N_38354);
and U39138 (N_39138,N_38820,N_38478);
and U39139 (N_39139,N_38369,N_38907);
xor U39140 (N_39140,N_38017,N_38678);
or U39141 (N_39141,N_38872,N_38357);
and U39142 (N_39142,N_38851,N_38994);
nand U39143 (N_39143,N_38626,N_38178);
xnor U39144 (N_39144,N_38091,N_38757);
or U39145 (N_39145,N_38821,N_38375);
xor U39146 (N_39146,N_38327,N_38401);
nand U39147 (N_39147,N_38045,N_38666);
or U39148 (N_39148,N_38488,N_38861);
xnor U39149 (N_39149,N_38629,N_38276);
or U39150 (N_39150,N_38699,N_38672);
nand U39151 (N_39151,N_38441,N_38001);
nand U39152 (N_39152,N_38391,N_38044);
nor U39153 (N_39153,N_38114,N_38931);
nand U39154 (N_39154,N_38054,N_38356);
or U39155 (N_39155,N_38103,N_38084);
nor U39156 (N_39156,N_38342,N_38445);
xor U39157 (N_39157,N_38040,N_38545);
nor U39158 (N_39158,N_38380,N_38275);
nand U39159 (N_39159,N_38684,N_38568);
or U39160 (N_39160,N_38145,N_38559);
xor U39161 (N_39161,N_38058,N_38890);
xnor U39162 (N_39162,N_38283,N_38961);
and U39163 (N_39163,N_38878,N_38787);
nand U39164 (N_39164,N_38135,N_38093);
and U39165 (N_39165,N_38260,N_38639);
nor U39166 (N_39166,N_38137,N_38378);
nand U39167 (N_39167,N_38254,N_38020);
or U39168 (N_39168,N_38694,N_38035);
and U39169 (N_39169,N_38937,N_38432);
nor U39170 (N_39170,N_38598,N_38476);
xnor U39171 (N_39171,N_38353,N_38214);
nand U39172 (N_39172,N_38006,N_38073);
nor U39173 (N_39173,N_38884,N_38295);
nand U39174 (N_39174,N_38105,N_38247);
nor U39175 (N_39175,N_38431,N_38519);
nor U39176 (N_39176,N_38552,N_38442);
and U39177 (N_39177,N_38854,N_38953);
and U39178 (N_39178,N_38226,N_38744);
or U39179 (N_39179,N_38352,N_38115);
xor U39180 (N_39180,N_38730,N_38171);
or U39181 (N_39181,N_38541,N_38156);
nor U39182 (N_39182,N_38903,N_38339);
xnor U39183 (N_39183,N_38896,N_38083);
xnor U39184 (N_39184,N_38587,N_38087);
nand U39185 (N_39185,N_38755,N_38670);
xnor U39186 (N_39186,N_38829,N_38316);
and U39187 (N_39187,N_38271,N_38089);
or U39188 (N_39188,N_38143,N_38109);
nand U39189 (N_39189,N_38608,N_38724);
nor U39190 (N_39190,N_38853,N_38995);
and U39191 (N_39191,N_38886,N_38981);
or U39192 (N_39192,N_38546,N_38584);
xor U39193 (N_39193,N_38862,N_38622);
and U39194 (N_39194,N_38219,N_38323);
or U39195 (N_39195,N_38223,N_38934);
nand U39196 (N_39196,N_38418,N_38673);
xor U39197 (N_39197,N_38444,N_38160);
and U39198 (N_39198,N_38983,N_38077);
and U39199 (N_39199,N_38313,N_38451);
nor U39200 (N_39200,N_38492,N_38649);
nor U39201 (N_39201,N_38529,N_38350);
xor U39202 (N_39202,N_38830,N_38681);
nand U39203 (N_39203,N_38392,N_38452);
and U39204 (N_39204,N_38456,N_38847);
or U39205 (N_39205,N_38660,N_38580);
and U39206 (N_39206,N_38997,N_38657);
nor U39207 (N_39207,N_38303,N_38701);
nor U39208 (N_39208,N_38117,N_38737);
and U39209 (N_39209,N_38758,N_38068);
xor U39210 (N_39210,N_38919,N_38406);
nor U39211 (N_39211,N_38414,N_38499);
or U39212 (N_39212,N_38146,N_38037);
or U39213 (N_39213,N_38586,N_38536);
or U39214 (N_39214,N_38071,N_38638);
nor U39215 (N_39215,N_38599,N_38162);
and U39216 (N_39216,N_38547,N_38565);
or U39217 (N_39217,N_38725,N_38992);
or U39218 (N_39218,N_38532,N_38769);
and U39219 (N_39219,N_38263,N_38078);
xnor U39220 (N_39220,N_38705,N_38617);
xor U39221 (N_39221,N_38879,N_38894);
xnor U39222 (N_39222,N_38504,N_38754);
or U39223 (N_39223,N_38876,N_38874);
and U39224 (N_39224,N_38819,N_38142);
or U39225 (N_39225,N_38557,N_38941);
nor U39226 (N_39226,N_38685,N_38197);
and U39227 (N_39227,N_38234,N_38297);
and U39228 (N_39228,N_38321,N_38453);
nor U39229 (N_39229,N_38422,N_38687);
or U39230 (N_39230,N_38258,N_38123);
nand U39231 (N_39231,N_38202,N_38549);
nor U39232 (N_39232,N_38059,N_38677);
or U39233 (N_39233,N_38487,N_38465);
xnor U39234 (N_39234,N_38280,N_38623);
xor U39235 (N_39235,N_38184,N_38222);
or U39236 (N_39236,N_38635,N_38505);
nand U39237 (N_39237,N_38916,N_38917);
or U39238 (N_39238,N_38891,N_38945);
nand U39239 (N_39239,N_38538,N_38319);
or U39240 (N_39240,N_38521,N_38960);
xor U39241 (N_39241,N_38383,N_38326);
xor U39242 (N_39242,N_38097,N_38625);
xor U39243 (N_39243,N_38533,N_38585);
and U39244 (N_39244,N_38591,N_38791);
nand U39245 (N_39245,N_38224,N_38273);
or U39246 (N_39246,N_38513,N_38053);
nor U39247 (N_39247,N_38172,N_38577);
nor U39248 (N_39248,N_38139,N_38449);
nor U39249 (N_39249,N_38329,N_38578);
nand U39250 (N_39250,N_38261,N_38195);
nand U39251 (N_39251,N_38088,N_38060);
or U39252 (N_39252,N_38090,N_38812);
xnor U39253 (N_39253,N_38736,N_38572);
nor U39254 (N_39254,N_38967,N_38738);
or U39255 (N_39255,N_38512,N_38604);
and U39256 (N_39256,N_38016,N_38494);
and U39257 (N_39257,N_38363,N_38417);
or U39258 (N_39258,N_38624,N_38510);
nor U39259 (N_39259,N_38030,N_38696);
nor U39260 (N_39260,N_38228,N_38688);
nand U39261 (N_39261,N_38808,N_38296);
xor U39262 (N_39262,N_38436,N_38050);
xor U39263 (N_39263,N_38731,N_38718);
xor U39264 (N_39264,N_38899,N_38897);
and U39265 (N_39265,N_38621,N_38804);
and U39266 (N_39266,N_38697,N_38468);
nand U39267 (N_39267,N_38307,N_38762);
and U39268 (N_39268,N_38509,N_38338);
and U39269 (N_39269,N_38750,N_38159);
xor U39270 (N_39270,N_38390,N_38593);
and U39271 (N_39271,N_38583,N_38373);
nand U39272 (N_39272,N_38080,N_38141);
and U39273 (N_39273,N_38480,N_38686);
and U39274 (N_39274,N_38927,N_38789);
and U39275 (N_39275,N_38211,N_38482);
nand U39276 (N_39276,N_38070,N_38000);
nand U39277 (N_39277,N_38232,N_38935);
xor U39278 (N_39278,N_38038,N_38643);
nor U39279 (N_39279,N_38550,N_38101);
nand U39280 (N_39280,N_38257,N_38753);
nor U39281 (N_39281,N_38479,N_38939);
and U39282 (N_39282,N_38704,N_38601);
xnor U39283 (N_39283,N_38570,N_38563);
nor U39284 (N_39284,N_38713,N_38126);
or U39285 (N_39285,N_38901,N_38998);
and U39286 (N_39286,N_38841,N_38842);
and U39287 (N_39287,N_38188,N_38185);
nand U39288 (N_39288,N_38241,N_38798);
and U39289 (N_39289,N_38291,N_38810);
nor U39290 (N_39290,N_38166,N_38285);
or U39291 (N_39291,N_38636,N_38827);
or U39292 (N_39292,N_38523,N_38244);
or U39293 (N_39293,N_38759,N_38064);
nand U39294 (N_39294,N_38169,N_38493);
and U39295 (N_39295,N_38402,N_38511);
nor U39296 (N_39296,N_38721,N_38619);
nand U39297 (N_39297,N_38880,N_38946);
and U39298 (N_39298,N_38975,N_38613);
xnor U39299 (N_39299,N_38397,N_38322);
and U39300 (N_39300,N_38364,N_38845);
and U39301 (N_39301,N_38485,N_38100);
xor U39302 (N_39302,N_38255,N_38707);
and U39303 (N_39303,N_38194,N_38936);
and U39304 (N_39304,N_38558,N_38785);
xor U39305 (N_39305,N_38999,N_38034);
nor U39306 (N_39306,N_38330,N_38489);
nand U39307 (N_39307,N_38949,N_38265);
nor U39308 (N_39308,N_38940,N_38554);
nor U39309 (N_39309,N_38706,N_38656);
and U39310 (N_39310,N_38500,N_38267);
and U39311 (N_39311,N_38119,N_38952);
and U39312 (N_39312,N_38534,N_38454);
or U39313 (N_39313,N_38264,N_38175);
or U39314 (N_39314,N_38978,N_38590);
xor U39315 (N_39315,N_38695,N_38920);
or U39316 (N_39316,N_38698,N_38426);
nor U39317 (N_39317,N_38314,N_38517);
or U39318 (N_39318,N_38419,N_38317);
nand U39319 (N_39319,N_38735,N_38531);
nand U39320 (N_39320,N_38199,N_38747);
nor U39321 (N_39321,N_38450,N_38046);
or U39322 (N_39322,N_38032,N_38859);
xor U39323 (N_39323,N_38661,N_38404);
and U39324 (N_39324,N_38116,N_38246);
and U39325 (N_39325,N_38474,N_38092);
nand U39326 (N_39326,N_38801,N_38370);
xor U39327 (N_39327,N_38388,N_38467);
nor U39328 (N_39328,N_38438,N_38320);
nor U39329 (N_39329,N_38455,N_38781);
nor U39330 (N_39330,N_38074,N_38009);
and U39331 (N_39331,N_38268,N_38144);
nor U39332 (N_39332,N_38096,N_38873);
and U39333 (N_39333,N_38348,N_38581);
xor U39334 (N_39334,N_38155,N_38662);
or U39335 (N_39335,N_38650,N_38973);
xnor U39336 (N_39336,N_38926,N_38425);
nor U39337 (N_39337,N_38807,N_38190);
nor U39338 (N_39338,N_38120,N_38732);
or U39339 (N_39339,N_38805,N_38760);
nor U39340 (N_39340,N_38292,N_38640);
nand U39341 (N_39341,N_38560,N_38405);
nor U39342 (N_39342,N_38113,N_38990);
nand U39343 (N_39343,N_38655,N_38318);
nand U39344 (N_39344,N_38932,N_38250);
xnor U39345 (N_39345,N_38710,N_38607);
nand U39346 (N_39346,N_38817,N_38023);
nor U39347 (N_39347,N_38871,N_38056);
or U39348 (N_39348,N_38130,N_38075);
nand U39349 (N_39349,N_38733,N_38900);
or U39350 (N_39350,N_38408,N_38957);
and U39351 (N_39351,N_38716,N_38203);
nand U39352 (N_39352,N_38239,N_38968);
xor U39353 (N_39353,N_38281,N_38768);
or U39354 (N_39354,N_38039,N_38770);
xor U39355 (N_39355,N_38620,N_38102);
nand U39356 (N_39356,N_38612,N_38852);
nand U39357 (N_39357,N_38514,N_38086);
and U39358 (N_39358,N_38229,N_38288);
nor U39359 (N_39359,N_38543,N_38602);
or U39360 (N_39360,N_38277,N_38520);
xor U39361 (N_39361,N_38793,N_38208);
xor U39362 (N_39362,N_38377,N_38714);
and U39363 (N_39363,N_38179,N_38381);
and U39364 (N_39364,N_38379,N_38382);
xnor U39365 (N_39365,N_38605,N_38469);
and U39366 (N_39366,N_38440,N_38386);
nor U39367 (N_39367,N_38631,N_38632);
nand U39368 (N_39368,N_38867,N_38098);
nor U39369 (N_39369,N_38969,N_38502);
nand U39370 (N_39370,N_38385,N_38189);
xnor U39371 (N_39371,N_38669,N_38384);
or U39372 (N_39372,N_38671,N_38589);
nand U39373 (N_39373,N_38518,N_38372);
nand U39374 (N_39374,N_38715,N_38042);
xnor U39375 (N_39375,N_38230,N_38484);
xor U39376 (N_39376,N_38421,N_38031);
and U39377 (N_39377,N_38933,N_38439);
xor U39378 (N_39378,N_38033,N_38561);
xnor U39379 (N_39379,N_38866,N_38865);
nand U39380 (N_39380,N_38956,N_38081);
xor U39381 (N_39381,N_38965,N_38227);
nor U39382 (N_39382,N_38911,N_38407);
nor U39383 (N_39383,N_38993,N_38739);
or U39384 (N_39384,N_38832,N_38200);
or U39385 (N_39385,N_38659,N_38248);
nand U39386 (N_39386,N_38844,N_38691);
and U39387 (N_39387,N_38245,N_38014);
or U39388 (N_39388,N_38788,N_38201);
and U39389 (N_39389,N_38958,N_38977);
xor U39390 (N_39390,N_38991,N_38412);
nand U39391 (N_39391,N_38122,N_38883);
or U39392 (N_39392,N_38795,N_38152);
nand U39393 (N_39393,N_38309,N_38121);
and U39394 (N_39394,N_38340,N_38892);
xnor U39395 (N_39395,N_38460,N_38516);
and U39396 (N_39396,N_38641,N_38740);
xor U39397 (N_39397,N_38816,N_38618);
nand U39398 (N_39398,N_38349,N_38217);
or U39399 (N_39399,N_38930,N_38361);
xnor U39400 (N_39400,N_38206,N_38002);
nand U39401 (N_39401,N_38818,N_38024);
nor U39402 (N_39402,N_38393,N_38887);
or U39403 (N_39403,N_38026,N_38496);
xor U39404 (N_39404,N_38712,N_38299);
or U39405 (N_39405,N_38302,N_38836);
or U39406 (N_39406,N_38204,N_38792);
and U39407 (N_39407,N_38653,N_38308);
nand U39408 (N_39408,N_38161,N_38221);
or U39409 (N_39409,N_38182,N_38556);
nor U39410 (N_39410,N_38574,N_38838);
nor U39411 (N_39411,N_38674,N_38399);
nand U39412 (N_39412,N_38196,N_38938);
nand U39413 (N_39413,N_38914,N_38651);
nor U39414 (N_39414,N_38849,N_38332);
nor U39415 (N_39415,N_38012,N_38877);
and U39416 (N_39416,N_38287,N_38215);
nand U39417 (N_39417,N_38306,N_38095);
nor U39418 (N_39418,N_38905,N_38954);
or U39419 (N_39419,N_38134,N_38424);
nor U39420 (N_39420,N_38630,N_38048);
nor U39421 (N_39421,N_38634,N_38067);
nor U39422 (N_39422,N_38177,N_38863);
xnor U39423 (N_39423,N_38592,N_38700);
nor U39424 (N_39424,N_38526,N_38429);
or U39425 (N_39425,N_38825,N_38163);
or U39426 (N_39426,N_38010,N_38237);
and U39427 (N_39427,N_38553,N_38708);
xnor U39428 (N_39428,N_38596,N_38835);
or U39429 (N_39429,N_38420,N_38497);
nor U39430 (N_39430,N_38328,N_38462);
and U39431 (N_39431,N_38881,N_38133);
or U39432 (N_39432,N_38437,N_38427);
xnor U39433 (N_39433,N_38243,N_38848);
and U39434 (N_39434,N_38767,N_38270);
and U39435 (N_39435,N_38471,N_38374);
or U39436 (N_39436,N_38335,N_38394);
nand U39437 (N_39437,N_38703,N_38491);
xor U39438 (N_39438,N_38398,N_38079);
or U39439 (N_39439,N_38573,N_38483);
and U39440 (N_39440,N_38569,N_38094);
nand U39441 (N_39441,N_38470,N_38921);
xnor U39442 (N_39442,N_38108,N_38780);
nor U39443 (N_39443,N_38582,N_38003);
and U39444 (N_39444,N_38775,N_38154);
xor U39445 (N_39445,N_38435,N_38606);
nor U39446 (N_39446,N_38337,N_38225);
and U39447 (N_39447,N_38654,N_38962);
or U39448 (N_39448,N_38007,N_38022);
or U39449 (N_39449,N_38477,N_38472);
nand U39450 (N_39450,N_38238,N_38942);
nand U39451 (N_39451,N_38542,N_38235);
and U39452 (N_39452,N_38782,N_38118);
nand U39453 (N_39453,N_38151,N_38610);
nand U39454 (N_39454,N_38525,N_38915);
and U39455 (N_39455,N_38692,N_38310);
or U39456 (N_39456,N_38895,N_38136);
xnor U39457 (N_39457,N_38765,N_38987);
nor U39458 (N_39458,N_38846,N_38982);
or U39459 (N_39459,N_38191,N_38220);
or U39460 (N_39460,N_38282,N_38658);
and U39461 (N_39461,N_38351,N_38786);
xor U39462 (N_39462,N_38723,N_38212);
or U39463 (N_39463,N_38341,N_38652);
and U39464 (N_39464,N_38315,N_38614);
nor U39465 (N_39465,N_38528,N_38828);
or U39466 (N_39466,N_38076,N_38875);
and U39467 (N_39467,N_38072,N_38893);
and U39468 (N_39468,N_38779,N_38996);
nor U39469 (N_39469,N_38734,N_38181);
or U39470 (N_39470,N_38005,N_38955);
nor U39471 (N_39471,N_38749,N_38908);
or U39472 (N_39472,N_38192,N_38771);
or U39473 (N_39473,N_38376,N_38928);
and U39474 (N_39474,N_38794,N_38475);
xor U39475 (N_39475,N_38069,N_38286);
nand U39476 (N_39476,N_38415,N_38355);
or U39477 (N_39477,N_38576,N_38943);
nor U39478 (N_39478,N_38764,N_38645);
and U39479 (N_39479,N_38486,N_38262);
nor U39480 (N_39480,N_38147,N_38806);
nand U39481 (N_39481,N_38057,N_38683);
nor U39482 (N_39482,N_38447,N_38802);
xor U39483 (N_39483,N_38367,N_38822);
nor U39484 (N_39484,N_38860,N_38540);
and U39485 (N_39485,N_38198,N_38925);
nor U39486 (N_39486,N_38389,N_38564);
nand U39487 (N_39487,N_38870,N_38013);
nor U39488 (N_39488,N_38888,N_38498);
nor U39489 (N_39489,N_38929,N_38889);
xnor U39490 (N_39490,N_38976,N_38766);
nand U39491 (N_39491,N_38790,N_38803);
nor U39492 (N_39492,N_38099,N_38742);
and U39493 (N_39493,N_38772,N_38676);
and U39494 (N_39494,N_38503,N_38049);
nor U39495 (N_39495,N_38843,N_38170);
nand U39496 (N_39496,N_38082,N_38646);
and U39497 (N_39497,N_38358,N_38409);
nor U39498 (N_39498,N_38416,N_38167);
xor U39499 (N_39499,N_38796,N_38609);
xnor U39500 (N_39500,N_38749,N_38776);
nand U39501 (N_39501,N_38823,N_38289);
or U39502 (N_39502,N_38709,N_38328);
xnor U39503 (N_39503,N_38914,N_38213);
or U39504 (N_39504,N_38532,N_38088);
xor U39505 (N_39505,N_38464,N_38275);
or U39506 (N_39506,N_38077,N_38620);
and U39507 (N_39507,N_38529,N_38647);
and U39508 (N_39508,N_38600,N_38373);
and U39509 (N_39509,N_38143,N_38898);
and U39510 (N_39510,N_38177,N_38820);
or U39511 (N_39511,N_38334,N_38479);
nand U39512 (N_39512,N_38259,N_38759);
nor U39513 (N_39513,N_38872,N_38938);
nand U39514 (N_39514,N_38409,N_38530);
nor U39515 (N_39515,N_38209,N_38776);
xnor U39516 (N_39516,N_38668,N_38895);
and U39517 (N_39517,N_38328,N_38746);
nand U39518 (N_39518,N_38868,N_38678);
nor U39519 (N_39519,N_38429,N_38676);
or U39520 (N_39520,N_38918,N_38275);
or U39521 (N_39521,N_38866,N_38354);
xnor U39522 (N_39522,N_38322,N_38187);
nand U39523 (N_39523,N_38263,N_38501);
xnor U39524 (N_39524,N_38495,N_38888);
and U39525 (N_39525,N_38977,N_38766);
or U39526 (N_39526,N_38568,N_38719);
xnor U39527 (N_39527,N_38127,N_38224);
xor U39528 (N_39528,N_38795,N_38642);
nand U39529 (N_39529,N_38346,N_38345);
and U39530 (N_39530,N_38817,N_38593);
xor U39531 (N_39531,N_38025,N_38337);
and U39532 (N_39532,N_38258,N_38516);
or U39533 (N_39533,N_38212,N_38206);
or U39534 (N_39534,N_38702,N_38226);
and U39535 (N_39535,N_38904,N_38736);
nand U39536 (N_39536,N_38816,N_38387);
xor U39537 (N_39537,N_38516,N_38422);
nand U39538 (N_39538,N_38635,N_38880);
or U39539 (N_39539,N_38762,N_38375);
or U39540 (N_39540,N_38425,N_38399);
xnor U39541 (N_39541,N_38095,N_38405);
nor U39542 (N_39542,N_38688,N_38997);
and U39543 (N_39543,N_38543,N_38231);
and U39544 (N_39544,N_38329,N_38958);
or U39545 (N_39545,N_38109,N_38535);
and U39546 (N_39546,N_38537,N_38354);
xor U39547 (N_39547,N_38116,N_38645);
nor U39548 (N_39548,N_38162,N_38832);
xor U39549 (N_39549,N_38479,N_38050);
xnor U39550 (N_39550,N_38427,N_38075);
nor U39551 (N_39551,N_38630,N_38121);
nand U39552 (N_39552,N_38288,N_38909);
or U39553 (N_39553,N_38650,N_38458);
nor U39554 (N_39554,N_38258,N_38141);
or U39555 (N_39555,N_38610,N_38617);
nor U39556 (N_39556,N_38853,N_38246);
nand U39557 (N_39557,N_38021,N_38427);
nor U39558 (N_39558,N_38247,N_38790);
nand U39559 (N_39559,N_38234,N_38993);
xnor U39560 (N_39560,N_38750,N_38731);
nand U39561 (N_39561,N_38245,N_38199);
nand U39562 (N_39562,N_38964,N_38677);
nand U39563 (N_39563,N_38963,N_38757);
or U39564 (N_39564,N_38329,N_38693);
nor U39565 (N_39565,N_38604,N_38232);
nand U39566 (N_39566,N_38958,N_38399);
nor U39567 (N_39567,N_38709,N_38014);
nor U39568 (N_39568,N_38182,N_38403);
and U39569 (N_39569,N_38256,N_38109);
nand U39570 (N_39570,N_38197,N_38395);
or U39571 (N_39571,N_38412,N_38933);
xnor U39572 (N_39572,N_38617,N_38633);
or U39573 (N_39573,N_38938,N_38028);
nand U39574 (N_39574,N_38817,N_38940);
and U39575 (N_39575,N_38960,N_38227);
and U39576 (N_39576,N_38163,N_38317);
or U39577 (N_39577,N_38642,N_38182);
or U39578 (N_39578,N_38087,N_38285);
and U39579 (N_39579,N_38603,N_38609);
xor U39580 (N_39580,N_38654,N_38714);
nand U39581 (N_39581,N_38736,N_38792);
and U39582 (N_39582,N_38409,N_38043);
xor U39583 (N_39583,N_38626,N_38897);
nor U39584 (N_39584,N_38572,N_38052);
and U39585 (N_39585,N_38148,N_38225);
or U39586 (N_39586,N_38070,N_38447);
xnor U39587 (N_39587,N_38815,N_38486);
nor U39588 (N_39588,N_38075,N_38720);
or U39589 (N_39589,N_38746,N_38181);
xor U39590 (N_39590,N_38085,N_38984);
nand U39591 (N_39591,N_38990,N_38777);
xnor U39592 (N_39592,N_38384,N_38970);
nor U39593 (N_39593,N_38461,N_38067);
nor U39594 (N_39594,N_38898,N_38696);
nand U39595 (N_39595,N_38984,N_38266);
xor U39596 (N_39596,N_38755,N_38675);
xnor U39597 (N_39597,N_38821,N_38824);
nand U39598 (N_39598,N_38668,N_38669);
or U39599 (N_39599,N_38733,N_38592);
and U39600 (N_39600,N_38573,N_38663);
and U39601 (N_39601,N_38051,N_38663);
nor U39602 (N_39602,N_38906,N_38009);
or U39603 (N_39603,N_38764,N_38941);
nor U39604 (N_39604,N_38945,N_38619);
nor U39605 (N_39605,N_38471,N_38992);
nand U39606 (N_39606,N_38983,N_38647);
or U39607 (N_39607,N_38318,N_38805);
xnor U39608 (N_39608,N_38127,N_38456);
nand U39609 (N_39609,N_38980,N_38547);
or U39610 (N_39610,N_38083,N_38513);
xnor U39611 (N_39611,N_38729,N_38706);
or U39612 (N_39612,N_38999,N_38286);
and U39613 (N_39613,N_38078,N_38265);
xor U39614 (N_39614,N_38205,N_38814);
and U39615 (N_39615,N_38623,N_38538);
and U39616 (N_39616,N_38361,N_38323);
xnor U39617 (N_39617,N_38492,N_38516);
or U39618 (N_39618,N_38034,N_38344);
or U39619 (N_39619,N_38613,N_38962);
xnor U39620 (N_39620,N_38265,N_38754);
xnor U39621 (N_39621,N_38015,N_38376);
xnor U39622 (N_39622,N_38347,N_38422);
nor U39623 (N_39623,N_38691,N_38943);
or U39624 (N_39624,N_38561,N_38657);
or U39625 (N_39625,N_38388,N_38762);
or U39626 (N_39626,N_38449,N_38458);
nor U39627 (N_39627,N_38642,N_38870);
and U39628 (N_39628,N_38028,N_38510);
nor U39629 (N_39629,N_38341,N_38886);
nor U39630 (N_39630,N_38028,N_38252);
and U39631 (N_39631,N_38325,N_38156);
nand U39632 (N_39632,N_38277,N_38941);
nor U39633 (N_39633,N_38301,N_38796);
nor U39634 (N_39634,N_38252,N_38191);
and U39635 (N_39635,N_38806,N_38117);
xnor U39636 (N_39636,N_38331,N_38335);
nor U39637 (N_39637,N_38937,N_38050);
xor U39638 (N_39638,N_38661,N_38129);
nand U39639 (N_39639,N_38387,N_38845);
nor U39640 (N_39640,N_38093,N_38463);
xor U39641 (N_39641,N_38254,N_38653);
nand U39642 (N_39642,N_38387,N_38940);
or U39643 (N_39643,N_38495,N_38648);
or U39644 (N_39644,N_38455,N_38665);
nand U39645 (N_39645,N_38166,N_38898);
and U39646 (N_39646,N_38447,N_38096);
xor U39647 (N_39647,N_38295,N_38226);
nand U39648 (N_39648,N_38432,N_38099);
nor U39649 (N_39649,N_38731,N_38413);
nor U39650 (N_39650,N_38966,N_38336);
or U39651 (N_39651,N_38545,N_38502);
and U39652 (N_39652,N_38964,N_38182);
nand U39653 (N_39653,N_38455,N_38200);
or U39654 (N_39654,N_38244,N_38867);
and U39655 (N_39655,N_38327,N_38599);
nor U39656 (N_39656,N_38795,N_38212);
xor U39657 (N_39657,N_38678,N_38217);
xnor U39658 (N_39658,N_38248,N_38736);
xnor U39659 (N_39659,N_38955,N_38313);
nor U39660 (N_39660,N_38640,N_38638);
or U39661 (N_39661,N_38273,N_38025);
nand U39662 (N_39662,N_38744,N_38208);
and U39663 (N_39663,N_38404,N_38431);
xnor U39664 (N_39664,N_38767,N_38578);
or U39665 (N_39665,N_38100,N_38812);
or U39666 (N_39666,N_38777,N_38911);
xor U39667 (N_39667,N_38213,N_38962);
nor U39668 (N_39668,N_38022,N_38922);
xor U39669 (N_39669,N_38434,N_38251);
and U39670 (N_39670,N_38020,N_38609);
and U39671 (N_39671,N_38928,N_38717);
and U39672 (N_39672,N_38095,N_38824);
nand U39673 (N_39673,N_38656,N_38333);
nor U39674 (N_39674,N_38134,N_38488);
nand U39675 (N_39675,N_38397,N_38806);
nor U39676 (N_39676,N_38839,N_38940);
and U39677 (N_39677,N_38480,N_38931);
nand U39678 (N_39678,N_38118,N_38131);
nor U39679 (N_39679,N_38478,N_38936);
or U39680 (N_39680,N_38065,N_38108);
and U39681 (N_39681,N_38750,N_38359);
or U39682 (N_39682,N_38920,N_38122);
and U39683 (N_39683,N_38631,N_38597);
and U39684 (N_39684,N_38688,N_38289);
or U39685 (N_39685,N_38198,N_38275);
or U39686 (N_39686,N_38130,N_38512);
and U39687 (N_39687,N_38955,N_38790);
and U39688 (N_39688,N_38796,N_38680);
xor U39689 (N_39689,N_38583,N_38356);
nand U39690 (N_39690,N_38922,N_38792);
nor U39691 (N_39691,N_38966,N_38551);
and U39692 (N_39692,N_38585,N_38406);
xnor U39693 (N_39693,N_38824,N_38515);
or U39694 (N_39694,N_38567,N_38523);
nand U39695 (N_39695,N_38011,N_38232);
or U39696 (N_39696,N_38496,N_38940);
or U39697 (N_39697,N_38157,N_38046);
and U39698 (N_39698,N_38770,N_38230);
and U39699 (N_39699,N_38324,N_38123);
or U39700 (N_39700,N_38308,N_38982);
xnor U39701 (N_39701,N_38350,N_38447);
nand U39702 (N_39702,N_38453,N_38733);
or U39703 (N_39703,N_38355,N_38942);
xnor U39704 (N_39704,N_38664,N_38969);
or U39705 (N_39705,N_38902,N_38132);
or U39706 (N_39706,N_38629,N_38191);
nor U39707 (N_39707,N_38691,N_38651);
nand U39708 (N_39708,N_38567,N_38915);
or U39709 (N_39709,N_38265,N_38613);
or U39710 (N_39710,N_38981,N_38608);
nand U39711 (N_39711,N_38619,N_38432);
or U39712 (N_39712,N_38825,N_38093);
nand U39713 (N_39713,N_38951,N_38274);
and U39714 (N_39714,N_38703,N_38531);
xor U39715 (N_39715,N_38246,N_38384);
nand U39716 (N_39716,N_38105,N_38303);
nor U39717 (N_39717,N_38417,N_38994);
xnor U39718 (N_39718,N_38806,N_38093);
xor U39719 (N_39719,N_38103,N_38718);
or U39720 (N_39720,N_38085,N_38661);
or U39721 (N_39721,N_38359,N_38981);
and U39722 (N_39722,N_38974,N_38719);
or U39723 (N_39723,N_38953,N_38496);
or U39724 (N_39724,N_38382,N_38606);
nand U39725 (N_39725,N_38588,N_38412);
nor U39726 (N_39726,N_38000,N_38801);
xnor U39727 (N_39727,N_38938,N_38615);
nand U39728 (N_39728,N_38115,N_38412);
nand U39729 (N_39729,N_38030,N_38245);
or U39730 (N_39730,N_38862,N_38972);
nand U39731 (N_39731,N_38181,N_38300);
nor U39732 (N_39732,N_38523,N_38593);
and U39733 (N_39733,N_38417,N_38582);
xnor U39734 (N_39734,N_38908,N_38148);
or U39735 (N_39735,N_38284,N_38937);
or U39736 (N_39736,N_38624,N_38507);
and U39737 (N_39737,N_38755,N_38194);
nor U39738 (N_39738,N_38776,N_38334);
nand U39739 (N_39739,N_38145,N_38324);
and U39740 (N_39740,N_38193,N_38937);
nand U39741 (N_39741,N_38162,N_38253);
nor U39742 (N_39742,N_38368,N_38218);
nor U39743 (N_39743,N_38671,N_38958);
and U39744 (N_39744,N_38141,N_38781);
xnor U39745 (N_39745,N_38821,N_38042);
or U39746 (N_39746,N_38420,N_38340);
nor U39747 (N_39747,N_38589,N_38501);
nor U39748 (N_39748,N_38727,N_38814);
and U39749 (N_39749,N_38645,N_38873);
or U39750 (N_39750,N_38245,N_38398);
and U39751 (N_39751,N_38178,N_38560);
and U39752 (N_39752,N_38509,N_38261);
nor U39753 (N_39753,N_38913,N_38385);
nand U39754 (N_39754,N_38768,N_38069);
xnor U39755 (N_39755,N_38751,N_38878);
and U39756 (N_39756,N_38830,N_38367);
and U39757 (N_39757,N_38081,N_38593);
and U39758 (N_39758,N_38648,N_38414);
nor U39759 (N_39759,N_38743,N_38117);
nand U39760 (N_39760,N_38345,N_38007);
nor U39761 (N_39761,N_38556,N_38545);
nor U39762 (N_39762,N_38053,N_38046);
xnor U39763 (N_39763,N_38292,N_38697);
nor U39764 (N_39764,N_38403,N_38378);
or U39765 (N_39765,N_38830,N_38725);
xnor U39766 (N_39766,N_38275,N_38932);
nor U39767 (N_39767,N_38757,N_38314);
nor U39768 (N_39768,N_38562,N_38761);
and U39769 (N_39769,N_38489,N_38074);
and U39770 (N_39770,N_38232,N_38308);
and U39771 (N_39771,N_38124,N_38736);
and U39772 (N_39772,N_38317,N_38655);
or U39773 (N_39773,N_38182,N_38727);
nand U39774 (N_39774,N_38724,N_38689);
xor U39775 (N_39775,N_38556,N_38637);
nor U39776 (N_39776,N_38367,N_38419);
or U39777 (N_39777,N_38920,N_38760);
xnor U39778 (N_39778,N_38263,N_38685);
or U39779 (N_39779,N_38098,N_38121);
nand U39780 (N_39780,N_38342,N_38333);
xnor U39781 (N_39781,N_38794,N_38034);
or U39782 (N_39782,N_38773,N_38625);
or U39783 (N_39783,N_38638,N_38423);
and U39784 (N_39784,N_38743,N_38780);
nor U39785 (N_39785,N_38595,N_38529);
xor U39786 (N_39786,N_38695,N_38369);
and U39787 (N_39787,N_38629,N_38409);
or U39788 (N_39788,N_38161,N_38756);
nand U39789 (N_39789,N_38632,N_38900);
nand U39790 (N_39790,N_38617,N_38605);
and U39791 (N_39791,N_38802,N_38973);
xnor U39792 (N_39792,N_38817,N_38445);
nor U39793 (N_39793,N_38825,N_38720);
nand U39794 (N_39794,N_38775,N_38963);
nand U39795 (N_39795,N_38614,N_38406);
nor U39796 (N_39796,N_38586,N_38249);
or U39797 (N_39797,N_38144,N_38081);
xnor U39798 (N_39798,N_38648,N_38598);
nor U39799 (N_39799,N_38106,N_38092);
nand U39800 (N_39800,N_38931,N_38637);
and U39801 (N_39801,N_38141,N_38481);
xor U39802 (N_39802,N_38894,N_38469);
nand U39803 (N_39803,N_38661,N_38508);
nand U39804 (N_39804,N_38524,N_38603);
or U39805 (N_39805,N_38084,N_38195);
nor U39806 (N_39806,N_38957,N_38575);
or U39807 (N_39807,N_38185,N_38405);
nor U39808 (N_39808,N_38535,N_38226);
nor U39809 (N_39809,N_38510,N_38776);
xnor U39810 (N_39810,N_38628,N_38085);
or U39811 (N_39811,N_38379,N_38371);
nand U39812 (N_39812,N_38125,N_38258);
and U39813 (N_39813,N_38913,N_38492);
and U39814 (N_39814,N_38188,N_38673);
or U39815 (N_39815,N_38401,N_38731);
and U39816 (N_39816,N_38338,N_38211);
and U39817 (N_39817,N_38813,N_38833);
or U39818 (N_39818,N_38155,N_38303);
nand U39819 (N_39819,N_38038,N_38841);
xor U39820 (N_39820,N_38761,N_38335);
nand U39821 (N_39821,N_38161,N_38344);
xor U39822 (N_39822,N_38711,N_38836);
or U39823 (N_39823,N_38222,N_38636);
nand U39824 (N_39824,N_38356,N_38125);
or U39825 (N_39825,N_38249,N_38606);
and U39826 (N_39826,N_38374,N_38817);
nor U39827 (N_39827,N_38304,N_38633);
nor U39828 (N_39828,N_38453,N_38107);
or U39829 (N_39829,N_38236,N_38313);
or U39830 (N_39830,N_38548,N_38516);
and U39831 (N_39831,N_38095,N_38609);
nand U39832 (N_39832,N_38280,N_38990);
nand U39833 (N_39833,N_38436,N_38313);
nor U39834 (N_39834,N_38700,N_38677);
or U39835 (N_39835,N_38177,N_38997);
xor U39836 (N_39836,N_38854,N_38947);
and U39837 (N_39837,N_38495,N_38714);
nand U39838 (N_39838,N_38077,N_38785);
xnor U39839 (N_39839,N_38003,N_38223);
nand U39840 (N_39840,N_38429,N_38021);
or U39841 (N_39841,N_38770,N_38155);
xnor U39842 (N_39842,N_38959,N_38451);
nand U39843 (N_39843,N_38426,N_38920);
xor U39844 (N_39844,N_38585,N_38617);
xor U39845 (N_39845,N_38980,N_38217);
xor U39846 (N_39846,N_38314,N_38587);
nand U39847 (N_39847,N_38118,N_38750);
xor U39848 (N_39848,N_38005,N_38597);
and U39849 (N_39849,N_38468,N_38182);
and U39850 (N_39850,N_38641,N_38247);
or U39851 (N_39851,N_38318,N_38018);
nand U39852 (N_39852,N_38041,N_38284);
nor U39853 (N_39853,N_38311,N_38683);
nand U39854 (N_39854,N_38719,N_38028);
xnor U39855 (N_39855,N_38564,N_38647);
nand U39856 (N_39856,N_38643,N_38554);
xor U39857 (N_39857,N_38139,N_38936);
and U39858 (N_39858,N_38461,N_38839);
nor U39859 (N_39859,N_38511,N_38852);
nand U39860 (N_39860,N_38234,N_38130);
or U39861 (N_39861,N_38740,N_38693);
xor U39862 (N_39862,N_38142,N_38042);
and U39863 (N_39863,N_38776,N_38408);
nor U39864 (N_39864,N_38844,N_38717);
nand U39865 (N_39865,N_38760,N_38665);
nand U39866 (N_39866,N_38820,N_38929);
nor U39867 (N_39867,N_38636,N_38249);
and U39868 (N_39868,N_38034,N_38427);
and U39869 (N_39869,N_38065,N_38124);
and U39870 (N_39870,N_38192,N_38785);
nand U39871 (N_39871,N_38810,N_38129);
nor U39872 (N_39872,N_38286,N_38024);
nor U39873 (N_39873,N_38870,N_38160);
nor U39874 (N_39874,N_38683,N_38205);
or U39875 (N_39875,N_38626,N_38973);
nand U39876 (N_39876,N_38110,N_38041);
nand U39877 (N_39877,N_38856,N_38980);
nor U39878 (N_39878,N_38061,N_38359);
or U39879 (N_39879,N_38667,N_38948);
xor U39880 (N_39880,N_38763,N_38936);
xnor U39881 (N_39881,N_38778,N_38299);
xnor U39882 (N_39882,N_38359,N_38139);
xor U39883 (N_39883,N_38809,N_38710);
nand U39884 (N_39884,N_38386,N_38979);
nor U39885 (N_39885,N_38360,N_38451);
and U39886 (N_39886,N_38122,N_38787);
xor U39887 (N_39887,N_38594,N_38698);
nand U39888 (N_39888,N_38471,N_38255);
xor U39889 (N_39889,N_38853,N_38474);
nand U39890 (N_39890,N_38899,N_38245);
nor U39891 (N_39891,N_38506,N_38788);
nand U39892 (N_39892,N_38918,N_38376);
or U39893 (N_39893,N_38045,N_38638);
nor U39894 (N_39894,N_38069,N_38231);
nand U39895 (N_39895,N_38748,N_38023);
or U39896 (N_39896,N_38384,N_38803);
and U39897 (N_39897,N_38089,N_38190);
or U39898 (N_39898,N_38502,N_38705);
or U39899 (N_39899,N_38808,N_38003);
nor U39900 (N_39900,N_38777,N_38914);
xnor U39901 (N_39901,N_38802,N_38711);
nand U39902 (N_39902,N_38208,N_38582);
nor U39903 (N_39903,N_38815,N_38042);
nor U39904 (N_39904,N_38253,N_38926);
nand U39905 (N_39905,N_38588,N_38141);
and U39906 (N_39906,N_38291,N_38911);
and U39907 (N_39907,N_38519,N_38467);
and U39908 (N_39908,N_38810,N_38247);
xor U39909 (N_39909,N_38595,N_38451);
nand U39910 (N_39910,N_38538,N_38910);
xor U39911 (N_39911,N_38867,N_38222);
xnor U39912 (N_39912,N_38238,N_38654);
and U39913 (N_39913,N_38859,N_38313);
xor U39914 (N_39914,N_38751,N_38896);
nor U39915 (N_39915,N_38549,N_38171);
nand U39916 (N_39916,N_38011,N_38893);
or U39917 (N_39917,N_38151,N_38788);
or U39918 (N_39918,N_38310,N_38902);
or U39919 (N_39919,N_38046,N_38147);
and U39920 (N_39920,N_38401,N_38776);
nor U39921 (N_39921,N_38549,N_38140);
nor U39922 (N_39922,N_38199,N_38614);
nor U39923 (N_39923,N_38706,N_38448);
nand U39924 (N_39924,N_38300,N_38304);
xnor U39925 (N_39925,N_38811,N_38934);
or U39926 (N_39926,N_38225,N_38607);
xnor U39927 (N_39927,N_38979,N_38744);
and U39928 (N_39928,N_38805,N_38710);
and U39929 (N_39929,N_38880,N_38553);
or U39930 (N_39930,N_38380,N_38794);
and U39931 (N_39931,N_38329,N_38038);
nor U39932 (N_39932,N_38822,N_38069);
nand U39933 (N_39933,N_38598,N_38779);
nand U39934 (N_39934,N_38031,N_38462);
nand U39935 (N_39935,N_38309,N_38803);
or U39936 (N_39936,N_38224,N_38415);
xor U39937 (N_39937,N_38029,N_38114);
nand U39938 (N_39938,N_38704,N_38205);
or U39939 (N_39939,N_38660,N_38270);
or U39940 (N_39940,N_38605,N_38989);
nand U39941 (N_39941,N_38827,N_38564);
xnor U39942 (N_39942,N_38853,N_38972);
nand U39943 (N_39943,N_38736,N_38669);
xor U39944 (N_39944,N_38588,N_38007);
nor U39945 (N_39945,N_38369,N_38730);
or U39946 (N_39946,N_38743,N_38059);
xor U39947 (N_39947,N_38920,N_38665);
nand U39948 (N_39948,N_38736,N_38309);
nand U39949 (N_39949,N_38785,N_38098);
or U39950 (N_39950,N_38595,N_38051);
nand U39951 (N_39951,N_38453,N_38241);
xor U39952 (N_39952,N_38016,N_38200);
or U39953 (N_39953,N_38213,N_38613);
and U39954 (N_39954,N_38196,N_38143);
and U39955 (N_39955,N_38123,N_38891);
or U39956 (N_39956,N_38645,N_38367);
or U39957 (N_39957,N_38068,N_38636);
and U39958 (N_39958,N_38875,N_38415);
nor U39959 (N_39959,N_38488,N_38430);
and U39960 (N_39960,N_38817,N_38904);
nand U39961 (N_39961,N_38515,N_38477);
nor U39962 (N_39962,N_38773,N_38499);
or U39963 (N_39963,N_38931,N_38482);
or U39964 (N_39964,N_38594,N_38021);
nand U39965 (N_39965,N_38801,N_38966);
or U39966 (N_39966,N_38335,N_38005);
nand U39967 (N_39967,N_38489,N_38213);
xnor U39968 (N_39968,N_38211,N_38523);
or U39969 (N_39969,N_38154,N_38361);
and U39970 (N_39970,N_38377,N_38129);
xor U39971 (N_39971,N_38969,N_38620);
nand U39972 (N_39972,N_38784,N_38711);
nor U39973 (N_39973,N_38054,N_38510);
and U39974 (N_39974,N_38150,N_38536);
nand U39975 (N_39975,N_38872,N_38934);
nor U39976 (N_39976,N_38914,N_38499);
and U39977 (N_39977,N_38421,N_38606);
or U39978 (N_39978,N_38704,N_38567);
nor U39979 (N_39979,N_38707,N_38581);
nor U39980 (N_39980,N_38837,N_38278);
nor U39981 (N_39981,N_38014,N_38029);
nor U39982 (N_39982,N_38351,N_38672);
or U39983 (N_39983,N_38161,N_38894);
xor U39984 (N_39984,N_38290,N_38324);
or U39985 (N_39985,N_38391,N_38257);
or U39986 (N_39986,N_38885,N_38557);
and U39987 (N_39987,N_38782,N_38870);
xor U39988 (N_39988,N_38198,N_38615);
nor U39989 (N_39989,N_38386,N_38391);
nand U39990 (N_39990,N_38498,N_38014);
xnor U39991 (N_39991,N_38561,N_38730);
xnor U39992 (N_39992,N_38746,N_38735);
or U39993 (N_39993,N_38789,N_38086);
or U39994 (N_39994,N_38334,N_38713);
or U39995 (N_39995,N_38308,N_38856);
and U39996 (N_39996,N_38556,N_38815);
xor U39997 (N_39997,N_38790,N_38650);
nand U39998 (N_39998,N_38360,N_38190);
nand U39999 (N_39999,N_38272,N_38936);
or U40000 (N_40000,N_39800,N_39369);
or U40001 (N_40001,N_39585,N_39043);
nor U40002 (N_40002,N_39162,N_39681);
nand U40003 (N_40003,N_39006,N_39498);
xnor U40004 (N_40004,N_39875,N_39699);
and U40005 (N_40005,N_39373,N_39047);
nand U40006 (N_40006,N_39330,N_39801);
xor U40007 (N_40007,N_39962,N_39327);
nand U40008 (N_40008,N_39821,N_39775);
xor U40009 (N_40009,N_39764,N_39956);
or U40010 (N_40010,N_39305,N_39634);
xnor U40011 (N_40011,N_39187,N_39514);
xnor U40012 (N_40012,N_39935,N_39156);
or U40013 (N_40013,N_39858,N_39131);
nand U40014 (N_40014,N_39721,N_39744);
xnor U40015 (N_40015,N_39667,N_39204);
nor U40016 (N_40016,N_39346,N_39135);
xnor U40017 (N_40017,N_39980,N_39575);
xnor U40018 (N_40018,N_39070,N_39948);
xor U40019 (N_40019,N_39524,N_39053);
xor U40020 (N_40020,N_39874,N_39146);
nand U40021 (N_40021,N_39640,N_39426);
nor U40022 (N_40022,N_39407,N_39519);
nand U40023 (N_40023,N_39415,N_39615);
nor U40024 (N_40024,N_39574,N_39352);
or U40025 (N_40025,N_39805,N_39753);
nand U40026 (N_40026,N_39291,N_39774);
nand U40027 (N_40027,N_39653,N_39378);
nand U40028 (N_40028,N_39724,N_39376);
nand U40029 (N_40029,N_39335,N_39927);
xor U40030 (N_40030,N_39032,N_39404);
nand U40031 (N_40031,N_39833,N_39629);
and U40032 (N_40032,N_39392,N_39234);
and U40033 (N_40033,N_39865,N_39123);
and U40034 (N_40034,N_39755,N_39087);
or U40035 (N_40035,N_39785,N_39528);
xor U40036 (N_40036,N_39590,N_39786);
xnor U40037 (N_40037,N_39567,N_39876);
nand U40038 (N_40038,N_39068,N_39175);
and U40039 (N_40039,N_39555,N_39861);
nor U40040 (N_40040,N_39757,N_39967);
nor U40041 (N_40041,N_39468,N_39516);
and U40042 (N_40042,N_39584,N_39160);
or U40043 (N_40043,N_39534,N_39961);
nand U40044 (N_40044,N_39414,N_39896);
or U40045 (N_40045,N_39826,N_39892);
nand U40046 (N_40046,N_39056,N_39224);
or U40047 (N_40047,N_39121,N_39023);
xor U40048 (N_40048,N_39010,N_39208);
and U40049 (N_40049,N_39400,N_39024);
and U40050 (N_40050,N_39088,N_39894);
nand U40051 (N_40051,N_39608,N_39676);
and U40052 (N_40052,N_39005,N_39211);
or U40053 (N_40053,N_39097,N_39069);
xor U40054 (N_40054,N_39958,N_39602);
nor U40055 (N_40055,N_39474,N_39030);
nand U40056 (N_40056,N_39491,N_39994);
and U40057 (N_40057,N_39003,N_39141);
or U40058 (N_40058,N_39500,N_39571);
nor U40059 (N_40059,N_39643,N_39758);
nand U40060 (N_40060,N_39132,N_39455);
xnor U40061 (N_40061,N_39192,N_39701);
xor U40062 (N_40062,N_39201,N_39067);
or U40063 (N_40063,N_39792,N_39260);
xor U40064 (N_40064,N_39209,N_39811);
xnor U40065 (N_40065,N_39720,N_39292);
or U40066 (N_40066,N_39521,N_39550);
and U40067 (N_40067,N_39014,N_39397);
and U40068 (N_40068,N_39173,N_39638);
or U40069 (N_40069,N_39463,N_39458);
or U40070 (N_40070,N_39381,N_39975);
and U40071 (N_40071,N_39679,N_39194);
nand U40072 (N_40072,N_39318,N_39706);
nor U40073 (N_40073,N_39154,N_39249);
nand U40074 (N_40074,N_39997,N_39625);
or U40075 (N_40075,N_39929,N_39022);
nor U40076 (N_40076,N_39839,N_39158);
nand U40077 (N_40077,N_39045,N_39347);
or U40078 (N_40078,N_39092,N_39512);
nand U40079 (N_40079,N_39081,N_39624);
and U40080 (N_40080,N_39112,N_39509);
and U40081 (N_40081,N_39915,N_39423);
or U40082 (N_40082,N_39960,N_39762);
or U40083 (N_40083,N_39340,N_39589);
nor U40084 (N_40084,N_39662,N_39663);
nand U40085 (N_40085,N_39227,N_39303);
and U40086 (N_40086,N_39499,N_39237);
nor U40087 (N_40087,N_39829,N_39502);
xor U40088 (N_40088,N_39274,N_39835);
and U40089 (N_40089,N_39287,N_39845);
xnor U40090 (N_40090,N_39772,N_39421);
or U40091 (N_40091,N_39887,N_39220);
nor U40092 (N_40092,N_39408,N_39425);
xnor U40093 (N_40093,N_39036,N_39661);
nor U40094 (N_40094,N_39333,N_39686);
and U40095 (N_40095,N_39129,N_39636);
nand U40096 (N_40096,N_39705,N_39825);
and U40097 (N_40097,N_39177,N_39137);
xor U40098 (N_40098,N_39280,N_39579);
and U40099 (N_40099,N_39497,N_39779);
nor U40100 (N_40100,N_39905,N_39196);
and U40101 (N_40101,N_39122,N_39647);
and U40102 (N_40102,N_39749,N_39941);
or U40103 (N_40103,N_39649,N_39691);
nor U40104 (N_40104,N_39612,N_39072);
or U40105 (N_40105,N_39853,N_39596);
nor U40106 (N_40106,N_39264,N_39044);
nor U40107 (N_40107,N_39664,N_39322);
xnor U40108 (N_40108,N_39405,N_39385);
xor U40109 (N_40109,N_39880,N_39374);
and U40110 (N_40110,N_39645,N_39553);
xor U40111 (N_40111,N_39102,N_39111);
xor U40112 (N_40112,N_39738,N_39592);
nand U40113 (N_40113,N_39242,N_39711);
nand U40114 (N_40114,N_39936,N_39859);
and U40115 (N_40115,N_39100,N_39058);
or U40116 (N_40116,N_39171,N_39221);
xor U40117 (N_40117,N_39362,N_39660);
and U40118 (N_40118,N_39933,N_39505);
and U40119 (N_40119,N_39120,N_39963);
nor U40120 (N_40120,N_39441,N_39708);
nor U40121 (N_40121,N_39114,N_39422);
xnor U40122 (N_40122,N_39968,N_39506);
nand U40123 (N_40123,N_39940,N_39982);
xnor U40124 (N_40124,N_39304,N_39763);
or U40125 (N_40125,N_39059,N_39034);
nand U40126 (N_40126,N_39259,N_39899);
or U40127 (N_40127,N_39680,N_39478);
nor U40128 (N_40128,N_39213,N_39206);
or U40129 (N_40129,N_39957,N_39804);
nor U40130 (N_40130,N_39168,N_39730);
xor U40131 (N_40131,N_39411,N_39151);
xor U40132 (N_40132,N_39586,N_39665);
nor U40133 (N_40133,N_39626,N_39153);
xnor U40134 (N_40134,N_39257,N_39564);
nand U40135 (N_40135,N_39906,N_39911);
or U40136 (N_40136,N_39517,N_39678);
xnor U40137 (N_40137,N_39566,N_39191);
nand U40138 (N_40138,N_39312,N_39394);
or U40139 (N_40139,N_39148,N_39820);
nand U40140 (N_40140,N_39934,N_39520);
or U40141 (N_40141,N_39469,N_39181);
xnor U40142 (N_40142,N_39562,N_39197);
and U40143 (N_40143,N_39082,N_39991);
nor U40144 (N_40144,N_39480,N_39818);
nor U40145 (N_40145,N_39704,N_39430);
xnor U40146 (N_40146,N_39637,N_39011);
xnor U40147 (N_40147,N_39025,N_39690);
xor U40148 (N_40148,N_39914,N_39782);
xor U40149 (N_40149,N_39573,N_39931);
nand U40150 (N_40150,N_39282,N_39989);
xor U40151 (N_40151,N_39557,N_39877);
nor U40152 (N_40152,N_39951,N_39273);
nand U40153 (N_40153,N_39379,N_39695);
nand U40154 (N_40154,N_39581,N_39712);
nand U40155 (N_40155,N_39071,N_39605);
xor U40156 (N_40156,N_39549,N_39570);
and U40157 (N_40157,N_39281,N_39113);
nand U40158 (N_40158,N_39286,N_39816);
and U40159 (N_40159,N_39552,N_39923);
nor U40160 (N_40160,N_39138,N_39115);
nor U40161 (N_40161,N_39255,N_39041);
nor U40162 (N_40162,N_39873,N_39313);
xnor U40163 (N_40163,N_39922,N_39364);
and U40164 (N_40164,N_39784,N_39739);
or U40165 (N_40165,N_39190,N_39306);
nor U40166 (N_40166,N_39604,N_39727);
nand U40167 (N_40167,N_39450,N_39078);
xor U40168 (N_40168,N_39470,N_39607);
xor U40169 (N_40169,N_39671,N_39079);
or U40170 (N_40170,N_39317,N_39236);
nand U40171 (N_40171,N_39103,N_39359);
nand U40172 (N_40172,N_39993,N_39830);
nand U40173 (N_40173,N_39673,N_39916);
nor U40174 (N_40174,N_39822,N_39366);
or U40175 (N_40175,N_39527,N_39717);
nor U40176 (N_40176,N_39345,N_39361);
and U40177 (N_40177,N_39371,N_39884);
xnor U40178 (N_40178,N_39928,N_39870);
nor U40179 (N_40179,N_39658,N_39326);
nor U40180 (N_40180,N_39895,N_39062);
or U40181 (N_40181,N_39108,N_39503);
xor U40182 (N_40182,N_39719,N_39203);
nor U40183 (N_40183,N_39453,N_39551);
xnor U40184 (N_40184,N_39620,N_39946);
nand U40185 (N_40185,N_39541,N_39294);
nand U40186 (N_40186,N_39283,N_39085);
xnor U40187 (N_40187,N_39560,N_39743);
nor U40188 (N_40188,N_39917,N_39457);
nor U40189 (N_40189,N_39879,N_39489);
or U40190 (N_40190,N_39756,N_39091);
nor U40191 (N_40191,N_39977,N_39587);
or U40192 (N_40192,N_39882,N_39554);
nor U40193 (N_40193,N_39561,N_39038);
xnor U40194 (N_40194,N_39331,N_39733);
and U40195 (N_40195,N_39613,N_39391);
nor U40196 (N_40196,N_39483,N_39716);
xnor U40197 (N_40197,N_39254,N_39429);
nand U40198 (N_40198,N_39693,N_39856);
xor U40199 (N_40199,N_39836,N_39995);
and U40200 (N_40200,N_39179,N_39261);
and U40201 (N_40201,N_39867,N_39382);
xor U40202 (N_40202,N_39631,N_39504);
and U40203 (N_40203,N_39913,N_39576);
nand U40204 (N_40204,N_39996,N_39169);
nand U40205 (N_40205,N_39768,N_39621);
nand U40206 (N_40206,N_39295,N_39563);
xor U40207 (N_40207,N_39271,N_39230);
and U40208 (N_40208,N_39066,N_39511);
nor U40209 (N_40209,N_39198,N_39903);
or U40210 (N_40210,N_39545,N_39599);
nand U40211 (N_40211,N_39380,N_39164);
or U40212 (N_40212,N_39614,N_39452);
nor U40213 (N_40213,N_39942,N_39692);
nor U40214 (N_40214,N_39226,N_39046);
and U40215 (N_40215,N_39101,N_39742);
nor U40216 (N_40216,N_39329,N_39760);
and U40217 (N_40217,N_39793,N_39881);
or U40218 (N_40218,N_39812,N_39428);
xnor U40219 (N_40219,N_39795,N_39205);
and U40220 (N_40220,N_39001,N_39950);
nand U40221 (N_40221,N_39464,N_39149);
or U40222 (N_40222,N_39752,N_39200);
and U40223 (N_40223,N_39855,N_39471);
or U40224 (N_40224,N_39598,N_39670);
and U40225 (N_40225,N_39969,N_39798);
nor U40226 (N_40226,N_39487,N_39180);
xor U40227 (N_40227,N_39183,N_39750);
nand U40228 (N_40228,N_39276,N_39508);
or U40229 (N_40229,N_39002,N_39709);
nand U40230 (N_40230,N_39998,N_39386);
nor U40231 (N_40231,N_39944,N_39336);
and U40232 (N_40232,N_39029,N_39529);
nand U40233 (N_40233,N_39096,N_39633);
nor U40234 (N_40234,N_39161,N_39488);
xnor U40235 (N_40235,N_39451,N_39398);
nand U40236 (N_40236,N_39650,N_39300);
xor U40237 (N_40237,N_39703,N_39815);
xor U40238 (N_40238,N_39819,N_39150);
nand U40239 (N_40239,N_39924,N_39250);
and U40240 (N_40240,N_39424,N_39432);
xnor U40241 (N_40241,N_39338,N_39533);
xor U40242 (N_40242,N_39492,N_39258);
xnor U40243 (N_40243,N_39178,N_39443);
and U40244 (N_40244,N_39435,N_39751);
nor U40245 (N_40245,N_39482,N_39279);
or U40246 (N_40246,N_39904,N_39710);
or U40247 (N_40247,N_39891,N_39272);
nor U40248 (N_40248,N_39182,N_39837);
nor U40249 (N_40249,N_39806,N_39808);
or U40250 (N_40250,N_39410,N_39965);
xor U40251 (N_40251,N_39908,N_39296);
and U40252 (N_40252,N_39669,N_39000);
nand U40253 (N_40253,N_39231,N_39442);
nor U40254 (N_40254,N_39142,N_39212);
xnor U40255 (N_40255,N_39729,N_39099);
nand U40256 (N_40256,N_39406,N_39239);
xor U40257 (N_40257,N_39810,N_39084);
xor U40258 (N_40258,N_39635,N_39093);
xnor U40259 (N_40259,N_39814,N_39732);
nor U40260 (N_40260,N_39128,N_39124);
nand U40261 (N_40261,N_39841,N_39544);
nor U40262 (N_40262,N_39897,N_39052);
or U40263 (N_40263,N_39696,N_39357);
xnor U40264 (N_40264,N_39513,N_39728);
or U40265 (N_40265,N_39207,N_39467);
or U40266 (N_40266,N_39921,N_39803);
or U40267 (N_40267,N_39064,N_39610);
and U40268 (N_40268,N_39736,N_39652);
nor U40269 (N_40269,N_39603,N_39518);
xor U40270 (N_40270,N_39438,N_39454);
and U40271 (N_40271,N_39990,N_39668);
nand U40272 (N_40272,N_39387,N_39321);
xor U40273 (N_40273,N_39004,N_39525);
xor U40274 (N_40274,N_39864,N_39086);
nand U40275 (N_40275,N_39912,N_39606);
nand U40276 (N_40276,N_39857,N_39367);
xor U40277 (N_40277,N_39689,N_39817);
xnor U40278 (N_40278,N_39697,N_39339);
nand U40279 (N_40279,N_39440,N_39163);
nor U40280 (N_40280,N_39403,N_39298);
nor U40281 (N_40281,N_39444,N_39308);
xnor U40282 (N_40282,N_39964,N_39523);
and U40283 (N_40283,N_39372,N_39813);
and U40284 (N_40284,N_39278,N_39215);
xnor U40285 (N_40285,N_39427,N_39832);
xor U40286 (N_40286,N_39290,N_39569);
xnor U40287 (N_40287,N_39125,N_39983);
or U40288 (N_40288,N_39332,N_39796);
or U40289 (N_40289,N_39787,N_39985);
xnor U40290 (N_40290,N_39495,N_39365);
or U40291 (N_40291,N_39019,N_39012);
or U40292 (N_40292,N_39399,N_39683);
or U40293 (N_40293,N_39018,N_39042);
xor U40294 (N_40294,N_39878,N_39789);
nand U40295 (N_40295,N_39119,N_39186);
and U40296 (N_40296,N_39218,N_39799);
xnor U40297 (N_40297,N_39389,N_39746);
or U40298 (N_40298,N_39953,N_39490);
or U40299 (N_40299,N_39838,N_39848);
nand U40300 (N_40300,N_39866,N_39401);
xnor U40301 (N_40301,N_39165,N_39077);
xnor U40302 (N_40302,N_39307,N_39228);
xor U40303 (N_40303,N_39472,N_39309);
nand U40304 (N_40304,N_39167,N_39243);
or U40305 (N_40305,N_39040,N_39981);
nand U40306 (N_40306,N_39823,N_39737);
nor U40307 (N_40307,N_39687,N_39767);
nor U40308 (N_40308,N_39639,N_39484);
or U40309 (N_40309,N_39354,N_39577);
nor U40310 (N_40310,N_39133,N_39824);
and U40311 (N_40311,N_39493,N_39140);
and U40312 (N_40312,N_39745,N_39334);
nand U40313 (N_40313,N_39431,N_39932);
nor U40314 (N_40314,N_39846,N_39754);
xnor U40315 (N_40315,N_39802,N_39349);
or U40316 (N_40316,N_39646,N_39247);
nand U40317 (N_40317,N_39535,N_39016);
xnor U40318 (N_40318,N_39597,N_39869);
and U40319 (N_40319,N_39642,N_39268);
nor U40320 (N_40320,N_39672,N_39350);
or U40321 (N_40321,N_39343,N_39199);
nor U40322 (N_40322,N_39157,N_39166);
nand U40323 (N_40323,N_39026,N_39644);
and U40324 (N_40324,N_39501,N_39110);
nor U40325 (N_40325,N_39972,N_39314);
nand U40326 (N_40326,N_39075,N_39434);
nor U40327 (N_40327,N_39766,N_39475);
xnor U40328 (N_40328,N_39588,N_39828);
xor U40329 (N_40329,N_39999,N_39959);
and U40330 (N_40330,N_39240,N_39297);
or U40331 (N_40331,N_39136,N_39104);
xor U40332 (N_40332,N_39548,N_39176);
nand U40333 (N_40333,N_39834,N_39460);
and U40334 (N_40334,N_39627,N_39542);
nand U40335 (N_40335,N_39061,N_39462);
nor U40336 (N_40336,N_39284,N_39035);
or U40337 (N_40337,N_39890,N_39285);
or U40338 (N_40338,N_39057,N_39252);
nor U40339 (N_40339,N_39437,N_39275);
and U40340 (N_40340,N_39143,N_39048);
and U40341 (N_40341,N_39074,N_39976);
nor U40342 (N_40342,N_39885,N_39147);
xor U40343 (N_40343,N_39609,N_39952);
or U40344 (N_40344,N_39033,N_39117);
xnor U40345 (N_40345,N_39531,N_39971);
nand U40346 (N_40346,N_39807,N_39685);
nand U40347 (N_40347,N_39390,N_39344);
nor U40348 (N_40348,N_39628,N_39898);
nand U40349 (N_40349,N_39355,N_39481);
or U40350 (N_40350,N_39725,N_39698);
or U40351 (N_40351,N_39193,N_39127);
or U40352 (N_40352,N_39189,N_39049);
nand U40353 (N_40353,N_39051,N_39844);
and U40354 (N_40354,N_39436,N_39174);
nand U40355 (N_40355,N_39417,N_39479);
and U40356 (N_40356,N_39532,N_39572);
xor U40357 (N_40357,N_39731,N_39778);
nand U40358 (N_40358,N_39447,N_39862);
nand U40359 (N_40359,N_39939,N_39740);
or U40360 (N_40360,N_39920,N_39184);
and U40361 (N_40361,N_39648,N_39328);
xnor U40362 (N_40362,N_39311,N_39776);
nand U40363 (N_40363,N_39797,N_39263);
xor U40364 (N_40364,N_39852,N_39393);
nor U40365 (N_40365,N_39970,N_39718);
and U40366 (N_40366,N_39515,N_39289);
nand U40367 (N_40367,N_39847,N_39055);
nand U40368 (N_40368,N_39269,N_39188);
and U40369 (N_40369,N_39210,N_39871);
and U40370 (N_40370,N_39031,N_39172);
nor U40371 (N_40371,N_39316,N_39159);
and U40372 (N_40372,N_39641,N_39780);
nand U40373 (N_40373,N_39507,N_39419);
xor U40374 (N_40374,N_39688,N_39765);
nor U40375 (N_40375,N_39761,N_39301);
nand U40376 (N_40376,N_39396,N_39013);
xor U40377 (N_40377,N_39677,N_39909);
nor U40378 (N_40378,N_39988,N_39409);
and U40379 (N_40379,N_39324,N_39109);
xnor U40380 (N_40380,N_39170,N_39539);
nand U40381 (N_40381,N_39674,N_39293);
and U40382 (N_40382,N_39145,N_39217);
nor U40383 (N_40383,N_39494,N_39565);
nor U40384 (N_40384,N_39863,N_39351);
nand U40385 (N_40385,N_39461,N_39039);
or U40386 (N_40386,N_39580,N_39134);
and U40387 (N_40387,N_39868,N_39849);
or U40388 (N_40388,N_39886,N_39219);
nor U40389 (N_40389,N_39526,N_39594);
nor U40390 (N_40390,N_39009,N_39547);
xnor U40391 (N_40391,N_39418,N_39530);
nor U40392 (N_40392,N_39028,N_39017);
xnor U40393 (N_40393,N_39007,N_39771);
nand U40394 (N_40394,N_39860,N_39232);
nand U40395 (N_40395,N_39256,N_39902);
xor U40396 (N_40396,N_39356,N_39233);
xor U40397 (N_40397,N_39439,N_39947);
and U40398 (N_40398,N_39595,N_39937);
xnor U40399 (N_40399,N_39684,N_39723);
nor U40400 (N_40400,N_39659,N_39593);
or U40401 (N_40401,N_39788,N_39954);
nand U40402 (N_40402,N_39558,N_39459);
or U40403 (N_40403,N_39496,N_39144);
and U40404 (N_40404,N_39600,N_39901);
xor U40405 (N_40405,N_39310,N_39358);
xnor U40406 (N_40406,N_39216,N_39449);
nand U40407 (N_40407,N_39850,N_39583);
and U40408 (N_40408,N_39370,N_39918);
nand U40409 (N_40409,N_39021,N_39888);
nand U40410 (N_40410,N_39543,N_39632);
xor U40411 (N_40411,N_39223,N_39783);
nor U40412 (N_40412,N_39770,N_39262);
or U40413 (N_40413,N_39476,N_39794);
or U40414 (N_40414,N_39466,N_39253);
xor U40415 (N_40415,N_39020,N_39473);
and U40416 (N_40416,N_39925,N_39065);
or U40417 (N_40417,N_39986,N_39773);
nand U40418 (N_40418,N_39656,N_39126);
nand U40419 (N_40419,N_39323,N_39202);
nand U40420 (N_40420,N_39267,N_39395);
nand U40421 (N_40421,N_39617,N_39225);
nor U40422 (N_40422,N_39368,N_39777);
nand U40423 (N_40423,N_39987,N_39682);
nor U40424 (N_40424,N_39106,N_39095);
nand U40425 (N_40425,N_39827,N_39277);
or U40426 (N_40426,N_39537,N_39889);
nor U40427 (N_40427,N_39843,N_39791);
nand U40428 (N_40428,N_39027,N_39465);
nand U40429 (N_40429,N_39556,N_39591);
nor U40430 (N_40430,N_39341,N_39416);
and U40431 (N_40431,N_39388,N_39651);
and U40432 (N_40432,N_39522,N_39089);
xor U40433 (N_40433,N_39966,N_39734);
or U40434 (N_40434,N_39342,N_39337);
nand U40435 (N_40435,N_39546,N_39616);
and U40436 (N_40436,N_39325,N_39130);
or U40437 (N_40437,N_39222,N_39266);
and U40438 (N_40438,N_39383,N_39402);
nand U40439 (N_40439,N_39722,N_39715);
nand U40440 (N_40440,N_39107,N_39938);
and U40441 (N_40441,N_39477,N_39118);
and U40442 (N_40442,N_39375,N_39657);
nand U40443 (N_40443,N_39116,N_39076);
xor U40444 (N_40444,N_39288,N_39883);
and U40445 (N_40445,N_39949,N_39155);
xnor U40446 (N_40446,N_39348,N_39973);
and U40447 (N_40447,N_39420,N_39666);
nor U40448 (N_40448,N_39245,N_39015);
or U40449 (N_40449,N_39781,N_39248);
xnor U40450 (N_40450,N_39265,N_39320);
xor U40451 (N_40451,N_39707,N_39578);
nand U40452 (N_40452,N_39630,N_39700);
or U40453 (N_40453,N_39360,N_39809);
nand U40454 (N_40454,N_39910,N_39675);
or U40455 (N_40455,N_39930,N_39105);
or U40456 (N_40456,N_39083,N_39741);
nand U40457 (N_40457,N_39060,N_39185);
or U40458 (N_40458,N_39448,N_39433);
and U40459 (N_40459,N_39456,N_39098);
nor U40460 (N_40460,N_39538,N_39054);
or U40461 (N_40461,N_39945,N_39008);
nor U40462 (N_40462,N_39377,N_39851);
nor U40463 (N_40463,N_39559,N_39050);
and U40464 (N_40464,N_39195,N_39979);
xnor U40465 (N_40465,N_39919,N_39713);
and U40466 (N_40466,N_39214,N_39790);
and U40467 (N_40467,N_39831,N_39943);
nor U40468 (N_40468,N_39747,N_39759);
or U40469 (N_40469,N_39139,N_39568);
xnor U40470 (N_40470,N_39978,N_39251);
nor U40471 (N_40471,N_39622,N_39611);
and U40472 (N_40472,N_39900,N_39984);
nor U40473 (N_40473,N_39363,N_39446);
and U40474 (N_40474,N_39299,N_39872);
and U40475 (N_40475,N_39842,N_39353);
xnor U40476 (N_40476,N_39241,N_39485);
nor U40477 (N_40477,N_39413,N_39080);
nand U40478 (N_40478,N_39238,N_39655);
nor U40479 (N_40479,N_39510,N_39384);
and U40480 (N_40480,N_39840,N_39769);
nand U40481 (N_40481,N_39854,N_39229);
or U40482 (N_40482,N_39235,N_39601);
xor U40483 (N_40483,N_39246,N_39037);
xnor U40484 (N_40484,N_39702,N_39926);
or U40485 (N_40485,N_39907,N_39992);
and U40486 (N_40486,N_39654,N_39748);
or U40487 (N_40487,N_39619,N_39714);
and U40488 (N_40488,N_39244,N_39315);
and U40489 (N_40489,N_39582,N_39445);
nand U40490 (N_40490,N_39486,N_39412);
nor U40491 (N_40491,N_39063,N_39536);
and U40492 (N_40492,N_39974,N_39152);
xnor U40493 (N_40493,N_39955,N_39090);
and U40494 (N_40494,N_39302,N_39694);
xnor U40495 (N_40495,N_39094,N_39073);
or U40496 (N_40496,N_39726,N_39270);
or U40497 (N_40497,N_39618,N_39623);
or U40498 (N_40498,N_39540,N_39319);
nor U40499 (N_40499,N_39735,N_39893);
or U40500 (N_40500,N_39940,N_39568);
nor U40501 (N_40501,N_39865,N_39465);
and U40502 (N_40502,N_39507,N_39791);
nor U40503 (N_40503,N_39555,N_39146);
xnor U40504 (N_40504,N_39498,N_39400);
xor U40505 (N_40505,N_39144,N_39479);
nand U40506 (N_40506,N_39855,N_39005);
nand U40507 (N_40507,N_39422,N_39785);
or U40508 (N_40508,N_39813,N_39759);
and U40509 (N_40509,N_39377,N_39072);
xor U40510 (N_40510,N_39093,N_39984);
xor U40511 (N_40511,N_39880,N_39044);
xnor U40512 (N_40512,N_39396,N_39131);
or U40513 (N_40513,N_39291,N_39058);
or U40514 (N_40514,N_39871,N_39256);
nand U40515 (N_40515,N_39437,N_39265);
nand U40516 (N_40516,N_39540,N_39743);
and U40517 (N_40517,N_39277,N_39704);
xnor U40518 (N_40518,N_39286,N_39649);
or U40519 (N_40519,N_39715,N_39932);
and U40520 (N_40520,N_39386,N_39657);
xnor U40521 (N_40521,N_39592,N_39078);
nand U40522 (N_40522,N_39131,N_39263);
xnor U40523 (N_40523,N_39384,N_39418);
xor U40524 (N_40524,N_39856,N_39039);
or U40525 (N_40525,N_39228,N_39557);
and U40526 (N_40526,N_39925,N_39251);
nand U40527 (N_40527,N_39175,N_39743);
and U40528 (N_40528,N_39771,N_39367);
or U40529 (N_40529,N_39278,N_39633);
xor U40530 (N_40530,N_39152,N_39773);
or U40531 (N_40531,N_39583,N_39023);
nand U40532 (N_40532,N_39823,N_39345);
xor U40533 (N_40533,N_39814,N_39194);
xor U40534 (N_40534,N_39990,N_39050);
and U40535 (N_40535,N_39887,N_39003);
or U40536 (N_40536,N_39676,N_39258);
nor U40537 (N_40537,N_39793,N_39129);
or U40538 (N_40538,N_39601,N_39757);
and U40539 (N_40539,N_39386,N_39216);
nand U40540 (N_40540,N_39771,N_39966);
xnor U40541 (N_40541,N_39162,N_39368);
xnor U40542 (N_40542,N_39628,N_39448);
xnor U40543 (N_40543,N_39794,N_39844);
and U40544 (N_40544,N_39260,N_39150);
or U40545 (N_40545,N_39158,N_39029);
and U40546 (N_40546,N_39455,N_39986);
nand U40547 (N_40547,N_39826,N_39616);
or U40548 (N_40548,N_39465,N_39490);
or U40549 (N_40549,N_39078,N_39767);
or U40550 (N_40550,N_39460,N_39370);
nor U40551 (N_40551,N_39556,N_39947);
or U40552 (N_40552,N_39517,N_39588);
and U40553 (N_40553,N_39859,N_39017);
nand U40554 (N_40554,N_39017,N_39789);
or U40555 (N_40555,N_39685,N_39667);
and U40556 (N_40556,N_39961,N_39899);
and U40557 (N_40557,N_39746,N_39016);
and U40558 (N_40558,N_39886,N_39742);
and U40559 (N_40559,N_39546,N_39127);
and U40560 (N_40560,N_39742,N_39179);
and U40561 (N_40561,N_39950,N_39017);
nor U40562 (N_40562,N_39956,N_39141);
nand U40563 (N_40563,N_39371,N_39507);
or U40564 (N_40564,N_39674,N_39570);
and U40565 (N_40565,N_39065,N_39178);
nand U40566 (N_40566,N_39191,N_39846);
and U40567 (N_40567,N_39680,N_39234);
xnor U40568 (N_40568,N_39305,N_39635);
nor U40569 (N_40569,N_39558,N_39653);
and U40570 (N_40570,N_39233,N_39660);
xnor U40571 (N_40571,N_39526,N_39403);
xor U40572 (N_40572,N_39721,N_39962);
nor U40573 (N_40573,N_39629,N_39923);
nand U40574 (N_40574,N_39574,N_39490);
nand U40575 (N_40575,N_39281,N_39800);
nand U40576 (N_40576,N_39201,N_39620);
nand U40577 (N_40577,N_39485,N_39690);
nand U40578 (N_40578,N_39346,N_39742);
xor U40579 (N_40579,N_39035,N_39065);
nand U40580 (N_40580,N_39370,N_39750);
xnor U40581 (N_40581,N_39345,N_39583);
and U40582 (N_40582,N_39315,N_39890);
and U40583 (N_40583,N_39632,N_39362);
xor U40584 (N_40584,N_39098,N_39925);
or U40585 (N_40585,N_39904,N_39368);
nand U40586 (N_40586,N_39456,N_39954);
or U40587 (N_40587,N_39487,N_39446);
xnor U40588 (N_40588,N_39158,N_39481);
and U40589 (N_40589,N_39415,N_39757);
or U40590 (N_40590,N_39128,N_39833);
nand U40591 (N_40591,N_39277,N_39553);
nand U40592 (N_40592,N_39889,N_39240);
xor U40593 (N_40593,N_39304,N_39499);
nor U40594 (N_40594,N_39942,N_39708);
nor U40595 (N_40595,N_39562,N_39938);
xnor U40596 (N_40596,N_39009,N_39124);
xnor U40597 (N_40597,N_39624,N_39901);
nor U40598 (N_40598,N_39562,N_39376);
xor U40599 (N_40599,N_39588,N_39014);
xor U40600 (N_40600,N_39293,N_39798);
nand U40601 (N_40601,N_39130,N_39646);
or U40602 (N_40602,N_39646,N_39430);
nor U40603 (N_40603,N_39199,N_39267);
and U40604 (N_40604,N_39487,N_39270);
and U40605 (N_40605,N_39963,N_39928);
and U40606 (N_40606,N_39401,N_39245);
and U40607 (N_40607,N_39055,N_39044);
nor U40608 (N_40608,N_39997,N_39458);
xor U40609 (N_40609,N_39168,N_39346);
nand U40610 (N_40610,N_39630,N_39563);
xor U40611 (N_40611,N_39020,N_39013);
or U40612 (N_40612,N_39050,N_39083);
xnor U40613 (N_40613,N_39438,N_39723);
nor U40614 (N_40614,N_39087,N_39724);
nand U40615 (N_40615,N_39783,N_39359);
nand U40616 (N_40616,N_39363,N_39034);
nand U40617 (N_40617,N_39930,N_39056);
xor U40618 (N_40618,N_39716,N_39685);
xor U40619 (N_40619,N_39806,N_39812);
xor U40620 (N_40620,N_39858,N_39030);
and U40621 (N_40621,N_39515,N_39136);
and U40622 (N_40622,N_39702,N_39413);
and U40623 (N_40623,N_39198,N_39373);
nand U40624 (N_40624,N_39541,N_39880);
and U40625 (N_40625,N_39405,N_39572);
xnor U40626 (N_40626,N_39819,N_39556);
nor U40627 (N_40627,N_39684,N_39776);
or U40628 (N_40628,N_39867,N_39834);
nand U40629 (N_40629,N_39512,N_39032);
and U40630 (N_40630,N_39625,N_39334);
nor U40631 (N_40631,N_39751,N_39289);
nand U40632 (N_40632,N_39663,N_39900);
nand U40633 (N_40633,N_39642,N_39623);
nand U40634 (N_40634,N_39758,N_39199);
nand U40635 (N_40635,N_39031,N_39806);
nand U40636 (N_40636,N_39018,N_39609);
nand U40637 (N_40637,N_39210,N_39228);
and U40638 (N_40638,N_39852,N_39889);
nor U40639 (N_40639,N_39639,N_39888);
or U40640 (N_40640,N_39735,N_39192);
nand U40641 (N_40641,N_39815,N_39500);
or U40642 (N_40642,N_39548,N_39393);
or U40643 (N_40643,N_39896,N_39510);
or U40644 (N_40644,N_39848,N_39362);
nor U40645 (N_40645,N_39126,N_39765);
nor U40646 (N_40646,N_39753,N_39643);
nand U40647 (N_40647,N_39493,N_39687);
and U40648 (N_40648,N_39818,N_39255);
and U40649 (N_40649,N_39193,N_39964);
and U40650 (N_40650,N_39260,N_39392);
and U40651 (N_40651,N_39053,N_39885);
xnor U40652 (N_40652,N_39201,N_39230);
and U40653 (N_40653,N_39062,N_39880);
nor U40654 (N_40654,N_39606,N_39719);
and U40655 (N_40655,N_39461,N_39233);
nand U40656 (N_40656,N_39416,N_39321);
and U40657 (N_40657,N_39305,N_39209);
nand U40658 (N_40658,N_39464,N_39379);
nor U40659 (N_40659,N_39060,N_39190);
and U40660 (N_40660,N_39617,N_39753);
and U40661 (N_40661,N_39865,N_39916);
and U40662 (N_40662,N_39920,N_39783);
or U40663 (N_40663,N_39552,N_39847);
and U40664 (N_40664,N_39568,N_39307);
nand U40665 (N_40665,N_39113,N_39620);
xnor U40666 (N_40666,N_39726,N_39763);
xor U40667 (N_40667,N_39176,N_39688);
or U40668 (N_40668,N_39058,N_39153);
or U40669 (N_40669,N_39227,N_39454);
or U40670 (N_40670,N_39947,N_39788);
xor U40671 (N_40671,N_39927,N_39316);
nand U40672 (N_40672,N_39350,N_39911);
and U40673 (N_40673,N_39896,N_39911);
nand U40674 (N_40674,N_39704,N_39336);
or U40675 (N_40675,N_39261,N_39753);
and U40676 (N_40676,N_39797,N_39754);
or U40677 (N_40677,N_39445,N_39883);
or U40678 (N_40678,N_39972,N_39194);
or U40679 (N_40679,N_39376,N_39900);
nand U40680 (N_40680,N_39242,N_39098);
nand U40681 (N_40681,N_39762,N_39438);
nor U40682 (N_40682,N_39809,N_39035);
or U40683 (N_40683,N_39562,N_39815);
or U40684 (N_40684,N_39109,N_39140);
or U40685 (N_40685,N_39375,N_39584);
or U40686 (N_40686,N_39557,N_39934);
and U40687 (N_40687,N_39349,N_39769);
xnor U40688 (N_40688,N_39338,N_39077);
and U40689 (N_40689,N_39794,N_39575);
xor U40690 (N_40690,N_39520,N_39603);
xnor U40691 (N_40691,N_39005,N_39475);
nor U40692 (N_40692,N_39020,N_39305);
nor U40693 (N_40693,N_39023,N_39566);
or U40694 (N_40694,N_39525,N_39070);
or U40695 (N_40695,N_39287,N_39994);
nor U40696 (N_40696,N_39595,N_39321);
nand U40697 (N_40697,N_39276,N_39300);
nand U40698 (N_40698,N_39859,N_39551);
and U40699 (N_40699,N_39372,N_39282);
nor U40700 (N_40700,N_39857,N_39982);
and U40701 (N_40701,N_39410,N_39891);
or U40702 (N_40702,N_39666,N_39350);
or U40703 (N_40703,N_39086,N_39339);
or U40704 (N_40704,N_39117,N_39638);
or U40705 (N_40705,N_39751,N_39076);
nand U40706 (N_40706,N_39156,N_39510);
xnor U40707 (N_40707,N_39765,N_39853);
nor U40708 (N_40708,N_39366,N_39691);
or U40709 (N_40709,N_39937,N_39023);
or U40710 (N_40710,N_39090,N_39380);
and U40711 (N_40711,N_39912,N_39624);
and U40712 (N_40712,N_39148,N_39303);
and U40713 (N_40713,N_39127,N_39618);
and U40714 (N_40714,N_39257,N_39851);
nor U40715 (N_40715,N_39434,N_39993);
xnor U40716 (N_40716,N_39581,N_39522);
xnor U40717 (N_40717,N_39069,N_39670);
nor U40718 (N_40718,N_39296,N_39580);
and U40719 (N_40719,N_39298,N_39962);
nand U40720 (N_40720,N_39492,N_39802);
xor U40721 (N_40721,N_39835,N_39056);
nor U40722 (N_40722,N_39533,N_39746);
nand U40723 (N_40723,N_39628,N_39401);
nand U40724 (N_40724,N_39800,N_39608);
and U40725 (N_40725,N_39777,N_39653);
or U40726 (N_40726,N_39696,N_39975);
and U40727 (N_40727,N_39510,N_39076);
nand U40728 (N_40728,N_39243,N_39372);
xnor U40729 (N_40729,N_39434,N_39043);
nor U40730 (N_40730,N_39031,N_39110);
nor U40731 (N_40731,N_39636,N_39756);
nand U40732 (N_40732,N_39387,N_39527);
xnor U40733 (N_40733,N_39275,N_39537);
xnor U40734 (N_40734,N_39313,N_39957);
nor U40735 (N_40735,N_39940,N_39437);
xnor U40736 (N_40736,N_39464,N_39421);
nand U40737 (N_40737,N_39957,N_39644);
nor U40738 (N_40738,N_39567,N_39940);
xor U40739 (N_40739,N_39992,N_39943);
nor U40740 (N_40740,N_39222,N_39973);
xor U40741 (N_40741,N_39756,N_39308);
nand U40742 (N_40742,N_39473,N_39295);
nand U40743 (N_40743,N_39244,N_39501);
nor U40744 (N_40744,N_39705,N_39708);
and U40745 (N_40745,N_39504,N_39234);
or U40746 (N_40746,N_39913,N_39513);
and U40747 (N_40747,N_39238,N_39605);
and U40748 (N_40748,N_39769,N_39896);
nor U40749 (N_40749,N_39597,N_39718);
or U40750 (N_40750,N_39033,N_39443);
and U40751 (N_40751,N_39006,N_39594);
and U40752 (N_40752,N_39244,N_39789);
nor U40753 (N_40753,N_39882,N_39703);
nand U40754 (N_40754,N_39403,N_39218);
nand U40755 (N_40755,N_39962,N_39679);
and U40756 (N_40756,N_39057,N_39261);
xor U40757 (N_40757,N_39363,N_39852);
nand U40758 (N_40758,N_39590,N_39947);
and U40759 (N_40759,N_39878,N_39804);
nand U40760 (N_40760,N_39938,N_39335);
xor U40761 (N_40761,N_39492,N_39450);
or U40762 (N_40762,N_39249,N_39097);
or U40763 (N_40763,N_39346,N_39916);
nand U40764 (N_40764,N_39084,N_39698);
xor U40765 (N_40765,N_39851,N_39115);
and U40766 (N_40766,N_39290,N_39329);
or U40767 (N_40767,N_39022,N_39129);
and U40768 (N_40768,N_39237,N_39964);
xnor U40769 (N_40769,N_39853,N_39096);
nand U40770 (N_40770,N_39152,N_39438);
xor U40771 (N_40771,N_39063,N_39133);
nor U40772 (N_40772,N_39937,N_39341);
or U40773 (N_40773,N_39616,N_39790);
or U40774 (N_40774,N_39952,N_39349);
nor U40775 (N_40775,N_39096,N_39766);
nor U40776 (N_40776,N_39954,N_39664);
or U40777 (N_40777,N_39083,N_39899);
nand U40778 (N_40778,N_39616,N_39356);
nor U40779 (N_40779,N_39128,N_39982);
or U40780 (N_40780,N_39751,N_39066);
nor U40781 (N_40781,N_39218,N_39763);
and U40782 (N_40782,N_39952,N_39759);
nand U40783 (N_40783,N_39672,N_39094);
nand U40784 (N_40784,N_39781,N_39612);
nand U40785 (N_40785,N_39286,N_39798);
nor U40786 (N_40786,N_39644,N_39990);
and U40787 (N_40787,N_39407,N_39135);
xnor U40788 (N_40788,N_39111,N_39212);
and U40789 (N_40789,N_39452,N_39807);
or U40790 (N_40790,N_39774,N_39271);
or U40791 (N_40791,N_39919,N_39856);
or U40792 (N_40792,N_39385,N_39020);
and U40793 (N_40793,N_39653,N_39421);
nor U40794 (N_40794,N_39828,N_39135);
nor U40795 (N_40795,N_39018,N_39692);
and U40796 (N_40796,N_39903,N_39905);
or U40797 (N_40797,N_39616,N_39269);
nand U40798 (N_40798,N_39004,N_39113);
nor U40799 (N_40799,N_39556,N_39474);
xor U40800 (N_40800,N_39026,N_39126);
xor U40801 (N_40801,N_39827,N_39012);
xor U40802 (N_40802,N_39175,N_39991);
xnor U40803 (N_40803,N_39645,N_39222);
and U40804 (N_40804,N_39246,N_39411);
nand U40805 (N_40805,N_39663,N_39212);
xor U40806 (N_40806,N_39391,N_39827);
xnor U40807 (N_40807,N_39276,N_39647);
and U40808 (N_40808,N_39884,N_39153);
and U40809 (N_40809,N_39168,N_39167);
or U40810 (N_40810,N_39634,N_39474);
nor U40811 (N_40811,N_39952,N_39333);
nand U40812 (N_40812,N_39919,N_39196);
xnor U40813 (N_40813,N_39191,N_39140);
nand U40814 (N_40814,N_39647,N_39272);
nor U40815 (N_40815,N_39479,N_39965);
nand U40816 (N_40816,N_39374,N_39518);
nor U40817 (N_40817,N_39973,N_39832);
or U40818 (N_40818,N_39849,N_39935);
nand U40819 (N_40819,N_39115,N_39934);
nor U40820 (N_40820,N_39137,N_39523);
xnor U40821 (N_40821,N_39767,N_39210);
nand U40822 (N_40822,N_39584,N_39910);
nand U40823 (N_40823,N_39996,N_39015);
or U40824 (N_40824,N_39624,N_39439);
nand U40825 (N_40825,N_39652,N_39147);
xor U40826 (N_40826,N_39261,N_39333);
and U40827 (N_40827,N_39742,N_39530);
xor U40828 (N_40828,N_39359,N_39871);
or U40829 (N_40829,N_39546,N_39147);
or U40830 (N_40830,N_39831,N_39850);
nand U40831 (N_40831,N_39940,N_39142);
nand U40832 (N_40832,N_39733,N_39118);
xor U40833 (N_40833,N_39581,N_39484);
nand U40834 (N_40834,N_39748,N_39931);
and U40835 (N_40835,N_39366,N_39579);
nor U40836 (N_40836,N_39461,N_39114);
and U40837 (N_40837,N_39219,N_39336);
or U40838 (N_40838,N_39134,N_39120);
and U40839 (N_40839,N_39743,N_39400);
nor U40840 (N_40840,N_39993,N_39112);
and U40841 (N_40841,N_39763,N_39802);
or U40842 (N_40842,N_39190,N_39123);
nor U40843 (N_40843,N_39884,N_39840);
nor U40844 (N_40844,N_39115,N_39316);
nor U40845 (N_40845,N_39010,N_39541);
or U40846 (N_40846,N_39944,N_39920);
nor U40847 (N_40847,N_39987,N_39545);
nor U40848 (N_40848,N_39332,N_39315);
and U40849 (N_40849,N_39351,N_39486);
or U40850 (N_40850,N_39389,N_39694);
xnor U40851 (N_40851,N_39683,N_39870);
xor U40852 (N_40852,N_39775,N_39851);
or U40853 (N_40853,N_39409,N_39408);
or U40854 (N_40854,N_39288,N_39402);
xor U40855 (N_40855,N_39826,N_39190);
or U40856 (N_40856,N_39921,N_39617);
and U40857 (N_40857,N_39032,N_39300);
xnor U40858 (N_40858,N_39691,N_39497);
xor U40859 (N_40859,N_39276,N_39356);
xnor U40860 (N_40860,N_39881,N_39890);
nor U40861 (N_40861,N_39306,N_39163);
and U40862 (N_40862,N_39969,N_39280);
xor U40863 (N_40863,N_39169,N_39737);
xnor U40864 (N_40864,N_39253,N_39660);
and U40865 (N_40865,N_39862,N_39028);
nor U40866 (N_40866,N_39954,N_39108);
nand U40867 (N_40867,N_39988,N_39168);
or U40868 (N_40868,N_39697,N_39125);
or U40869 (N_40869,N_39689,N_39032);
xnor U40870 (N_40870,N_39548,N_39792);
nor U40871 (N_40871,N_39184,N_39220);
or U40872 (N_40872,N_39396,N_39316);
nor U40873 (N_40873,N_39665,N_39741);
nor U40874 (N_40874,N_39070,N_39500);
xor U40875 (N_40875,N_39358,N_39312);
or U40876 (N_40876,N_39456,N_39595);
nand U40877 (N_40877,N_39467,N_39047);
nand U40878 (N_40878,N_39550,N_39147);
and U40879 (N_40879,N_39710,N_39226);
nor U40880 (N_40880,N_39589,N_39720);
and U40881 (N_40881,N_39330,N_39988);
or U40882 (N_40882,N_39628,N_39376);
and U40883 (N_40883,N_39837,N_39435);
nor U40884 (N_40884,N_39981,N_39705);
nand U40885 (N_40885,N_39753,N_39791);
nand U40886 (N_40886,N_39350,N_39994);
or U40887 (N_40887,N_39561,N_39487);
nor U40888 (N_40888,N_39327,N_39328);
nor U40889 (N_40889,N_39055,N_39371);
xor U40890 (N_40890,N_39271,N_39200);
nand U40891 (N_40891,N_39279,N_39704);
or U40892 (N_40892,N_39849,N_39394);
or U40893 (N_40893,N_39542,N_39292);
and U40894 (N_40894,N_39615,N_39783);
nor U40895 (N_40895,N_39655,N_39176);
nor U40896 (N_40896,N_39080,N_39829);
xor U40897 (N_40897,N_39585,N_39556);
or U40898 (N_40898,N_39210,N_39668);
or U40899 (N_40899,N_39711,N_39787);
or U40900 (N_40900,N_39297,N_39005);
xor U40901 (N_40901,N_39044,N_39158);
nor U40902 (N_40902,N_39204,N_39322);
xnor U40903 (N_40903,N_39853,N_39720);
nand U40904 (N_40904,N_39779,N_39054);
nor U40905 (N_40905,N_39754,N_39778);
and U40906 (N_40906,N_39629,N_39578);
and U40907 (N_40907,N_39880,N_39240);
xnor U40908 (N_40908,N_39270,N_39334);
and U40909 (N_40909,N_39907,N_39244);
nor U40910 (N_40910,N_39536,N_39329);
and U40911 (N_40911,N_39220,N_39243);
nor U40912 (N_40912,N_39741,N_39116);
nand U40913 (N_40913,N_39826,N_39970);
and U40914 (N_40914,N_39754,N_39893);
nand U40915 (N_40915,N_39885,N_39488);
nand U40916 (N_40916,N_39192,N_39563);
xor U40917 (N_40917,N_39406,N_39467);
xor U40918 (N_40918,N_39800,N_39186);
and U40919 (N_40919,N_39519,N_39900);
xor U40920 (N_40920,N_39856,N_39464);
xnor U40921 (N_40921,N_39912,N_39734);
or U40922 (N_40922,N_39809,N_39308);
and U40923 (N_40923,N_39511,N_39768);
nor U40924 (N_40924,N_39882,N_39230);
nor U40925 (N_40925,N_39066,N_39332);
nor U40926 (N_40926,N_39137,N_39928);
nand U40927 (N_40927,N_39896,N_39524);
nor U40928 (N_40928,N_39872,N_39688);
or U40929 (N_40929,N_39040,N_39207);
or U40930 (N_40930,N_39842,N_39501);
xnor U40931 (N_40931,N_39335,N_39833);
nor U40932 (N_40932,N_39052,N_39335);
or U40933 (N_40933,N_39104,N_39342);
nor U40934 (N_40934,N_39850,N_39213);
xor U40935 (N_40935,N_39145,N_39670);
nor U40936 (N_40936,N_39475,N_39220);
nor U40937 (N_40937,N_39694,N_39740);
xnor U40938 (N_40938,N_39317,N_39152);
xnor U40939 (N_40939,N_39343,N_39925);
xor U40940 (N_40940,N_39205,N_39901);
xor U40941 (N_40941,N_39554,N_39547);
xor U40942 (N_40942,N_39910,N_39648);
xnor U40943 (N_40943,N_39633,N_39531);
nand U40944 (N_40944,N_39560,N_39046);
xor U40945 (N_40945,N_39570,N_39353);
or U40946 (N_40946,N_39642,N_39717);
nor U40947 (N_40947,N_39525,N_39221);
and U40948 (N_40948,N_39870,N_39279);
xnor U40949 (N_40949,N_39717,N_39295);
xor U40950 (N_40950,N_39262,N_39509);
nand U40951 (N_40951,N_39804,N_39142);
nor U40952 (N_40952,N_39256,N_39831);
or U40953 (N_40953,N_39387,N_39930);
nor U40954 (N_40954,N_39765,N_39403);
or U40955 (N_40955,N_39434,N_39629);
nand U40956 (N_40956,N_39698,N_39723);
or U40957 (N_40957,N_39603,N_39236);
or U40958 (N_40958,N_39622,N_39310);
or U40959 (N_40959,N_39411,N_39277);
nor U40960 (N_40960,N_39908,N_39481);
xor U40961 (N_40961,N_39884,N_39094);
xor U40962 (N_40962,N_39900,N_39033);
nor U40963 (N_40963,N_39188,N_39053);
nor U40964 (N_40964,N_39503,N_39377);
and U40965 (N_40965,N_39628,N_39701);
xor U40966 (N_40966,N_39193,N_39126);
nor U40967 (N_40967,N_39109,N_39114);
and U40968 (N_40968,N_39043,N_39696);
nor U40969 (N_40969,N_39586,N_39229);
nand U40970 (N_40970,N_39025,N_39394);
nand U40971 (N_40971,N_39121,N_39672);
nor U40972 (N_40972,N_39898,N_39630);
xnor U40973 (N_40973,N_39697,N_39761);
xor U40974 (N_40974,N_39465,N_39364);
and U40975 (N_40975,N_39652,N_39746);
nor U40976 (N_40976,N_39123,N_39630);
or U40977 (N_40977,N_39058,N_39507);
nand U40978 (N_40978,N_39739,N_39843);
and U40979 (N_40979,N_39566,N_39932);
nand U40980 (N_40980,N_39694,N_39422);
or U40981 (N_40981,N_39927,N_39512);
xor U40982 (N_40982,N_39374,N_39999);
xnor U40983 (N_40983,N_39367,N_39193);
nor U40984 (N_40984,N_39618,N_39649);
nor U40985 (N_40985,N_39932,N_39936);
or U40986 (N_40986,N_39957,N_39529);
or U40987 (N_40987,N_39152,N_39927);
nor U40988 (N_40988,N_39513,N_39860);
xor U40989 (N_40989,N_39566,N_39467);
nor U40990 (N_40990,N_39950,N_39300);
or U40991 (N_40991,N_39535,N_39118);
or U40992 (N_40992,N_39365,N_39845);
nor U40993 (N_40993,N_39559,N_39435);
nand U40994 (N_40994,N_39338,N_39508);
and U40995 (N_40995,N_39908,N_39637);
and U40996 (N_40996,N_39396,N_39442);
xor U40997 (N_40997,N_39233,N_39939);
nand U40998 (N_40998,N_39660,N_39320);
xnor U40999 (N_40999,N_39899,N_39297);
or U41000 (N_41000,N_40785,N_40010);
and U41001 (N_41001,N_40444,N_40170);
nor U41002 (N_41002,N_40939,N_40161);
and U41003 (N_41003,N_40841,N_40833);
and U41004 (N_41004,N_40539,N_40373);
or U41005 (N_41005,N_40307,N_40320);
xnor U41006 (N_41006,N_40817,N_40204);
xnor U41007 (N_41007,N_40150,N_40225);
and U41008 (N_41008,N_40366,N_40583);
or U41009 (N_41009,N_40657,N_40134);
nand U41010 (N_41010,N_40387,N_40547);
and U41011 (N_41011,N_40753,N_40760);
and U41012 (N_41012,N_40698,N_40358);
xor U41013 (N_41013,N_40850,N_40523);
nor U41014 (N_41014,N_40035,N_40721);
or U41015 (N_41015,N_40432,N_40412);
xor U41016 (N_41016,N_40233,N_40506);
or U41017 (N_41017,N_40559,N_40402);
and U41018 (N_41018,N_40864,N_40232);
or U41019 (N_41019,N_40828,N_40933);
xnor U41020 (N_41020,N_40812,N_40878);
and U41021 (N_41021,N_40025,N_40143);
nand U41022 (N_41022,N_40857,N_40778);
or U41023 (N_41023,N_40991,N_40574);
xor U41024 (N_41024,N_40069,N_40431);
nor U41025 (N_41025,N_40199,N_40997);
or U41026 (N_41026,N_40724,N_40228);
or U41027 (N_41027,N_40052,N_40784);
or U41028 (N_41028,N_40490,N_40832);
nor U41029 (N_41029,N_40231,N_40931);
xor U41030 (N_41030,N_40118,N_40382);
nand U41031 (N_41031,N_40397,N_40588);
nand U41032 (N_41032,N_40208,N_40972);
or U41033 (N_41033,N_40398,N_40461);
and U41034 (N_41034,N_40867,N_40889);
xnor U41035 (N_41035,N_40486,N_40517);
nand U41036 (N_41036,N_40745,N_40219);
and U41037 (N_41037,N_40028,N_40562);
nand U41038 (N_41038,N_40108,N_40148);
nand U41039 (N_41039,N_40942,N_40755);
nor U41040 (N_41040,N_40827,N_40625);
nand U41041 (N_41041,N_40503,N_40576);
and U41042 (N_41042,N_40502,N_40626);
or U41043 (N_41043,N_40835,N_40883);
xnor U41044 (N_41044,N_40314,N_40280);
xnor U41045 (N_41045,N_40844,N_40239);
nand U41046 (N_41046,N_40141,N_40904);
and U41047 (N_41047,N_40560,N_40212);
nor U41048 (N_41048,N_40943,N_40317);
or U41049 (N_41049,N_40075,N_40121);
nor U41050 (N_41050,N_40369,N_40874);
or U41051 (N_41051,N_40650,N_40473);
nand U41052 (N_41052,N_40282,N_40123);
nand U41053 (N_41053,N_40954,N_40762);
nand U41054 (N_41054,N_40306,N_40554);
nand U41055 (N_41055,N_40303,N_40852);
or U41056 (N_41056,N_40663,N_40532);
xor U41057 (N_41057,N_40132,N_40862);
xor U41058 (N_41058,N_40460,N_40405);
and U41059 (N_41059,N_40315,N_40816);
nand U41060 (N_41060,N_40815,N_40185);
nor U41061 (N_41061,N_40799,N_40484);
xnor U41062 (N_41062,N_40428,N_40088);
and U41063 (N_41063,N_40814,N_40423);
nand U41064 (N_41064,N_40795,N_40806);
nand U41065 (N_41065,N_40530,N_40772);
nor U41066 (N_41066,N_40377,N_40313);
nand U41067 (N_41067,N_40858,N_40868);
xnor U41068 (N_41068,N_40359,N_40528);
or U41069 (N_41069,N_40468,N_40579);
and U41070 (N_41070,N_40585,N_40009);
xor U41071 (N_41071,N_40736,N_40617);
xnor U41072 (N_41072,N_40916,N_40876);
and U41073 (N_41073,N_40129,N_40362);
nor U41074 (N_41074,N_40008,N_40630);
nor U41075 (N_41075,N_40986,N_40634);
xnor U41076 (N_41076,N_40341,N_40122);
and U41077 (N_41077,N_40016,N_40589);
or U41078 (N_41078,N_40743,N_40462);
nand U41079 (N_41079,N_40384,N_40356);
xor U41080 (N_41080,N_40826,N_40352);
and U41081 (N_41081,N_40168,N_40869);
xnor U41082 (N_41082,N_40422,N_40598);
and U41083 (N_41083,N_40913,N_40558);
xor U41084 (N_41084,N_40919,N_40987);
or U41085 (N_41085,N_40408,N_40443);
or U41086 (N_41086,N_40990,N_40970);
nand U41087 (N_41087,N_40304,N_40037);
nor U41088 (N_41088,N_40266,N_40284);
nand U41089 (N_41089,N_40770,N_40066);
or U41090 (N_41090,N_40151,N_40848);
or U41091 (N_41091,N_40995,N_40071);
or U41092 (N_41092,N_40810,N_40363);
xor U41093 (N_41093,N_40768,N_40985);
xnor U41094 (N_41094,N_40636,N_40386);
xnor U41095 (N_41095,N_40555,N_40556);
xnor U41096 (N_41096,N_40774,N_40701);
and U41097 (N_41097,N_40205,N_40156);
nand U41098 (N_41098,N_40163,N_40251);
xnor U41099 (N_41099,N_40569,N_40209);
nand U41100 (N_41100,N_40514,N_40116);
and U41101 (N_41101,N_40090,N_40063);
and U41102 (N_41102,N_40808,N_40064);
and U41103 (N_41103,N_40800,N_40409);
xor U41104 (N_41104,N_40780,N_40566);
xnor U41105 (N_41105,N_40181,N_40087);
nor U41106 (N_41106,N_40061,N_40334);
xor U41107 (N_41107,N_40323,N_40477);
nand U41108 (N_41108,N_40710,N_40880);
or U41109 (N_41109,N_40550,N_40279);
nand U41110 (N_41110,N_40689,N_40048);
or U41111 (N_41111,N_40714,N_40411);
and U41112 (N_41112,N_40330,N_40081);
xnor U41113 (N_41113,N_40746,N_40045);
nor U41114 (N_41114,N_40012,N_40975);
nand U41115 (N_41115,N_40082,N_40407);
and U41116 (N_41116,N_40096,N_40716);
nand U41117 (N_41117,N_40672,N_40343);
nor U41118 (N_41118,N_40637,N_40103);
nand U41119 (N_41119,N_40024,N_40529);
nor U41120 (N_41120,N_40115,N_40447);
nand U41121 (N_41121,N_40038,N_40573);
or U41122 (N_41122,N_40624,N_40659);
xnor U41123 (N_41123,N_40840,N_40979);
or U41124 (N_41124,N_40202,N_40821);
nor U41125 (N_41125,N_40178,N_40699);
nor U41126 (N_41126,N_40033,N_40182);
nand U41127 (N_41127,N_40922,N_40452);
nand U41128 (N_41128,N_40142,N_40733);
and U41129 (N_41129,N_40434,N_40516);
xnor U41130 (N_41130,N_40830,N_40571);
or U41131 (N_41131,N_40929,N_40507);
nor U41132 (N_41132,N_40807,N_40882);
and U41133 (N_41133,N_40581,N_40060);
and U41134 (N_41134,N_40145,N_40348);
nand U41135 (N_41135,N_40759,N_40368);
or U41136 (N_41136,N_40458,N_40819);
xnor U41137 (N_41137,N_40504,N_40091);
xor U41138 (N_41138,N_40053,N_40195);
xnor U41139 (N_41139,N_40522,N_40027);
nor U41140 (N_41140,N_40109,N_40645);
nand U41141 (N_41141,N_40898,N_40180);
nand U41142 (N_41142,N_40691,N_40842);
xnor U41143 (N_41143,N_40793,N_40139);
and U41144 (N_41144,N_40325,N_40511);
nor U41145 (N_41145,N_40544,N_40453);
nor U41146 (N_41146,N_40921,N_40633);
and U41147 (N_41147,N_40597,N_40247);
or U41148 (N_41148,N_40336,N_40809);
nor U41149 (N_41149,N_40958,N_40196);
or U41150 (N_41150,N_40305,N_40289);
nand U41151 (N_41151,N_40584,N_40160);
xor U41152 (N_41152,N_40338,N_40272);
nand U41153 (N_41153,N_40962,N_40687);
nand U41154 (N_41154,N_40870,N_40321);
and U41155 (N_41155,N_40273,N_40354);
or U41156 (N_41156,N_40041,N_40927);
nand U41157 (N_41157,N_40189,N_40527);
nor U41158 (N_41158,N_40102,N_40389);
and U41159 (N_41159,N_40283,N_40892);
or U41160 (N_41160,N_40641,N_40437);
nand U41161 (N_41161,N_40073,N_40946);
nor U41162 (N_41162,N_40187,N_40183);
or U41163 (N_41163,N_40992,N_40393);
nor U41164 (N_41164,N_40104,N_40934);
nor U41165 (N_41165,N_40909,N_40744);
nor U41166 (N_41166,N_40619,N_40474);
xnor U41167 (N_41167,N_40899,N_40254);
xor U41168 (N_41168,N_40007,N_40629);
or U41169 (N_41169,N_40243,N_40798);
nand U41170 (N_41170,N_40551,N_40157);
nor U41171 (N_41171,N_40312,N_40639);
nor U41172 (N_41172,N_40615,N_40030);
or U41173 (N_41173,N_40476,N_40302);
nand U41174 (N_41174,N_40964,N_40895);
or U41175 (N_41175,N_40329,N_40153);
or U41176 (N_41176,N_40955,N_40824);
or U41177 (N_41177,N_40738,N_40531);
and U41178 (N_41178,N_40385,N_40847);
nor U41179 (N_41179,N_40250,N_40885);
nand U41180 (N_41180,N_40241,N_40335);
nor U41181 (N_41181,N_40860,N_40059);
xnor U41182 (N_41182,N_40996,N_40519);
nor U41183 (N_41183,N_40133,N_40940);
nor U41184 (N_41184,N_40649,N_40553);
nand U41185 (N_41185,N_40968,N_40427);
nor U41186 (N_41186,N_40238,N_40752);
nand U41187 (N_41187,N_40074,N_40717);
nor U41188 (N_41188,N_40999,N_40804);
nor U41189 (N_41189,N_40601,N_40072);
nor U41190 (N_41190,N_40667,N_40119);
xnor U41191 (N_41191,N_40740,N_40177);
xor U41192 (N_41192,N_40246,N_40342);
nand U41193 (N_41193,N_40011,N_40548);
nand U41194 (N_41194,N_40983,N_40401);
nor U41195 (N_41195,N_40887,N_40891);
and U41196 (N_41196,N_40686,N_40269);
and U41197 (N_41197,N_40570,N_40612);
nor U41198 (N_41198,N_40318,N_40230);
nand U41199 (N_41199,N_40498,N_40879);
nor U41200 (N_41200,N_40062,N_40166);
xnor U41201 (N_41201,N_40974,N_40781);
xnor U41202 (N_41202,N_40322,N_40831);
nand U41203 (N_41203,N_40274,N_40252);
or U41204 (N_41204,N_40056,N_40608);
and U41205 (N_41205,N_40897,N_40789);
nand U41206 (N_41206,N_40413,N_40920);
xor U41207 (N_41207,N_40677,N_40614);
nor U41208 (N_41208,N_40355,N_40101);
or U41209 (N_41209,N_40357,N_40154);
nor U41210 (N_41210,N_40005,N_40396);
or U41211 (N_41211,N_40813,N_40478);
or U41212 (N_41212,N_40515,N_40100);
and U41213 (N_41213,N_40333,N_40543);
xor U41214 (N_41214,N_40855,N_40894);
or U41215 (N_41215,N_40068,N_40644);
or U41216 (N_41216,N_40167,N_40327);
nand U41217 (N_41217,N_40802,N_40026);
or U41218 (N_41218,N_40747,N_40711);
xor U41219 (N_41219,N_40656,N_40803);
xor U41220 (N_41220,N_40552,N_40094);
nand U41221 (N_41221,N_40372,N_40492);
and U41222 (N_41222,N_40928,N_40537);
xor U41223 (N_41223,N_40620,N_40877);
and U41224 (N_41224,N_40905,N_40300);
xor U41225 (N_41225,N_40521,N_40337);
and U41226 (N_41226,N_40915,N_40345);
xnor U41227 (N_41227,N_40147,N_40399);
and U41228 (N_41228,N_40198,N_40930);
xnor U41229 (N_41229,N_40705,N_40594);
nand U41230 (N_41230,N_40932,N_40582);
or U41231 (N_41231,N_40077,N_40192);
nand U41232 (N_41232,N_40875,N_40445);
nand U41233 (N_41233,N_40339,N_40797);
nor U41234 (N_41234,N_40114,N_40169);
nor U41235 (N_41235,N_40264,N_40741);
nand U41236 (N_41236,N_40380,N_40410);
and U41237 (N_41237,N_40859,N_40281);
xor U41238 (N_41238,N_40414,N_40046);
or U41239 (N_41239,N_40873,N_40051);
nor U41240 (N_41240,N_40765,N_40678);
nor U41241 (N_41241,N_40456,N_40117);
nand U41242 (N_41242,N_40568,N_40349);
and U41243 (N_41243,N_40001,N_40015);
nor U41244 (N_41244,N_40839,N_40378);
or U41245 (N_41245,N_40771,N_40896);
nor U41246 (N_41246,N_40846,N_40646);
and U41247 (N_41247,N_40618,N_40376);
nor U41248 (N_41248,N_40949,N_40790);
nor U41249 (N_41249,N_40065,N_40777);
xnor U41250 (N_41250,N_40144,N_40076);
and U41251 (N_41251,N_40311,N_40863);
nand U41252 (N_41252,N_40365,N_40188);
or U41253 (N_41253,N_40638,N_40956);
or U41254 (N_41254,N_40725,N_40600);
xnor U41255 (N_41255,N_40165,N_40079);
nand U41256 (N_41256,N_40006,N_40497);
xor U41257 (N_41257,N_40957,N_40845);
xnor U41258 (N_41258,N_40483,N_40912);
nand U41259 (N_41259,N_40206,N_40660);
xor U41260 (N_41260,N_40487,N_40057);
xor U41261 (N_41261,N_40328,N_40702);
nor U41262 (N_41262,N_40331,N_40494);
or U41263 (N_41263,N_40695,N_40734);
nand U41264 (N_41264,N_40655,N_40666);
or U41265 (N_41265,N_40587,N_40018);
and U41266 (N_41266,N_40764,N_40856);
or U41267 (N_41267,N_40671,N_40379);
or U41268 (N_41268,N_40351,N_40616);
nand U41269 (N_41269,N_40207,N_40332);
or U41270 (N_41270,N_40610,N_40316);
nand U41271 (N_41271,N_40938,N_40261);
and U41272 (N_41272,N_40713,N_40464);
nand U41273 (N_41273,N_40174,N_40567);
xor U41274 (N_41274,N_40276,N_40155);
nand U41275 (N_41275,N_40640,N_40977);
and U41276 (N_41276,N_40124,N_40766);
and U41277 (N_41277,N_40643,N_40715);
nand U41278 (N_41278,N_40682,N_40164);
or U41279 (N_41279,N_40138,N_40093);
nand U41280 (N_41280,N_40361,N_40112);
xor U41281 (N_41281,N_40805,N_40838);
nor U41282 (N_41282,N_40843,N_40684);
or U41283 (N_41283,N_40210,N_40286);
xor U41284 (N_41284,N_40299,N_40936);
and U41285 (N_41285,N_40203,N_40392);
nor U41286 (N_41286,N_40110,N_40425);
nand U41287 (N_41287,N_40673,N_40240);
and U41288 (N_41288,N_40439,N_40287);
nor U41289 (N_41289,N_40888,N_40265);
or U41290 (N_41290,N_40245,N_40084);
xnor U41291 (N_41291,N_40665,N_40820);
nor U41292 (N_41292,N_40326,N_40495);
nand U41293 (N_41293,N_40267,N_40653);
and U41294 (N_41294,N_40963,N_40647);
and U41295 (N_41295,N_40095,N_40099);
xor U41296 (N_41296,N_40149,N_40395);
nand U41297 (N_41297,N_40706,N_40535);
nor U41298 (N_41298,N_40602,N_40757);
nor U41299 (N_41299,N_40125,N_40186);
xor U41300 (N_41300,N_40262,N_40500);
xnor U41301 (N_41301,N_40089,N_40466);
and U41302 (N_41302,N_40222,N_40036);
xnor U41303 (N_41303,N_40541,N_40034);
xnor U41304 (N_41304,N_40324,N_40982);
or U41305 (N_41305,N_40236,N_40690);
nand U41306 (N_41306,N_40669,N_40903);
or U41307 (N_41307,N_40923,N_40749);
and U41308 (N_41308,N_40175,N_40967);
or U41309 (N_41309,N_40591,N_40989);
nor U41310 (N_41310,N_40849,N_40438);
xnor U41311 (N_41311,N_40998,N_40390);
or U41312 (N_41312,N_40201,N_40911);
xnor U41313 (N_41313,N_40295,N_40463);
xnor U41314 (N_41314,N_40216,N_40910);
and U41315 (N_41315,N_40621,N_40501);
xnor U41316 (N_41316,N_40694,N_40563);
or U41317 (N_41317,N_40811,N_40049);
and U41318 (N_41318,N_40127,N_40491);
nor U41319 (N_41319,N_40421,N_40436);
nor U41320 (N_41320,N_40249,N_40681);
nand U41321 (N_41321,N_40945,N_40596);
nor U41322 (N_41322,N_40459,N_40966);
nor U41323 (N_41323,N_40680,N_40586);
or U41324 (N_41324,N_40263,N_40538);
nor U41325 (N_41325,N_40416,N_40851);
nor U41326 (N_41326,N_40173,N_40561);
and U41327 (N_41327,N_40572,N_40176);
nand U41328 (N_41328,N_40426,N_40465);
nor U41329 (N_41329,N_40661,N_40993);
xnor U41330 (N_41330,N_40244,N_40914);
and U41331 (N_41331,N_40190,N_40105);
or U41332 (N_41332,N_40592,N_40722);
xnor U41333 (N_41333,N_40769,N_40773);
and U41334 (N_41334,N_40854,N_40391);
xor U41335 (N_41335,N_40235,N_40257);
nand U41336 (N_41336,N_40723,N_40424);
nor U41337 (N_41337,N_40685,N_40603);
nor U41338 (N_41338,N_40374,N_40294);
and U41339 (N_41339,N_40924,N_40613);
and U41340 (N_41340,N_40525,N_40679);
nor U41341 (N_41341,N_40131,N_40120);
and U41342 (N_41342,N_40978,N_40524);
nand U41343 (N_41343,N_40253,N_40788);
xnor U41344 (N_41344,N_40260,N_40042);
or U41345 (N_41345,N_40215,N_40783);
and U41346 (N_41346,N_40482,N_40834);
nand U41347 (N_41347,N_40013,N_40433);
xor U41348 (N_41348,N_40505,N_40435);
xnor U41349 (N_41349,N_40727,N_40092);
xor U41350 (N_41350,N_40418,N_40565);
nor U41351 (N_41351,N_40900,N_40292);
nor U41352 (N_41352,N_40980,N_40350);
xnor U41353 (N_41353,N_40836,N_40111);
xor U41354 (N_41354,N_40726,N_40308);
and U41355 (N_41355,N_40575,N_40298);
and U41356 (N_41356,N_40627,N_40906);
xor U41357 (N_41357,N_40782,N_40775);
and U41358 (N_41358,N_40429,N_40730);
and U41359 (N_41359,N_40526,N_40837);
nand U41360 (N_41360,N_40578,N_40654);
nand U41361 (N_41361,N_40622,N_40184);
xnor U41362 (N_41362,N_40440,N_40002);
nor U41363 (N_41363,N_40632,N_40213);
nand U41364 (N_41364,N_40381,N_40595);
nand U41365 (N_41365,N_40031,N_40590);
or U41366 (N_41366,N_40748,N_40277);
and U41367 (N_41367,N_40676,N_40004);
nor U41368 (N_41368,N_40022,N_40128);
and U41369 (N_41369,N_40017,N_40969);
and U41370 (N_41370,N_40224,N_40564);
nand U41371 (N_41371,N_40536,N_40137);
nand U41372 (N_41372,N_40703,N_40750);
nand U41373 (N_41373,N_40960,N_40364);
xor U41374 (N_41374,N_40829,N_40309);
nand U41375 (N_41375,N_40822,N_40540);
nor U41376 (N_41376,N_40794,N_40097);
nand U41377 (N_41377,N_40388,N_40475);
xnor U41378 (N_41378,N_40040,N_40021);
or U41379 (N_41379,N_40448,N_40683);
nand U41380 (N_41380,N_40512,N_40605);
and U41381 (N_41381,N_40193,N_40801);
or U41382 (N_41382,N_40607,N_40948);
xnor U41383 (N_41383,N_40712,N_40179);
xor U41384 (N_41384,N_40787,N_40126);
nand U41385 (N_41385,N_40344,N_40080);
or U41386 (N_41386,N_40481,N_40054);
nor U41387 (N_41387,N_40729,N_40973);
nor U41388 (N_41388,N_40454,N_40696);
xor U41389 (N_41389,N_40796,N_40083);
nor U41390 (N_41390,N_40200,N_40234);
and U41391 (N_41391,N_40893,N_40020);
nor U41392 (N_41392,N_40107,N_40908);
nand U41393 (N_41393,N_40499,N_40085);
and U41394 (N_41394,N_40420,N_40242);
xor U41395 (N_41395,N_40709,N_40533);
nand U41396 (N_41396,N_40670,N_40197);
nor U41397 (N_41397,N_40606,N_40078);
and U41398 (N_41398,N_40394,N_40296);
or U41399 (N_41399,N_40098,N_40278);
nand U41400 (N_41400,N_40707,N_40375);
nand U41401 (N_41401,N_40951,N_40662);
nor U41402 (N_41402,N_40140,N_40223);
nand U41403 (N_41403,N_40471,N_40965);
and U41404 (N_41404,N_40470,N_40546);
nand U41405 (N_41405,N_40791,N_40518);
or U41406 (N_41406,N_40545,N_40767);
or U41407 (N_41407,N_40886,N_40952);
or U41408 (N_41408,N_40872,N_40367);
nor U41409 (N_41409,N_40675,N_40430);
nor U41410 (N_41410,N_40229,N_40902);
or U41411 (N_41411,N_40534,N_40510);
and U41412 (N_41412,N_40070,N_40731);
nor U41413 (N_41413,N_40728,N_40441);
and U41414 (N_41414,N_40959,N_40258);
or U41415 (N_41415,N_40971,N_40704);
nor U41416 (N_41416,N_40214,N_40248);
xor U41417 (N_41417,N_40668,N_40457);
nand U41418 (N_41418,N_40310,N_40158);
nand U41419 (N_41419,N_40635,N_40937);
nand U41420 (N_41420,N_40029,N_40086);
nor U41421 (N_41421,N_40818,N_40981);
nor U41422 (N_41422,N_40271,N_40370);
or U41423 (N_41423,N_40135,N_40000);
and U41424 (N_41424,N_40623,N_40693);
xor U41425 (N_41425,N_40146,N_40628);
or U41426 (N_41426,N_40754,N_40479);
xor U41427 (N_41427,N_40419,N_40043);
or U41428 (N_41428,N_40211,N_40651);
and U41429 (N_41429,N_40648,N_40944);
nor U41430 (N_41430,N_40019,N_40050);
nor U41431 (N_41431,N_40925,N_40631);
nand U41432 (N_41432,N_40067,N_40270);
or U41433 (N_41433,N_40493,N_40058);
nand U41434 (N_41434,N_40871,N_40226);
nor U41435 (N_41435,N_40918,N_40599);
nand U41436 (N_41436,N_40935,N_40756);
and U41437 (N_41437,N_40488,N_40988);
nand U41438 (N_41438,N_40218,N_40917);
or U41439 (N_41439,N_40984,N_40301);
and U41440 (N_41440,N_40268,N_40825);
nand U41441 (N_41441,N_40901,N_40737);
or U41442 (N_41442,N_40947,N_40580);
or U41443 (N_41443,N_40881,N_40792);
and U41444 (N_41444,N_40823,N_40346);
and U41445 (N_41445,N_40865,N_40758);
nand U41446 (N_41446,N_40604,N_40285);
or U41447 (N_41447,N_40130,N_40542);
nand U41448 (N_41448,N_40941,N_40255);
and U41449 (N_41449,N_40557,N_40469);
nor U41450 (N_41450,N_40417,N_40776);
nor U41451 (N_41451,N_40489,N_40761);
nor U41452 (N_41452,N_40159,N_40735);
and U41453 (N_41453,N_40191,N_40220);
and U41454 (N_41454,N_40288,N_40861);
or U41455 (N_41455,N_40853,N_40513);
xor U41456 (N_41456,N_40472,N_40194);
xor U41457 (N_41457,N_40319,N_40976);
nor U41458 (N_41458,N_40446,N_40779);
and U41459 (N_41459,N_40496,N_40485);
xor U41460 (N_41460,N_40742,N_40577);
xnor U41461 (N_41461,N_40259,N_40652);
nand U41462 (N_41462,N_40047,N_40450);
or U41463 (N_41463,N_40113,N_40961);
or U41464 (N_41464,N_40039,N_40720);
nor U41465 (N_41465,N_40926,N_40297);
xor U41466 (N_41466,N_40275,N_40032);
and U41467 (N_41467,N_40014,N_40293);
nor U41468 (N_41468,N_40044,N_40291);
or U41469 (N_41469,N_40611,N_40953);
xnor U41470 (N_41470,N_40415,N_40593);
xnor U41471 (N_41471,N_40371,N_40347);
or U41472 (N_41472,N_40340,N_40674);
and U41473 (N_41473,N_40403,N_40406);
xnor U41474 (N_41474,N_40136,N_40509);
or U41475 (N_41475,N_40383,N_40162);
nor U41476 (N_41476,N_40688,N_40106);
xor U41477 (N_41477,N_40451,N_40055);
and U41478 (N_41478,N_40023,N_40697);
and U41479 (N_41479,N_40890,N_40290);
nor U41480 (N_41480,N_40449,N_40467);
nand U41481 (N_41481,N_40152,N_40786);
xnor U41482 (N_41482,N_40763,N_40549);
nor U41483 (N_41483,N_40480,N_40609);
nor U41484 (N_41484,N_40719,N_40664);
and U41485 (N_41485,N_40884,N_40256);
nand U41486 (N_41486,N_40732,N_40950);
or U41487 (N_41487,N_40237,N_40172);
nand U41488 (N_41488,N_40718,N_40708);
xnor U41489 (N_41489,N_40400,N_40994);
or U41490 (N_41490,N_40227,N_40360);
or U41491 (N_41491,N_40751,N_40642);
nor U41492 (N_41492,N_40739,N_40455);
or U41493 (N_41493,N_40866,N_40907);
nor U41494 (N_41494,N_40700,N_40520);
nor U41495 (N_41495,N_40692,N_40658);
xnor U41496 (N_41496,N_40171,N_40353);
and U41497 (N_41497,N_40508,N_40003);
xor U41498 (N_41498,N_40404,N_40442);
xnor U41499 (N_41499,N_40221,N_40217);
xor U41500 (N_41500,N_40350,N_40783);
nand U41501 (N_41501,N_40905,N_40971);
nand U41502 (N_41502,N_40002,N_40660);
nor U41503 (N_41503,N_40939,N_40865);
or U41504 (N_41504,N_40658,N_40753);
xnor U41505 (N_41505,N_40180,N_40233);
nand U41506 (N_41506,N_40884,N_40192);
nand U41507 (N_41507,N_40247,N_40086);
and U41508 (N_41508,N_40730,N_40243);
nand U41509 (N_41509,N_40577,N_40233);
and U41510 (N_41510,N_40732,N_40631);
xnor U41511 (N_41511,N_40377,N_40203);
nor U41512 (N_41512,N_40636,N_40814);
and U41513 (N_41513,N_40620,N_40258);
and U41514 (N_41514,N_40594,N_40843);
nor U41515 (N_41515,N_40366,N_40530);
nor U41516 (N_41516,N_40720,N_40707);
nor U41517 (N_41517,N_40911,N_40378);
and U41518 (N_41518,N_40460,N_40698);
nand U41519 (N_41519,N_40763,N_40433);
xor U41520 (N_41520,N_40919,N_40349);
or U41521 (N_41521,N_40278,N_40378);
xor U41522 (N_41522,N_40217,N_40250);
nand U41523 (N_41523,N_40506,N_40686);
xnor U41524 (N_41524,N_40619,N_40888);
and U41525 (N_41525,N_40651,N_40312);
nand U41526 (N_41526,N_40035,N_40982);
nor U41527 (N_41527,N_40231,N_40631);
or U41528 (N_41528,N_40190,N_40125);
xnor U41529 (N_41529,N_40805,N_40799);
nand U41530 (N_41530,N_40280,N_40888);
xor U41531 (N_41531,N_40000,N_40129);
nand U41532 (N_41532,N_40920,N_40645);
or U41533 (N_41533,N_40282,N_40280);
xor U41534 (N_41534,N_40449,N_40127);
or U41535 (N_41535,N_40031,N_40847);
xnor U41536 (N_41536,N_40069,N_40288);
or U41537 (N_41537,N_40697,N_40048);
xnor U41538 (N_41538,N_40137,N_40884);
nand U41539 (N_41539,N_40392,N_40913);
nand U41540 (N_41540,N_40148,N_40397);
nor U41541 (N_41541,N_40683,N_40297);
xnor U41542 (N_41542,N_40100,N_40880);
nand U41543 (N_41543,N_40991,N_40815);
xnor U41544 (N_41544,N_40494,N_40611);
nor U41545 (N_41545,N_40201,N_40894);
nand U41546 (N_41546,N_40578,N_40554);
and U41547 (N_41547,N_40894,N_40390);
xor U41548 (N_41548,N_40518,N_40554);
nor U41549 (N_41549,N_40095,N_40303);
and U41550 (N_41550,N_40451,N_40416);
xor U41551 (N_41551,N_40091,N_40361);
and U41552 (N_41552,N_40845,N_40097);
and U41553 (N_41553,N_40112,N_40075);
or U41554 (N_41554,N_40394,N_40430);
xor U41555 (N_41555,N_40183,N_40076);
nand U41556 (N_41556,N_40936,N_40061);
nor U41557 (N_41557,N_40803,N_40634);
and U41558 (N_41558,N_40248,N_40413);
or U41559 (N_41559,N_40133,N_40691);
xor U41560 (N_41560,N_40630,N_40445);
or U41561 (N_41561,N_40807,N_40078);
or U41562 (N_41562,N_40376,N_40303);
xor U41563 (N_41563,N_40707,N_40059);
or U41564 (N_41564,N_40778,N_40134);
and U41565 (N_41565,N_40267,N_40678);
and U41566 (N_41566,N_40846,N_40987);
nor U41567 (N_41567,N_40744,N_40010);
nor U41568 (N_41568,N_40246,N_40799);
or U41569 (N_41569,N_40746,N_40878);
or U41570 (N_41570,N_40987,N_40724);
nand U41571 (N_41571,N_40498,N_40713);
or U41572 (N_41572,N_40811,N_40611);
xor U41573 (N_41573,N_40792,N_40317);
nand U41574 (N_41574,N_40133,N_40277);
or U41575 (N_41575,N_40709,N_40731);
nand U41576 (N_41576,N_40279,N_40638);
and U41577 (N_41577,N_40897,N_40667);
nand U41578 (N_41578,N_40581,N_40659);
or U41579 (N_41579,N_40147,N_40023);
xnor U41580 (N_41580,N_40501,N_40379);
or U41581 (N_41581,N_40200,N_40873);
and U41582 (N_41582,N_40205,N_40384);
or U41583 (N_41583,N_40581,N_40450);
xor U41584 (N_41584,N_40866,N_40821);
xor U41585 (N_41585,N_40719,N_40645);
xnor U41586 (N_41586,N_40998,N_40827);
and U41587 (N_41587,N_40895,N_40040);
nor U41588 (N_41588,N_40006,N_40829);
and U41589 (N_41589,N_40388,N_40681);
and U41590 (N_41590,N_40662,N_40128);
or U41591 (N_41591,N_40392,N_40905);
nand U41592 (N_41592,N_40548,N_40426);
and U41593 (N_41593,N_40283,N_40551);
nand U41594 (N_41594,N_40444,N_40782);
xnor U41595 (N_41595,N_40194,N_40314);
xnor U41596 (N_41596,N_40429,N_40347);
nand U41597 (N_41597,N_40571,N_40304);
nor U41598 (N_41598,N_40258,N_40397);
or U41599 (N_41599,N_40365,N_40190);
nand U41600 (N_41600,N_40214,N_40068);
nand U41601 (N_41601,N_40056,N_40524);
nand U41602 (N_41602,N_40108,N_40316);
nor U41603 (N_41603,N_40964,N_40764);
nor U41604 (N_41604,N_40869,N_40661);
nor U41605 (N_41605,N_40949,N_40226);
and U41606 (N_41606,N_40304,N_40978);
nor U41607 (N_41607,N_40042,N_40962);
and U41608 (N_41608,N_40252,N_40714);
or U41609 (N_41609,N_40701,N_40244);
nand U41610 (N_41610,N_40604,N_40660);
xnor U41611 (N_41611,N_40985,N_40049);
xnor U41612 (N_41612,N_40595,N_40253);
or U41613 (N_41613,N_40010,N_40759);
nand U41614 (N_41614,N_40488,N_40342);
nand U41615 (N_41615,N_40678,N_40009);
xor U41616 (N_41616,N_40744,N_40992);
and U41617 (N_41617,N_40225,N_40432);
or U41618 (N_41618,N_40210,N_40216);
nand U41619 (N_41619,N_40108,N_40930);
nor U41620 (N_41620,N_40157,N_40329);
nand U41621 (N_41621,N_40530,N_40589);
and U41622 (N_41622,N_40650,N_40242);
xor U41623 (N_41623,N_40770,N_40619);
nor U41624 (N_41624,N_40155,N_40160);
xnor U41625 (N_41625,N_40675,N_40637);
nand U41626 (N_41626,N_40024,N_40816);
and U41627 (N_41627,N_40802,N_40998);
nor U41628 (N_41628,N_40649,N_40300);
and U41629 (N_41629,N_40328,N_40648);
xnor U41630 (N_41630,N_40482,N_40801);
nand U41631 (N_41631,N_40741,N_40795);
and U41632 (N_41632,N_40438,N_40319);
nor U41633 (N_41633,N_40143,N_40912);
or U41634 (N_41634,N_40279,N_40191);
and U41635 (N_41635,N_40236,N_40881);
xor U41636 (N_41636,N_40734,N_40366);
and U41637 (N_41637,N_40435,N_40661);
or U41638 (N_41638,N_40022,N_40284);
and U41639 (N_41639,N_40202,N_40506);
and U41640 (N_41640,N_40561,N_40514);
or U41641 (N_41641,N_40150,N_40882);
or U41642 (N_41642,N_40028,N_40775);
xor U41643 (N_41643,N_40907,N_40346);
or U41644 (N_41644,N_40681,N_40591);
nand U41645 (N_41645,N_40159,N_40247);
or U41646 (N_41646,N_40594,N_40120);
and U41647 (N_41647,N_40880,N_40218);
or U41648 (N_41648,N_40782,N_40931);
nor U41649 (N_41649,N_40246,N_40174);
and U41650 (N_41650,N_40248,N_40616);
nor U41651 (N_41651,N_40196,N_40514);
and U41652 (N_41652,N_40554,N_40566);
and U41653 (N_41653,N_40598,N_40087);
nor U41654 (N_41654,N_40309,N_40787);
nor U41655 (N_41655,N_40693,N_40139);
nand U41656 (N_41656,N_40338,N_40946);
nand U41657 (N_41657,N_40953,N_40886);
nand U41658 (N_41658,N_40499,N_40563);
and U41659 (N_41659,N_40965,N_40777);
and U41660 (N_41660,N_40440,N_40327);
nor U41661 (N_41661,N_40297,N_40566);
nor U41662 (N_41662,N_40081,N_40486);
or U41663 (N_41663,N_40373,N_40086);
xnor U41664 (N_41664,N_40750,N_40049);
or U41665 (N_41665,N_40792,N_40937);
or U41666 (N_41666,N_40407,N_40406);
xnor U41667 (N_41667,N_40997,N_40648);
xor U41668 (N_41668,N_40985,N_40355);
or U41669 (N_41669,N_40713,N_40443);
and U41670 (N_41670,N_40579,N_40788);
nand U41671 (N_41671,N_40444,N_40651);
nor U41672 (N_41672,N_40893,N_40357);
and U41673 (N_41673,N_40067,N_40015);
or U41674 (N_41674,N_40106,N_40582);
nor U41675 (N_41675,N_40951,N_40085);
nand U41676 (N_41676,N_40575,N_40761);
xnor U41677 (N_41677,N_40804,N_40340);
nand U41678 (N_41678,N_40399,N_40639);
xor U41679 (N_41679,N_40293,N_40677);
and U41680 (N_41680,N_40819,N_40616);
xor U41681 (N_41681,N_40138,N_40892);
and U41682 (N_41682,N_40641,N_40441);
or U41683 (N_41683,N_40617,N_40349);
or U41684 (N_41684,N_40898,N_40912);
nand U41685 (N_41685,N_40452,N_40695);
nor U41686 (N_41686,N_40620,N_40004);
nor U41687 (N_41687,N_40735,N_40639);
xor U41688 (N_41688,N_40563,N_40605);
and U41689 (N_41689,N_40328,N_40744);
and U41690 (N_41690,N_40062,N_40177);
or U41691 (N_41691,N_40932,N_40282);
or U41692 (N_41692,N_40946,N_40348);
or U41693 (N_41693,N_40035,N_40610);
nand U41694 (N_41694,N_40532,N_40496);
nand U41695 (N_41695,N_40744,N_40190);
xor U41696 (N_41696,N_40165,N_40923);
and U41697 (N_41697,N_40249,N_40513);
and U41698 (N_41698,N_40981,N_40780);
and U41699 (N_41699,N_40124,N_40853);
or U41700 (N_41700,N_40292,N_40604);
and U41701 (N_41701,N_40997,N_40240);
xor U41702 (N_41702,N_40390,N_40119);
or U41703 (N_41703,N_40507,N_40301);
or U41704 (N_41704,N_40671,N_40433);
nor U41705 (N_41705,N_40649,N_40416);
xnor U41706 (N_41706,N_40010,N_40100);
and U41707 (N_41707,N_40256,N_40800);
or U41708 (N_41708,N_40254,N_40468);
nand U41709 (N_41709,N_40469,N_40844);
or U41710 (N_41710,N_40024,N_40231);
nand U41711 (N_41711,N_40738,N_40870);
and U41712 (N_41712,N_40529,N_40100);
xnor U41713 (N_41713,N_40740,N_40020);
nor U41714 (N_41714,N_40279,N_40778);
nand U41715 (N_41715,N_40060,N_40585);
nor U41716 (N_41716,N_40738,N_40211);
and U41717 (N_41717,N_40099,N_40852);
nor U41718 (N_41718,N_40345,N_40557);
nor U41719 (N_41719,N_40657,N_40229);
xor U41720 (N_41720,N_40993,N_40674);
and U41721 (N_41721,N_40565,N_40636);
or U41722 (N_41722,N_40069,N_40180);
nand U41723 (N_41723,N_40644,N_40591);
xnor U41724 (N_41724,N_40505,N_40785);
nand U41725 (N_41725,N_40477,N_40288);
xnor U41726 (N_41726,N_40451,N_40526);
xor U41727 (N_41727,N_40630,N_40944);
and U41728 (N_41728,N_40093,N_40789);
or U41729 (N_41729,N_40400,N_40048);
xor U41730 (N_41730,N_40105,N_40882);
or U41731 (N_41731,N_40770,N_40700);
nand U41732 (N_41732,N_40369,N_40287);
nand U41733 (N_41733,N_40526,N_40890);
nand U41734 (N_41734,N_40160,N_40473);
xnor U41735 (N_41735,N_40983,N_40294);
nor U41736 (N_41736,N_40161,N_40713);
nand U41737 (N_41737,N_40970,N_40422);
and U41738 (N_41738,N_40136,N_40518);
and U41739 (N_41739,N_40727,N_40135);
and U41740 (N_41740,N_40296,N_40680);
or U41741 (N_41741,N_40119,N_40724);
nor U41742 (N_41742,N_40340,N_40978);
or U41743 (N_41743,N_40267,N_40658);
and U41744 (N_41744,N_40061,N_40105);
and U41745 (N_41745,N_40394,N_40513);
nand U41746 (N_41746,N_40193,N_40304);
xnor U41747 (N_41747,N_40441,N_40367);
nand U41748 (N_41748,N_40891,N_40201);
xor U41749 (N_41749,N_40121,N_40062);
xor U41750 (N_41750,N_40247,N_40514);
and U41751 (N_41751,N_40200,N_40381);
xor U41752 (N_41752,N_40620,N_40164);
and U41753 (N_41753,N_40271,N_40501);
or U41754 (N_41754,N_40468,N_40685);
or U41755 (N_41755,N_40937,N_40351);
xor U41756 (N_41756,N_40798,N_40119);
and U41757 (N_41757,N_40912,N_40348);
and U41758 (N_41758,N_40906,N_40246);
and U41759 (N_41759,N_40388,N_40595);
and U41760 (N_41760,N_40056,N_40068);
nand U41761 (N_41761,N_40673,N_40965);
nor U41762 (N_41762,N_40848,N_40649);
nor U41763 (N_41763,N_40314,N_40477);
xnor U41764 (N_41764,N_40563,N_40578);
or U41765 (N_41765,N_40453,N_40858);
xnor U41766 (N_41766,N_40258,N_40666);
nor U41767 (N_41767,N_40992,N_40713);
and U41768 (N_41768,N_40931,N_40412);
xor U41769 (N_41769,N_40417,N_40393);
nand U41770 (N_41770,N_40138,N_40356);
and U41771 (N_41771,N_40490,N_40140);
nand U41772 (N_41772,N_40409,N_40555);
or U41773 (N_41773,N_40415,N_40606);
nor U41774 (N_41774,N_40110,N_40218);
nand U41775 (N_41775,N_40010,N_40863);
nand U41776 (N_41776,N_40440,N_40008);
nand U41777 (N_41777,N_40402,N_40035);
and U41778 (N_41778,N_40386,N_40207);
and U41779 (N_41779,N_40627,N_40401);
and U41780 (N_41780,N_40461,N_40959);
xor U41781 (N_41781,N_40089,N_40917);
nand U41782 (N_41782,N_40352,N_40012);
nor U41783 (N_41783,N_40785,N_40308);
nand U41784 (N_41784,N_40335,N_40833);
or U41785 (N_41785,N_40425,N_40775);
nand U41786 (N_41786,N_40694,N_40845);
nand U41787 (N_41787,N_40565,N_40639);
nor U41788 (N_41788,N_40211,N_40595);
and U41789 (N_41789,N_40439,N_40897);
nor U41790 (N_41790,N_40656,N_40117);
xnor U41791 (N_41791,N_40352,N_40036);
nand U41792 (N_41792,N_40940,N_40648);
xnor U41793 (N_41793,N_40446,N_40600);
nor U41794 (N_41794,N_40729,N_40811);
xor U41795 (N_41795,N_40278,N_40074);
or U41796 (N_41796,N_40601,N_40781);
and U41797 (N_41797,N_40994,N_40581);
nand U41798 (N_41798,N_40363,N_40122);
and U41799 (N_41799,N_40917,N_40144);
nor U41800 (N_41800,N_40147,N_40865);
xor U41801 (N_41801,N_40499,N_40756);
nand U41802 (N_41802,N_40972,N_40836);
and U41803 (N_41803,N_40604,N_40099);
or U41804 (N_41804,N_40266,N_40406);
or U41805 (N_41805,N_40850,N_40769);
xor U41806 (N_41806,N_40600,N_40704);
nor U41807 (N_41807,N_40637,N_40173);
xnor U41808 (N_41808,N_40968,N_40413);
and U41809 (N_41809,N_40572,N_40427);
and U41810 (N_41810,N_40741,N_40737);
nand U41811 (N_41811,N_40172,N_40440);
nand U41812 (N_41812,N_40162,N_40960);
xnor U41813 (N_41813,N_40771,N_40104);
nor U41814 (N_41814,N_40759,N_40787);
or U41815 (N_41815,N_40900,N_40007);
xnor U41816 (N_41816,N_40789,N_40182);
nand U41817 (N_41817,N_40410,N_40810);
or U41818 (N_41818,N_40261,N_40880);
nor U41819 (N_41819,N_40066,N_40247);
or U41820 (N_41820,N_40926,N_40527);
and U41821 (N_41821,N_40897,N_40233);
and U41822 (N_41822,N_40488,N_40578);
nor U41823 (N_41823,N_40204,N_40779);
nor U41824 (N_41824,N_40675,N_40655);
and U41825 (N_41825,N_40918,N_40436);
xor U41826 (N_41826,N_40414,N_40784);
and U41827 (N_41827,N_40129,N_40777);
xnor U41828 (N_41828,N_40141,N_40444);
nand U41829 (N_41829,N_40177,N_40259);
and U41830 (N_41830,N_40518,N_40707);
and U41831 (N_41831,N_40997,N_40399);
nand U41832 (N_41832,N_40151,N_40194);
and U41833 (N_41833,N_40952,N_40019);
nand U41834 (N_41834,N_40842,N_40757);
nand U41835 (N_41835,N_40135,N_40028);
nor U41836 (N_41836,N_40387,N_40602);
or U41837 (N_41837,N_40491,N_40992);
nand U41838 (N_41838,N_40849,N_40299);
and U41839 (N_41839,N_40984,N_40798);
and U41840 (N_41840,N_40917,N_40568);
xor U41841 (N_41841,N_40480,N_40315);
or U41842 (N_41842,N_40651,N_40755);
nand U41843 (N_41843,N_40656,N_40725);
xnor U41844 (N_41844,N_40817,N_40220);
nor U41845 (N_41845,N_40335,N_40897);
nand U41846 (N_41846,N_40853,N_40286);
nor U41847 (N_41847,N_40578,N_40631);
nor U41848 (N_41848,N_40955,N_40832);
nand U41849 (N_41849,N_40514,N_40893);
xnor U41850 (N_41850,N_40363,N_40513);
nand U41851 (N_41851,N_40664,N_40942);
or U41852 (N_41852,N_40951,N_40579);
xor U41853 (N_41853,N_40898,N_40361);
or U41854 (N_41854,N_40141,N_40537);
nor U41855 (N_41855,N_40003,N_40371);
xor U41856 (N_41856,N_40381,N_40776);
or U41857 (N_41857,N_40179,N_40226);
or U41858 (N_41858,N_40750,N_40339);
xnor U41859 (N_41859,N_40410,N_40553);
nor U41860 (N_41860,N_40602,N_40144);
nor U41861 (N_41861,N_40773,N_40852);
nand U41862 (N_41862,N_40512,N_40931);
nand U41863 (N_41863,N_40989,N_40308);
or U41864 (N_41864,N_40352,N_40730);
xnor U41865 (N_41865,N_40958,N_40761);
and U41866 (N_41866,N_40838,N_40694);
or U41867 (N_41867,N_40176,N_40817);
xnor U41868 (N_41868,N_40269,N_40293);
or U41869 (N_41869,N_40825,N_40442);
or U41870 (N_41870,N_40790,N_40002);
xor U41871 (N_41871,N_40184,N_40400);
nor U41872 (N_41872,N_40735,N_40391);
xnor U41873 (N_41873,N_40356,N_40543);
and U41874 (N_41874,N_40108,N_40565);
or U41875 (N_41875,N_40547,N_40651);
or U41876 (N_41876,N_40660,N_40066);
and U41877 (N_41877,N_40799,N_40563);
and U41878 (N_41878,N_40273,N_40836);
and U41879 (N_41879,N_40847,N_40452);
or U41880 (N_41880,N_40480,N_40289);
nor U41881 (N_41881,N_40077,N_40135);
and U41882 (N_41882,N_40509,N_40790);
xnor U41883 (N_41883,N_40959,N_40912);
xor U41884 (N_41884,N_40529,N_40211);
nor U41885 (N_41885,N_40373,N_40635);
nand U41886 (N_41886,N_40947,N_40744);
nor U41887 (N_41887,N_40855,N_40729);
nand U41888 (N_41888,N_40928,N_40345);
xor U41889 (N_41889,N_40816,N_40813);
or U41890 (N_41890,N_40321,N_40386);
xnor U41891 (N_41891,N_40442,N_40890);
or U41892 (N_41892,N_40332,N_40368);
nor U41893 (N_41893,N_40938,N_40561);
or U41894 (N_41894,N_40832,N_40472);
nand U41895 (N_41895,N_40231,N_40396);
nor U41896 (N_41896,N_40890,N_40456);
xnor U41897 (N_41897,N_40620,N_40475);
xnor U41898 (N_41898,N_40571,N_40945);
or U41899 (N_41899,N_40703,N_40402);
xnor U41900 (N_41900,N_40665,N_40088);
and U41901 (N_41901,N_40539,N_40450);
xnor U41902 (N_41902,N_40874,N_40813);
nor U41903 (N_41903,N_40614,N_40753);
and U41904 (N_41904,N_40551,N_40293);
xnor U41905 (N_41905,N_40321,N_40559);
xnor U41906 (N_41906,N_40904,N_40791);
nor U41907 (N_41907,N_40940,N_40543);
or U41908 (N_41908,N_40089,N_40036);
and U41909 (N_41909,N_40630,N_40932);
nor U41910 (N_41910,N_40822,N_40414);
and U41911 (N_41911,N_40488,N_40144);
nand U41912 (N_41912,N_40587,N_40562);
nand U41913 (N_41913,N_40016,N_40097);
nand U41914 (N_41914,N_40677,N_40839);
or U41915 (N_41915,N_40053,N_40843);
nor U41916 (N_41916,N_40564,N_40362);
nand U41917 (N_41917,N_40703,N_40456);
and U41918 (N_41918,N_40479,N_40182);
nor U41919 (N_41919,N_40847,N_40007);
xnor U41920 (N_41920,N_40900,N_40793);
or U41921 (N_41921,N_40059,N_40789);
nand U41922 (N_41922,N_40120,N_40225);
and U41923 (N_41923,N_40621,N_40881);
and U41924 (N_41924,N_40799,N_40088);
nor U41925 (N_41925,N_40743,N_40009);
nand U41926 (N_41926,N_40390,N_40519);
nor U41927 (N_41927,N_40500,N_40167);
nand U41928 (N_41928,N_40002,N_40283);
nor U41929 (N_41929,N_40446,N_40755);
xor U41930 (N_41930,N_40786,N_40675);
xor U41931 (N_41931,N_40902,N_40235);
or U41932 (N_41932,N_40408,N_40466);
xnor U41933 (N_41933,N_40052,N_40057);
or U41934 (N_41934,N_40370,N_40358);
or U41935 (N_41935,N_40166,N_40945);
nor U41936 (N_41936,N_40346,N_40249);
nand U41937 (N_41937,N_40685,N_40381);
xor U41938 (N_41938,N_40698,N_40580);
nand U41939 (N_41939,N_40056,N_40520);
and U41940 (N_41940,N_40438,N_40901);
nand U41941 (N_41941,N_40620,N_40122);
nor U41942 (N_41942,N_40635,N_40774);
and U41943 (N_41943,N_40818,N_40978);
or U41944 (N_41944,N_40732,N_40786);
or U41945 (N_41945,N_40602,N_40458);
and U41946 (N_41946,N_40392,N_40338);
xor U41947 (N_41947,N_40668,N_40734);
and U41948 (N_41948,N_40946,N_40435);
nand U41949 (N_41949,N_40220,N_40153);
xnor U41950 (N_41950,N_40167,N_40495);
or U41951 (N_41951,N_40775,N_40266);
nor U41952 (N_41952,N_40927,N_40567);
xor U41953 (N_41953,N_40158,N_40611);
xor U41954 (N_41954,N_40176,N_40976);
xnor U41955 (N_41955,N_40271,N_40260);
or U41956 (N_41956,N_40495,N_40294);
nand U41957 (N_41957,N_40979,N_40916);
or U41958 (N_41958,N_40892,N_40846);
and U41959 (N_41959,N_40930,N_40245);
nand U41960 (N_41960,N_40062,N_40482);
nand U41961 (N_41961,N_40474,N_40061);
or U41962 (N_41962,N_40887,N_40200);
and U41963 (N_41963,N_40550,N_40000);
or U41964 (N_41964,N_40348,N_40312);
nor U41965 (N_41965,N_40814,N_40978);
xnor U41966 (N_41966,N_40503,N_40578);
or U41967 (N_41967,N_40796,N_40711);
or U41968 (N_41968,N_40100,N_40026);
xnor U41969 (N_41969,N_40736,N_40786);
and U41970 (N_41970,N_40828,N_40782);
xor U41971 (N_41971,N_40396,N_40252);
or U41972 (N_41972,N_40426,N_40185);
nand U41973 (N_41973,N_40060,N_40386);
and U41974 (N_41974,N_40053,N_40065);
nor U41975 (N_41975,N_40639,N_40977);
or U41976 (N_41976,N_40869,N_40716);
nor U41977 (N_41977,N_40236,N_40943);
nand U41978 (N_41978,N_40492,N_40453);
nor U41979 (N_41979,N_40811,N_40778);
xor U41980 (N_41980,N_40070,N_40901);
nor U41981 (N_41981,N_40121,N_40307);
or U41982 (N_41982,N_40163,N_40801);
xor U41983 (N_41983,N_40418,N_40608);
xor U41984 (N_41984,N_40774,N_40256);
or U41985 (N_41985,N_40787,N_40937);
and U41986 (N_41986,N_40395,N_40958);
or U41987 (N_41987,N_40805,N_40090);
nor U41988 (N_41988,N_40591,N_40599);
xor U41989 (N_41989,N_40074,N_40404);
nand U41990 (N_41990,N_40331,N_40472);
and U41991 (N_41991,N_40418,N_40458);
xor U41992 (N_41992,N_40111,N_40259);
and U41993 (N_41993,N_40339,N_40247);
and U41994 (N_41994,N_40567,N_40145);
or U41995 (N_41995,N_40673,N_40599);
nand U41996 (N_41996,N_40989,N_40045);
and U41997 (N_41997,N_40040,N_40990);
xor U41998 (N_41998,N_40875,N_40690);
or U41999 (N_41999,N_40255,N_40850);
xnor U42000 (N_42000,N_41495,N_41794);
or U42001 (N_42001,N_41944,N_41526);
and U42002 (N_42002,N_41324,N_41383);
xnor U42003 (N_42003,N_41965,N_41616);
nand U42004 (N_42004,N_41350,N_41121);
xnor U42005 (N_42005,N_41893,N_41129);
xnor U42006 (N_42006,N_41870,N_41068);
or U42007 (N_42007,N_41499,N_41478);
or U42008 (N_42008,N_41813,N_41020);
or U42009 (N_42009,N_41030,N_41178);
or U42010 (N_42010,N_41697,N_41017);
and U42011 (N_42011,N_41329,N_41958);
nor U42012 (N_42012,N_41467,N_41149);
or U42013 (N_42013,N_41942,N_41130);
and U42014 (N_42014,N_41554,N_41483);
nand U42015 (N_42015,N_41657,N_41821);
xnor U42016 (N_42016,N_41994,N_41216);
nand U42017 (N_42017,N_41161,N_41909);
nand U42018 (N_42018,N_41079,N_41264);
nand U42019 (N_42019,N_41168,N_41112);
nor U42020 (N_42020,N_41640,N_41023);
or U42021 (N_42021,N_41583,N_41285);
xor U42022 (N_42022,N_41096,N_41947);
or U42023 (N_42023,N_41214,N_41408);
xnor U42024 (N_42024,N_41425,N_41533);
nor U42025 (N_42025,N_41781,N_41065);
and U42026 (N_42026,N_41253,N_41557);
nand U42027 (N_42027,N_41160,N_41268);
xnor U42028 (N_42028,N_41798,N_41258);
and U42029 (N_42029,N_41931,N_41793);
xnor U42030 (N_42030,N_41566,N_41035);
or U42031 (N_42031,N_41341,N_41036);
nand U42032 (N_42032,N_41191,N_41379);
xnor U42033 (N_42033,N_41703,N_41937);
and U42034 (N_42034,N_41126,N_41935);
nand U42035 (N_42035,N_41818,N_41704);
nor U42036 (N_42036,N_41599,N_41570);
xor U42037 (N_42037,N_41820,N_41580);
nor U42038 (N_42038,N_41282,N_41915);
nor U42039 (N_42039,N_41644,N_41155);
xnor U42040 (N_42040,N_41122,N_41418);
or U42041 (N_42041,N_41680,N_41267);
xor U42042 (N_42042,N_41313,N_41249);
nand U42043 (N_42043,N_41359,N_41104);
nor U42044 (N_42044,N_41838,N_41535);
xnor U42045 (N_42045,N_41611,N_41349);
nor U42046 (N_42046,N_41770,N_41028);
and U42047 (N_42047,N_41466,N_41945);
and U42048 (N_42048,N_41801,N_41338);
or U42049 (N_42049,N_41992,N_41360);
and U42050 (N_42050,N_41627,N_41345);
xor U42051 (N_42051,N_41973,N_41077);
xnor U42052 (N_42052,N_41560,N_41142);
or U42053 (N_42053,N_41508,N_41118);
or U42054 (N_42054,N_41553,N_41760);
and U42055 (N_42055,N_41853,N_41825);
xnor U42056 (N_42056,N_41783,N_41343);
and U42057 (N_42057,N_41854,N_41391);
xor U42058 (N_42058,N_41691,N_41746);
nand U42059 (N_42059,N_41876,N_41990);
nor U42060 (N_42060,N_41731,N_41806);
nor U42061 (N_42061,N_41624,N_41366);
or U42062 (N_42062,N_41940,N_41843);
or U42063 (N_42063,N_41355,N_41339);
and U42064 (N_42064,N_41320,N_41445);
xor U42065 (N_42065,N_41153,N_41358);
xnor U42066 (N_42066,N_41658,N_41518);
or U42067 (N_42067,N_41710,N_41219);
xor U42068 (N_42068,N_41163,N_41974);
nand U42069 (N_42069,N_41397,N_41812);
nand U42070 (N_42070,N_41913,N_41110);
nand U42071 (N_42071,N_41986,N_41503);
or U42072 (N_42072,N_41674,N_41239);
or U42073 (N_42073,N_41089,N_41552);
nor U42074 (N_42074,N_41098,N_41735);
or U42075 (N_42075,N_41486,N_41026);
and U42076 (N_42076,N_41839,N_41524);
nand U42077 (N_42077,N_41449,N_41882);
or U42078 (N_42078,N_41493,N_41582);
nand U42079 (N_42079,N_41227,N_41659);
nor U42080 (N_42080,N_41435,N_41759);
nor U42081 (N_42081,N_41861,N_41701);
xor U42082 (N_42082,N_41137,N_41771);
xnor U42083 (N_42083,N_41021,N_41747);
or U42084 (N_42084,N_41632,N_41978);
and U42085 (N_42085,N_41459,N_41082);
nor U42086 (N_42086,N_41594,N_41862);
nor U42087 (N_42087,N_41590,N_41544);
xor U42088 (N_42088,N_41167,N_41979);
xor U42089 (N_42089,N_41361,N_41591);
nand U42090 (N_42090,N_41943,N_41393);
nand U42091 (N_42091,N_41502,N_41099);
nand U42092 (N_42092,N_41381,N_41846);
or U42093 (N_42093,N_41917,N_41673);
nand U42094 (N_42094,N_41421,N_41369);
xnor U42095 (N_42095,N_41817,N_41384);
nand U42096 (N_42096,N_41071,N_41884);
and U42097 (N_42097,N_41165,N_41936);
nor U42098 (N_42098,N_41215,N_41956);
xnor U42099 (N_42099,N_41631,N_41934);
or U42100 (N_42100,N_41795,N_41211);
nor U42101 (N_42101,N_41698,N_41728);
nand U42102 (N_42102,N_41787,N_41744);
nand U42103 (N_42103,N_41908,N_41724);
nand U42104 (N_42104,N_41709,N_41378);
nand U42105 (N_42105,N_41789,N_41038);
nand U42106 (N_42106,N_41683,N_41436);
and U42107 (N_42107,N_41173,N_41602);
xnor U42108 (N_42108,N_41629,N_41612);
or U42109 (N_42109,N_41070,N_41265);
or U42110 (N_42110,N_41233,N_41454);
or U42111 (N_42111,N_41625,N_41831);
nor U42112 (N_42112,N_41278,N_41274);
nor U42113 (N_42113,N_41133,N_41596);
or U42114 (N_42114,N_41891,N_41837);
xnor U42115 (N_42115,N_41729,N_41883);
or U42116 (N_42116,N_41567,N_41504);
nand U42117 (N_42117,N_41643,N_41573);
xnor U42118 (N_42118,N_41194,N_41323);
xor U42119 (N_42119,N_41392,N_41585);
or U42120 (N_42120,N_41808,N_41311);
or U42121 (N_42121,N_41456,N_41575);
nand U42122 (N_42122,N_41388,N_41604);
or U42123 (N_42123,N_41677,N_41881);
or U42124 (N_42124,N_41962,N_41321);
xor U42125 (N_42125,N_41540,N_41461);
and U42126 (N_42126,N_41353,N_41059);
xnor U42127 (N_42127,N_41765,N_41874);
or U42128 (N_42128,N_41957,N_41827);
and U42129 (N_42129,N_41308,N_41333);
nand U42130 (N_42130,N_41052,N_41492);
xnor U42131 (N_42131,N_41251,N_41772);
or U42132 (N_42132,N_41487,N_41911);
and U42133 (N_42133,N_41696,N_41042);
and U42134 (N_42134,N_41675,N_41548);
nand U42135 (N_42135,N_41715,N_41780);
or U42136 (N_42136,N_41334,N_41342);
nand U42137 (N_42137,N_41288,N_41754);
xor U42138 (N_42138,N_41745,N_41694);
and U42139 (N_42139,N_41272,N_41471);
or U42140 (N_42140,N_41901,N_41152);
nand U42141 (N_42141,N_41062,N_41100);
nor U42142 (N_42142,N_41287,N_41016);
nor U42143 (N_42143,N_41719,N_41046);
nor U42144 (N_42144,N_41234,N_41900);
nand U42145 (N_42145,N_41971,N_41564);
xor U42146 (N_42146,N_41791,N_41107);
xnor U42147 (N_42147,N_41725,N_41286);
and U42148 (N_42148,N_41245,N_41872);
xnor U42149 (N_42149,N_41409,N_41140);
and U42150 (N_42150,N_41444,N_41983);
nand U42151 (N_42151,N_41396,N_41182);
nand U42152 (N_42152,N_41574,N_41183);
or U42153 (N_42153,N_41693,N_41948);
or U42154 (N_42154,N_41921,N_41148);
and U42155 (N_42155,N_41664,N_41739);
or U42156 (N_42156,N_41006,N_41886);
or U42157 (N_42157,N_41880,N_41032);
xnor U42158 (N_42158,N_41143,N_41075);
nor U42159 (N_42159,N_41447,N_41097);
nor U42160 (N_42160,N_41768,N_41617);
xnor U42161 (N_42161,N_41555,N_41476);
or U42162 (N_42162,N_41919,N_41998);
xnor U42163 (N_42163,N_41738,N_41687);
or U42164 (N_42164,N_41316,N_41201);
or U42165 (N_42165,N_41231,N_41949);
or U42166 (N_42166,N_41225,N_41722);
and U42167 (N_42167,N_41465,N_41667);
nand U42168 (N_42168,N_41346,N_41755);
nand U42169 (N_42169,N_41815,N_41297);
nor U42170 (N_42170,N_41000,N_41666);
nor U42171 (N_42171,N_41022,N_41619);
or U42172 (N_42172,N_41576,N_41996);
xnor U42173 (N_42173,N_41377,N_41069);
nand U42174 (N_42174,N_41930,N_41312);
or U42175 (N_42175,N_41162,N_41690);
or U42176 (N_42176,N_41926,N_41198);
nand U42177 (N_42177,N_41967,N_41106);
xnor U42178 (N_42178,N_41423,N_41654);
xnor U42179 (N_42179,N_41189,N_41319);
nor U42180 (N_42180,N_41185,N_41115);
nor U42181 (N_42181,N_41105,N_41980);
and U42182 (N_42182,N_41601,N_41382);
nor U42183 (N_42183,N_41752,N_41792);
or U42184 (N_42184,N_41404,N_41330);
or U42185 (N_42185,N_41784,N_41174);
nor U42186 (N_42186,N_41048,N_41802);
xor U42187 (N_42187,N_41685,N_41261);
or U42188 (N_42188,N_41322,N_41761);
nand U42189 (N_42189,N_41788,N_41209);
and U42190 (N_42190,N_41850,N_41037);
and U42191 (N_42191,N_41141,N_41108);
and U42192 (N_42192,N_41428,N_41136);
and U42193 (N_42193,N_41277,N_41672);
and U42194 (N_42194,N_41623,N_41295);
nand U42195 (N_42195,N_41630,N_41542);
nand U42196 (N_42196,N_41208,N_41840);
nor U42197 (N_42197,N_41269,N_41117);
nand U42198 (N_42198,N_41205,N_41064);
nand U42199 (N_42199,N_41804,N_41426);
and U42200 (N_42200,N_41797,N_41844);
or U42201 (N_42201,N_41340,N_41531);
xnor U42202 (N_42202,N_41912,N_41712);
nand U42203 (N_42203,N_41733,N_41859);
nor U42204 (N_42204,N_41561,N_41955);
xor U42205 (N_42205,N_41448,N_41608);
or U42206 (N_42206,N_41109,N_41364);
nor U42207 (N_42207,N_41647,N_41475);
or U42208 (N_42208,N_41641,N_41520);
and U42209 (N_42209,N_41873,N_41635);
and U42210 (N_42210,N_41681,N_41088);
or U42211 (N_42211,N_41541,N_41488);
or U42212 (N_42212,N_41939,N_41145);
xnor U42213 (N_42213,N_41595,N_41250);
or U42214 (N_42214,N_41648,N_41529);
or U42215 (N_42215,N_41453,N_41362);
nand U42216 (N_42216,N_41634,N_41443);
and U42217 (N_42217,N_41519,N_41603);
nand U42218 (N_42218,N_41645,N_41695);
and U42219 (N_42219,N_41925,N_41777);
and U42220 (N_42220,N_41179,N_41546);
and U42221 (N_42221,N_41841,N_41197);
or U42222 (N_42222,N_41730,N_41609);
nor U42223 (N_42223,N_41462,N_41228);
and U42224 (N_42224,N_41757,N_41271);
or U42225 (N_42225,N_41014,N_41981);
or U42226 (N_42226,N_41906,N_41442);
nand U42227 (N_42227,N_41127,N_41828);
nor U42228 (N_42228,N_41663,N_41887);
nand U42229 (N_42229,N_41325,N_41440);
nor U42230 (N_42230,N_41896,N_41852);
nor U42231 (N_42231,N_41721,N_41385);
nand U42232 (N_42232,N_41816,N_41221);
and U42233 (N_42233,N_41004,N_41970);
nand U42234 (N_42234,N_41671,N_41417);
or U42235 (N_42235,N_41550,N_41232);
or U42236 (N_42236,N_41489,N_41434);
xnor U42237 (N_42237,N_41537,N_41424);
nor U42238 (N_42238,N_41318,N_41154);
xor U42239 (N_42239,N_41805,N_41705);
or U42240 (N_42240,N_41774,N_41276);
and U42241 (N_42241,N_41914,N_41003);
xor U42242 (N_42242,N_41008,N_41830);
and U42243 (N_42243,N_41933,N_41146);
nor U42244 (N_42244,N_41950,N_41598);
or U42245 (N_42245,N_41243,N_41241);
nand U42246 (N_42246,N_41438,N_41019);
and U42247 (N_42247,N_41995,N_41170);
nand U42248 (N_42248,N_41422,N_41063);
xnor U42249 (N_42249,N_41646,N_41199);
or U42250 (N_42250,N_41875,N_41164);
xnor U42251 (N_42251,N_41414,N_41090);
xnor U42252 (N_42252,N_41969,N_41545);
xor U42253 (N_42253,N_41707,N_41855);
xor U42254 (N_42254,N_41833,N_41336);
xnor U42255 (N_42255,N_41758,N_41002);
xnor U42256 (N_42256,N_41289,N_41354);
nand U42257 (N_42257,N_41651,N_41348);
nor U42258 (N_42258,N_41190,N_41015);
nand U42259 (N_42259,N_41718,N_41655);
or U42260 (N_42260,N_41702,N_41521);
xnor U42261 (N_42261,N_41051,N_41894);
and U42262 (N_42262,N_41558,N_41866);
nor U42263 (N_42263,N_41571,N_41281);
or U42264 (N_42264,N_41296,N_41773);
nor U42265 (N_42265,N_41670,N_41290);
and U42266 (N_42266,N_41387,N_41976);
and U42267 (N_42267,N_41776,N_41514);
and U42268 (N_42268,N_41723,N_41903);
nand U42269 (N_42269,N_41613,N_41073);
nand U42270 (N_42270,N_41280,N_41058);
xor U42271 (N_42271,N_41357,N_41522);
nor U42272 (N_42272,N_41748,N_41700);
or U42273 (N_42273,N_41736,N_41864);
xor U42274 (N_42274,N_41260,N_41551);
xor U42275 (N_42275,N_41890,N_41961);
and U42276 (N_42276,N_41351,N_41213);
xor U42277 (N_42277,N_41181,N_41605);
nand U42278 (N_42278,N_41224,N_41916);
or U42279 (N_42279,N_41223,N_41317);
nor U42280 (N_42280,N_41819,N_41033);
nand U42281 (N_42281,N_41229,N_41398);
xor U42282 (N_42282,N_41203,N_41653);
xor U42283 (N_42283,N_41867,N_41273);
and U42284 (N_42284,N_41158,N_41649);
nand U42285 (N_42285,N_41457,N_41547);
or U42286 (N_42286,N_41132,N_41041);
or U42287 (N_42287,N_41138,N_41468);
or U42288 (N_42288,N_41490,N_41084);
and U42289 (N_42289,N_41188,N_41885);
nand U42290 (N_42290,N_41898,N_41579);
xor U42291 (N_42291,N_41055,N_41991);
or U42292 (N_42292,N_41220,N_41530);
and U42293 (N_42293,N_41678,N_41309);
nor U42294 (N_42294,N_41403,N_41628);
or U42295 (N_42295,N_41202,N_41923);
and U42296 (N_42296,N_41863,N_41727);
nand U42297 (N_42297,N_41860,N_41217);
nor U42298 (N_42298,N_41186,N_41699);
nor U42299 (N_42299,N_41822,N_41266);
nor U42300 (N_42300,N_41650,N_41275);
xnor U42301 (N_42301,N_41834,N_41989);
xnor U42302 (N_42302,N_41218,N_41235);
or U42303 (N_42303,N_41686,N_41399);
and U42304 (N_42304,N_41907,N_41175);
or U42305 (N_42305,N_41169,N_41123);
xnor U42306 (N_42306,N_41512,N_41248);
or U42307 (N_42307,N_41389,N_41314);
nand U42308 (N_42308,N_41067,N_41714);
nor U42309 (N_42309,N_41257,N_41877);
nand U42310 (N_42310,N_41419,N_41741);
and U42311 (N_42311,N_41786,N_41928);
nand U42312 (N_42312,N_41993,N_41053);
xnor U42313 (N_42313,N_41606,N_41057);
nand U42314 (N_42314,N_41597,N_41195);
xnor U42315 (N_42315,N_41676,N_41386);
nand U42316 (N_42316,N_41256,N_41511);
or U42317 (N_42317,N_41543,N_41684);
and U42318 (N_42318,N_41826,N_41929);
or U42319 (N_42319,N_41299,N_41559);
or U42320 (N_42320,N_41525,N_41412);
nor U42321 (N_42321,N_41708,N_41011);
xnor U42322 (N_42322,N_41018,N_41706);
or U42323 (N_42323,N_41782,N_41103);
and U42324 (N_42324,N_41230,N_41614);
xor U42325 (N_42325,N_41306,N_41966);
nand U42326 (N_42326,N_41507,N_41865);
or U42327 (N_42327,N_41785,N_41124);
nor U42328 (N_42328,N_41013,N_41963);
and U42329 (N_42329,N_41135,N_41842);
nor U42330 (N_42330,N_41044,N_41307);
nand U42331 (N_42331,N_41892,N_41536);
nand U42332 (N_42332,N_41618,N_41607);
nor U42333 (N_42333,N_41086,N_41172);
nor U42334 (N_42334,N_41851,N_41402);
and U42335 (N_42335,N_41807,N_41331);
xor U42336 (N_42336,N_41610,N_41128);
nand U42337 (N_42337,N_41437,N_41473);
or U42338 (N_42338,N_41415,N_41577);
or U42339 (N_42339,N_41941,N_41439);
and U42340 (N_42340,N_41085,N_41156);
nand U42341 (N_42341,N_41458,N_41327);
xnor U42342 (N_42342,N_41572,N_41147);
nand U42343 (N_42343,N_41775,N_41193);
nor U42344 (N_42344,N_41455,N_41056);
xor U42345 (N_42345,N_41192,N_41588);
and U42346 (N_42346,N_41238,N_41661);
nor U42347 (N_42347,N_41120,N_41692);
and U42348 (N_42348,N_41380,N_41005);
or U42349 (N_42349,N_41938,N_41102);
xnor U42350 (N_42350,N_41332,N_41034);
or U42351 (N_42351,N_41868,N_41497);
xor U42352 (N_42352,N_41751,N_41593);
xor U42353 (N_42353,N_41997,N_41375);
and U42354 (N_42354,N_41074,N_41335);
nand U42355 (N_42355,N_41116,N_41410);
xnor U42356 (N_42356,N_41626,N_41637);
or U42357 (N_42357,N_41711,N_41113);
nor U42358 (N_42358,N_41263,N_41451);
nand U42359 (N_42359,N_41304,N_41960);
nand U42360 (N_42360,N_41592,N_41920);
or U42361 (N_42361,N_41226,N_41726);
nor U42362 (N_42362,N_41298,N_41857);
xor U42363 (N_42363,N_41095,N_41254);
nand U42364 (N_42364,N_41578,N_41762);
or U42365 (N_42365,N_41985,N_41420);
or U42366 (N_42366,N_41310,N_41569);
nand U42367 (N_42367,N_41328,N_41395);
and U42368 (N_42368,N_41049,N_41452);
xnor U42369 (N_42369,N_41878,N_41742);
xor U42370 (N_42370,N_41946,N_41959);
nor U42371 (N_42371,N_41469,N_41463);
nand U42372 (N_42372,N_41144,N_41480);
and U42373 (N_42373,N_41134,N_41713);
nor U42374 (N_42374,N_41356,N_41847);
or U42375 (N_42375,N_41769,N_41212);
nand U42376 (N_42376,N_41516,N_41433);
and U42377 (N_42377,N_41347,N_41427);
nand U42378 (N_42378,N_41363,N_41581);
xnor U42379 (N_42379,N_41157,N_41093);
or U42380 (N_42380,N_41888,N_41236);
nor U42381 (N_42381,N_41027,N_41092);
and U42382 (N_42382,N_41968,N_41600);
nand U42383 (N_42383,N_41045,N_41527);
nor U42384 (N_42384,N_41125,N_41244);
and U42385 (N_42385,N_41720,N_41829);
xnor U42386 (N_42386,N_41371,N_41688);
nand U42387 (N_42387,N_41464,N_41210);
nor U42388 (N_42388,N_41879,N_41301);
nor U42389 (N_42389,N_41897,N_41589);
nand U42390 (N_42390,N_41796,N_41679);
and U42391 (N_42391,N_41977,N_41528);
nor U42392 (N_42392,N_41753,N_41496);
or U42393 (N_42393,N_41491,N_41662);
nand U42394 (N_42394,N_41562,N_41639);
xnor U42395 (N_42395,N_41012,N_41368);
and U42396 (N_42396,N_41856,N_41450);
nor U42397 (N_42397,N_41622,N_41061);
nand U42398 (N_42398,N_41823,N_41344);
nand U42399 (N_42399,N_41902,N_41895);
nand U42400 (N_42400,N_41337,N_41506);
nor U42401 (N_42401,N_41087,N_41764);
nor U42402 (N_42402,N_41638,N_41665);
and U42403 (N_42403,N_41482,N_41252);
nor U42404 (N_42404,N_41066,N_41636);
nand U42405 (N_42405,N_41446,N_41689);
nor U42406 (N_42406,N_41766,N_41054);
nand U42407 (N_42407,N_41166,N_41501);
nor U42408 (N_42408,N_41171,N_41242);
xnor U42409 (N_42409,N_41740,N_41565);
nor U42410 (N_42410,N_41405,N_41204);
nor U42411 (N_42411,N_41119,N_41905);
nor U42412 (N_42412,N_41159,N_41050);
and U42413 (N_42413,N_41372,N_41932);
nor U42414 (N_42414,N_41401,N_41367);
or U42415 (N_42415,N_41656,N_41262);
xnor U42416 (N_42416,N_41407,N_41150);
or U42417 (N_42417,N_41951,N_41669);
nand U42418 (N_42418,N_41889,N_41539);
nor U42419 (N_42419,N_41294,N_41400);
xnor U42420 (N_42420,N_41799,N_41394);
and U42421 (N_42421,N_41176,N_41039);
and U42422 (N_42422,N_41767,N_41832);
nand U42423 (N_42423,N_41481,N_41431);
or U42424 (N_42424,N_41029,N_41479);
or U42425 (N_42425,N_41305,N_41984);
and U42426 (N_42426,N_41460,N_41472);
nor U42427 (N_42427,N_41682,N_41101);
and U42428 (N_42428,N_41899,N_41790);
nor U42429 (N_42429,N_41810,N_41432);
or U42430 (N_42430,N_41292,N_41568);
or U42431 (N_42431,N_41259,N_41836);
and U42432 (N_42432,N_41809,N_41081);
xor U42433 (N_42433,N_41009,N_41078);
nand U42434 (N_42434,N_41114,N_41513);
or U42435 (N_42435,N_41556,N_41352);
nor U42436 (N_42436,N_41953,N_41734);
nand U42437 (N_42437,N_41083,N_41534);
nor U42438 (N_42438,N_41811,N_41315);
and U42439 (N_42439,N_41982,N_41291);
or U42440 (N_42440,N_41184,N_41500);
nor U42441 (N_42441,N_41131,N_41177);
nand U42442 (N_42442,N_41494,N_41716);
and U42443 (N_42443,N_41279,N_41411);
and U42444 (N_42444,N_41376,N_41523);
nand U42445 (N_42445,N_41076,N_41633);
and U42446 (N_42446,N_41988,N_41302);
or U42447 (N_42447,N_41532,N_41918);
xor U42448 (N_42448,N_41749,N_41406);
or U42449 (N_42449,N_41848,N_41952);
xnor U42450 (N_42450,N_41779,N_41047);
xnor U42451 (N_42451,N_41660,N_41270);
xnor U42452 (N_42452,N_41756,N_41237);
xor U42453 (N_42453,N_41080,N_41668);
and U42454 (N_42454,N_41510,N_41975);
xor U42455 (N_42455,N_41835,N_41586);
or U42456 (N_42456,N_41470,N_41001);
and U42457 (N_42457,N_41743,N_41430);
nand U42458 (N_42458,N_41031,N_41007);
or U42459 (N_42459,N_41849,N_41927);
xor U42460 (N_42460,N_41326,N_41538);
or U42461 (N_42461,N_41365,N_41615);
or U42462 (N_42462,N_41222,N_41814);
or U42463 (N_42463,N_41111,N_41300);
nor U42464 (N_42464,N_41800,N_41498);
nand U42465 (N_42465,N_41924,N_41187);
nand U42466 (N_42466,N_41778,N_41416);
or U42467 (N_42467,N_41732,N_41010);
xnor U42468 (N_42468,N_41139,N_41206);
xnor U42469 (N_42469,N_41255,N_41858);
nand U42470 (N_42470,N_41374,N_41845);
xor U42471 (N_42471,N_41196,N_41485);
and U42472 (N_42472,N_41750,N_41441);
and U42473 (N_42473,N_41474,N_41025);
and U42474 (N_42474,N_41515,N_41390);
and U42475 (N_42475,N_41094,N_41517);
xnor U42476 (N_42476,N_41869,N_41207);
nor U42477 (N_42477,N_41043,N_41293);
or U42478 (N_42478,N_41151,N_41737);
or U42479 (N_42479,N_41987,N_41072);
xnor U42480 (N_42480,N_41284,N_41803);
or U42481 (N_42481,N_41240,N_41972);
xnor U42482 (N_42482,N_41373,N_41247);
nor U42483 (N_42483,N_41954,N_41040);
or U42484 (N_42484,N_41717,N_41091);
or U42485 (N_42485,N_41910,N_41587);
and U42486 (N_42486,N_41620,N_41824);
nor U42487 (N_42487,N_41642,N_41922);
nor U42488 (N_42488,N_41652,N_41549);
and U42489 (N_42489,N_41563,N_41477);
and U42490 (N_42490,N_41484,N_41584);
nand U42491 (N_42491,N_41246,N_41964);
xnor U42492 (N_42492,N_41283,N_41024);
nand U42493 (N_42493,N_41509,N_41429);
nor U42494 (N_42494,N_41370,N_41871);
nor U42495 (N_42495,N_41621,N_41763);
xor U42496 (N_42496,N_41060,N_41904);
nand U42497 (N_42497,N_41303,N_41505);
nor U42498 (N_42498,N_41413,N_41200);
nor U42499 (N_42499,N_41999,N_41180);
nor U42500 (N_42500,N_41426,N_41727);
xnor U42501 (N_42501,N_41542,N_41824);
nor U42502 (N_42502,N_41008,N_41875);
or U42503 (N_42503,N_41986,N_41379);
xnor U42504 (N_42504,N_41438,N_41025);
xor U42505 (N_42505,N_41077,N_41909);
nor U42506 (N_42506,N_41974,N_41060);
nor U42507 (N_42507,N_41517,N_41943);
or U42508 (N_42508,N_41758,N_41646);
nand U42509 (N_42509,N_41019,N_41585);
and U42510 (N_42510,N_41469,N_41363);
xor U42511 (N_42511,N_41676,N_41460);
nor U42512 (N_42512,N_41334,N_41654);
and U42513 (N_42513,N_41059,N_41551);
nand U42514 (N_42514,N_41878,N_41483);
or U42515 (N_42515,N_41379,N_41946);
and U42516 (N_42516,N_41186,N_41167);
and U42517 (N_42517,N_41677,N_41365);
or U42518 (N_42518,N_41402,N_41736);
and U42519 (N_42519,N_41762,N_41623);
and U42520 (N_42520,N_41932,N_41962);
nand U42521 (N_42521,N_41832,N_41308);
xnor U42522 (N_42522,N_41628,N_41738);
and U42523 (N_42523,N_41560,N_41112);
or U42524 (N_42524,N_41857,N_41909);
and U42525 (N_42525,N_41305,N_41951);
and U42526 (N_42526,N_41279,N_41889);
or U42527 (N_42527,N_41899,N_41266);
nand U42528 (N_42528,N_41652,N_41875);
or U42529 (N_42529,N_41742,N_41686);
xor U42530 (N_42530,N_41517,N_41889);
xor U42531 (N_42531,N_41692,N_41750);
xor U42532 (N_42532,N_41116,N_41696);
or U42533 (N_42533,N_41832,N_41361);
nor U42534 (N_42534,N_41468,N_41644);
and U42535 (N_42535,N_41507,N_41286);
or U42536 (N_42536,N_41607,N_41043);
nor U42537 (N_42537,N_41238,N_41613);
nor U42538 (N_42538,N_41042,N_41147);
or U42539 (N_42539,N_41833,N_41859);
or U42540 (N_42540,N_41492,N_41923);
nor U42541 (N_42541,N_41105,N_41359);
and U42542 (N_42542,N_41012,N_41229);
xnor U42543 (N_42543,N_41973,N_41489);
nor U42544 (N_42544,N_41019,N_41828);
nand U42545 (N_42545,N_41510,N_41106);
nand U42546 (N_42546,N_41012,N_41949);
and U42547 (N_42547,N_41367,N_41746);
and U42548 (N_42548,N_41115,N_41750);
or U42549 (N_42549,N_41117,N_41771);
and U42550 (N_42550,N_41694,N_41788);
or U42551 (N_42551,N_41793,N_41620);
xnor U42552 (N_42552,N_41494,N_41434);
and U42553 (N_42553,N_41603,N_41259);
nor U42554 (N_42554,N_41401,N_41974);
nor U42555 (N_42555,N_41927,N_41944);
nand U42556 (N_42556,N_41419,N_41779);
nand U42557 (N_42557,N_41774,N_41825);
or U42558 (N_42558,N_41303,N_41985);
and U42559 (N_42559,N_41292,N_41672);
xnor U42560 (N_42560,N_41007,N_41349);
nand U42561 (N_42561,N_41475,N_41222);
and U42562 (N_42562,N_41746,N_41888);
nand U42563 (N_42563,N_41356,N_41858);
nand U42564 (N_42564,N_41916,N_41550);
or U42565 (N_42565,N_41798,N_41651);
xor U42566 (N_42566,N_41719,N_41550);
xnor U42567 (N_42567,N_41191,N_41071);
and U42568 (N_42568,N_41526,N_41774);
xor U42569 (N_42569,N_41281,N_41644);
nand U42570 (N_42570,N_41726,N_41983);
nand U42571 (N_42571,N_41145,N_41943);
or U42572 (N_42572,N_41109,N_41925);
xnor U42573 (N_42573,N_41235,N_41600);
or U42574 (N_42574,N_41930,N_41240);
or U42575 (N_42575,N_41221,N_41247);
and U42576 (N_42576,N_41570,N_41987);
or U42577 (N_42577,N_41729,N_41357);
nand U42578 (N_42578,N_41999,N_41109);
xnor U42579 (N_42579,N_41025,N_41904);
xnor U42580 (N_42580,N_41847,N_41481);
or U42581 (N_42581,N_41883,N_41855);
nand U42582 (N_42582,N_41431,N_41050);
or U42583 (N_42583,N_41875,N_41039);
nand U42584 (N_42584,N_41822,N_41179);
xnor U42585 (N_42585,N_41867,N_41377);
nor U42586 (N_42586,N_41684,N_41282);
xor U42587 (N_42587,N_41140,N_41489);
and U42588 (N_42588,N_41742,N_41624);
xor U42589 (N_42589,N_41101,N_41869);
xnor U42590 (N_42590,N_41473,N_41852);
nor U42591 (N_42591,N_41315,N_41468);
nand U42592 (N_42592,N_41116,N_41603);
and U42593 (N_42593,N_41459,N_41206);
nor U42594 (N_42594,N_41156,N_41487);
nand U42595 (N_42595,N_41211,N_41387);
or U42596 (N_42596,N_41908,N_41464);
nor U42597 (N_42597,N_41217,N_41319);
and U42598 (N_42598,N_41584,N_41602);
xor U42599 (N_42599,N_41044,N_41112);
nand U42600 (N_42600,N_41924,N_41376);
xnor U42601 (N_42601,N_41825,N_41148);
nand U42602 (N_42602,N_41250,N_41355);
nand U42603 (N_42603,N_41354,N_41682);
nand U42604 (N_42604,N_41766,N_41725);
nor U42605 (N_42605,N_41159,N_41524);
xnor U42606 (N_42606,N_41862,N_41984);
xor U42607 (N_42607,N_41553,N_41868);
xor U42608 (N_42608,N_41672,N_41171);
and U42609 (N_42609,N_41890,N_41357);
xnor U42610 (N_42610,N_41938,N_41210);
nand U42611 (N_42611,N_41957,N_41208);
or U42612 (N_42612,N_41285,N_41061);
nand U42613 (N_42613,N_41069,N_41086);
and U42614 (N_42614,N_41957,N_41475);
and U42615 (N_42615,N_41976,N_41182);
and U42616 (N_42616,N_41397,N_41135);
or U42617 (N_42617,N_41901,N_41694);
nand U42618 (N_42618,N_41885,N_41769);
nand U42619 (N_42619,N_41357,N_41094);
nor U42620 (N_42620,N_41064,N_41699);
and U42621 (N_42621,N_41247,N_41631);
or U42622 (N_42622,N_41839,N_41732);
xnor U42623 (N_42623,N_41716,N_41871);
xor U42624 (N_42624,N_41870,N_41387);
or U42625 (N_42625,N_41253,N_41134);
nand U42626 (N_42626,N_41371,N_41801);
and U42627 (N_42627,N_41380,N_41925);
nor U42628 (N_42628,N_41346,N_41005);
nand U42629 (N_42629,N_41734,N_41442);
nor U42630 (N_42630,N_41848,N_41970);
and U42631 (N_42631,N_41750,N_41194);
nor U42632 (N_42632,N_41515,N_41916);
nand U42633 (N_42633,N_41093,N_41516);
and U42634 (N_42634,N_41743,N_41247);
or U42635 (N_42635,N_41228,N_41028);
nand U42636 (N_42636,N_41423,N_41551);
xor U42637 (N_42637,N_41036,N_41597);
xnor U42638 (N_42638,N_41883,N_41861);
and U42639 (N_42639,N_41811,N_41795);
nand U42640 (N_42640,N_41796,N_41208);
xor U42641 (N_42641,N_41969,N_41261);
and U42642 (N_42642,N_41835,N_41973);
xnor U42643 (N_42643,N_41612,N_41909);
or U42644 (N_42644,N_41328,N_41163);
xnor U42645 (N_42645,N_41994,N_41194);
nand U42646 (N_42646,N_41658,N_41774);
or U42647 (N_42647,N_41737,N_41419);
or U42648 (N_42648,N_41551,N_41211);
and U42649 (N_42649,N_41987,N_41004);
nand U42650 (N_42650,N_41335,N_41728);
xor U42651 (N_42651,N_41124,N_41237);
nor U42652 (N_42652,N_41452,N_41676);
xor U42653 (N_42653,N_41105,N_41375);
and U42654 (N_42654,N_41667,N_41171);
nor U42655 (N_42655,N_41109,N_41816);
nand U42656 (N_42656,N_41912,N_41366);
and U42657 (N_42657,N_41178,N_41569);
or U42658 (N_42658,N_41940,N_41670);
or U42659 (N_42659,N_41067,N_41815);
nor U42660 (N_42660,N_41850,N_41962);
and U42661 (N_42661,N_41849,N_41907);
or U42662 (N_42662,N_41082,N_41117);
nor U42663 (N_42663,N_41686,N_41612);
nor U42664 (N_42664,N_41864,N_41296);
xnor U42665 (N_42665,N_41921,N_41044);
and U42666 (N_42666,N_41382,N_41076);
or U42667 (N_42667,N_41143,N_41064);
nand U42668 (N_42668,N_41543,N_41437);
and U42669 (N_42669,N_41825,N_41107);
and U42670 (N_42670,N_41843,N_41172);
and U42671 (N_42671,N_41332,N_41848);
and U42672 (N_42672,N_41609,N_41528);
or U42673 (N_42673,N_41751,N_41865);
or U42674 (N_42674,N_41201,N_41225);
nor U42675 (N_42675,N_41387,N_41856);
nor U42676 (N_42676,N_41134,N_41248);
nor U42677 (N_42677,N_41326,N_41140);
and U42678 (N_42678,N_41973,N_41934);
xnor U42679 (N_42679,N_41228,N_41370);
xnor U42680 (N_42680,N_41310,N_41758);
or U42681 (N_42681,N_41575,N_41530);
xnor U42682 (N_42682,N_41004,N_41259);
nand U42683 (N_42683,N_41109,N_41827);
or U42684 (N_42684,N_41822,N_41188);
or U42685 (N_42685,N_41213,N_41431);
nand U42686 (N_42686,N_41204,N_41628);
and U42687 (N_42687,N_41154,N_41269);
and U42688 (N_42688,N_41652,N_41844);
xnor U42689 (N_42689,N_41957,N_41109);
or U42690 (N_42690,N_41870,N_41848);
xor U42691 (N_42691,N_41450,N_41654);
nand U42692 (N_42692,N_41765,N_41605);
nor U42693 (N_42693,N_41822,N_41129);
nand U42694 (N_42694,N_41672,N_41388);
nand U42695 (N_42695,N_41057,N_41952);
xnor U42696 (N_42696,N_41273,N_41511);
or U42697 (N_42697,N_41287,N_41059);
nand U42698 (N_42698,N_41702,N_41724);
and U42699 (N_42699,N_41154,N_41477);
nor U42700 (N_42700,N_41878,N_41956);
nand U42701 (N_42701,N_41200,N_41189);
nand U42702 (N_42702,N_41298,N_41947);
xnor U42703 (N_42703,N_41991,N_41544);
and U42704 (N_42704,N_41712,N_41335);
nor U42705 (N_42705,N_41189,N_41386);
and U42706 (N_42706,N_41893,N_41048);
or U42707 (N_42707,N_41400,N_41771);
and U42708 (N_42708,N_41611,N_41931);
and U42709 (N_42709,N_41412,N_41905);
nand U42710 (N_42710,N_41716,N_41984);
xor U42711 (N_42711,N_41277,N_41409);
and U42712 (N_42712,N_41238,N_41957);
nor U42713 (N_42713,N_41521,N_41610);
and U42714 (N_42714,N_41535,N_41645);
nor U42715 (N_42715,N_41250,N_41829);
xnor U42716 (N_42716,N_41557,N_41626);
and U42717 (N_42717,N_41230,N_41897);
or U42718 (N_42718,N_41869,N_41119);
xor U42719 (N_42719,N_41555,N_41093);
and U42720 (N_42720,N_41958,N_41742);
nand U42721 (N_42721,N_41377,N_41043);
nor U42722 (N_42722,N_41855,N_41854);
nand U42723 (N_42723,N_41741,N_41994);
nor U42724 (N_42724,N_41583,N_41024);
nor U42725 (N_42725,N_41758,N_41678);
or U42726 (N_42726,N_41023,N_41641);
nand U42727 (N_42727,N_41286,N_41732);
or U42728 (N_42728,N_41345,N_41364);
nor U42729 (N_42729,N_41252,N_41435);
nor U42730 (N_42730,N_41133,N_41208);
nand U42731 (N_42731,N_41391,N_41760);
xor U42732 (N_42732,N_41225,N_41315);
or U42733 (N_42733,N_41536,N_41329);
nor U42734 (N_42734,N_41764,N_41747);
and U42735 (N_42735,N_41176,N_41513);
and U42736 (N_42736,N_41171,N_41154);
or U42737 (N_42737,N_41231,N_41603);
nor U42738 (N_42738,N_41692,N_41771);
or U42739 (N_42739,N_41399,N_41488);
nor U42740 (N_42740,N_41422,N_41355);
nand U42741 (N_42741,N_41088,N_41193);
nor U42742 (N_42742,N_41568,N_41791);
nor U42743 (N_42743,N_41411,N_41608);
or U42744 (N_42744,N_41078,N_41643);
nand U42745 (N_42745,N_41560,N_41915);
xor U42746 (N_42746,N_41390,N_41286);
or U42747 (N_42747,N_41034,N_41691);
or U42748 (N_42748,N_41332,N_41062);
or U42749 (N_42749,N_41006,N_41732);
and U42750 (N_42750,N_41956,N_41949);
or U42751 (N_42751,N_41008,N_41357);
nor U42752 (N_42752,N_41559,N_41261);
nor U42753 (N_42753,N_41458,N_41056);
and U42754 (N_42754,N_41059,N_41064);
nor U42755 (N_42755,N_41277,N_41833);
and U42756 (N_42756,N_41974,N_41655);
nand U42757 (N_42757,N_41110,N_41633);
xnor U42758 (N_42758,N_41665,N_41706);
nor U42759 (N_42759,N_41364,N_41631);
nor U42760 (N_42760,N_41195,N_41829);
xnor U42761 (N_42761,N_41871,N_41251);
or U42762 (N_42762,N_41372,N_41920);
nor U42763 (N_42763,N_41595,N_41871);
nor U42764 (N_42764,N_41973,N_41773);
nand U42765 (N_42765,N_41285,N_41807);
or U42766 (N_42766,N_41257,N_41840);
or U42767 (N_42767,N_41881,N_41728);
xnor U42768 (N_42768,N_41316,N_41176);
and U42769 (N_42769,N_41182,N_41472);
xor U42770 (N_42770,N_41073,N_41958);
xnor U42771 (N_42771,N_41280,N_41462);
nand U42772 (N_42772,N_41574,N_41961);
and U42773 (N_42773,N_41125,N_41357);
nor U42774 (N_42774,N_41992,N_41561);
nand U42775 (N_42775,N_41322,N_41173);
or U42776 (N_42776,N_41231,N_41465);
xor U42777 (N_42777,N_41784,N_41480);
and U42778 (N_42778,N_41829,N_41590);
nand U42779 (N_42779,N_41572,N_41421);
nand U42780 (N_42780,N_41108,N_41407);
or U42781 (N_42781,N_41946,N_41505);
nor U42782 (N_42782,N_41268,N_41332);
and U42783 (N_42783,N_41949,N_41562);
xnor U42784 (N_42784,N_41290,N_41665);
or U42785 (N_42785,N_41636,N_41396);
and U42786 (N_42786,N_41487,N_41114);
xor U42787 (N_42787,N_41214,N_41351);
or U42788 (N_42788,N_41917,N_41000);
nand U42789 (N_42789,N_41889,N_41526);
or U42790 (N_42790,N_41225,N_41819);
xnor U42791 (N_42791,N_41671,N_41099);
xor U42792 (N_42792,N_41799,N_41898);
nand U42793 (N_42793,N_41258,N_41768);
nand U42794 (N_42794,N_41209,N_41419);
xnor U42795 (N_42795,N_41393,N_41026);
nand U42796 (N_42796,N_41012,N_41662);
xnor U42797 (N_42797,N_41168,N_41428);
xnor U42798 (N_42798,N_41497,N_41025);
and U42799 (N_42799,N_41586,N_41530);
nor U42800 (N_42800,N_41549,N_41893);
or U42801 (N_42801,N_41152,N_41133);
nor U42802 (N_42802,N_41714,N_41881);
and U42803 (N_42803,N_41652,N_41806);
nor U42804 (N_42804,N_41994,N_41086);
and U42805 (N_42805,N_41099,N_41312);
nor U42806 (N_42806,N_41265,N_41199);
and U42807 (N_42807,N_41203,N_41148);
or U42808 (N_42808,N_41206,N_41931);
nand U42809 (N_42809,N_41089,N_41762);
or U42810 (N_42810,N_41415,N_41364);
nand U42811 (N_42811,N_41331,N_41989);
or U42812 (N_42812,N_41071,N_41447);
and U42813 (N_42813,N_41920,N_41130);
nor U42814 (N_42814,N_41877,N_41901);
nand U42815 (N_42815,N_41046,N_41841);
nor U42816 (N_42816,N_41453,N_41092);
or U42817 (N_42817,N_41934,N_41483);
nand U42818 (N_42818,N_41519,N_41405);
xor U42819 (N_42819,N_41538,N_41837);
nor U42820 (N_42820,N_41090,N_41064);
nand U42821 (N_42821,N_41890,N_41912);
or U42822 (N_42822,N_41659,N_41397);
nor U42823 (N_42823,N_41765,N_41749);
and U42824 (N_42824,N_41706,N_41175);
nor U42825 (N_42825,N_41249,N_41592);
or U42826 (N_42826,N_41174,N_41431);
nand U42827 (N_42827,N_41664,N_41117);
nand U42828 (N_42828,N_41253,N_41088);
and U42829 (N_42829,N_41575,N_41765);
or U42830 (N_42830,N_41275,N_41239);
or U42831 (N_42831,N_41792,N_41433);
or U42832 (N_42832,N_41431,N_41758);
and U42833 (N_42833,N_41038,N_41745);
xor U42834 (N_42834,N_41806,N_41541);
xnor U42835 (N_42835,N_41832,N_41046);
and U42836 (N_42836,N_41285,N_41814);
and U42837 (N_42837,N_41308,N_41776);
nor U42838 (N_42838,N_41100,N_41512);
or U42839 (N_42839,N_41981,N_41358);
xnor U42840 (N_42840,N_41643,N_41792);
and U42841 (N_42841,N_41958,N_41046);
xnor U42842 (N_42842,N_41775,N_41042);
nand U42843 (N_42843,N_41443,N_41092);
or U42844 (N_42844,N_41566,N_41444);
nor U42845 (N_42845,N_41441,N_41159);
nand U42846 (N_42846,N_41203,N_41028);
xnor U42847 (N_42847,N_41713,N_41628);
nand U42848 (N_42848,N_41415,N_41147);
nor U42849 (N_42849,N_41313,N_41546);
and U42850 (N_42850,N_41484,N_41556);
xor U42851 (N_42851,N_41907,N_41754);
nand U42852 (N_42852,N_41196,N_41488);
xor U42853 (N_42853,N_41091,N_41474);
nand U42854 (N_42854,N_41264,N_41073);
xnor U42855 (N_42855,N_41135,N_41123);
nand U42856 (N_42856,N_41079,N_41917);
or U42857 (N_42857,N_41501,N_41121);
nor U42858 (N_42858,N_41611,N_41824);
and U42859 (N_42859,N_41466,N_41853);
nand U42860 (N_42860,N_41559,N_41804);
nand U42861 (N_42861,N_41043,N_41343);
or U42862 (N_42862,N_41750,N_41106);
and U42863 (N_42863,N_41444,N_41739);
xor U42864 (N_42864,N_41660,N_41026);
and U42865 (N_42865,N_41341,N_41062);
nor U42866 (N_42866,N_41285,N_41730);
and U42867 (N_42867,N_41100,N_41397);
or U42868 (N_42868,N_41967,N_41054);
or U42869 (N_42869,N_41806,N_41229);
or U42870 (N_42870,N_41260,N_41486);
and U42871 (N_42871,N_41999,N_41214);
or U42872 (N_42872,N_41502,N_41704);
and U42873 (N_42873,N_41206,N_41601);
nand U42874 (N_42874,N_41102,N_41223);
xnor U42875 (N_42875,N_41389,N_41189);
xnor U42876 (N_42876,N_41623,N_41258);
nand U42877 (N_42877,N_41219,N_41378);
or U42878 (N_42878,N_41380,N_41281);
and U42879 (N_42879,N_41805,N_41606);
and U42880 (N_42880,N_41175,N_41266);
or U42881 (N_42881,N_41941,N_41335);
or U42882 (N_42882,N_41900,N_41369);
nor U42883 (N_42883,N_41167,N_41160);
or U42884 (N_42884,N_41588,N_41824);
and U42885 (N_42885,N_41267,N_41223);
or U42886 (N_42886,N_41376,N_41319);
and U42887 (N_42887,N_41989,N_41667);
xor U42888 (N_42888,N_41714,N_41134);
xnor U42889 (N_42889,N_41803,N_41745);
nor U42890 (N_42890,N_41773,N_41471);
and U42891 (N_42891,N_41050,N_41460);
nor U42892 (N_42892,N_41530,N_41465);
nor U42893 (N_42893,N_41468,N_41601);
nor U42894 (N_42894,N_41077,N_41042);
and U42895 (N_42895,N_41253,N_41303);
xnor U42896 (N_42896,N_41153,N_41150);
nand U42897 (N_42897,N_41231,N_41180);
nor U42898 (N_42898,N_41324,N_41089);
or U42899 (N_42899,N_41897,N_41722);
xnor U42900 (N_42900,N_41360,N_41513);
nand U42901 (N_42901,N_41380,N_41202);
and U42902 (N_42902,N_41334,N_41918);
nor U42903 (N_42903,N_41575,N_41203);
or U42904 (N_42904,N_41158,N_41011);
nor U42905 (N_42905,N_41064,N_41506);
nand U42906 (N_42906,N_41282,N_41034);
nand U42907 (N_42907,N_41799,N_41868);
nand U42908 (N_42908,N_41840,N_41692);
xor U42909 (N_42909,N_41070,N_41345);
nor U42910 (N_42910,N_41541,N_41634);
nor U42911 (N_42911,N_41387,N_41379);
nor U42912 (N_42912,N_41946,N_41809);
xnor U42913 (N_42913,N_41254,N_41790);
xnor U42914 (N_42914,N_41026,N_41554);
xnor U42915 (N_42915,N_41725,N_41431);
or U42916 (N_42916,N_41174,N_41889);
and U42917 (N_42917,N_41979,N_41279);
or U42918 (N_42918,N_41921,N_41095);
nor U42919 (N_42919,N_41948,N_41238);
nand U42920 (N_42920,N_41765,N_41164);
nor U42921 (N_42921,N_41293,N_41852);
or U42922 (N_42922,N_41395,N_41185);
or U42923 (N_42923,N_41724,N_41548);
nand U42924 (N_42924,N_41139,N_41164);
and U42925 (N_42925,N_41978,N_41439);
nand U42926 (N_42926,N_41219,N_41619);
and U42927 (N_42927,N_41265,N_41072);
nand U42928 (N_42928,N_41938,N_41161);
xor U42929 (N_42929,N_41298,N_41081);
xor U42930 (N_42930,N_41109,N_41647);
nor U42931 (N_42931,N_41696,N_41139);
nor U42932 (N_42932,N_41261,N_41752);
nand U42933 (N_42933,N_41460,N_41773);
and U42934 (N_42934,N_41329,N_41375);
nand U42935 (N_42935,N_41519,N_41836);
nor U42936 (N_42936,N_41437,N_41525);
nand U42937 (N_42937,N_41137,N_41794);
nand U42938 (N_42938,N_41149,N_41058);
nand U42939 (N_42939,N_41792,N_41975);
and U42940 (N_42940,N_41249,N_41780);
and U42941 (N_42941,N_41812,N_41859);
nor U42942 (N_42942,N_41979,N_41633);
and U42943 (N_42943,N_41872,N_41140);
nand U42944 (N_42944,N_41966,N_41783);
nand U42945 (N_42945,N_41756,N_41809);
nor U42946 (N_42946,N_41193,N_41850);
nand U42947 (N_42947,N_41015,N_41544);
xnor U42948 (N_42948,N_41371,N_41539);
nor U42949 (N_42949,N_41951,N_41565);
nor U42950 (N_42950,N_41641,N_41551);
nor U42951 (N_42951,N_41195,N_41521);
xor U42952 (N_42952,N_41093,N_41607);
xor U42953 (N_42953,N_41611,N_41251);
nand U42954 (N_42954,N_41892,N_41618);
or U42955 (N_42955,N_41135,N_41424);
or U42956 (N_42956,N_41232,N_41066);
or U42957 (N_42957,N_41328,N_41309);
xnor U42958 (N_42958,N_41164,N_41633);
or U42959 (N_42959,N_41440,N_41747);
nand U42960 (N_42960,N_41898,N_41550);
xor U42961 (N_42961,N_41676,N_41506);
nor U42962 (N_42962,N_41623,N_41897);
nor U42963 (N_42963,N_41781,N_41240);
or U42964 (N_42964,N_41188,N_41043);
or U42965 (N_42965,N_41441,N_41644);
xor U42966 (N_42966,N_41019,N_41367);
or U42967 (N_42967,N_41473,N_41557);
or U42968 (N_42968,N_41479,N_41513);
nand U42969 (N_42969,N_41301,N_41393);
nand U42970 (N_42970,N_41140,N_41398);
nand U42971 (N_42971,N_41790,N_41031);
nand U42972 (N_42972,N_41821,N_41473);
xnor U42973 (N_42973,N_41671,N_41420);
xor U42974 (N_42974,N_41547,N_41343);
nor U42975 (N_42975,N_41538,N_41136);
and U42976 (N_42976,N_41860,N_41738);
nor U42977 (N_42977,N_41860,N_41613);
and U42978 (N_42978,N_41962,N_41820);
or U42979 (N_42979,N_41730,N_41573);
nand U42980 (N_42980,N_41198,N_41340);
xnor U42981 (N_42981,N_41426,N_41608);
nand U42982 (N_42982,N_41194,N_41869);
nor U42983 (N_42983,N_41890,N_41196);
or U42984 (N_42984,N_41866,N_41404);
and U42985 (N_42985,N_41241,N_41490);
nand U42986 (N_42986,N_41010,N_41173);
nand U42987 (N_42987,N_41915,N_41458);
xor U42988 (N_42988,N_41071,N_41642);
xnor U42989 (N_42989,N_41350,N_41294);
and U42990 (N_42990,N_41320,N_41190);
or U42991 (N_42991,N_41745,N_41548);
nor U42992 (N_42992,N_41980,N_41161);
nor U42993 (N_42993,N_41118,N_41642);
nor U42994 (N_42994,N_41173,N_41067);
and U42995 (N_42995,N_41250,N_41067);
or U42996 (N_42996,N_41247,N_41739);
or U42997 (N_42997,N_41752,N_41075);
nand U42998 (N_42998,N_41302,N_41507);
nor U42999 (N_42999,N_41483,N_41706);
and U43000 (N_43000,N_42465,N_42639);
nand U43001 (N_43001,N_42916,N_42103);
nand U43002 (N_43002,N_42901,N_42526);
and U43003 (N_43003,N_42585,N_42056);
nor U43004 (N_43004,N_42407,N_42166);
nand U43005 (N_43005,N_42837,N_42392);
nor U43006 (N_43006,N_42836,N_42927);
and U43007 (N_43007,N_42224,N_42621);
nand U43008 (N_43008,N_42134,N_42949);
or U43009 (N_43009,N_42084,N_42905);
xnor U43010 (N_43010,N_42842,N_42334);
xnor U43011 (N_43011,N_42571,N_42098);
nor U43012 (N_43012,N_42113,N_42488);
and U43013 (N_43013,N_42999,N_42705);
nor U43014 (N_43014,N_42427,N_42071);
nor U43015 (N_43015,N_42373,N_42294);
and U43016 (N_43016,N_42269,N_42934);
or U43017 (N_43017,N_42142,N_42893);
or U43018 (N_43018,N_42514,N_42300);
nand U43019 (N_43019,N_42727,N_42401);
or U43020 (N_43020,N_42509,N_42438);
or U43021 (N_43021,N_42039,N_42760);
nand U43022 (N_43022,N_42755,N_42674);
and U43023 (N_43023,N_42771,N_42910);
and U43024 (N_43024,N_42603,N_42960);
xnor U43025 (N_43025,N_42770,N_42829);
xor U43026 (N_43026,N_42006,N_42447);
nor U43027 (N_43027,N_42521,N_42956);
xnor U43028 (N_43028,N_42767,N_42408);
nand U43029 (N_43029,N_42076,N_42761);
nor U43030 (N_43030,N_42917,N_42497);
and U43031 (N_43031,N_42498,N_42951);
and U43032 (N_43032,N_42321,N_42278);
nor U43033 (N_43033,N_42965,N_42024);
xor U43034 (N_43034,N_42840,N_42087);
nor U43035 (N_43035,N_42788,N_42764);
nand U43036 (N_43036,N_42969,N_42993);
nor U43037 (N_43037,N_42979,N_42012);
and U43038 (N_43038,N_42726,N_42703);
and U43039 (N_43039,N_42768,N_42099);
or U43040 (N_43040,N_42240,N_42141);
xnor U43041 (N_43041,N_42400,N_42594);
nor U43042 (N_43042,N_42077,N_42534);
nor U43043 (N_43043,N_42417,N_42452);
nor U43044 (N_43044,N_42994,N_42816);
nor U43045 (N_43045,N_42130,N_42347);
xnor U43046 (N_43046,N_42894,N_42777);
xnor U43047 (N_43047,N_42353,N_42185);
or U43048 (N_43048,N_42237,N_42030);
nand U43049 (N_43049,N_42838,N_42535);
xor U43050 (N_43050,N_42355,N_42468);
or U43051 (N_43051,N_42093,N_42343);
or U43052 (N_43052,N_42647,N_42462);
nand U43053 (N_43053,N_42614,N_42293);
nand U43054 (N_43054,N_42065,N_42987);
and U43055 (N_43055,N_42439,N_42698);
or U43056 (N_43056,N_42389,N_42435);
and U43057 (N_43057,N_42442,N_42358);
xor U43058 (N_43058,N_42558,N_42940);
nand U43059 (N_43059,N_42425,N_42069);
nor U43060 (N_43060,N_42072,N_42298);
xnor U43061 (N_43061,N_42644,N_42413);
nor U43062 (N_43062,N_42483,N_42181);
or U43063 (N_43063,N_42158,N_42105);
nor U43064 (N_43064,N_42376,N_42932);
nor U43065 (N_43065,N_42653,N_42988);
xor U43066 (N_43066,N_42020,N_42210);
and U43067 (N_43067,N_42544,N_42792);
nand U43068 (N_43068,N_42375,N_42441);
nor U43069 (N_43069,N_42820,N_42980);
xnor U43070 (N_43070,N_42649,N_42051);
nand U43071 (N_43071,N_42067,N_42868);
nand U43072 (N_43072,N_42952,N_42902);
or U43073 (N_43073,N_42057,N_42464);
nor U43074 (N_43074,N_42776,N_42361);
xor U43075 (N_43075,N_42001,N_42944);
xor U43076 (N_43076,N_42615,N_42522);
xor U43077 (N_43077,N_42708,N_42195);
xnor U43078 (N_43078,N_42244,N_42446);
nor U43079 (N_43079,N_42756,N_42814);
xor U43080 (N_43080,N_42915,N_42505);
nor U43081 (N_43081,N_42660,N_42149);
and U43082 (N_43082,N_42551,N_42564);
or U43083 (N_43083,N_42774,N_42196);
or U43084 (N_43084,N_42909,N_42096);
or U43085 (N_43085,N_42707,N_42312);
and U43086 (N_43086,N_42168,N_42011);
nand U43087 (N_43087,N_42429,N_42613);
and U43088 (N_43088,N_42961,N_42699);
xnor U43089 (N_43089,N_42262,N_42877);
nand U43090 (N_43090,N_42007,N_42207);
and U43091 (N_43091,N_42570,N_42587);
nor U43092 (N_43092,N_42914,N_42741);
xnor U43093 (N_43093,N_42199,N_42907);
and U43094 (N_43094,N_42454,N_42068);
nand U43095 (N_43095,N_42518,N_42476);
nand U43096 (N_43096,N_42605,N_42136);
and U43097 (N_43097,N_42747,N_42265);
nand U43098 (N_43098,N_42947,N_42608);
nor U43099 (N_43099,N_42460,N_42310);
nor U43100 (N_43100,N_42888,N_42664);
nor U43101 (N_43101,N_42694,N_42859);
nor U43102 (N_43102,N_42044,N_42139);
or U43103 (N_43103,N_42931,N_42268);
or U43104 (N_43104,N_42701,N_42306);
xnor U43105 (N_43105,N_42780,N_42754);
or U43106 (N_43106,N_42576,N_42709);
and U43107 (N_43107,N_42272,N_42824);
or U43108 (N_43108,N_42396,N_42283);
or U43109 (N_43109,N_42617,N_42881);
nand U43110 (N_43110,N_42669,N_42147);
or U43111 (N_43111,N_42911,N_42882);
and U43112 (N_43112,N_42804,N_42304);
nor U43113 (N_43113,N_42192,N_42493);
and U43114 (N_43114,N_42981,N_42871);
or U43115 (N_43115,N_42088,N_42878);
nand U43116 (N_43116,N_42217,N_42630);
nand U43117 (N_43117,N_42772,N_42696);
xnor U43118 (N_43118,N_42364,N_42081);
or U43119 (N_43119,N_42242,N_42140);
xnor U43120 (N_43120,N_42326,N_42656);
nand U43121 (N_43121,N_42216,N_42582);
and U43122 (N_43122,N_42880,N_42299);
xor U43123 (N_43123,N_42249,N_42561);
xor U43124 (N_43124,N_42611,N_42174);
or U43125 (N_43125,N_42177,N_42331);
xnor U43126 (N_43126,N_42229,N_42054);
nand U43127 (N_43127,N_42205,N_42636);
nor U43128 (N_43128,N_42945,N_42720);
nor U43129 (N_43129,N_42398,N_42338);
and U43130 (N_43130,N_42155,N_42038);
nand U43131 (N_43131,N_42208,N_42463);
xor U43132 (N_43132,N_42284,N_42854);
or U43133 (N_43133,N_42110,N_42367);
xor U43134 (N_43134,N_42697,N_42519);
or U43135 (N_43135,N_42973,N_42743);
nand U43136 (N_43136,N_42554,N_42808);
nor U43137 (N_43137,N_42371,N_42520);
and U43138 (N_43138,N_42264,N_42586);
nor U43139 (N_43139,N_42975,N_42752);
xnor U43140 (N_43140,N_42287,N_42750);
and U43141 (N_43141,N_42512,N_42557);
or U43142 (N_43142,N_42145,N_42380);
nand U43143 (N_43143,N_42692,N_42785);
or U43144 (N_43144,N_42496,N_42926);
or U43145 (N_43145,N_42059,N_42797);
nor U43146 (N_43146,N_42307,N_42173);
nand U43147 (N_43147,N_42675,N_42393);
xor U43148 (N_43148,N_42434,N_42964);
and U43149 (N_43149,N_42959,N_42886);
or U43150 (N_43150,N_42957,N_42676);
nand U43151 (N_43151,N_42252,N_42146);
nor U43152 (N_43152,N_42507,N_42455);
or U43153 (N_43153,N_42948,N_42029);
and U43154 (N_43154,N_42009,N_42451);
nand U43155 (N_43155,N_42555,N_42853);
or U43156 (N_43156,N_42480,N_42976);
and U43157 (N_43157,N_42157,N_42598);
and U43158 (N_43158,N_42045,N_42835);
or U43159 (N_43159,N_42308,N_42341);
nand U43160 (N_43160,N_42623,N_42085);
nand U43161 (N_43161,N_42690,N_42101);
nand U43162 (N_43162,N_42550,N_42037);
and U43163 (N_43163,N_42672,N_42289);
or U43164 (N_43164,N_42572,N_42494);
or U43165 (N_43165,N_42120,N_42935);
nand U43166 (N_43166,N_42748,N_42728);
and U43167 (N_43167,N_42167,N_42958);
nor U43168 (N_43168,N_42805,N_42612);
and U43169 (N_43169,N_42688,N_42230);
nand U43170 (N_43170,N_42796,N_42740);
nor U43171 (N_43171,N_42083,N_42744);
xor U43172 (N_43172,N_42271,N_42047);
and U43173 (N_43173,N_42722,N_42857);
nand U43174 (N_43174,N_42938,N_42547);
xor U43175 (N_43175,N_42263,N_42991);
xnor U43176 (N_43176,N_42161,N_42388);
and U43177 (N_43177,N_42872,N_42875);
xnor U43178 (N_43178,N_42015,N_42220);
and U43179 (N_43179,N_42831,N_42937);
and U43180 (N_43180,N_42682,N_42552);
nand U43181 (N_43181,N_42259,N_42667);
or U43182 (N_43182,N_42052,N_42869);
xnor U43183 (N_43183,N_42784,N_42543);
nand U43184 (N_43184,N_42811,N_42733);
xor U43185 (N_43185,N_42243,N_42590);
and U43186 (N_43186,N_42686,N_42365);
xor U43187 (N_43187,N_42266,N_42445);
xor U43188 (N_43188,N_42848,N_42503);
or U43189 (N_43189,N_42529,N_42459);
and U43190 (N_43190,N_42953,N_42635);
or U43191 (N_43191,N_42972,N_42563);
nor U43192 (N_43192,N_42511,N_42584);
or U43193 (N_43193,N_42896,N_42286);
nor U43194 (N_43194,N_42346,N_42383);
nor U43195 (N_43195,N_42486,N_42276);
or U43196 (N_43196,N_42599,N_42183);
xor U43197 (N_43197,N_42390,N_42016);
xnor U43198 (N_43198,N_42179,N_42348);
xor U43199 (N_43199,N_42864,N_42345);
xnor U43200 (N_43200,N_42601,N_42583);
or U43201 (N_43201,N_42092,N_42638);
and U43202 (N_43202,N_42395,N_42654);
and U43203 (N_43203,N_42420,N_42484);
nand U43204 (N_43204,N_42971,N_42763);
nand U43205 (N_43205,N_42625,N_42899);
and U43206 (N_43206,N_42954,N_42022);
xnor U43207 (N_43207,N_42187,N_42714);
nand U43208 (N_43208,N_42409,N_42135);
and U43209 (N_43209,N_42873,N_42034);
xnor U43210 (N_43210,N_42236,N_42565);
nor U43211 (N_43211,N_42382,N_42549);
and U43212 (N_43212,N_42156,N_42591);
nand U43213 (N_43213,N_42821,N_42721);
nand U43214 (N_43214,N_42789,N_42658);
nand U43215 (N_43215,N_42049,N_42327);
or U43216 (N_43216,N_42121,N_42247);
and U43217 (N_43217,N_42381,N_42523);
and U43218 (N_43218,N_42983,N_42801);
xnor U43219 (N_43219,N_42324,N_42372);
or U43220 (N_43220,N_42004,N_42320);
or U43221 (N_43221,N_42366,N_42079);
nor U43222 (N_43222,N_42448,N_42432);
xor U43223 (N_43223,N_42074,N_42679);
xnor U43224 (N_43224,N_42596,N_42280);
or U43225 (N_43225,N_42642,N_42423);
nor U43226 (N_43226,N_42443,N_42203);
nor U43227 (N_43227,N_42295,N_42719);
and U43228 (N_43228,N_42633,N_42627);
nor U43229 (N_43229,N_42604,N_42212);
nand U43230 (N_43230,N_42489,N_42080);
nor U43231 (N_43231,N_42405,N_42211);
or U43232 (N_43232,N_42680,N_42610);
nand U43233 (N_43233,N_42370,N_42170);
or U43234 (N_43234,N_42033,N_42867);
nand U43235 (N_43235,N_42863,N_42990);
or U43236 (N_43236,N_42791,N_42702);
or U43237 (N_43237,N_42732,N_42759);
nand U43238 (N_43238,N_42691,N_42333);
and U43239 (N_43239,N_42193,N_42807);
nand U43240 (N_43240,N_42089,N_42330);
and U43241 (N_43241,N_42884,N_42645);
and U43242 (N_43242,N_42362,N_42578);
or U43243 (N_43243,N_42533,N_42678);
or U43244 (N_43244,N_42502,N_42412);
and U43245 (N_43245,N_42318,N_42270);
nor U43246 (N_43246,N_42588,N_42941);
and U43247 (N_43247,N_42643,N_42773);
or U43248 (N_43248,N_42053,N_42234);
nand U43249 (N_43249,N_42078,N_42695);
or U43250 (N_43250,N_42828,N_42670);
xnor U43251 (N_43251,N_42782,N_42580);
nand U43252 (N_43252,N_42111,N_42525);
nor U43253 (N_43253,N_42325,N_42499);
or U43254 (N_43254,N_42086,N_42100);
nor U43255 (N_43255,N_42624,N_42036);
or U43256 (N_43256,N_42303,N_42946);
xnor U43257 (N_43257,N_42787,N_42753);
and U43258 (N_43258,N_42713,N_42568);
nand U43259 (N_43259,N_42123,N_42176);
or U43260 (N_43260,N_42860,N_42449);
or U43261 (N_43261,N_42119,N_42479);
nor U43262 (N_43262,N_42538,N_42023);
and U43263 (N_43263,N_42492,N_42742);
nor U43264 (N_43264,N_42921,N_42977);
nand U43265 (N_43265,N_42474,N_42666);
or U43266 (N_43266,N_42651,N_42920);
nor U43267 (N_43267,N_42819,N_42215);
and U43268 (N_43268,N_42000,N_42481);
and U43269 (N_43269,N_42404,N_42410);
nor U43270 (N_43270,N_42221,N_42715);
or U43271 (N_43271,N_42731,N_42717);
nand U43272 (N_43272,N_42524,N_42553);
nor U43273 (N_43273,N_42144,N_42609);
or U43274 (N_43274,N_42094,N_42340);
xor U43275 (N_43275,N_42218,N_42018);
nand U43276 (N_43276,N_42560,N_42995);
or U43277 (N_43277,N_42491,N_42440);
or U43278 (N_43278,N_42936,N_42718);
or U43279 (N_43279,N_42391,N_42962);
or U43280 (N_43280,N_42904,N_42430);
nand U43281 (N_43281,N_42495,N_42040);
or U43282 (N_43282,N_42852,N_42124);
and U43283 (N_43283,N_42273,N_42632);
nand U43284 (N_43284,N_42329,N_42540);
nor U43285 (N_43285,N_42301,N_42851);
xnor U43286 (N_43286,N_42515,N_42267);
nor U43287 (N_43287,N_42206,N_42803);
and U43288 (N_43288,N_42794,N_42209);
nor U43289 (N_43289,N_42548,N_42245);
xnor U43290 (N_43290,N_42339,N_42433);
xnor U43291 (N_43291,N_42966,N_42516);
or U43292 (N_43292,N_42924,N_42150);
nand U43293 (N_43293,N_42189,N_42845);
and U43294 (N_43294,N_42062,N_42403);
xnor U43295 (N_43295,N_42027,N_42444);
nand U43296 (N_43296,N_42198,N_42475);
or U43297 (N_43297,N_42416,N_42188);
nand U43298 (N_43298,N_42929,N_42885);
nand U43299 (N_43299,N_42032,N_42169);
nor U43300 (N_43300,N_42201,N_42257);
or U43301 (N_43301,N_42665,N_42302);
and U43302 (N_43302,N_42017,N_42351);
or U43303 (N_43303,N_42827,N_42014);
nor U43304 (N_43304,N_42757,N_42335);
nand U43305 (N_43305,N_42737,N_42222);
nor U43306 (N_43306,N_42182,N_42275);
xnor U43307 (N_43307,N_42323,N_42419);
xnor U43308 (N_43308,N_42214,N_42456);
nand U43309 (N_43309,N_42528,N_42013);
and U43310 (N_43310,N_42527,N_42274);
nor U43311 (N_43311,N_42640,N_42809);
and U43312 (N_43312,N_42883,N_42781);
and U43313 (N_43313,N_42704,N_42746);
xor U43314 (N_43314,N_42626,N_42127);
nor U43315 (N_43315,N_42411,N_42865);
and U43316 (N_43316,N_42659,N_42279);
xor U43317 (N_43317,N_42133,N_42231);
xor U43318 (N_43318,N_42517,N_42890);
or U43319 (N_43319,N_42928,N_42629);
and U43320 (N_43320,N_42115,N_42681);
nand U43321 (N_43321,N_42470,N_42839);
nand U43322 (N_43322,N_42313,N_42125);
or U43323 (N_43323,N_42414,N_42542);
and U43324 (N_43324,N_42736,N_42876);
or U43325 (N_43325,N_42683,N_42200);
and U43326 (N_43326,N_42379,N_42620);
xor U43327 (N_43327,N_42126,N_42309);
xor U43328 (N_43328,N_42246,N_42058);
xor U43329 (N_43329,N_42426,N_42104);
nor U43330 (N_43330,N_42344,N_42858);
or U43331 (N_43331,N_42422,N_42290);
nor U43332 (N_43332,N_42261,N_42394);
or U43333 (N_43333,N_42655,N_42870);
xor U43334 (N_43334,N_42943,N_42490);
or U43335 (N_43335,N_42843,N_42634);
or U43336 (N_43336,N_42356,N_42833);
or U43337 (N_43337,N_42700,N_42874);
xor U43338 (N_43338,N_42043,N_42729);
nor U43339 (N_43339,N_42415,N_42897);
nand U43340 (N_43340,N_42162,N_42175);
nor U43341 (N_43341,N_42569,N_42559);
nand U43342 (N_43342,N_42288,N_42765);
and U43343 (N_43343,N_42895,N_42315);
or U43344 (N_43344,N_42311,N_42637);
nor U43345 (N_43345,N_42473,N_42779);
xor U43346 (N_43346,N_42606,N_42090);
and U43347 (N_43347,N_42850,N_42424);
nand U43348 (N_43348,N_42671,N_42122);
nand U43349 (N_43349,N_42360,N_42292);
xor U43350 (N_43350,N_42129,N_42725);
and U43351 (N_43351,N_42735,N_42532);
nor U43352 (N_43352,N_42592,N_42641);
nor U43353 (N_43353,N_42546,N_42689);
nor U43354 (N_43354,N_42855,N_42378);
nor U43355 (N_43355,N_42005,N_42107);
nand U43356 (N_43356,N_42912,N_42762);
and U43357 (N_43357,N_42577,N_42834);
nor U43358 (N_43358,N_42469,N_42930);
nand U43359 (N_43359,N_42806,N_42710);
and U43360 (N_43360,N_42368,N_42028);
and U43361 (N_43361,N_42766,N_42813);
xnor U43362 (N_43362,N_42758,N_42992);
or U43363 (N_43363,N_42091,N_42114);
or U43364 (N_43364,N_42841,N_42457);
xnor U43365 (N_43365,N_42508,N_42970);
nand U43366 (N_43366,N_42437,N_42233);
and U43367 (N_43367,N_42661,N_42963);
or U43368 (N_43368,N_42048,N_42482);
or U43369 (N_43369,N_42418,N_42073);
and U43370 (N_43370,N_42600,N_42628);
or U43371 (N_43371,N_42618,N_42539);
or U43372 (N_43372,N_42137,N_42802);
or U43373 (N_43373,N_42530,N_42402);
xnor U43374 (N_43374,N_42219,N_42238);
nand U43375 (N_43375,N_42567,N_42783);
and U43376 (N_43376,N_42984,N_42428);
or U43377 (N_43377,N_42436,N_42172);
and U43378 (N_43378,N_42685,N_42461);
and U43379 (N_43379,N_42749,N_42154);
and U43380 (N_43380,N_42003,N_42450);
nand U43381 (N_43381,N_42466,N_42019);
xor U43382 (N_43382,N_42844,N_42745);
nor U43383 (N_43383,N_42186,N_42989);
and U43384 (N_43384,N_42866,N_42102);
xor U43385 (N_43385,N_42232,N_42202);
xor U43386 (N_43386,N_42723,N_42734);
or U43387 (N_43387,N_42562,N_42662);
nand U43388 (N_43388,N_42925,N_42021);
xor U43389 (N_43389,N_42041,N_42684);
xnor U43390 (N_43390,N_42008,N_42861);
xor U43391 (N_43391,N_42297,N_42374);
nand U43392 (N_43392,N_42223,N_42349);
nand U43393 (N_43393,N_42035,N_42248);
and U43394 (N_43394,N_42291,N_42163);
and U43395 (N_43395,N_42055,N_42846);
nor U43396 (N_43396,N_42541,N_42918);
nor U43397 (N_43397,N_42317,N_42227);
nor U43398 (N_43398,N_42974,N_42652);
xnor U43399 (N_43399,N_42256,N_42900);
or U43400 (N_43400,N_42369,N_42898);
nor U43401 (N_43401,N_42471,N_42545);
nor U43402 (N_43402,N_42328,N_42128);
xnor U43403 (N_43403,N_42285,N_42026);
and U43404 (N_43404,N_42108,N_42913);
xnor U43405 (N_43405,N_42357,N_42143);
xor U43406 (N_43406,N_42847,N_42254);
xnor U43407 (N_43407,N_42810,N_42922);
and U43408 (N_43408,N_42397,N_42118);
nor U43409 (N_43409,N_42849,N_42751);
and U43410 (N_43410,N_42165,N_42453);
nor U43411 (N_43411,N_42738,N_42431);
or U43412 (N_43412,N_42574,N_42923);
or U43413 (N_43413,N_42967,N_42010);
nor U43414 (N_43414,N_42892,N_42812);
and U43415 (N_43415,N_42472,N_42504);
and U43416 (N_43416,N_42190,N_42650);
and U43417 (N_43417,N_42501,N_42506);
or U43418 (N_43418,N_42399,N_42180);
and U43419 (N_43419,N_42677,N_42706);
nand U43420 (N_43420,N_42536,N_42421);
and U43421 (N_43421,N_42573,N_42354);
nor U43422 (N_43422,N_42191,N_42800);
nand U43423 (N_43423,N_42826,N_42064);
or U43424 (N_43424,N_42194,N_42385);
and U43425 (N_43425,N_42891,N_42815);
and U43426 (N_43426,N_42082,N_42031);
nor U43427 (N_43427,N_42386,N_42939);
or U43428 (N_43428,N_42769,N_42817);
nand U43429 (N_43429,N_42790,N_42566);
or U43430 (N_43430,N_42458,N_42500);
nand U43431 (N_43431,N_42322,N_42225);
nor U43432 (N_43432,N_42942,N_42314);
and U43433 (N_43433,N_42204,N_42968);
nor U43434 (N_43434,N_42619,N_42097);
nand U43435 (N_43435,N_42985,N_42879);
and U43436 (N_43436,N_42595,N_42159);
nand U43437 (N_43437,N_42138,N_42795);
nand U43438 (N_43438,N_42657,N_42887);
nand U43439 (N_43439,N_42616,N_42998);
and U43440 (N_43440,N_42352,N_42213);
and U43441 (N_43441,N_42152,N_42342);
nand U43442 (N_43442,N_42116,N_42117);
nor U43443 (N_43443,N_42978,N_42002);
xnor U43444 (N_43444,N_42332,N_42646);
and U43445 (N_43445,N_42477,N_42799);
nor U43446 (N_43446,N_42337,N_42982);
nand U43447 (N_43447,N_42579,N_42239);
xor U43448 (N_43448,N_42487,N_42387);
nor U43449 (N_43449,N_42226,N_42050);
xnor U43450 (N_43450,N_42319,N_42406);
nand U43451 (N_43451,N_42822,N_42823);
nand U43452 (N_43452,N_42336,N_42862);
and U43453 (N_43453,N_42997,N_42607);
xnor U43454 (N_43454,N_42250,N_42818);
and U43455 (N_43455,N_42631,N_42950);
nor U43456 (N_43456,N_42160,N_42485);
and U43457 (N_43457,N_42687,N_42258);
nor U43458 (N_43458,N_42589,N_42075);
xnor U43459 (N_43459,N_42106,N_42171);
nor U43460 (N_43460,N_42253,N_42131);
or U43461 (N_43461,N_42063,N_42070);
nand U43462 (N_43462,N_42793,N_42919);
xor U43463 (N_43463,N_42668,N_42712);
xor U43464 (N_43464,N_42739,N_42673);
xor U43465 (N_43465,N_42153,N_42363);
xnor U43466 (N_43466,N_42663,N_42716);
nand U43467 (N_43467,N_42537,N_42575);
nor U43468 (N_43468,N_42648,N_42830);
and U43469 (N_43469,N_42148,N_42622);
xnor U43470 (N_43470,N_42350,N_42377);
and U43471 (N_43471,N_42908,N_42132);
or U43472 (N_43472,N_42060,N_42832);
and U43473 (N_43473,N_42933,N_42711);
and U43474 (N_43474,N_42906,N_42281);
nand U43475 (N_43475,N_42693,N_42109);
xnor U43476 (N_43476,N_42095,N_42581);
and U43477 (N_43477,N_42856,N_42025);
and U43478 (N_43478,N_42778,N_42467);
and U43479 (N_43479,N_42798,N_42282);
or U43480 (N_43480,N_42597,N_42251);
nor U43481 (N_43481,N_42316,N_42889);
and U43482 (N_43482,N_42197,N_42384);
and U43483 (N_43483,N_42112,N_42602);
nor U43484 (N_43484,N_42478,N_42178);
nand U43485 (N_43485,N_42510,N_42730);
xnor U43486 (N_43486,N_42184,N_42724);
and U43487 (N_43487,N_42296,N_42061);
and U43488 (N_43488,N_42241,N_42164);
nand U43489 (N_43489,N_42066,N_42825);
nand U43490 (N_43490,N_42955,N_42531);
and U43491 (N_43491,N_42513,N_42228);
xor U43492 (N_43492,N_42046,N_42042);
xor U43493 (N_43493,N_42260,N_42255);
or U43494 (N_43494,N_42986,N_42305);
or U43495 (N_43495,N_42903,N_42556);
or U43496 (N_43496,N_42786,N_42996);
nand U43497 (N_43497,N_42593,N_42151);
or U43498 (N_43498,N_42277,N_42775);
xor U43499 (N_43499,N_42359,N_42235);
nor U43500 (N_43500,N_42617,N_42743);
nand U43501 (N_43501,N_42410,N_42932);
nand U43502 (N_43502,N_42538,N_42645);
xnor U43503 (N_43503,N_42053,N_42454);
xnor U43504 (N_43504,N_42122,N_42797);
and U43505 (N_43505,N_42087,N_42145);
and U43506 (N_43506,N_42236,N_42220);
xor U43507 (N_43507,N_42557,N_42726);
nor U43508 (N_43508,N_42556,N_42016);
nand U43509 (N_43509,N_42531,N_42264);
xnor U43510 (N_43510,N_42984,N_42128);
nand U43511 (N_43511,N_42098,N_42862);
or U43512 (N_43512,N_42257,N_42724);
or U43513 (N_43513,N_42812,N_42841);
and U43514 (N_43514,N_42442,N_42622);
xor U43515 (N_43515,N_42202,N_42763);
or U43516 (N_43516,N_42395,N_42026);
nand U43517 (N_43517,N_42395,N_42366);
or U43518 (N_43518,N_42290,N_42381);
xor U43519 (N_43519,N_42490,N_42741);
or U43520 (N_43520,N_42610,N_42770);
xor U43521 (N_43521,N_42984,N_42704);
xor U43522 (N_43522,N_42569,N_42283);
nor U43523 (N_43523,N_42681,N_42191);
nand U43524 (N_43524,N_42503,N_42163);
or U43525 (N_43525,N_42130,N_42270);
nand U43526 (N_43526,N_42149,N_42094);
or U43527 (N_43527,N_42208,N_42574);
nand U43528 (N_43528,N_42770,N_42193);
nand U43529 (N_43529,N_42361,N_42104);
or U43530 (N_43530,N_42523,N_42697);
nor U43531 (N_43531,N_42885,N_42615);
or U43532 (N_43532,N_42167,N_42441);
xnor U43533 (N_43533,N_42856,N_42252);
nand U43534 (N_43534,N_42691,N_42715);
or U43535 (N_43535,N_42985,N_42091);
nor U43536 (N_43536,N_42630,N_42793);
or U43537 (N_43537,N_42457,N_42640);
and U43538 (N_43538,N_42453,N_42582);
nand U43539 (N_43539,N_42078,N_42137);
nand U43540 (N_43540,N_42675,N_42078);
or U43541 (N_43541,N_42034,N_42708);
and U43542 (N_43542,N_42827,N_42172);
or U43543 (N_43543,N_42032,N_42325);
nand U43544 (N_43544,N_42667,N_42904);
or U43545 (N_43545,N_42281,N_42133);
xnor U43546 (N_43546,N_42854,N_42587);
nand U43547 (N_43547,N_42051,N_42471);
xnor U43548 (N_43548,N_42217,N_42990);
xnor U43549 (N_43549,N_42046,N_42449);
nor U43550 (N_43550,N_42051,N_42396);
xor U43551 (N_43551,N_42917,N_42748);
xnor U43552 (N_43552,N_42135,N_42012);
or U43553 (N_43553,N_42730,N_42028);
nand U43554 (N_43554,N_42381,N_42451);
nor U43555 (N_43555,N_42415,N_42937);
or U43556 (N_43556,N_42641,N_42589);
nor U43557 (N_43557,N_42029,N_42926);
or U43558 (N_43558,N_42677,N_42959);
nor U43559 (N_43559,N_42567,N_42853);
nor U43560 (N_43560,N_42255,N_42427);
or U43561 (N_43561,N_42043,N_42135);
nor U43562 (N_43562,N_42205,N_42953);
or U43563 (N_43563,N_42646,N_42884);
nor U43564 (N_43564,N_42579,N_42940);
xnor U43565 (N_43565,N_42926,N_42427);
xnor U43566 (N_43566,N_42332,N_42257);
or U43567 (N_43567,N_42110,N_42752);
nand U43568 (N_43568,N_42183,N_42827);
nor U43569 (N_43569,N_42406,N_42767);
or U43570 (N_43570,N_42609,N_42572);
and U43571 (N_43571,N_42273,N_42278);
nor U43572 (N_43572,N_42305,N_42517);
and U43573 (N_43573,N_42519,N_42386);
and U43574 (N_43574,N_42042,N_42226);
or U43575 (N_43575,N_42996,N_42749);
and U43576 (N_43576,N_42042,N_42212);
nor U43577 (N_43577,N_42149,N_42784);
and U43578 (N_43578,N_42002,N_42529);
or U43579 (N_43579,N_42127,N_42344);
or U43580 (N_43580,N_42556,N_42572);
nand U43581 (N_43581,N_42972,N_42350);
nor U43582 (N_43582,N_42256,N_42683);
nand U43583 (N_43583,N_42364,N_42293);
xor U43584 (N_43584,N_42792,N_42354);
nand U43585 (N_43585,N_42985,N_42664);
and U43586 (N_43586,N_42169,N_42341);
or U43587 (N_43587,N_42725,N_42373);
and U43588 (N_43588,N_42479,N_42806);
and U43589 (N_43589,N_42743,N_42598);
nand U43590 (N_43590,N_42101,N_42367);
and U43591 (N_43591,N_42988,N_42628);
nand U43592 (N_43592,N_42038,N_42173);
and U43593 (N_43593,N_42603,N_42285);
xnor U43594 (N_43594,N_42505,N_42324);
xor U43595 (N_43595,N_42097,N_42126);
and U43596 (N_43596,N_42486,N_42024);
nand U43597 (N_43597,N_42624,N_42905);
or U43598 (N_43598,N_42213,N_42017);
and U43599 (N_43599,N_42804,N_42895);
xor U43600 (N_43600,N_42800,N_42054);
nand U43601 (N_43601,N_42589,N_42626);
or U43602 (N_43602,N_42988,N_42225);
xor U43603 (N_43603,N_42436,N_42959);
nor U43604 (N_43604,N_42039,N_42381);
nand U43605 (N_43605,N_42898,N_42657);
xnor U43606 (N_43606,N_42574,N_42087);
nand U43607 (N_43607,N_42236,N_42717);
xor U43608 (N_43608,N_42122,N_42176);
and U43609 (N_43609,N_42455,N_42432);
nor U43610 (N_43610,N_42508,N_42692);
and U43611 (N_43611,N_42752,N_42295);
or U43612 (N_43612,N_42659,N_42762);
and U43613 (N_43613,N_42723,N_42233);
and U43614 (N_43614,N_42941,N_42864);
nor U43615 (N_43615,N_42180,N_42859);
and U43616 (N_43616,N_42574,N_42764);
xnor U43617 (N_43617,N_42480,N_42894);
and U43618 (N_43618,N_42408,N_42178);
xor U43619 (N_43619,N_42578,N_42780);
nand U43620 (N_43620,N_42027,N_42557);
xor U43621 (N_43621,N_42882,N_42555);
and U43622 (N_43622,N_42609,N_42295);
nor U43623 (N_43623,N_42001,N_42543);
nor U43624 (N_43624,N_42928,N_42718);
nor U43625 (N_43625,N_42626,N_42357);
or U43626 (N_43626,N_42395,N_42791);
and U43627 (N_43627,N_42827,N_42593);
nand U43628 (N_43628,N_42603,N_42033);
nor U43629 (N_43629,N_42641,N_42071);
nor U43630 (N_43630,N_42902,N_42848);
nand U43631 (N_43631,N_42715,N_42756);
or U43632 (N_43632,N_42343,N_42289);
xnor U43633 (N_43633,N_42945,N_42928);
or U43634 (N_43634,N_42882,N_42741);
nand U43635 (N_43635,N_42000,N_42583);
and U43636 (N_43636,N_42620,N_42120);
nand U43637 (N_43637,N_42882,N_42463);
xnor U43638 (N_43638,N_42445,N_42206);
and U43639 (N_43639,N_42470,N_42592);
and U43640 (N_43640,N_42424,N_42608);
nor U43641 (N_43641,N_42309,N_42147);
xor U43642 (N_43642,N_42841,N_42276);
nand U43643 (N_43643,N_42845,N_42784);
and U43644 (N_43644,N_42166,N_42234);
or U43645 (N_43645,N_42933,N_42344);
nand U43646 (N_43646,N_42040,N_42467);
or U43647 (N_43647,N_42494,N_42430);
or U43648 (N_43648,N_42601,N_42188);
and U43649 (N_43649,N_42204,N_42924);
xnor U43650 (N_43650,N_42507,N_42534);
nand U43651 (N_43651,N_42638,N_42661);
and U43652 (N_43652,N_42101,N_42059);
nor U43653 (N_43653,N_42918,N_42397);
or U43654 (N_43654,N_42478,N_42630);
nand U43655 (N_43655,N_42021,N_42605);
and U43656 (N_43656,N_42897,N_42430);
and U43657 (N_43657,N_42114,N_42491);
xor U43658 (N_43658,N_42458,N_42389);
nor U43659 (N_43659,N_42691,N_42272);
nand U43660 (N_43660,N_42692,N_42418);
xnor U43661 (N_43661,N_42265,N_42616);
and U43662 (N_43662,N_42963,N_42560);
nor U43663 (N_43663,N_42041,N_42967);
or U43664 (N_43664,N_42645,N_42238);
nor U43665 (N_43665,N_42261,N_42536);
or U43666 (N_43666,N_42746,N_42075);
nor U43667 (N_43667,N_42962,N_42083);
nand U43668 (N_43668,N_42807,N_42138);
xnor U43669 (N_43669,N_42342,N_42341);
or U43670 (N_43670,N_42067,N_42737);
nand U43671 (N_43671,N_42943,N_42507);
xor U43672 (N_43672,N_42778,N_42436);
xor U43673 (N_43673,N_42231,N_42910);
or U43674 (N_43674,N_42432,N_42986);
and U43675 (N_43675,N_42155,N_42289);
xnor U43676 (N_43676,N_42168,N_42391);
nor U43677 (N_43677,N_42034,N_42382);
or U43678 (N_43678,N_42984,N_42992);
xnor U43679 (N_43679,N_42961,N_42591);
nor U43680 (N_43680,N_42986,N_42008);
and U43681 (N_43681,N_42354,N_42672);
nor U43682 (N_43682,N_42289,N_42817);
xnor U43683 (N_43683,N_42594,N_42106);
nand U43684 (N_43684,N_42689,N_42936);
or U43685 (N_43685,N_42618,N_42950);
or U43686 (N_43686,N_42504,N_42973);
and U43687 (N_43687,N_42956,N_42945);
or U43688 (N_43688,N_42498,N_42920);
nor U43689 (N_43689,N_42605,N_42048);
nand U43690 (N_43690,N_42063,N_42123);
xor U43691 (N_43691,N_42411,N_42684);
nand U43692 (N_43692,N_42411,N_42028);
xor U43693 (N_43693,N_42822,N_42141);
nor U43694 (N_43694,N_42744,N_42598);
nand U43695 (N_43695,N_42717,N_42706);
xor U43696 (N_43696,N_42214,N_42774);
nand U43697 (N_43697,N_42288,N_42033);
nor U43698 (N_43698,N_42207,N_42815);
and U43699 (N_43699,N_42435,N_42964);
xnor U43700 (N_43700,N_42124,N_42574);
or U43701 (N_43701,N_42026,N_42569);
xnor U43702 (N_43702,N_42484,N_42108);
or U43703 (N_43703,N_42583,N_42697);
nand U43704 (N_43704,N_42657,N_42548);
nor U43705 (N_43705,N_42559,N_42089);
or U43706 (N_43706,N_42191,N_42809);
or U43707 (N_43707,N_42580,N_42166);
xor U43708 (N_43708,N_42421,N_42360);
nor U43709 (N_43709,N_42619,N_42812);
xnor U43710 (N_43710,N_42908,N_42385);
xor U43711 (N_43711,N_42847,N_42308);
nand U43712 (N_43712,N_42544,N_42239);
nand U43713 (N_43713,N_42419,N_42181);
nand U43714 (N_43714,N_42103,N_42164);
and U43715 (N_43715,N_42304,N_42100);
or U43716 (N_43716,N_42247,N_42278);
nor U43717 (N_43717,N_42792,N_42237);
nor U43718 (N_43718,N_42643,N_42128);
nor U43719 (N_43719,N_42421,N_42723);
nand U43720 (N_43720,N_42530,N_42627);
nor U43721 (N_43721,N_42725,N_42602);
xor U43722 (N_43722,N_42495,N_42140);
nor U43723 (N_43723,N_42630,N_42014);
nor U43724 (N_43724,N_42273,N_42317);
nor U43725 (N_43725,N_42327,N_42311);
nand U43726 (N_43726,N_42017,N_42187);
xor U43727 (N_43727,N_42831,N_42401);
nand U43728 (N_43728,N_42432,N_42454);
nor U43729 (N_43729,N_42474,N_42595);
nand U43730 (N_43730,N_42793,N_42214);
nand U43731 (N_43731,N_42725,N_42369);
or U43732 (N_43732,N_42597,N_42454);
nand U43733 (N_43733,N_42687,N_42451);
and U43734 (N_43734,N_42198,N_42197);
nor U43735 (N_43735,N_42837,N_42994);
xor U43736 (N_43736,N_42449,N_42574);
or U43737 (N_43737,N_42822,N_42251);
or U43738 (N_43738,N_42813,N_42328);
nand U43739 (N_43739,N_42859,N_42495);
xnor U43740 (N_43740,N_42794,N_42490);
nor U43741 (N_43741,N_42061,N_42272);
or U43742 (N_43742,N_42952,N_42879);
or U43743 (N_43743,N_42589,N_42538);
or U43744 (N_43744,N_42377,N_42815);
nand U43745 (N_43745,N_42925,N_42851);
xor U43746 (N_43746,N_42328,N_42321);
xnor U43747 (N_43747,N_42041,N_42830);
xnor U43748 (N_43748,N_42806,N_42678);
nor U43749 (N_43749,N_42376,N_42131);
nor U43750 (N_43750,N_42887,N_42567);
or U43751 (N_43751,N_42588,N_42993);
or U43752 (N_43752,N_42491,N_42963);
or U43753 (N_43753,N_42985,N_42371);
nor U43754 (N_43754,N_42360,N_42716);
nand U43755 (N_43755,N_42876,N_42716);
xnor U43756 (N_43756,N_42559,N_42877);
nor U43757 (N_43757,N_42219,N_42852);
or U43758 (N_43758,N_42267,N_42037);
xnor U43759 (N_43759,N_42128,N_42712);
nor U43760 (N_43760,N_42956,N_42952);
or U43761 (N_43761,N_42762,N_42648);
or U43762 (N_43762,N_42887,N_42750);
and U43763 (N_43763,N_42344,N_42058);
or U43764 (N_43764,N_42581,N_42750);
nor U43765 (N_43765,N_42334,N_42724);
or U43766 (N_43766,N_42312,N_42241);
nor U43767 (N_43767,N_42581,N_42101);
and U43768 (N_43768,N_42278,N_42644);
nand U43769 (N_43769,N_42330,N_42662);
or U43770 (N_43770,N_42448,N_42467);
xor U43771 (N_43771,N_42639,N_42653);
or U43772 (N_43772,N_42826,N_42440);
nand U43773 (N_43773,N_42513,N_42477);
or U43774 (N_43774,N_42200,N_42312);
and U43775 (N_43775,N_42110,N_42698);
nand U43776 (N_43776,N_42767,N_42312);
or U43777 (N_43777,N_42304,N_42480);
or U43778 (N_43778,N_42543,N_42776);
or U43779 (N_43779,N_42286,N_42609);
xnor U43780 (N_43780,N_42553,N_42887);
and U43781 (N_43781,N_42684,N_42937);
and U43782 (N_43782,N_42885,N_42841);
or U43783 (N_43783,N_42469,N_42133);
nor U43784 (N_43784,N_42356,N_42031);
and U43785 (N_43785,N_42241,N_42496);
nor U43786 (N_43786,N_42013,N_42279);
or U43787 (N_43787,N_42555,N_42957);
or U43788 (N_43788,N_42539,N_42193);
and U43789 (N_43789,N_42933,N_42805);
or U43790 (N_43790,N_42460,N_42217);
xor U43791 (N_43791,N_42123,N_42480);
nand U43792 (N_43792,N_42420,N_42793);
and U43793 (N_43793,N_42210,N_42524);
or U43794 (N_43794,N_42573,N_42879);
nor U43795 (N_43795,N_42702,N_42871);
nand U43796 (N_43796,N_42842,N_42070);
nand U43797 (N_43797,N_42170,N_42361);
xor U43798 (N_43798,N_42201,N_42508);
or U43799 (N_43799,N_42732,N_42199);
xnor U43800 (N_43800,N_42198,N_42104);
and U43801 (N_43801,N_42776,N_42924);
or U43802 (N_43802,N_42975,N_42248);
nor U43803 (N_43803,N_42690,N_42820);
xnor U43804 (N_43804,N_42009,N_42127);
nand U43805 (N_43805,N_42941,N_42023);
or U43806 (N_43806,N_42001,N_42674);
and U43807 (N_43807,N_42772,N_42524);
or U43808 (N_43808,N_42551,N_42487);
xnor U43809 (N_43809,N_42972,N_42066);
xor U43810 (N_43810,N_42750,N_42618);
nor U43811 (N_43811,N_42307,N_42411);
and U43812 (N_43812,N_42590,N_42425);
and U43813 (N_43813,N_42566,N_42621);
or U43814 (N_43814,N_42221,N_42799);
nand U43815 (N_43815,N_42290,N_42944);
nand U43816 (N_43816,N_42689,N_42717);
nor U43817 (N_43817,N_42095,N_42223);
and U43818 (N_43818,N_42659,N_42292);
nand U43819 (N_43819,N_42945,N_42841);
and U43820 (N_43820,N_42495,N_42535);
and U43821 (N_43821,N_42327,N_42512);
nor U43822 (N_43822,N_42152,N_42622);
xnor U43823 (N_43823,N_42617,N_42843);
or U43824 (N_43824,N_42499,N_42106);
nor U43825 (N_43825,N_42765,N_42874);
or U43826 (N_43826,N_42867,N_42025);
or U43827 (N_43827,N_42501,N_42424);
nor U43828 (N_43828,N_42005,N_42318);
xnor U43829 (N_43829,N_42518,N_42712);
or U43830 (N_43830,N_42810,N_42240);
nand U43831 (N_43831,N_42202,N_42321);
nor U43832 (N_43832,N_42007,N_42942);
or U43833 (N_43833,N_42344,N_42148);
nor U43834 (N_43834,N_42686,N_42118);
and U43835 (N_43835,N_42963,N_42676);
nand U43836 (N_43836,N_42228,N_42414);
nor U43837 (N_43837,N_42543,N_42177);
nor U43838 (N_43838,N_42578,N_42392);
xor U43839 (N_43839,N_42585,N_42826);
xor U43840 (N_43840,N_42429,N_42187);
nand U43841 (N_43841,N_42884,N_42403);
nand U43842 (N_43842,N_42060,N_42960);
or U43843 (N_43843,N_42985,N_42431);
or U43844 (N_43844,N_42206,N_42499);
and U43845 (N_43845,N_42280,N_42750);
and U43846 (N_43846,N_42063,N_42618);
nand U43847 (N_43847,N_42346,N_42435);
nor U43848 (N_43848,N_42082,N_42783);
or U43849 (N_43849,N_42168,N_42156);
nand U43850 (N_43850,N_42315,N_42455);
nor U43851 (N_43851,N_42118,N_42345);
nor U43852 (N_43852,N_42943,N_42753);
nor U43853 (N_43853,N_42754,N_42314);
and U43854 (N_43854,N_42780,N_42589);
or U43855 (N_43855,N_42392,N_42516);
nand U43856 (N_43856,N_42313,N_42668);
xor U43857 (N_43857,N_42156,N_42101);
and U43858 (N_43858,N_42407,N_42494);
nor U43859 (N_43859,N_42190,N_42488);
and U43860 (N_43860,N_42251,N_42948);
and U43861 (N_43861,N_42390,N_42477);
nor U43862 (N_43862,N_42242,N_42474);
nor U43863 (N_43863,N_42136,N_42599);
or U43864 (N_43864,N_42856,N_42950);
xor U43865 (N_43865,N_42715,N_42736);
xnor U43866 (N_43866,N_42076,N_42393);
nand U43867 (N_43867,N_42191,N_42403);
xor U43868 (N_43868,N_42195,N_42966);
nand U43869 (N_43869,N_42093,N_42149);
nor U43870 (N_43870,N_42394,N_42165);
nor U43871 (N_43871,N_42082,N_42795);
nand U43872 (N_43872,N_42554,N_42387);
and U43873 (N_43873,N_42403,N_42484);
nor U43874 (N_43874,N_42831,N_42562);
xor U43875 (N_43875,N_42988,N_42459);
nor U43876 (N_43876,N_42857,N_42313);
nor U43877 (N_43877,N_42497,N_42104);
nor U43878 (N_43878,N_42936,N_42984);
or U43879 (N_43879,N_42413,N_42940);
nand U43880 (N_43880,N_42689,N_42132);
xor U43881 (N_43881,N_42673,N_42314);
nand U43882 (N_43882,N_42863,N_42284);
or U43883 (N_43883,N_42876,N_42388);
and U43884 (N_43884,N_42515,N_42501);
or U43885 (N_43885,N_42536,N_42643);
xnor U43886 (N_43886,N_42995,N_42793);
or U43887 (N_43887,N_42589,N_42852);
and U43888 (N_43888,N_42618,N_42048);
nand U43889 (N_43889,N_42005,N_42524);
nor U43890 (N_43890,N_42482,N_42804);
nand U43891 (N_43891,N_42122,N_42460);
xnor U43892 (N_43892,N_42132,N_42471);
xor U43893 (N_43893,N_42400,N_42401);
or U43894 (N_43894,N_42948,N_42531);
and U43895 (N_43895,N_42932,N_42657);
xnor U43896 (N_43896,N_42963,N_42822);
xnor U43897 (N_43897,N_42152,N_42514);
nor U43898 (N_43898,N_42750,N_42190);
nor U43899 (N_43899,N_42495,N_42369);
xor U43900 (N_43900,N_42753,N_42408);
nand U43901 (N_43901,N_42816,N_42309);
nand U43902 (N_43902,N_42963,N_42435);
xnor U43903 (N_43903,N_42821,N_42967);
nand U43904 (N_43904,N_42740,N_42726);
and U43905 (N_43905,N_42690,N_42733);
and U43906 (N_43906,N_42307,N_42950);
nor U43907 (N_43907,N_42121,N_42272);
nor U43908 (N_43908,N_42007,N_42573);
nand U43909 (N_43909,N_42098,N_42766);
and U43910 (N_43910,N_42699,N_42337);
or U43911 (N_43911,N_42945,N_42460);
nor U43912 (N_43912,N_42696,N_42510);
and U43913 (N_43913,N_42072,N_42703);
or U43914 (N_43914,N_42855,N_42734);
nand U43915 (N_43915,N_42776,N_42060);
nand U43916 (N_43916,N_42893,N_42197);
nor U43917 (N_43917,N_42461,N_42398);
or U43918 (N_43918,N_42678,N_42685);
xor U43919 (N_43919,N_42129,N_42150);
nand U43920 (N_43920,N_42802,N_42029);
nor U43921 (N_43921,N_42012,N_42653);
nand U43922 (N_43922,N_42410,N_42360);
nand U43923 (N_43923,N_42176,N_42024);
and U43924 (N_43924,N_42096,N_42462);
and U43925 (N_43925,N_42256,N_42912);
nor U43926 (N_43926,N_42800,N_42944);
and U43927 (N_43927,N_42087,N_42726);
nor U43928 (N_43928,N_42912,N_42759);
xor U43929 (N_43929,N_42607,N_42740);
nand U43930 (N_43930,N_42674,N_42306);
nor U43931 (N_43931,N_42473,N_42505);
xor U43932 (N_43932,N_42060,N_42676);
and U43933 (N_43933,N_42035,N_42836);
nand U43934 (N_43934,N_42448,N_42932);
or U43935 (N_43935,N_42378,N_42806);
nor U43936 (N_43936,N_42969,N_42087);
or U43937 (N_43937,N_42871,N_42905);
nand U43938 (N_43938,N_42137,N_42534);
xnor U43939 (N_43939,N_42581,N_42610);
xnor U43940 (N_43940,N_42708,N_42485);
xnor U43941 (N_43941,N_42432,N_42534);
or U43942 (N_43942,N_42110,N_42716);
or U43943 (N_43943,N_42036,N_42521);
and U43944 (N_43944,N_42417,N_42451);
and U43945 (N_43945,N_42460,N_42021);
nand U43946 (N_43946,N_42102,N_42883);
or U43947 (N_43947,N_42457,N_42938);
nor U43948 (N_43948,N_42451,N_42954);
and U43949 (N_43949,N_42052,N_42532);
nor U43950 (N_43950,N_42202,N_42656);
xor U43951 (N_43951,N_42821,N_42898);
nor U43952 (N_43952,N_42127,N_42001);
xor U43953 (N_43953,N_42963,N_42249);
nor U43954 (N_43954,N_42739,N_42991);
and U43955 (N_43955,N_42344,N_42334);
xnor U43956 (N_43956,N_42066,N_42609);
nor U43957 (N_43957,N_42630,N_42269);
xnor U43958 (N_43958,N_42162,N_42734);
and U43959 (N_43959,N_42548,N_42467);
xnor U43960 (N_43960,N_42176,N_42368);
xor U43961 (N_43961,N_42196,N_42334);
nand U43962 (N_43962,N_42803,N_42061);
nand U43963 (N_43963,N_42718,N_42571);
and U43964 (N_43964,N_42707,N_42239);
xnor U43965 (N_43965,N_42612,N_42585);
nor U43966 (N_43966,N_42253,N_42154);
nand U43967 (N_43967,N_42779,N_42101);
nand U43968 (N_43968,N_42154,N_42896);
and U43969 (N_43969,N_42985,N_42012);
xor U43970 (N_43970,N_42363,N_42529);
xor U43971 (N_43971,N_42385,N_42168);
xor U43972 (N_43972,N_42636,N_42291);
nand U43973 (N_43973,N_42087,N_42152);
nand U43974 (N_43974,N_42333,N_42056);
and U43975 (N_43975,N_42383,N_42914);
xor U43976 (N_43976,N_42828,N_42636);
nor U43977 (N_43977,N_42259,N_42664);
or U43978 (N_43978,N_42359,N_42532);
and U43979 (N_43979,N_42130,N_42202);
xor U43980 (N_43980,N_42088,N_42146);
xnor U43981 (N_43981,N_42531,N_42810);
nand U43982 (N_43982,N_42789,N_42907);
or U43983 (N_43983,N_42391,N_42268);
nand U43984 (N_43984,N_42257,N_42149);
and U43985 (N_43985,N_42235,N_42279);
or U43986 (N_43986,N_42955,N_42514);
or U43987 (N_43987,N_42020,N_42689);
or U43988 (N_43988,N_42473,N_42224);
nand U43989 (N_43989,N_42342,N_42426);
and U43990 (N_43990,N_42198,N_42418);
xnor U43991 (N_43991,N_42811,N_42599);
and U43992 (N_43992,N_42831,N_42131);
and U43993 (N_43993,N_42548,N_42590);
and U43994 (N_43994,N_42489,N_42079);
nand U43995 (N_43995,N_42611,N_42904);
nand U43996 (N_43996,N_42420,N_42670);
nand U43997 (N_43997,N_42933,N_42221);
xor U43998 (N_43998,N_42967,N_42881);
nor U43999 (N_43999,N_42284,N_42970);
or U44000 (N_44000,N_43105,N_43045);
nor U44001 (N_44001,N_43622,N_43933);
xor U44002 (N_44002,N_43230,N_43974);
or U44003 (N_44003,N_43624,N_43885);
xor U44004 (N_44004,N_43957,N_43113);
and U44005 (N_44005,N_43056,N_43851);
nor U44006 (N_44006,N_43138,N_43188);
and U44007 (N_44007,N_43048,N_43371);
nand U44008 (N_44008,N_43554,N_43961);
or U44009 (N_44009,N_43035,N_43540);
nor U44010 (N_44010,N_43183,N_43812);
and U44011 (N_44011,N_43835,N_43758);
nor U44012 (N_44012,N_43970,N_43353);
and U44013 (N_44013,N_43460,N_43401);
xor U44014 (N_44014,N_43538,N_43017);
nor U44015 (N_44015,N_43517,N_43997);
nor U44016 (N_44016,N_43968,N_43432);
and U44017 (N_44017,N_43626,N_43595);
or U44018 (N_44018,N_43257,N_43918);
or U44019 (N_44019,N_43549,N_43139);
xor U44020 (N_44020,N_43450,N_43261);
xnor U44021 (N_44021,N_43842,N_43561);
nor U44022 (N_44022,N_43516,N_43518);
nor U44023 (N_44023,N_43982,N_43279);
xnor U44024 (N_44024,N_43576,N_43133);
nor U44025 (N_44025,N_43030,N_43180);
nand U44026 (N_44026,N_43775,N_43154);
nor U44027 (N_44027,N_43208,N_43715);
nand U44028 (N_44028,N_43800,N_43345);
xnor U44029 (N_44029,N_43234,N_43370);
and U44030 (N_44030,N_43550,N_43224);
xor U44031 (N_44031,N_43608,N_43284);
nand U44032 (N_44032,N_43741,N_43125);
or U44033 (N_44033,N_43567,N_43060);
nand U44034 (N_44034,N_43011,N_43987);
or U44035 (N_44035,N_43860,N_43900);
nor U44036 (N_44036,N_43973,N_43667);
nor U44037 (N_44037,N_43964,N_43843);
nand U44038 (N_44038,N_43110,N_43569);
and U44039 (N_44039,N_43912,N_43196);
nor U44040 (N_44040,N_43453,N_43470);
and U44041 (N_44041,N_43124,N_43876);
nand U44042 (N_44042,N_43445,N_43132);
or U44043 (N_44043,N_43648,N_43267);
nand U44044 (N_44044,N_43384,N_43927);
nand U44045 (N_44045,N_43128,N_43808);
nand U44046 (N_44046,N_43013,N_43350);
and U44047 (N_44047,N_43523,N_43740);
nand U44048 (N_44048,N_43661,N_43087);
nand U44049 (N_44049,N_43612,N_43332);
nand U44050 (N_44050,N_43820,N_43906);
nand U44051 (N_44051,N_43066,N_43857);
nand U44052 (N_44052,N_43738,N_43072);
and U44053 (N_44053,N_43680,N_43043);
xor U44054 (N_44054,N_43844,N_43037);
or U44055 (N_44055,N_43052,N_43577);
and U44056 (N_44056,N_43111,N_43962);
xor U44057 (N_44057,N_43354,N_43519);
or U44058 (N_44058,N_43006,N_43206);
and U44059 (N_44059,N_43046,N_43794);
and U44060 (N_44060,N_43644,N_43995);
or U44061 (N_44061,N_43493,N_43325);
nor U44062 (N_44062,N_43189,N_43647);
and U44063 (N_44063,N_43764,N_43483);
nor U44064 (N_44064,N_43559,N_43818);
or U44065 (N_44065,N_43593,N_43191);
or U44066 (N_44066,N_43454,N_43223);
nand U44067 (N_44067,N_43341,N_43496);
nor U44068 (N_44068,N_43263,N_43435);
or U44069 (N_44069,N_43788,N_43057);
xnor U44070 (N_44070,N_43225,N_43536);
or U44071 (N_44071,N_43699,N_43032);
and U44072 (N_44072,N_43815,N_43753);
nand U44073 (N_44073,N_43481,N_43803);
and U44074 (N_44074,N_43780,N_43513);
nor U44075 (N_44075,N_43728,N_43638);
and U44076 (N_44076,N_43976,N_43315);
nand U44077 (N_44077,N_43200,N_43346);
and U44078 (N_44078,N_43362,N_43763);
xnor U44079 (N_44079,N_43091,N_43235);
xor U44080 (N_44080,N_43027,N_43630);
or U44081 (N_44081,N_43601,N_43387);
xnor U44082 (N_44082,N_43155,N_43299);
nand U44083 (N_44083,N_43891,N_43243);
or U44084 (N_44084,N_43821,N_43283);
xnor U44085 (N_44085,N_43427,N_43932);
nand U44086 (N_44086,N_43621,N_43302);
nand U44087 (N_44087,N_43407,N_43244);
and U44088 (N_44088,N_43931,N_43543);
nor U44089 (N_44089,N_43233,N_43792);
and U44090 (N_44090,N_43116,N_43218);
nor U44091 (N_44091,N_43149,N_43745);
nand U44092 (N_44092,N_43374,N_43285);
nand U44093 (N_44093,N_43838,N_43683);
nand U44094 (N_44094,N_43656,N_43102);
xor U44095 (N_44095,N_43980,N_43022);
xor U44096 (N_44096,N_43688,N_43399);
or U44097 (N_44097,N_43573,N_43274);
or U44098 (N_44098,N_43433,N_43489);
nand U44099 (N_44099,N_43028,N_43364);
nand U44100 (N_44100,N_43804,N_43190);
xnor U44101 (N_44101,N_43222,N_43275);
or U44102 (N_44102,N_43660,N_43337);
xnor U44103 (N_44103,N_43682,N_43205);
xor U44104 (N_44104,N_43239,N_43446);
nor U44105 (N_44105,N_43025,N_43534);
and U44106 (N_44106,N_43319,N_43499);
nand U44107 (N_44107,N_43107,N_43329);
nor U44108 (N_44108,N_43007,N_43358);
and U44109 (N_44109,N_43907,N_43198);
nand U44110 (N_44110,N_43458,N_43684);
or U44111 (N_44111,N_43823,N_43634);
nand U44112 (N_44112,N_43054,N_43181);
xnor U44113 (N_44113,N_43743,N_43877);
nor U44114 (N_44114,N_43598,N_43734);
and U44115 (N_44115,N_43395,N_43179);
xor U44116 (N_44116,N_43153,N_43557);
and U44117 (N_44117,N_43207,N_43832);
nand U44118 (N_44118,N_43195,N_43761);
nand U44119 (N_44119,N_43672,N_43747);
nor U44120 (N_44120,N_43340,N_43449);
or U44121 (N_44121,N_43563,N_43485);
nand U44122 (N_44122,N_43178,N_43530);
xor U44123 (N_44123,N_43498,N_43651);
or U44124 (N_44124,N_43021,N_43342);
and U44125 (N_44125,N_43751,N_43548);
and U44126 (N_44126,N_43442,N_43256);
and U44127 (N_44127,N_43571,N_43073);
nand U44128 (N_44128,N_43952,N_43905);
nand U44129 (N_44129,N_43533,N_43824);
or U44130 (N_44130,N_43739,N_43303);
nor U44131 (N_44131,N_43650,N_43908);
xor U44132 (N_44132,N_43024,N_43038);
and U44133 (N_44133,N_43524,N_43948);
nor U44134 (N_44134,N_43730,N_43100);
and U44135 (N_44135,N_43171,N_43448);
or U44136 (N_44136,N_43055,N_43400);
xor U44137 (N_44137,N_43286,N_43926);
nor U44138 (N_44138,N_43270,N_43566);
xor U44139 (N_44139,N_43978,N_43609);
nand U44140 (N_44140,N_43381,N_43920);
nor U44141 (N_44141,N_43430,N_43999);
or U44142 (N_44142,N_43542,N_43570);
and U44143 (N_44143,N_43685,N_43152);
or U44144 (N_44144,N_43439,N_43018);
or U44145 (N_44145,N_43781,N_43831);
nand U44146 (N_44146,N_43503,N_43151);
nor U44147 (N_44147,N_43867,N_43238);
xnor U44148 (N_44148,N_43869,N_43847);
nand U44149 (N_44149,N_43690,N_43164);
nand U44150 (N_44150,N_43994,N_43093);
nand U44151 (N_44151,N_43452,N_43115);
nor U44152 (N_44152,N_43352,N_43242);
or U44153 (N_44153,N_43520,N_43936);
xor U44154 (N_44154,N_43720,N_43960);
xor U44155 (N_44155,N_43491,N_43776);
nand U44156 (N_44156,N_43922,N_43036);
xnor U44157 (N_44157,N_43532,N_43678);
xnor U44158 (N_44158,N_43273,N_43785);
nand U44159 (N_44159,N_43258,N_43810);
nor U44160 (N_44160,N_43417,N_43801);
nor U44161 (N_44161,N_43248,N_43950);
and U44162 (N_44162,N_43604,N_43406);
and U44163 (N_44163,N_43975,N_43185);
nand U44164 (N_44164,N_43515,N_43061);
or U44165 (N_44165,N_43335,N_43240);
nand U44166 (N_44166,N_43969,N_43292);
and U44167 (N_44167,N_43797,N_43632);
xor U44168 (N_44168,N_43296,N_43276);
nand U44169 (N_44169,N_43689,N_43714);
nand U44170 (N_44170,N_43393,N_43361);
nand U44171 (N_44171,N_43090,N_43348);
nand U44172 (N_44172,N_43378,N_43098);
nand U44173 (N_44173,N_43527,N_43886);
and U44174 (N_44174,N_43713,N_43985);
and U44175 (N_44175,N_43349,N_43799);
or U44176 (N_44176,N_43160,N_43881);
xor U44177 (N_44177,N_43252,N_43526);
and U44178 (N_44178,N_43809,N_43525);
nand U44179 (N_44179,N_43016,N_43311);
nor U44180 (N_44180,N_43039,N_43676);
nand U44181 (N_44181,N_43408,N_43404);
nand U44182 (N_44182,N_43459,N_43707);
xnor U44183 (N_44183,N_43723,N_43537);
or U44184 (N_44184,N_43574,N_43594);
and U44185 (N_44185,N_43053,N_43615);
nand U44186 (N_44186,N_43255,N_43042);
and U44187 (N_44187,N_43123,N_43162);
xnor U44188 (N_44188,N_43210,N_43323);
xnor U44189 (N_44189,N_43122,N_43423);
nand U44190 (N_44190,N_43898,N_43896);
or U44191 (N_44191,N_43836,N_43883);
xor U44192 (N_44192,N_43865,N_43431);
nor U44193 (N_44193,N_43783,N_43703);
and U44194 (N_44194,N_43318,N_43941);
or U44195 (N_44195,N_43635,N_43589);
nand U44196 (N_44196,N_43500,N_43558);
or U44197 (N_44197,N_43760,N_43373);
xnor U44198 (N_44198,N_43888,N_43071);
nand U44199 (N_44199,N_43597,N_43646);
xor U44200 (N_44200,N_43878,N_43009);
and U44201 (N_44201,N_43848,N_43958);
nor U44202 (N_44202,N_43471,N_43484);
xnor U44203 (N_44203,N_43586,N_43778);
and U44204 (N_44204,N_43953,N_43089);
and U44205 (N_44205,N_43663,N_43963);
or U44206 (N_44206,N_43117,N_43031);
and U44207 (N_44207,N_43861,N_43592);
nor U44208 (N_44208,N_43456,N_43895);
or U44209 (N_44209,N_43157,N_43590);
xor U44210 (N_44210,N_43165,N_43547);
and U44211 (N_44211,N_43509,N_43405);
or U44212 (N_44212,N_43451,N_43686);
or U44213 (N_44213,N_43610,N_43972);
or U44214 (N_44214,N_43677,N_43514);
nor U44215 (N_44215,N_43717,N_43029);
nand U44216 (N_44216,N_43790,N_43575);
nand U44217 (N_44217,N_43119,N_43217);
or U44218 (N_44218,N_43000,N_43382);
nor U44219 (N_44219,N_43864,N_43879);
or U44220 (N_44220,N_43347,N_43560);
xor U44221 (N_44221,N_43137,N_43837);
xor U44222 (N_44222,N_43892,N_43159);
or U44223 (N_44223,N_43639,N_43001);
nand U44224 (N_44224,N_43623,N_43786);
xnor U44225 (N_44225,N_43902,N_43981);
and U44226 (N_44226,N_43856,N_43033);
and U44227 (N_44227,N_43120,N_43236);
xnor U44228 (N_44228,N_43587,N_43288);
or U44229 (N_44229,N_43805,N_43546);
nand U44230 (N_44230,N_43817,N_43965);
xor U44231 (N_44231,N_43736,N_43194);
xor U44232 (N_44232,N_43798,N_43356);
and U44233 (N_44233,N_43203,N_43913);
nor U44234 (N_44234,N_43437,N_43897);
or U44235 (N_44235,N_43331,N_43398);
nor U44236 (N_44236,N_43840,N_43658);
and U44237 (N_44237,N_43187,N_43814);
nand U44238 (N_44238,N_43394,N_43939);
and U44239 (N_44239,N_43182,N_43979);
or U44240 (N_44240,N_43923,N_43784);
nand U44241 (N_44241,N_43625,N_43099);
nor U44242 (N_44242,N_43641,N_43619);
nor U44243 (N_44243,N_43079,N_43146);
or U44244 (N_44244,N_43993,N_43330);
nand U44245 (N_44245,N_43849,N_43725);
nand U44246 (N_44246,N_43887,N_43167);
or U44247 (N_44247,N_43868,N_43403);
xor U44248 (N_44248,N_43556,N_43919);
nor U44249 (N_44249,N_43769,N_43578);
or U44250 (N_44250,N_43768,N_43679);
xor U44251 (N_44251,N_43938,N_43260);
nor U44252 (N_44252,N_43825,N_43946);
nor U44253 (N_44253,N_43213,N_43705);
nor U44254 (N_44254,N_43322,N_43893);
xnor U44255 (N_44255,N_43562,N_43476);
nor U44256 (N_44256,N_43301,N_43724);
and U44257 (N_44257,N_43568,N_43305);
nand U44258 (N_44258,N_43482,N_43265);
xnor U44259 (N_44259,N_43507,N_43718);
xor U44260 (N_44260,N_43280,N_43565);
nor U44261 (N_44261,N_43637,N_43695);
or U44262 (N_44262,N_43771,N_43426);
nand U44263 (N_44263,N_43461,N_43034);
nor U44264 (N_44264,N_43614,N_43246);
nand U44265 (N_44265,N_43068,N_43748);
and U44266 (N_44266,N_43700,N_43872);
or U44267 (N_44267,N_43492,N_43334);
nand U44268 (N_44268,N_43416,N_43343);
nor U44269 (N_44269,N_43959,N_43134);
or U44270 (N_44270,N_43304,N_43464);
xnor U44271 (N_44271,N_43620,N_43522);
nand U44272 (N_44272,N_43954,N_43062);
and U44273 (N_44273,N_43161,N_43924);
and U44274 (N_44274,N_43226,N_43219);
nor U44275 (N_44275,N_43126,N_43854);
nand U44276 (N_44276,N_43521,N_43441);
xor U44277 (N_44277,N_43067,N_43177);
nor U44278 (N_44278,N_43019,N_43990);
nand U44279 (N_44279,N_43584,N_43074);
and U44280 (N_44280,N_43793,N_43142);
xnor U44281 (N_44281,N_43147,N_43465);
nor U44282 (N_44282,N_43163,N_43169);
nand U44283 (N_44283,N_43173,N_43511);
or U44284 (N_44284,N_43654,N_43585);
nand U44285 (N_44285,N_43468,N_43581);
nor U44286 (N_44286,N_43106,N_43752);
or U44287 (N_44287,N_43135,N_43497);
xor U44288 (N_44288,N_43710,N_43321);
nand U44289 (N_44289,N_43469,N_43086);
and U44290 (N_44290,N_43429,N_43859);
or U44291 (N_44291,N_43834,N_43649);
nand U44292 (N_44292,N_43731,N_43657);
xnor U44293 (N_44293,N_43702,N_43040);
nor U44294 (N_44294,N_43297,N_43773);
nor U44295 (N_44295,N_43064,N_43419);
or U44296 (N_44296,N_43708,N_43186);
nor U44297 (N_44297,N_43653,N_43541);
and U44298 (N_44298,N_43420,N_43599);
nor U44299 (N_44299,N_43313,N_43050);
xnor U44300 (N_44300,N_43691,N_43505);
or U44301 (N_44301,N_43366,N_43145);
xor U44302 (N_44302,N_43827,N_43044);
and U44303 (N_44303,N_43228,N_43262);
nor U44304 (N_44304,N_43490,N_43192);
nor U44305 (N_44305,N_43320,N_43076);
or U44306 (N_44306,N_43121,N_43618);
and U44307 (N_44307,N_43884,N_43508);
nor U44308 (N_44308,N_43457,N_43291);
or U44309 (N_44309,N_43967,N_43212);
nor U44310 (N_44310,N_43069,N_43360);
or U44311 (N_44311,N_43202,N_43108);
or U44312 (N_44312,N_43041,N_43921);
nand U44313 (N_44313,N_43855,N_43298);
and U44314 (N_44314,N_43669,N_43328);
nand U44315 (N_44315,N_43277,N_43531);
or U44316 (N_44316,N_43294,N_43026);
nand U44317 (N_44317,N_43097,N_43081);
nor U44318 (N_44318,N_43380,N_43983);
or U44319 (N_44319,N_43455,N_43310);
or U44320 (N_44320,N_43480,N_43940);
nor U44321 (N_44321,N_43813,N_43101);
xor U44322 (N_44322,N_43986,N_43357);
and U44323 (N_44323,N_43487,N_43992);
and U44324 (N_44324,N_43338,N_43909);
nand U44325 (N_44325,N_43766,N_43796);
xnor U44326 (N_44326,N_43424,N_43698);
xor U44327 (N_44327,N_43929,N_43627);
nor U44328 (N_44328,N_43379,N_43237);
xnor U44329 (N_44329,N_43103,N_43600);
and U44330 (N_44330,N_43949,N_43479);
or U44331 (N_44331,N_43529,N_43158);
and U44332 (N_44332,N_43616,N_43966);
or U44333 (N_44333,N_43716,N_43080);
xnor U44334 (N_44334,N_43065,N_43652);
xor U44335 (N_44335,N_43308,N_43726);
nand U44336 (N_44336,N_43984,N_43383);
and U44337 (N_44337,N_43211,N_43247);
nand U44338 (N_44338,N_43579,N_43673);
and U44339 (N_44339,N_43670,N_43118);
or U44340 (N_44340,N_43369,N_43392);
nor U44341 (N_44341,N_43324,N_43942);
or U44342 (N_44342,N_43853,N_43944);
or U44343 (N_44343,N_43735,N_43882);
or U44344 (N_44344,N_43862,N_43762);
and U44345 (N_44345,N_43774,N_43681);
xnor U44346 (N_44346,N_43082,N_43359);
xnor U44347 (N_44347,N_43693,N_43306);
or U44348 (N_44348,N_43588,N_43870);
and U44349 (N_44349,N_43023,N_43339);
or U44350 (N_44350,N_43282,N_43839);
xor U44351 (N_44351,N_43414,N_43826);
nor U44352 (N_44352,N_43271,N_43757);
xnor U44353 (N_44353,N_43692,N_43910);
or U44354 (N_44354,N_43628,N_43396);
and U44355 (N_44355,N_43911,N_43436);
or U44356 (N_44356,N_43174,N_43943);
or U44357 (N_44357,N_43737,N_43789);
xnor U44358 (N_44358,N_43372,N_43596);
nor U44359 (N_44359,N_43004,N_43659);
or U44360 (N_44360,N_43486,N_43863);
and U44361 (N_44361,N_43755,N_43020);
nand U44362 (N_44362,N_43894,N_43934);
nand U44363 (N_44363,N_43201,N_43216);
and U44364 (N_44364,N_43421,N_43742);
or U44365 (N_44365,N_43197,N_43841);
nand U44366 (N_44366,N_43049,N_43150);
nand U44367 (N_44367,N_43871,N_43591);
or U44368 (N_44368,N_43114,N_43309);
or U44369 (N_44369,N_43925,N_43807);
or U44370 (N_44370,N_43172,N_43156);
xor U44371 (N_44371,N_43607,N_43259);
xor U44372 (N_44372,N_43991,N_43336);
or U44373 (N_44373,N_43719,N_43890);
or U44374 (N_44374,N_43996,N_43665);
and U44375 (N_44375,N_43687,N_43051);
xor U44376 (N_44376,N_43444,N_43852);
or U44377 (N_44377,N_43377,N_43175);
or U44378 (N_44378,N_43643,N_43209);
nand U44379 (N_44379,N_43935,N_43367);
and U44380 (N_44380,N_43666,N_43830);
and U44381 (N_44381,N_43333,N_43148);
xor U44382 (N_44382,N_43129,N_43088);
nand U44383 (N_44383,N_43750,N_43951);
nor U44384 (N_44384,N_43928,N_43010);
nand U44385 (N_44385,N_43096,N_43312);
nand U44386 (N_44386,N_43409,N_43552);
nand U44387 (N_44387,N_43440,N_43811);
xor U44388 (N_44388,N_43822,N_43866);
nor U44389 (N_44389,N_43502,N_43300);
or U44390 (N_44390,N_43386,N_43447);
or U44391 (N_44391,N_43903,N_43014);
xnor U44392 (N_44392,N_43916,N_43389);
nand U44393 (N_44393,N_43008,N_43316);
nand U44394 (N_44394,N_43795,N_43845);
xnor U44395 (N_44395,N_43744,N_43415);
nor U44396 (N_44396,N_43095,N_43402);
xor U44397 (N_44397,N_43711,N_43241);
nor U44398 (N_44398,N_43528,N_43988);
nand U44399 (N_44399,N_43144,N_43215);
nor U44400 (N_44400,N_43281,N_43474);
or U44401 (N_44401,N_43729,N_43112);
nand U44402 (N_44402,N_43221,N_43606);
and U44403 (N_44403,N_43278,N_43874);
nor U44404 (N_44404,N_43229,N_43477);
and U44405 (N_44405,N_43858,N_43472);
and U44406 (N_44406,N_43184,N_43955);
nand U44407 (N_44407,N_43140,N_43272);
nor U44408 (N_44408,N_43582,N_43756);
nand U44409 (N_44409,N_43880,N_43268);
or U44410 (N_44410,N_43251,N_43553);
nand U44411 (N_44411,N_43344,N_43914);
and U44412 (N_44412,N_43782,N_43015);
nor U44413 (N_44413,N_43494,N_43058);
or U44414 (N_44414,N_43722,N_43617);
xor U44415 (N_44415,N_43603,N_43231);
and U44416 (N_44416,N_43662,N_43754);
nand U44417 (N_44417,N_43873,N_43697);
or U44418 (N_44418,N_43204,N_43410);
xnor U44419 (N_44419,N_43136,N_43443);
and U44420 (N_44420,N_43668,N_43674);
or U44421 (N_44421,N_43463,N_43168);
or U44422 (N_44422,N_43506,N_43307);
nor U44423 (N_44423,N_43732,N_43193);
or U44424 (N_44424,N_43078,N_43478);
xnor U44425 (N_44425,N_43629,N_43535);
nor U44426 (N_44426,N_43696,N_43438);
or U44427 (N_44427,N_43390,N_43249);
nand U44428 (N_44428,N_43413,N_43539);
xor U44429 (N_44429,N_43411,N_43850);
and U44430 (N_44430,N_43351,N_43376);
nand U44431 (N_44431,N_43293,N_43326);
and U44432 (N_44432,N_43232,N_43388);
nand U44433 (N_44433,N_43846,N_43901);
xnor U44434 (N_44434,N_43545,N_43564);
nor U44435 (N_44435,N_43462,N_43806);
nor U44436 (N_44436,N_43613,N_43937);
nand U44437 (N_44437,N_43675,N_43904);
or U44438 (N_44438,N_43130,N_43504);
xnor U44439 (N_44439,N_43645,N_43363);
and U44440 (N_44440,N_43802,N_43572);
nand U44441 (N_44441,N_43706,N_43269);
nor U44442 (N_44442,N_43671,N_43290);
nor U44443 (N_44443,N_43250,N_43544);
xor U44444 (N_44444,N_43664,N_43495);
xnor U44445 (N_44445,N_43109,N_43214);
xnor U44446 (N_44446,N_43131,N_43295);
or U44447 (N_44447,N_43829,N_43059);
xnor U44448 (N_44448,N_43428,N_43727);
or U44449 (N_44449,N_43989,N_43759);
or U44450 (N_44450,N_43875,N_43166);
xor U44451 (N_44451,N_43083,N_43749);
or U44452 (N_44452,N_43501,N_43475);
xor U44453 (N_44453,N_43510,N_43085);
or U44454 (N_44454,N_43003,N_43767);
xor U44455 (N_44455,N_43791,N_43075);
xor U44456 (N_44456,N_43012,N_43104);
or U44457 (N_44457,N_43746,N_43473);
nor U44458 (N_44458,N_43816,N_43287);
xor U44459 (N_44459,N_43220,N_43998);
and U44460 (N_44460,N_43092,N_43170);
and U44461 (N_44461,N_43327,N_43289);
xnor U44462 (N_44462,N_43712,N_43945);
nand U44463 (N_44463,N_43047,N_43772);
nor U44464 (N_44464,N_43245,N_43787);
xor U44465 (N_44465,N_43412,N_43956);
and U44466 (N_44466,N_43694,N_43094);
or U44467 (N_44467,N_43077,N_43397);
xnor U44468 (N_44468,N_43733,N_43930);
nand U44469 (N_44469,N_43947,N_43779);
nor U44470 (N_44470,N_43611,N_43434);
xnor U44471 (N_44471,N_43070,N_43709);
or U44472 (N_44472,N_43602,N_43005);
and U44473 (N_44473,N_43143,N_43467);
xor U44474 (N_44474,N_43899,N_43375);
nor U44475 (N_44475,N_43917,N_43317);
nor U44476 (N_44476,N_43254,N_43889);
nor U44477 (N_44477,N_43355,N_43580);
nand U44478 (N_44478,N_43199,N_43770);
or U44479 (N_44479,N_43176,N_43512);
or U44480 (N_44480,N_43127,N_43642);
nand U44481 (N_44481,N_43425,N_43551);
nor U44482 (N_44482,N_43368,N_43063);
or U44483 (N_44483,N_43253,N_43701);
xor U44484 (N_44484,N_43365,N_43977);
xnor U44485 (N_44485,N_43819,N_43314);
or U44486 (N_44486,N_43141,N_43828);
and U44487 (N_44487,N_43765,N_43488);
nor U44488 (N_44488,N_43631,N_43227);
xor U44489 (N_44489,N_43583,N_43633);
or U44490 (N_44490,N_43640,N_43915);
and U44491 (N_44491,N_43002,N_43264);
nand U44492 (N_44492,N_43704,N_43636);
nor U44493 (N_44493,N_43418,N_43385);
xor U44494 (N_44494,N_43971,N_43266);
nand U44495 (N_44495,N_43466,N_43833);
nor U44496 (N_44496,N_43605,N_43391);
xor U44497 (N_44497,N_43777,N_43084);
or U44498 (N_44498,N_43721,N_43422);
and U44499 (N_44499,N_43555,N_43655);
or U44500 (N_44500,N_43248,N_43097);
nor U44501 (N_44501,N_43450,N_43648);
xnor U44502 (N_44502,N_43052,N_43676);
xnor U44503 (N_44503,N_43162,N_43187);
nor U44504 (N_44504,N_43436,N_43943);
xnor U44505 (N_44505,N_43293,N_43922);
nor U44506 (N_44506,N_43842,N_43490);
nor U44507 (N_44507,N_43044,N_43843);
nand U44508 (N_44508,N_43158,N_43344);
nand U44509 (N_44509,N_43546,N_43572);
nor U44510 (N_44510,N_43156,N_43175);
or U44511 (N_44511,N_43962,N_43475);
and U44512 (N_44512,N_43075,N_43971);
or U44513 (N_44513,N_43507,N_43174);
nor U44514 (N_44514,N_43469,N_43821);
xor U44515 (N_44515,N_43233,N_43661);
nor U44516 (N_44516,N_43982,N_43795);
or U44517 (N_44517,N_43820,N_43750);
and U44518 (N_44518,N_43323,N_43408);
xor U44519 (N_44519,N_43133,N_43878);
nor U44520 (N_44520,N_43484,N_43672);
or U44521 (N_44521,N_43783,N_43388);
nor U44522 (N_44522,N_43491,N_43355);
xnor U44523 (N_44523,N_43862,N_43230);
xnor U44524 (N_44524,N_43482,N_43780);
or U44525 (N_44525,N_43912,N_43132);
xor U44526 (N_44526,N_43818,N_43386);
or U44527 (N_44527,N_43860,N_43103);
nand U44528 (N_44528,N_43892,N_43499);
and U44529 (N_44529,N_43987,N_43630);
nand U44530 (N_44530,N_43937,N_43122);
and U44531 (N_44531,N_43854,N_43919);
nor U44532 (N_44532,N_43568,N_43953);
and U44533 (N_44533,N_43325,N_43177);
xnor U44534 (N_44534,N_43657,N_43554);
nand U44535 (N_44535,N_43627,N_43886);
nand U44536 (N_44536,N_43627,N_43041);
nand U44537 (N_44537,N_43972,N_43213);
and U44538 (N_44538,N_43936,N_43025);
and U44539 (N_44539,N_43551,N_43834);
or U44540 (N_44540,N_43772,N_43751);
and U44541 (N_44541,N_43318,N_43528);
nand U44542 (N_44542,N_43844,N_43032);
or U44543 (N_44543,N_43711,N_43879);
or U44544 (N_44544,N_43289,N_43897);
nor U44545 (N_44545,N_43193,N_43174);
xnor U44546 (N_44546,N_43016,N_43509);
nand U44547 (N_44547,N_43589,N_43365);
nor U44548 (N_44548,N_43547,N_43532);
xor U44549 (N_44549,N_43744,N_43215);
xnor U44550 (N_44550,N_43758,N_43060);
nand U44551 (N_44551,N_43900,N_43684);
xnor U44552 (N_44552,N_43369,N_43017);
xor U44553 (N_44553,N_43321,N_43536);
and U44554 (N_44554,N_43620,N_43035);
or U44555 (N_44555,N_43041,N_43168);
nor U44556 (N_44556,N_43318,N_43413);
xnor U44557 (N_44557,N_43548,N_43901);
or U44558 (N_44558,N_43490,N_43117);
and U44559 (N_44559,N_43365,N_43785);
xor U44560 (N_44560,N_43294,N_43518);
nand U44561 (N_44561,N_43848,N_43172);
xnor U44562 (N_44562,N_43981,N_43267);
or U44563 (N_44563,N_43822,N_43496);
or U44564 (N_44564,N_43938,N_43409);
or U44565 (N_44565,N_43688,N_43922);
xor U44566 (N_44566,N_43687,N_43279);
nor U44567 (N_44567,N_43945,N_43289);
nand U44568 (N_44568,N_43440,N_43325);
or U44569 (N_44569,N_43561,N_43662);
nand U44570 (N_44570,N_43882,N_43472);
and U44571 (N_44571,N_43285,N_43556);
nand U44572 (N_44572,N_43348,N_43610);
xnor U44573 (N_44573,N_43482,N_43223);
and U44574 (N_44574,N_43184,N_43931);
and U44575 (N_44575,N_43055,N_43892);
nor U44576 (N_44576,N_43373,N_43110);
nor U44577 (N_44577,N_43432,N_43372);
nand U44578 (N_44578,N_43810,N_43194);
nor U44579 (N_44579,N_43993,N_43960);
or U44580 (N_44580,N_43645,N_43931);
or U44581 (N_44581,N_43446,N_43881);
or U44582 (N_44582,N_43367,N_43144);
and U44583 (N_44583,N_43070,N_43086);
xor U44584 (N_44584,N_43057,N_43472);
xor U44585 (N_44585,N_43124,N_43050);
nand U44586 (N_44586,N_43572,N_43083);
nand U44587 (N_44587,N_43821,N_43490);
and U44588 (N_44588,N_43805,N_43752);
xnor U44589 (N_44589,N_43682,N_43313);
nand U44590 (N_44590,N_43160,N_43788);
or U44591 (N_44591,N_43441,N_43306);
or U44592 (N_44592,N_43662,N_43680);
nand U44593 (N_44593,N_43302,N_43221);
or U44594 (N_44594,N_43646,N_43944);
or U44595 (N_44595,N_43641,N_43511);
or U44596 (N_44596,N_43415,N_43764);
and U44597 (N_44597,N_43733,N_43418);
or U44598 (N_44598,N_43372,N_43028);
or U44599 (N_44599,N_43167,N_43718);
xnor U44600 (N_44600,N_43639,N_43764);
or U44601 (N_44601,N_43989,N_43296);
or U44602 (N_44602,N_43299,N_43258);
nor U44603 (N_44603,N_43972,N_43781);
xor U44604 (N_44604,N_43906,N_43034);
nand U44605 (N_44605,N_43931,N_43488);
xor U44606 (N_44606,N_43413,N_43937);
nor U44607 (N_44607,N_43544,N_43984);
nand U44608 (N_44608,N_43244,N_43723);
and U44609 (N_44609,N_43543,N_43332);
nand U44610 (N_44610,N_43073,N_43767);
xnor U44611 (N_44611,N_43989,N_43289);
and U44612 (N_44612,N_43683,N_43982);
nor U44613 (N_44613,N_43656,N_43335);
and U44614 (N_44614,N_43340,N_43719);
xnor U44615 (N_44615,N_43172,N_43147);
nand U44616 (N_44616,N_43410,N_43611);
xor U44617 (N_44617,N_43055,N_43874);
or U44618 (N_44618,N_43633,N_43301);
nand U44619 (N_44619,N_43461,N_43096);
xor U44620 (N_44620,N_43231,N_43033);
nor U44621 (N_44621,N_43566,N_43426);
and U44622 (N_44622,N_43575,N_43665);
nor U44623 (N_44623,N_43780,N_43245);
xor U44624 (N_44624,N_43403,N_43027);
nand U44625 (N_44625,N_43646,N_43126);
nor U44626 (N_44626,N_43664,N_43168);
and U44627 (N_44627,N_43957,N_43787);
and U44628 (N_44628,N_43581,N_43042);
or U44629 (N_44629,N_43131,N_43362);
nand U44630 (N_44630,N_43003,N_43018);
nand U44631 (N_44631,N_43933,N_43524);
nand U44632 (N_44632,N_43659,N_43870);
nand U44633 (N_44633,N_43557,N_43953);
and U44634 (N_44634,N_43329,N_43471);
nand U44635 (N_44635,N_43257,N_43333);
nor U44636 (N_44636,N_43016,N_43767);
nor U44637 (N_44637,N_43349,N_43750);
nor U44638 (N_44638,N_43529,N_43938);
nor U44639 (N_44639,N_43414,N_43478);
nor U44640 (N_44640,N_43642,N_43774);
nand U44641 (N_44641,N_43311,N_43634);
nor U44642 (N_44642,N_43651,N_43363);
nor U44643 (N_44643,N_43568,N_43240);
xor U44644 (N_44644,N_43470,N_43682);
or U44645 (N_44645,N_43822,N_43043);
nor U44646 (N_44646,N_43879,N_43635);
and U44647 (N_44647,N_43565,N_43302);
and U44648 (N_44648,N_43100,N_43285);
xor U44649 (N_44649,N_43557,N_43998);
nand U44650 (N_44650,N_43041,N_43448);
nor U44651 (N_44651,N_43697,N_43342);
nor U44652 (N_44652,N_43924,N_43847);
xnor U44653 (N_44653,N_43581,N_43191);
nor U44654 (N_44654,N_43067,N_43342);
xnor U44655 (N_44655,N_43440,N_43976);
or U44656 (N_44656,N_43223,N_43604);
and U44657 (N_44657,N_43283,N_43800);
and U44658 (N_44658,N_43739,N_43814);
nor U44659 (N_44659,N_43488,N_43697);
or U44660 (N_44660,N_43790,N_43023);
nor U44661 (N_44661,N_43602,N_43029);
nand U44662 (N_44662,N_43837,N_43541);
nor U44663 (N_44663,N_43529,N_43902);
nor U44664 (N_44664,N_43098,N_43109);
xor U44665 (N_44665,N_43337,N_43102);
nand U44666 (N_44666,N_43971,N_43367);
nor U44667 (N_44667,N_43050,N_43241);
nand U44668 (N_44668,N_43028,N_43593);
nand U44669 (N_44669,N_43062,N_43201);
or U44670 (N_44670,N_43500,N_43878);
nor U44671 (N_44671,N_43155,N_43772);
nand U44672 (N_44672,N_43128,N_43026);
and U44673 (N_44673,N_43290,N_43986);
nor U44674 (N_44674,N_43979,N_43037);
nand U44675 (N_44675,N_43426,N_43833);
xnor U44676 (N_44676,N_43640,N_43723);
nand U44677 (N_44677,N_43896,N_43146);
nand U44678 (N_44678,N_43687,N_43990);
xnor U44679 (N_44679,N_43058,N_43902);
xnor U44680 (N_44680,N_43443,N_43890);
nand U44681 (N_44681,N_43604,N_43640);
nor U44682 (N_44682,N_43498,N_43446);
or U44683 (N_44683,N_43489,N_43083);
xnor U44684 (N_44684,N_43316,N_43304);
and U44685 (N_44685,N_43608,N_43253);
nor U44686 (N_44686,N_43443,N_43727);
nor U44687 (N_44687,N_43572,N_43408);
xnor U44688 (N_44688,N_43609,N_43418);
or U44689 (N_44689,N_43259,N_43267);
nor U44690 (N_44690,N_43440,N_43019);
or U44691 (N_44691,N_43078,N_43447);
nand U44692 (N_44692,N_43535,N_43305);
and U44693 (N_44693,N_43436,N_43438);
xor U44694 (N_44694,N_43300,N_43623);
and U44695 (N_44695,N_43960,N_43154);
or U44696 (N_44696,N_43215,N_43374);
or U44697 (N_44697,N_43793,N_43590);
or U44698 (N_44698,N_43049,N_43977);
nand U44699 (N_44699,N_43662,N_43995);
nor U44700 (N_44700,N_43731,N_43270);
nand U44701 (N_44701,N_43897,N_43132);
nor U44702 (N_44702,N_43364,N_43424);
xor U44703 (N_44703,N_43893,N_43094);
or U44704 (N_44704,N_43952,N_43333);
and U44705 (N_44705,N_43015,N_43421);
xnor U44706 (N_44706,N_43442,N_43066);
nor U44707 (N_44707,N_43511,N_43009);
xor U44708 (N_44708,N_43945,N_43755);
xor U44709 (N_44709,N_43944,N_43436);
nor U44710 (N_44710,N_43502,N_43963);
nand U44711 (N_44711,N_43958,N_43702);
and U44712 (N_44712,N_43799,N_43035);
nor U44713 (N_44713,N_43633,N_43051);
nand U44714 (N_44714,N_43273,N_43936);
nand U44715 (N_44715,N_43841,N_43086);
or U44716 (N_44716,N_43826,N_43092);
or U44717 (N_44717,N_43938,N_43255);
xor U44718 (N_44718,N_43727,N_43875);
xnor U44719 (N_44719,N_43770,N_43643);
nor U44720 (N_44720,N_43535,N_43224);
or U44721 (N_44721,N_43612,N_43400);
and U44722 (N_44722,N_43281,N_43638);
nor U44723 (N_44723,N_43712,N_43012);
or U44724 (N_44724,N_43386,N_43663);
or U44725 (N_44725,N_43667,N_43112);
xor U44726 (N_44726,N_43986,N_43177);
xnor U44727 (N_44727,N_43050,N_43309);
nand U44728 (N_44728,N_43854,N_43700);
or U44729 (N_44729,N_43458,N_43683);
and U44730 (N_44730,N_43305,N_43778);
or U44731 (N_44731,N_43556,N_43212);
xnor U44732 (N_44732,N_43239,N_43044);
or U44733 (N_44733,N_43338,N_43980);
xor U44734 (N_44734,N_43278,N_43204);
and U44735 (N_44735,N_43786,N_43736);
nand U44736 (N_44736,N_43572,N_43652);
xnor U44737 (N_44737,N_43645,N_43924);
nor U44738 (N_44738,N_43042,N_43843);
nor U44739 (N_44739,N_43865,N_43777);
or U44740 (N_44740,N_43745,N_43988);
and U44741 (N_44741,N_43007,N_43295);
nor U44742 (N_44742,N_43400,N_43821);
xor U44743 (N_44743,N_43554,N_43601);
nor U44744 (N_44744,N_43986,N_43819);
nand U44745 (N_44745,N_43690,N_43316);
and U44746 (N_44746,N_43963,N_43885);
and U44747 (N_44747,N_43992,N_43978);
or U44748 (N_44748,N_43203,N_43457);
nor U44749 (N_44749,N_43837,N_43330);
nor U44750 (N_44750,N_43914,N_43064);
nor U44751 (N_44751,N_43830,N_43524);
xor U44752 (N_44752,N_43702,N_43453);
nand U44753 (N_44753,N_43771,N_43950);
nand U44754 (N_44754,N_43419,N_43764);
nand U44755 (N_44755,N_43772,N_43480);
xnor U44756 (N_44756,N_43224,N_43218);
or U44757 (N_44757,N_43460,N_43547);
nor U44758 (N_44758,N_43019,N_43681);
and U44759 (N_44759,N_43533,N_43063);
nor U44760 (N_44760,N_43186,N_43477);
nor U44761 (N_44761,N_43360,N_43991);
or U44762 (N_44762,N_43652,N_43925);
nor U44763 (N_44763,N_43752,N_43147);
or U44764 (N_44764,N_43665,N_43912);
and U44765 (N_44765,N_43172,N_43540);
and U44766 (N_44766,N_43950,N_43503);
nand U44767 (N_44767,N_43673,N_43942);
xor U44768 (N_44768,N_43169,N_43903);
or U44769 (N_44769,N_43340,N_43872);
nand U44770 (N_44770,N_43112,N_43411);
nor U44771 (N_44771,N_43182,N_43953);
and U44772 (N_44772,N_43374,N_43549);
and U44773 (N_44773,N_43963,N_43805);
and U44774 (N_44774,N_43092,N_43767);
or U44775 (N_44775,N_43110,N_43626);
nand U44776 (N_44776,N_43422,N_43927);
and U44777 (N_44777,N_43595,N_43049);
and U44778 (N_44778,N_43521,N_43092);
nor U44779 (N_44779,N_43337,N_43117);
nand U44780 (N_44780,N_43457,N_43811);
or U44781 (N_44781,N_43907,N_43137);
nand U44782 (N_44782,N_43650,N_43827);
nand U44783 (N_44783,N_43902,N_43280);
nor U44784 (N_44784,N_43295,N_43363);
nor U44785 (N_44785,N_43914,N_43101);
xnor U44786 (N_44786,N_43525,N_43854);
xor U44787 (N_44787,N_43155,N_43179);
nor U44788 (N_44788,N_43178,N_43776);
xor U44789 (N_44789,N_43216,N_43849);
xor U44790 (N_44790,N_43026,N_43526);
and U44791 (N_44791,N_43714,N_43566);
nor U44792 (N_44792,N_43991,N_43066);
nor U44793 (N_44793,N_43477,N_43943);
xnor U44794 (N_44794,N_43848,N_43157);
and U44795 (N_44795,N_43931,N_43377);
nand U44796 (N_44796,N_43509,N_43334);
and U44797 (N_44797,N_43470,N_43895);
xnor U44798 (N_44798,N_43029,N_43479);
nand U44799 (N_44799,N_43713,N_43915);
xor U44800 (N_44800,N_43254,N_43074);
or U44801 (N_44801,N_43976,N_43356);
or U44802 (N_44802,N_43814,N_43881);
nor U44803 (N_44803,N_43633,N_43153);
nor U44804 (N_44804,N_43707,N_43098);
xor U44805 (N_44805,N_43059,N_43585);
or U44806 (N_44806,N_43343,N_43559);
and U44807 (N_44807,N_43579,N_43931);
and U44808 (N_44808,N_43020,N_43690);
nor U44809 (N_44809,N_43498,N_43568);
nand U44810 (N_44810,N_43096,N_43514);
nand U44811 (N_44811,N_43063,N_43967);
and U44812 (N_44812,N_43976,N_43114);
and U44813 (N_44813,N_43677,N_43203);
or U44814 (N_44814,N_43956,N_43318);
nor U44815 (N_44815,N_43541,N_43701);
and U44816 (N_44816,N_43150,N_43358);
nand U44817 (N_44817,N_43188,N_43526);
xnor U44818 (N_44818,N_43362,N_43523);
and U44819 (N_44819,N_43740,N_43787);
nand U44820 (N_44820,N_43079,N_43230);
nand U44821 (N_44821,N_43541,N_43778);
nor U44822 (N_44822,N_43654,N_43694);
nor U44823 (N_44823,N_43894,N_43177);
and U44824 (N_44824,N_43038,N_43864);
nor U44825 (N_44825,N_43246,N_43574);
nand U44826 (N_44826,N_43304,N_43586);
nor U44827 (N_44827,N_43037,N_43835);
or U44828 (N_44828,N_43184,N_43276);
nand U44829 (N_44829,N_43258,N_43797);
or U44830 (N_44830,N_43555,N_43977);
or U44831 (N_44831,N_43895,N_43730);
nand U44832 (N_44832,N_43338,N_43315);
nand U44833 (N_44833,N_43092,N_43094);
xor U44834 (N_44834,N_43223,N_43739);
and U44835 (N_44835,N_43047,N_43926);
nand U44836 (N_44836,N_43597,N_43768);
nand U44837 (N_44837,N_43365,N_43653);
xnor U44838 (N_44838,N_43800,N_43447);
nand U44839 (N_44839,N_43294,N_43468);
and U44840 (N_44840,N_43042,N_43238);
nor U44841 (N_44841,N_43482,N_43028);
and U44842 (N_44842,N_43930,N_43457);
or U44843 (N_44843,N_43057,N_43557);
nand U44844 (N_44844,N_43533,N_43632);
and U44845 (N_44845,N_43990,N_43895);
or U44846 (N_44846,N_43887,N_43873);
xnor U44847 (N_44847,N_43279,N_43648);
nand U44848 (N_44848,N_43354,N_43689);
nor U44849 (N_44849,N_43540,N_43282);
nor U44850 (N_44850,N_43150,N_43428);
nand U44851 (N_44851,N_43402,N_43250);
and U44852 (N_44852,N_43310,N_43643);
nor U44853 (N_44853,N_43398,N_43760);
xor U44854 (N_44854,N_43463,N_43531);
nand U44855 (N_44855,N_43757,N_43851);
nor U44856 (N_44856,N_43883,N_43988);
nor U44857 (N_44857,N_43777,N_43508);
nor U44858 (N_44858,N_43474,N_43044);
and U44859 (N_44859,N_43392,N_43628);
or U44860 (N_44860,N_43431,N_43286);
and U44861 (N_44861,N_43973,N_43326);
nor U44862 (N_44862,N_43034,N_43193);
and U44863 (N_44863,N_43514,N_43477);
nand U44864 (N_44864,N_43580,N_43296);
nand U44865 (N_44865,N_43185,N_43802);
and U44866 (N_44866,N_43777,N_43111);
or U44867 (N_44867,N_43120,N_43054);
xor U44868 (N_44868,N_43461,N_43788);
or U44869 (N_44869,N_43737,N_43906);
or U44870 (N_44870,N_43035,N_43636);
nand U44871 (N_44871,N_43465,N_43984);
or U44872 (N_44872,N_43294,N_43786);
nand U44873 (N_44873,N_43643,N_43975);
or U44874 (N_44874,N_43271,N_43302);
nand U44875 (N_44875,N_43631,N_43968);
nor U44876 (N_44876,N_43890,N_43517);
and U44877 (N_44877,N_43168,N_43534);
xor U44878 (N_44878,N_43535,N_43557);
nand U44879 (N_44879,N_43731,N_43071);
or U44880 (N_44880,N_43389,N_43950);
xor U44881 (N_44881,N_43182,N_43787);
nor U44882 (N_44882,N_43194,N_43921);
xnor U44883 (N_44883,N_43290,N_43305);
or U44884 (N_44884,N_43857,N_43174);
or U44885 (N_44885,N_43785,N_43840);
xor U44886 (N_44886,N_43059,N_43013);
or U44887 (N_44887,N_43073,N_43800);
and U44888 (N_44888,N_43264,N_43079);
nor U44889 (N_44889,N_43152,N_43536);
nor U44890 (N_44890,N_43233,N_43091);
and U44891 (N_44891,N_43828,N_43250);
nor U44892 (N_44892,N_43689,N_43801);
nand U44893 (N_44893,N_43393,N_43371);
or U44894 (N_44894,N_43027,N_43994);
nor U44895 (N_44895,N_43833,N_43202);
or U44896 (N_44896,N_43729,N_43544);
xor U44897 (N_44897,N_43778,N_43470);
or U44898 (N_44898,N_43568,N_43196);
or U44899 (N_44899,N_43798,N_43115);
xnor U44900 (N_44900,N_43917,N_43885);
nor U44901 (N_44901,N_43276,N_43028);
nor U44902 (N_44902,N_43588,N_43622);
nand U44903 (N_44903,N_43982,N_43145);
nor U44904 (N_44904,N_43967,N_43057);
nor U44905 (N_44905,N_43132,N_43531);
and U44906 (N_44906,N_43452,N_43435);
nand U44907 (N_44907,N_43996,N_43510);
and U44908 (N_44908,N_43605,N_43865);
nor U44909 (N_44909,N_43742,N_43616);
nand U44910 (N_44910,N_43512,N_43569);
and U44911 (N_44911,N_43620,N_43651);
nor U44912 (N_44912,N_43327,N_43533);
nand U44913 (N_44913,N_43268,N_43831);
nand U44914 (N_44914,N_43571,N_43289);
and U44915 (N_44915,N_43511,N_43555);
nand U44916 (N_44916,N_43618,N_43450);
nand U44917 (N_44917,N_43462,N_43712);
or U44918 (N_44918,N_43431,N_43167);
or U44919 (N_44919,N_43663,N_43803);
xnor U44920 (N_44920,N_43046,N_43723);
xor U44921 (N_44921,N_43152,N_43236);
or U44922 (N_44922,N_43359,N_43577);
nor U44923 (N_44923,N_43676,N_43076);
or U44924 (N_44924,N_43727,N_43738);
nor U44925 (N_44925,N_43483,N_43985);
xor U44926 (N_44926,N_43158,N_43451);
or U44927 (N_44927,N_43304,N_43465);
nand U44928 (N_44928,N_43591,N_43834);
nor U44929 (N_44929,N_43746,N_43689);
and U44930 (N_44930,N_43573,N_43105);
xor U44931 (N_44931,N_43415,N_43290);
or U44932 (N_44932,N_43205,N_43749);
and U44933 (N_44933,N_43507,N_43141);
nand U44934 (N_44934,N_43496,N_43694);
xor U44935 (N_44935,N_43389,N_43681);
and U44936 (N_44936,N_43967,N_43336);
nand U44937 (N_44937,N_43368,N_43110);
and U44938 (N_44938,N_43389,N_43012);
or U44939 (N_44939,N_43301,N_43400);
or U44940 (N_44940,N_43189,N_43724);
nor U44941 (N_44941,N_43312,N_43247);
xor U44942 (N_44942,N_43858,N_43788);
xnor U44943 (N_44943,N_43981,N_43868);
or U44944 (N_44944,N_43303,N_43320);
nand U44945 (N_44945,N_43669,N_43344);
and U44946 (N_44946,N_43768,N_43670);
or U44947 (N_44947,N_43288,N_43870);
nor U44948 (N_44948,N_43369,N_43621);
nand U44949 (N_44949,N_43273,N_43056);
nand U44950 (N_44950,N_43550,N_43112);
and U44951 (N_44951,N_43017,N_43007);
nand U44952 (N_44952,N_43020,N_43325);
and U44953 (N_44953,N_43358,N_43573);
xor U44954 (N_44954,N_43529,N_43700);
nand U44955 (N_44955,N_43040,N_43102);
or U44956 (N_44956,N_43848,N_43400);
and U44957 (N_44957,N_43471,N_43231);
nand U44958 (N_44958,N_43185,N_43120);
and U44959 (N_44959,N_43510,N_43689);
or U44960 (N_44960,N_43163,N_43152);
xnor U44961 (N_44961,N_43175,N_43284);
nor U44962 (N_44962,N_43190,N_43506);
or U44963 (N_44963,N_43990,N_43906);
and U44964 (N_44964,N_43164,N_43752);
nor U44965 (N_44965,N_43746,N_43574);
and U44966 (N_44966,N_43186,N_43584);
xnor U44967 (N_44967,N_43301,N_43529);
xnor U44968 (N_44968,N_43042,N_43643);
nand U44969 (N_44969,N_43650,N_43817);
and U44970 (N_44970,N_43578,N_43890);
xor U44971 (N_44971,N_43458,N_43293);
nor U44972 (N_44972,N_43728,N_43289);
or U44973 (N_44973,N_43847,N_43948);
or U44974 (N_44974,N_43185,N_43438);
xnor U44975 (N_44975,N_43974,N_43314);
nand U44976 (N_44976,N_43912,N_43734);
nor U44977 (N_44977,N_43555,N_43673);
nand U44978 (N_44978,N_43654,N_43949);
and U44979 (N_44979,N_43661,N_43083);
xnor U44980 (N_44980,N_43645,N_43675);
nor U44981 (N_44981,N_43897,N_43381);
or U44982 (N_44982,N_43905,N_43476);
nor U44983 (N_44983,N_43747,N_43778);
and U44984 (N_44984,N_43813,N_43648);
or U44985 (N_44985,N_43357,N_43245);
or U44986 (N_44986,N_43898,N_43019);
and U44987 (N_44987,N_43985,N_43583);
xnor U44988 (N_44988,N_43528,N_43100);
nand U44989 (N_44989,N_43054,N_43188);
and U44990 (N_44990,N_43550,N_43606);
and U44991 (N_44991,N_43285,N_43194);
nor U44992 (N_44992,N_43620,N_43684);
and U44993 (N_44993,N_43386,N_43541);
xor U44994 (N_44994,N_43383,N_43114);
nor U44995 (N_44995,N_43371,N_43224);
and U44996 (N_44996,N_43000,N_43586);
nor U44997 (N_44997,N_43068,N_43855);
nor U44998 (N_44998,N_43300,N_43477);
xnor U44999 (N_44999,N_43367,N_43970);
nand U45000 (N_45000,N_44318,N_44647);
nand U45001 (N_45001,N_44144,N_44189);
or U45002 (N_45002,N_44671,N_44152);
nand U45003 (N_45003,N_44995,N_44358);
nor U45004 (N_45004,N_44524,N_44748);
and U45005 (N_45005,N_44233,N_44076);
nor U45006 (N_45006,N_44057,N_44040);
nor U45007 (N_45007,N_44117,N_44330);
xor U45008 (N_45008,N_44405,N_44396);
nor U45009 (N_45009,N_44506,N_44537);
xnor U45010 (N_45010,N_44978,N_44250);
nor U45011 (N_45011,N_44719,N_44617);
nor U45012 (N_45012,N_44101,N_44648);
nor U45013 (N_45013,N_44734,N_44116);
and U45014 (N_45014,N_44413,N_44077);
or U45015 (N_45015,N_44469,N_44522);
nand U45016 (N_45016,N_44147,N_44319);
nand U45017 (N_45017,N_44324,N_44168);
and U45018 (N_45018,N_44482,N_44620);
xor U45019 (N_45019,N_44520,N_44030);
nand U45020 (N_45020,N_44155,N_44247);
nand U45021 (N_45021,N_44206,N_44765);
xnor U45022 (N_45022,N_44234,N_44756);
and U45023 (N_45023,N_44894,N_44228);
and U45024 (N_45024,N_44998,N_44463);
or U45025 (N_45025,N_44024,N_44665);
xnor U45026 (N_45026,N_44010,N_44928);
and U45027 (N_45027,N_44181,N_44270);
and U45028 (N_45028,N_44606,N_44218);
nand U45029 (N_45029,N_44246,N_44174);
xnor U45030 (N_45030,N_44422,N_44832);
nand U45031 (N_45031,N_44530,N_44162);
and U45032 (N_45032,N_44037,N_44738);
xor U45033 (N_45033,N_44811,N_44699);
and U45034 (N_45034,N_44380,N_44193);
and U45035 (N_45035,N_44643,N_44248);
xor U45036 (N_45036,N_44572,N_44382);
or U45037 (N_45037,N_44477,N_44223);
and U45038 (N_45038,N_44865,N_44093);
or U45039 (N_45039,N_44498,N_44690);
and U45040 (N_45040,N_44133,N_44088);
or U45041 (N_45041,N_44547,N_44489);
and U45042 (N_45042,N_44053,N_44979);
and U45043 (N_45043,N_44169,N_44458);
or U45044 (N_45044,N_44946,N_44373);
and U45045 (N_45045,N_44304,N_44586);
nand U45046 (N_45046,N_44518,N_44553);
nand U45047 (N_45047,N_44360,N_44187);
and U45048 (N_45048,N_44215,N_44836);
and U45049 (N_45049,N_44752,N_44940);
or U45050 (N_45050,N_44350,N_44416);
and U45051 (N_45051,N_44106,N_44723);
xor U45052 (N_45052,N_44342,N_44074);
and U45053 (N_45053,N_44801,N_44633);
or U45054 (N_45054,N_44161,N_44164);
nand U45055 (N_45055,N_44200,N_44800);
and U45056 (N_45056,N_44341,N_44126);
and U45057 (N_45057,N_44789,N_44676);
xnor U45058 (N_45058,N_44100,N_44343);
nor U45059 (N_45059,N_44531,N_44172);
and U45060 (N_45060,N_44579,N_44225);
xnor U45061 (N_45061,N_44207,N_44558);
xor U45062 (N_45062,N_44793,N_44542);
nor U45063 (N_45063,N_44700,N_44039);
nor U45064 (N_45064,N_44662,N_44301);
nand U45065 (N_45065,N_44792,N_44903);
xnor U45066 (N_45066,N_44230,N_44298);
and U45067 (N_45067,N_44483,N_44698);
or U45068 (N_45068,N_44922,N_44115);
nor U45069 (N_45069,N_44853,N_44761);
or U45070 (N_45070,N_44994,N_44610);
nand U45071 (N_45071,N_44476,N_44597);
nand U45072 (N_45072,N_44290,N_44732);
and U45073 (N_45073,N_44292,N_44226);
nand U45074 (N_45074,N_44136,N_44593);
xnor U45075 (N_45075,N_44452,N_44663);
and U45076 (N_45076,N_44316,N_44964);
xor U45077 (N_45077,N_44658,N_44878);
nor U45078 (N_45078,N_44959,N_44485);
and U45079 (N_45079,N_44950,N_44760);
xnor U45080 (N_45080,N_44650,N_44481);
or U45081 (N_45081,N_44592,N_44019);
nand U45082 (N_45082,N_44145,N_44807);
or U45083 (N_45083,N_44988,N_44159);
nand U45084 (N_45084,N_44001,N_44598);
or U45085 (N_45085,N_44219,N_44367);
xnor U45086 (N_45086,N_44656,N_44016);
nor U45087 (N_45087,N_44939,N_44747);
or U45088 (N_45088,N_44575,N_44990);
nand U45089 (N_45089,N_44720,N_44945);
xnor U45090 (N_45090,N_44997,N_44550);
and U45091 (N_45091,N_44075,N_44173);
and U45092 (N_45092,N_44495,N_44546);
nand U45093 (N_45093,N_44086,N_44651);
nand U45094 (N_45094,N_44139,N_44308);
xor U45095 (N_45095,N_44254,N_44914);
and U45096 (N_45096,N_44261,N_44385);
or U45097 (N_45097,N_44724,N_44376);
xor U45098 (N_45098,N_44119,N_44599);
nor U45099 (N_45099,N_44791,N_44839);
xor U45100 (N_45100,N_44241,N_44260);
and U45101 (N_45101,N_44653,N_44695);
xor U45102 (N_45102,N_44783,N_44762);
and U45103 (N_45103,N_44066,N_44677);
xnor U45104 (N_45104,N_44491,N_44114);
nor U45105 (N_45105,N_44786,N_44099);
nand U45106 (N_45106,N_44089,N_44927);
xnor U45107 (N_45107,N_44602,N_44862);
nand U45108 (N_45108,N_44977,N_44408);
or U45109 (N_45109,N_44779,N_44932);
nor U45110 (N_45110,N_44737,N_44838);
xor U45111 (N_45111,N_44435,N_44591);
nand U45112 (N_45112,N_44420,N_44920);
nand U45113 (N_45113,N_44965,N_44814);
xor U45114 (N_45114,N_44211,N_44992);
or U45115 (N_45115,N_44632,N_44044);
nor U45116 (N_45116,N_44852,N_44041);
xor U45117 (N_45117,N_44837,N_44455);
nor U45118 (N_45118,N_44600,N_44180);
nor U45119 (N_45119,N_44401,N_44845);
xnor U45120 (N_45120,N_44735,N_44028);
nand U45121 (N_45121,N_44901,N_44571);
and U45122 (N_45122,N_44440,N_44208);
nor U45123 (N_45123,N_44130,N_44742);
nor U45124 (N_45124,N_44038,N_44691);
xnor U45125 (N_45125,N_44210,N_44081);
and U45126 (N_45126,N_44909,N_44962);
nand U45127 (N_45127,N_44666,N_44657);
nor U45128 (N_45128,N_44743,N_44778);
nand U45129 (N_45129,N_44830,N_44252);
xnor U45130 (N_45130,N_44192,N_44340);
and U45131 (N_45131,N_44841,N_44107);
xor U45132 (N_45132,N_44834,N_44683);
or U45133 (N_45133,N_44564,N_44014);
or U45134 (N_45134,N_44003,N_44733);
nand U45135 (N_45135,N_44154,N_44880);
or U45136 (N_45136,N_44584,N_44124);
nor U45137 (N_45137,N_44644,N_44623);
and U45138 (N_45138,N_44980,N_44127);
xor U45139 (N_45139,N_44869,N_44848);
or U45140 (N_45140,N_44462,N_44718);
and U45141 (N_45141,N_44394,N_44635);
nor U45142 (N_45142,N_44976,N_44631);
xor U45143 (N_45143,N_44025,N_44335);
xor U45144 (N_45144,N_44796,N_44366);
nand U45145 (N_45145,N_44359,N_44943);
or U45146 (N_45146,N_44872,N_44924);
xnor U45147 (N_45147,N_44344,N_44365);
nand U45148 (N_45148,N_44326,N_44113);
or U45149 (N_45149,N_44804,N_44567);
xnor U45150 (N_45150,N_44955,N_44842);
xor U45151 (N_45151,N_44538,N_44797);
nor U45152 (N_45152,N_44312,N_44999);
xnor U45153 (N_45153,N_44479,N_44142);
and U45154 (N_45154,N_44274,N_44926);
or U45155 (N_45155,N_44242,N_44516);
xor U45156 (N_45156,N_44062,N_44393);
nand U45157 (N_45157,N_44555,N_44151);
nand U45158 (N_45158,N_44026,N_44276);
and U45159 (N_45159,N_44919,N_44397);
xor U45160 (N_45160,N_44654,N_44815);
nand U45161 (N_45161,N_44209,N_44311);
nor U45162 (N_45162,N_44672,N_44574);
xnor U45163 (N_45163,N_44160,N_44710);
and U45164 (N_45164,N_44492,N_44005);
nor U45165 (N_45165,N_44649,N_44176);
and U45166 (N_45166,N_44661,N_44355);
or U45167 (N_45167,N_44437,N_44079);
or U45168 (N_45168,N_44889,N_44256);
nor U45169 (N_45169,N_44320,N_44750);
nor U45170 (N_45170,N_44613,N_44787);
nand U45171 (N_45171,N_44973,N_44509);
and U45172 (N_45172,N_44892,N_44629);
nand U45173 (N_45173,N_44897,N_44125);
xor U45174 (N_45174,N_44194,N_44182);
or U45175 (N_45175,N_44887,N_44785);
nand U45176 (N_45176,N_44006,N_44507);
nor U45177 (N_45177,N_44430,N_44543);
nor U45178 (N_45178,N_44493,N_44601);
and U45179 (N_45179,N_44561,N_44614);
nand U45180 (N_45180,N_44011,N_44626);
nand U45181 (N_45181,N_44327,N_44983);
nand U45182 (N_45182,N_44707,N_44056);
and U45183 (N_45183,N_44560,N_44953);
nor U45184 (N_45184,N_44638,N_44122);
nand U45185 (N_45185,N_44729,N_44465);
xor U45186 (N_45186,N_44353,N_44863);
nor U45187 (N_45187,N_44891,N_44278);
xnor U45188 (N_45188,N_44501,N_44906);
or U45189 (N_45189,N_44552,N_44907);
nor U45190 (N_45190,N_44705,N_44717);
nor U45191 (N_45191,N_44406,N_44480);
or U45192 (N_45192,N_44767,N_44032);
nand U45193 (N_45193,N_44963,N_44156);
nand U45194 (N_45194,N_44378,N_44583);
nand U45195 (N_45195,N_44213,N_44621);
and U45196 (N_45196,N_44535,N_44947);
xnor U45197 (N_45197,N_44232,N_44387);
xor U45198 (N_45198,N_44725,N_44364);
nand U45199 (N_45199,N_44305,N_44694);
nor U45200 (N_45200,N_44461,N_44426);
or U45201 (N_45201,N_44871,N_44751);
nor U45202 (N_45202,N_44287,N_44050);
and U45203 (N_45203,N_44867,N_44948);
nor U45204 (N_45204,N_44466,N_44083);
or U45205 (N_45205,N_44589,N_44428);
nor U45206 (N_45206,N_44445,N_44612);
and U45207 (N_45207,N_44730,N_44027);
or U45208 (N_45208,N_44904,N_44214);
xnor U45209 (N_45209,N_44447,N_44294);
or U45210 (N_45210,N_44436,N_44628);
or U45211 (N_45211,N_44968,N_44494);
nor U45212 (N_45212,N_44701,N_44146);
nand U45213 (N_45213,N_44398,N_44059);
nor U45214 (N_45214,N_44110,N_44389);
xor U45215 (N_45215,N_44630,N_44286);
or U45216 (N_45216,N_44165,N_44457);
and U45217 (N_45217,N_44070,N_44098);
and U45218 (N_45218,N_44134,N_44686);
xnor U45219 (N_45219,N_44639,N_44956);
or U45220 (N_45220,N_44131,N_44285);
or U45221 (N_45221,N_44021,N_44798);
nor U45222 (N_45222,N_44105,N_44936);
nor U45223 (N_45223,N_44684,N_44714);
and U45224 (N_45224,N_44822,N_44108);
xnor U45225 (N_45225,N_44949,N_44033);
xor U45226 (N_45226,N_44064,N_44883);
or U45227 (N_45227,N_44712,N_44379);
nand U45228 (N_45228,N_44636,N_44879);
nand U45229 (N_45229,N_44351,N_44605);
xnor U45230 (N_45230,N_44138,N_44771);
or U45231 (N_45231,N_44381,N_44890);
nand U45232 (N_45232,N_44082,N_44736);
nand U45233 (N_45233,N_44450,N_44921);
nand U45234 (N_45234,N_44374,N_44840);
xor U45235 (N_45235,N_44915,N_44177);
and U45236 (N_45236,N_44236,N_44054);
xnor U45237 (N_45237,N_44669,N_44681);
and U45238 (N_45238,N_44345,N_44212);
nor U45239 (N_45239,N_44923,N_44938);
and U45240 (N_45240,N_44627,N_44338);
and U45241 (N_45241,N_44049,N_44846);
xnor U45242 (N_45242,N_44012,N_44908);
nand U45243 (N_45243,N_44859,N_44309);
xnor U45244 (N_45244,N_44467,N_44284);
nor U45245 (N_45245,N_44989,N_44487);
and U45246 (N_45246,N_44618,N_44410);
xnor U45247 (N_45247,N_44442,N_44143);
and U45248 (N_45248,N_44642,N_44521);
nor U45249 (N_45249,N_44198,N_44149);
and U45250 (N_45250,N_44809,N_44664);
or U45251 (N_45251,N_44795,N_44267);
nand U45252 (N_45252,N_44952,N_44478);
nand U45253 (N_45253,N_44148,N_44348);
nand U45254 (N_45254,N_44414,N_44910);
nor U45255 (N_45255,N_44877,N_44063);
and U45256 (N_45256,N_44870,N_44817);
or U45257 (N_45257,N_44625,N_44585);
and U45258 (N_45258,N_44587,N_44087);
nand U45259 (N_45259,N_44982,N_44931);
nor U45260 (N_45260,N_44641,N_44363);
xor U45261 (N_45261,N_44323,N_44015);
and U45262 (N_45262,N_44185,N_44170);
and U45263 (N_45263,N_44140,N_44166);
and U45264 (N_45264,N_44991,N_44511);
xor U45265 (N_45265,N_44757,N_44317);
nand U45266 (N_45266,N_44523,N_44881);
nor U45267 (N_45267,N_44655,N_44559);
xor U45268 (N_45268,N_44969,N_44217);
or U45269 (N_45269,N_44824,N_44526);
nor U45270 (N_45270,N_44570,N_44425);
nand U45271 (N_45271,N_44244,N_44268);
or U45272 (N_45272,N_44504,N_44061);
nand U45273 (N_45273,N_44510,N_44277);
xnor U45274 (N_45274,N_44532,N_44678);
or U45275 (N_45275,N_44418,N_44329);
or U45276 (N_45276,N_44595,N_44569);
and U45277 (N_45277,N_44580,N_44084);
nand U45278 (N_45278,N_44831,N_44749);
nor U45279 (N_45279,N_44768,N_44067);
or U45280 (N_45280,N_44545,N_44820);
and U45281 (N_45281,N_44687,N_44847);
xor U45282 (N_45282,N_44337,N_44893);
nor U45283 (N_45283,N_44864,N_44446);
xnor U45284 (N_45284,N_44716,N_44473);
xnor U45285 (N_45285,N_44873,N_44415);
xnor U45286 (N_45286,N_44310,N_44744);
nand U45287 (N_45287,N_44899,N_44812);
xnor U45288 (N_45288,N_44529,N_44412);
or U45289 (N_45289,N_44933,N_44400);
and U45290 (N_45290,N_44854,N_44433);
and U45291 (N_45291,N_44755,N_44935);
nor U45292 (N_45292,N_44539,N_44390);
nor U45293 (N_45293,N_44157,N_44417);
and U45294 (N_45294,N_44637,N_44557);
and U45295 (N_45295,N_44307,N_44388);
nor U45296 (N_45296,N_44175,N_44409);
xor U45297 (N_45297,N_44566,N_44085);
xor U45298 (N_45298,N_44191,N_44243);
xnor U45299 (N_45299,N_44281,N_44231);
and U45300 (N_45300,N_44505,N_44104);
nand U45301 (N_45301,N_44985,N_44758);
nor U45302 (N_45302,N_44150,N_44451);
nor U45303 (N_45303,N_44395,N_44803);
or U45304 (N_45304,N_44265,N_44224);
xnor U45305 (N_45305,N_44431,N_44017);
nor U45306 (N_45306,N_44513,N_44645);
and U45307 (N_45307,N_44322,N_44332);
nand U45308 (N_45308,N_44667,N_44715);
or U45309 (N_45309,N_44993,N_44788);
or U45310 (N_45310,N_44096,N_44488);
xor U45311 (N_45311,N_44556,N_44456);
and U45312 (N_45312,N_44986,N_44886);
xnor U45313 (N_45313,N_44336,N_44590);
and U45314 (N_45314,N_44253,N_44685);
nor U45315 (N_45315,N_44929,N_44582);
or U45316 (N_45316,N_44065,N_44153);
nand U45317 (N_45317,N_44764,N_44196);
xor U45318 (N_45318,N_44474,N_44448);
nand U45319 (N_45319,N_44023,N_44975);
and U45320 (N_45320,N_44484,N_44090);
xnor U45321 (N_45321,N_44711,N_44709);
and U45322 (N_45322,N_44073,N_44441);
xor U45323 (N_45323,N_44372,N_44679);
or U45324 (N_45324,N_44726,N_44634);
xnor U45325 (N_45325,N_44313,N_44438);
nand U45326 (N_45326,N_44369,N_44300);
xnor U45327 (N_45327,N_44565,N_44449);
xor U45328 (N_45328,N_44759,N_44371);
nor U45329 (N_45329,N_44549,N_44594);
and U45330 (N_45330,N_44043,N_44728);
and U45331 (N_45331,N_44519,N_44497);
xnor U45332 (N_45332,N_44652,N_44263);
nand U45333 (N_45333,N_44454,N_44884);
nor U45334 (N_45334,N_44399,N_44377);
nor U45335 (N_45335,N_44689,N_44052);
or U45336 (N_45336,N_44607,N_44905);
and U45337 (N_45337,N_44129,N_44802);
nor U45338 (N_45338,N_44283,N_44239);
nand U45339 (N_45339,N_44051,N_44609);
xor U45340 (N_45340,N_44971,N_44296);
and U45341 (N_45341,N_44293,N_44325);
xor U45342 (N_45342,N_44770,N_44045);
nand U45343 (N_45343,N_44913,N_44704);
or U45344 (N_45344,N_44900,N_44235);
nand U45345 (N_45345,N_44825,N_44002);
and U45346 (N_45346,N_44816,N_44996);
xnor U45347 (N_45347,N_44183,N_44222);
or U45348 (N_45348,N_44141,N_44111);
xnor U45349 (N_45349,N_44706,N_44974);
and U45350 (N_45350,N_44799,N_44930);
nand U45351 (N_45351,N_44944,N_44895);
xor U45352 (N_45352,N_44368,N_44184);
xnor U45353 (N_45353,N_44693,N_44271);
xnor U45354 (N_45354,N_44048,N_44500);
or U45355 (N_45355,N_44918,N_44357);
nand U45356 (N_45356,N_44876,N_44429);
or U45357 (N_45357,N_44000,N_44911);
nor U45358 (N_45358,N_44453,N_44525);
and U45359 (N_45359,N_44958,N_44275);
nor U45360 (N_45360,N_44502,N_44273);
or U45361 (N_45361,N_44121,N_44128);
nand U45362 (N_45362,N_44856,N_44272);
nand U45363 (N_45363,N_44740,N_44444);
nor U45364 (N_45364,N_44713,N_44981);
and U45365 (N_45365,N_44540,N_44216);
nand U45366 (N_45366,N_44527,N_44611);
or U45367 (N_45367,N_44533,N_44741);
nand U45368 (N_45368,N_44432,N_44282);
nor U45369 (N_45369,N_44072,N_44823);
or U45370 (N_45370,N_44898,N_44925);
nor U45371 (N_45371,N_44424,N_44069);
xor U45372 (N_45372,N_44548,N_44407);
or U45373 (N_45373,N_44616,N_44813);
xnor U45374 (N_45374,N_44375,N_44861);
and U45375 (N_45375,N_44238,N_44035);
xor U45376 (N_45376,N_44882,N_44468);
nor U45377 (N_45377,N_44339,N_44046);
xnor U45378 (N_45378,N_44934,N_44123);
nand U45379 (N_45379,N_44781,N_44776);
or U45380 (N_45380,N_44186,N_44362);
nand U45381 (N_45381,N_44008,N_44068);
xor U45382 (N_45382,N_44221,N_44179);
or U45383 (N_45383,N_44843,N_44640);
nor U45384 (N_45384,N_44581,N_44660);
nor U45385 (N_45385,N_44347,N_44554);
xor U45386 (N_45386,N_44203,N_44708);
xnor U45387 (N_45387,N_44471,N_44851);
or U45388 (N_45388,N_44503,N_44849);
xnor U45389 (N_45389,N_44608,N_44774);
and U45390 (N_45390,N_44916,N_44427);
xnor U45391 (N_45391,N_44470,N_44303);
nand U45392 (N_45392,N_44171,N_44888);
or U45393 (N_45393,N_44361,N_44858);
nor U45394 (N_45394,N_44205,N_44004);
or U45395 (N_45395,N_44821,N_44551);
nand U45396 (N_45396,N_44229,N_44103);
and U45397 (N_45397,N_44257,N_44334);
nand U45398 (N_45398,N_44135,N_44178);
nand U45399 (N_45399,N_44967,N_44829);
nor U45400 (N_45400,N_44109,N_44541);
nand U45401 (N_45401,N_44443,N_44528);
nand U45402 (N_45402,N_44951,N_44259);
nand U45403 (N_45403,N_44423,N_44810);
nand U45404 (N_45404,N_44163,N_44769);
or U45405 (N_45405,N_44835,N_44806);
nor U45406 (N_45406,N_44578,N_44315);
xor U45407 (N_45407,N_44603,N_44295);
xor U45408 (N_45408,N_44078,N_44688);
xnor U45409 (N_45409,N_44120,N_44302);
nor U45410 (N_45410,N_44102,N_44808);
xnor U45411 (N_45411,N_44352,N_44490);
xor U45412 (N_45412,N_44370,N_44622);
and U45413 (N_45413,N_44333,N_44860);
nor U45414 (N_45414,N_44091,N_44960);
and U45415 (N_45415,N_44702,N_44464);
xor U45416 (N_45416,N_44721,N_44987);
nor U45417 (N_45417,N_44646,N_44201);
nand U45418 (N_45418,N_44659,N_44753);
nor U45419 (N_45419,N_44346,N_44512);
nand U45420 (N_45420,N_44670,N_44668);
nor U45421 (N_45421,N_44696,N_44034);
or U45422 (N_45422,N_44972,N_44514);
or U45423 (N_45423,N_44288,N_44619);
or U45424 (N_45424,N_44197,N_44460);
xor U45425 (N_45425,N_44961,N_44047);
xnor U45426 (N_45426,N_44746,N_44739);
and U45427 (N_45427,N_44885,N_44404);
nand U45428 (N_45428,N_44917,N_44245);
and U45429 (N_45429,N_44703,N_44029);
nand U45430 (N_45430,N_44615,N_44722);
nor U45431 (N_45431,N_44060,N_44496);
or U45432 (N_45432,N_44596,N_44158);
nand U45433 (N_45433,N_44515,N_44790);
and U45434 (N_45434,N_44055,N_44459);
xnor U45435 (N_45435,N_44673,N_44818);
xnor U45436 (N_45436,N_44354,N_44167);
nor U45437 (N_45437,N_44279,N_44384);
and U45438 (N_45438,N_44970,N_44269);
nand U45439 (N_45439,N_44349,N_44280);
and U45440 (N_45440,N_44604,N_44321);
and U45441 (N_45441,N_44763,N_44577);
nand U45442 (N_45442,N_44486,N_44402);
nand U45443 (N_45443,N_44007,N_44264);
or U45444 (N_45444,N_44289,N_44777);
and U45445 (N_45445,N_44745,N_44874);
nand U45446 (N_45446,N_44563,N_44866);
and U45447 (N_45447,N_44118,N_44896);
nand U45448 (N_45448,N_44020,N_44071);
and U45449 (N_45449,N_44844,N_44692);
nor U45450 (N_45450,N_44775,N_44772);
nand U45451 (N_45451,N_44266,N_44042);
nor U45452 (N_45452,N_44544,N_44536);
xnor U45453 (N_45453,N_44568,N_44680);
xnor U45454 (N_45454,N_44697,N_44875);
or U45455 (N_45455,N_44199,N_44195);
and U45456 (N_45456,N_44112,N_44573);
xor U45457 (N_45457,N_44328,N_44828);
nand U45458 (N_45458,N_44833,N_44782);
or U45459 (N_45459,N_44826,N_44237);
nor U45460 (N_45460,N_44827,N_44499);
or U45461 (N_45461,N_44434,N_44754);
nor U45462 (N_45462,N_44857,N_44391);
nor U45463 (N_45463,N_44262,N_44240);
and U45464 (N_45464,N_44674,N_44356);
nor U45465 (N_45465,N_44475,N_44411);
nor U45466 (N_45466,N_44058,N_44291);
xor U45467 (N_45467,N_44137,N_44095);
and U45468 (N_45468,N_44941,N_44624);
or U45469 (N_45469,N_44258,N_44784);
or U45470 (N_45470,N_44682,N_44780);
nor U45471 (N_45471,N_44013,N_44386);
nand U45472 (N_45472,N_44092,N_44009);
xor U45473 (N_45473,N_44534,N_44472);
xor U45474 (N_45474,N_44022,N_44675);
xnor U45475 (N_45475,N_44227,N_44392);
xnor U45476 (N_45476,N_44576,N_44255);
nand U45477 (N_45477,N_44031,N_44942);
or U45478 (N_45478,N_44132,N_44202);
nor U45479 (N_45479,N_44819,N_44855);
and U45480 (N_45480,N_44080,N_44018);
and U45481 (N_45481,N_44036,N_44421);
nor U45482 (N_45482,N_44508,N_44902);
xor U45483 (N_45483,N_44805,N_44957);
or U45484 (N_45484,N_44188,N_44297);
or U45485 (N_45485,N_44850,N_44419);
and U45486 (N_45486,N_44251,N_44439);
xnor U45487 (N_45487,N_44984,N_44727);
nand U45488 (N_45488,N_44299,N_44097);
and U45489 (N_45489,N_44588,N_44249);
nor U45490 (N_45490,N_44094,N_44937);
nand U45491 (N_45491,N_44383,N_44403);
xor U45492 (N_45492,N_44331,N_44306);
nor U45493 (N_45493,N_44562,N_44966);
nand U45494 (N_45494,N_44773,N_44912);
nor U45495 (N_45495,N_44204,N_44220);
and U45496 (N_45496,N_44731,N_44766);
xnor U45497 (N_45497,N_44954,N_44868);
nor U45498 (N_45498,N_44517,N_44794);
nor U45499 (N_45499,N_44314,N_44190);
xor U45500 (N_45500,N_44719,N_44052);
and U45501 (N_45501,N_44210,N_44504);
and U45502 (N_45502,N_44468,N_44485);
nor U45503 (N_45503,N_44680,N_44522);
nor U45504 (N_45504,N_44711,N_44915);
nor U45505 (N_45505,N_44474,N_44597);
or U45506 (N_45506,N_44628,N_44054);
xor U45507 (N_45507,N_44531,N_44424);
xor U45508 (N_45508,N_44573,N_44554);
or U45509 (N_45509,N_44483,N_44874);
or U45510 (N_45510,N_44039,N_44337);
or U45511 (N_45511,N_44109,N_44098);
nand U45512 (N_45512,N_44599,N_44539);
xor U45513 (N_45513,N_44406,N_44639);
nor U45514 (N_45514,N_44954,N_44944);
or U45515 (N_45515,N_44299,N_44766);
nand U45516 (N_45516,N_44168,N_44050);
and U45517 (N_45517,N_44792,N_44537);
or U45518 (N_45518,N_44777,N_44908);
nor U45519 (N_45519,N_44117,N_44552);
xnor U45520 (N_45520,N_44977,N_44107);
xor U45521 (N_45521,N_44796,N_44671);
or U45522 (N_45522,N_44174,N_44977);
xor U45523 (N_45523,N_44314,N_44318);
xnor U45524 (N_45524,N_44426,N_44813);
and U45525 (N_45525,N_44948,N_44929);
or U45526 (N_45526,N_44219,N_44342);
and U45527 (N_45527,N_44776,N_44449);
and U45528 (N_45528,N_44918,N_44440);
nand U45529 (N_45529,N_44510,N_44975);
xnor U45530 (N_45530,N_44405,N_44647);
xor U45531 (N_45531,N_44971,N_44760);
nand U45532 (N_45532,N_44892,N_44062);
nand U45533 (N_45533,N_44385,N_44012);
and U45534 (N_45534,N_44953,N_44592);
nand U45535 (N_45535,N_44038,N_44255);
or U45536 (N_45536,N_44433,N_44310);
nand U45537 (N_45537,N_44034,N_44337);
nor U45538 (N_45538,N_44984,N_44379);
and U45539 (N_45539,N_44490,N_44811);
nor U45540 (N_45540,N_44352,N_44683);
nor U45541 (N_45541,N_44250,N_44565);
nand U45542 (N_45542,N_44374,N_44170);
xnor U45543 (N_45543,N_44818,N_44514);
nor U45544 (N_45544,N_44938,N_44986);
or U45545 (N_45545,N_44377,N_44338);
or U45546 (N_45546,N_44277,N_44730);
xor U45547 (N_45547,N_44549,N_44242);
nand U45548 (N_45548,N_44062,N_44806);
and U45549 (N_45549,N_44885,N_44828);
and U45550 (N_45550,N_44270,N_44074);
and U45551 (N_45551,N_44776,N_44833);
or U45552 (N_45552,N_44377,N_44925);
nor U45553 (N_45553,N_44142,N_44741);
xor U45554 (N_45554,N_44828,N_44148);
nand U45555 (N_45555,N_44203,N_44320);
or U45556 (N_45556,N_44399,N_44604);
nand U45557 (N_45557,N_44649,N_44276);
and U45558 (N_45558,N_44101,N_44600);
or U45559 (N_45559,N_44938,N_44603);
or U45560 (N_45560,N_44553,N_44001);
nand U45561 (N_45561,N_44299,N_44212);
nand U45562 (N_45562,N_44330,N_44871);
nand U45563 (N_45563,N_44833,N_44829);
nor U45564 (N_45564,N_44838,N_44541);
xor U45565 (N_45565,N_44979,N_44395);
and U45566 (N_45566,N_44329,N_44380);
xnor U45567 (N_45567,N_44260,N_44367);
or U45568 (N_45568,N_44381,N_44169);
or U45569 (N_45569,N_44748,N_44876);
nand U45570 (N_45570,N_44595,N_44944);
or U45571 (N_45571,N_44110,N_44907);
and U45572 (N_45572,N_44651,N_44922);
xnor U45573 (N_45573,N_44486,N_44032);
or U45574 (N_45574,N_44930,N_44232);
and U45575 (N_45575,N_44861,N_44184);
nor U45576 (N_45576,N_44202,N_44700);
nand U45577 (N_45577,N_44662,N_44944);
xor U45578 (N_45578,N_44390,N_44576);
or U45579 (N_45579,N_44378,N_44599);
nor U45580 (N_45580,N_44561,N_44384);
or U45581 (N_45581,N_44022,N_44366);
nor U45582 (N_45582,N_44738,N_44444);
xor U45583 (N_45583,N_44954,N_44542);
nor U45584 (N_45584,N_44489,N_44392);
nor U45585 (N_45585,N_44917,N_44186);
xor U45586 (N_45586,N_44352,N_44515);
xnor U45587 (N_45587,N_44565,N_44459);
or U45588 (N_45588,N_44594,N_44302);
and U45589 (N_45589,N_44631,N_44297);
or U45590 (N_45590,N_44286,N_44130);
or U45591 (N_45591,N_44830,N_44716);
nor U45592 (N_45592,N_44383,N_44373);
nand U45593 (N_45593,N_44012,N_44158);
xnor U45594 (N_45594,N_44217,N_44847);
and U45595 (N_45595,N_44584,N_44049);
or U45596 (N_45596,N_44249,N_44488);
xnor U45597 (N_45597,N_44541,N_44359);
and U45598 (N_45598,N_44304,N_44366);
nand U45599 (N_45599,N_44151,N_44710);
or U45600 (N_45600,N_44830,N_44158);
nor U45601 (N_45601,N_44594,N_44556);
nor U45602 (N_45602,N_44915,N_44716);
and U45603 (N_45603,N_44421,N_44434);
or U45604 (N_45604,N_44522,N_44247);
nor U45605 (N_45605,N_44594,N_44643);
xor U45606 (N_45606,N_44798,N_44032);
and U45607 (N_45607,N_44434,N_44715);
xor U45608 (N_45608,N_44484,N_44917);
xor U45609 (N_45609,N_44779,N_44006);
or U45610 (N_45610,N_44815,N_44539);
nor U45611 (N_45611,N_44406,N_44591);
or U45612 (N_45612,N_44591,N_44819);
nor U45613 (N_45613,N_44574,N_44157);
and U45614 (N_45614,N_44096,N_44600);
xor U45615 (N_45615,N_44616,N_44569);
nor U45616 (N_45616,N_44490,N_44266);
xnor U45617 (N_45617,N_44526,N_44608);
nand U45618 (N_45618,N_44603,N_44240);
xor U45619 (N_45619,N_44932,N_44231);
and U45620 (N_45620,N_44409,N_44250);
or U45621 (N_45621,N_44953,N_44323);
and U45622 (N_45622,N_44738,N_44039);
and U45623 (N_45623,N_44202,N_44522);
xor U45624 (N_45624,N_44250,N_44750);
xnor U45625 (N_45625,N_44316,N_44362);
or U45626 (N_45626,N_44506,N_44872);
or U45627 (N_45627,N_44977,N_44334);
xor U45628 (N_45628,N_44543,N_44987);
nand U45629 (N_45629,N_44196,N_44194);
and U45630 (N_45630,N_44875,N_44208);
xnor U45631 (N_45631,N_44905,N_44725);
or U45632 (N_45632,N_44070,N_44792);
or U45633 (N_45633,N_44037,N_44494);
nor U45634 (N_45634,N_44375,N_44026);
nand U45635 (N_45635,N_44281,N_44916);
nand U45636 (N_45636,N_44837,N_44028);
or U45637 (N_45637,N_44916,N_44393);
or U45638 (N_45638,N_44124,N_44656);
or U45639 (N_45639,N_44078,N_44473);
or U45640 (N_45640,N_44410,N_44972);
and U45641 (N_45641,N_44836,N_44433);
nand U45642 (N_45642,N_44292,N_44606);
xor U45643 (N_45643,N_44401,N_44010);
and U45644 (N_45644,N_44763,N_44700);
nor U45645 (N_45645,N_44682,N_44613);
and U45646 (N_45646,N_44568,N_44009);
nor U45647 (N_45647,N_44892,N_44075);
and U45648 (N_45648,N_44786,N_44156);
nor U45649 (N_45649,N_44201,N_44809);
nor U45650 (N_45650,N_44793,N_44289);
or U45651 (N_45651,N_44192,N_44193);
and U45652 (N_45652,N_44771,N_44736);
nor U45653 (N_45653,N_44261,N_44841);
nand U45654 (N_45654,N_44510,N_44959);
or U45655 (N_45655,N_44164,N_44813);
or U45656 (N_45656,N_44980,N_44421);
nor U45657 (N_45657,N_44427,N_44236);
and U45658 (N_45658,N_44904,N_44335);
or U45659 (N_45659,N_44436,N_44773);
xor U45660 (N_45660,N_44996,N_44257);
nor U45661 (N_45661,N_44994,N_44342);
xnor U45662 (N_45662,N_44012,N_44234);
or U45663 (N_45663,N_44238,N_44319);
nor U45664 (N_45664,N_44534,N_44888);
nand U45665 (N_45665,N_44989,N_44158);
and U45666 (N_45666,N_44405,N_44735);
or U45667 (N_45667,N_44253,N_44862);
nor U45668 (N_45668,N_44629,N_44995);
nand U45669 (N_45669,N_44242,N_44095);
or U45670 (N_45670,N_44799,N_44697);
or U45671 (N_45671,N_44174,N_44871);
nand U45672 (N_45672,N_44468,N_44919);
nand U45673 (N_45673,N_44252,N_44509);
xnor U45674 (N_45674,N_44475,N_44539);
or U45675 (N_45675,N_44885,N_44941);
or U45676 (N_45676,N_44696,N_44115);
or U45677 (N_45677,N_44209,N_44318);
or U45678 (N_45678,N_44110,N_44754);
nor U45679 (N_45679,N_44958,N_44541);
nor U45680 (N_45680,N_44365,N_44965);
and U45681 (N_45681,N_44476,N_44396);
xor U45682 (N_45682,N_44971,N_44805);
nor U45683 (N_45683,N_44016,N_44363);
xnor U45684 (N_45684,N_44369,N_44715);
nand U45685 (N_45685,N_44690,N_44771);
xnor U45686 (N_45686,N_44036,N_44308);
and U45687 (N_45687,N_44397,N_44053);
xnor U45688 (N_45688,N_44366,N_44678);
nor U45689 (N_45689,N_44876,N_44421);
or U45690 (N_45690,N_44203,N_44570);
nand U45691 (N_45691,N_44350,N_44194);
and U45692 (N_45692,N_44562,N_44051);
or U45693 (N_45693,N_44118,N_44639);
and U45694 (N_45694,N_44517,N_44460);
nand U45695 (N_45695,N_44516,N_44446);
and U45696 (N_45696,N_44683,N_44280);
or U45697 (N_45697,N_44702,N_44430);
xor U45698 (N_45698,N_44940,N_44070);
nor U45699 (N_45699,N_44304,N_44422);
or U45700 (N_45700,N_44113,N_44947);
nand U45701 (N_45701,N_44836,N_44715);
and U45702 (N_45702,N_44354,N_44472);
nor U45703 (N_45703,N_44205,N_44234);
xnor U45704 (N_45704,N_44470,N_44297);
or U45705 (N_45705,N_44153,N_44225);
nor U45706 (N_45706,N_44565,N_44230);
xnor U45707 (N_45707,N_44583,N_44576);
or U45708 (N_45708,N_44863,N_44645);
nand U45709 (N_45709,N_44785,N_44236);
nor U45710 (N_45710,N_44760,N_44406);
and U45711 (N_45711,N_44644,N_44033);
nor U45712 (N_45712,N_44654,N_44632);
xor U45713 (N_45713,N_44101,N_44677);
nand U45714 (N_45714,N_44950,N_44715);
xor U45715 (N_45715,N_44510,N_44701);
xor U45716 (N_45716,N_44183,N_44693);
nand U45717 (N_45717,N_44075,N_44186);
nand U45718 (N_45718,N_44445,N_44420);
or U45719 (N_45719,N_44877,N_44445);
or U45720 (N_45720,N_44134,N_44065);
or U45721 (N_45721,N_44134,N_44428);
nor U45722 (N_45722,N_44193,N_44340);
and U45723 (N_45723,N_44666,N_44946);
or U45724 (N_45724,N_44032,N_44837);
nor U45725 (N_45725,N_44424,N_44874);
or U45726 (N_45726,N_44536,N_44987);
xnor U45727 (N_45727,N_44522,N_44379);
nand U45728 (N_45728,N_44669,N_44770);
nor U45729 (N_45729,N_44451,N_44326);
nor U45730 (N_45730,N_44752,N_44600);
xor U45731 (N_45731,N_44481,N_44183);
and U45732 (N_45732,N_44248,N_44339);
and U45733 (N_45733,N_44694,N_44192);
and U45734 (N_45734,N_44824,N_44186);
or U45735 (N_45735,N_44463,N_44596);
nor U45736 (N_45736,N_44989,N_44777);
xnor U45737 (N_45737,N_44651,N_44399);
and U45738 (N_45738,N_44733,N_44250);
nand U45739 (N_45739,N_44981,N_44541);
xor U45740 (N_45740,N_44190,N_44480);
nand U45741 (N_45741,N_44823,N_44174);
and U45742 (N_45742,N_44596,N_44132);
nand U45743 (N_45743,N_44505,N_44955);
nand U45744 (N_45744,N_44613,N_44485);
nand U45745 (N_45745,N_44592,N_44491);
nand U45746 (N_45746,N_44193,N_44544);
xor U45747 (N_45747,N_44043,N_44097);
and U45748 (N_45748,N_44192,N_44336);
nor U45749 (N_45749,N_44329,N_44992);
xnor U45750 (N_45750,N_44063,N_44314);
nand U45751 (N_45751,N_44345,N_44757);
nor U45752 (N_45752,N_44522,N_44558);
nor U45753 (N_45753,N_44105,N_44727);
nor U45754 (N_45754,N_44895,N_44663);
and U45755 (N_45755,N_44258,N_44832);
and U45756 (N_45756,N_44636,N_44990);
nor U45757 (N_45757,N_44341,N_44209);
xnor U45758 (N_45758,N_44952,N_44240);
nor U45759 (N_45759,N_44404,N_44409);
xor U45760 (N_45760,N_44220,N_44079);
xnor U45761 (N_45761,N_44432,N_44113);
and U45762 (N_45762,N_44436,N_44802);
nand U45763 (N_45763,N_44890,N_44365);
or U45764 (N_45764,N_44337,N_44460);
nor U45765 (N_45765,N_44283,N_44209);
nand U45766 (N_45766,N_44572,N_44810);
and U45767 (N_45767,N_44384,N_44608);
and U45768 (N_45768,N_44192,N_44139);
and U45769 (N_45769,N_44270,N_44703);
xnor U45770 (N_45770,N_44026,N_44146);
and U45771 (N_45771,N_44464,N_44355);
or U45772 (N_45772,N_44836,N_44490);
xor U45773 (N_45773,N_44328,N_44883);
nor U45774 (N_45774,N_44003,N_44985);
nor U45775 (N_45775,N_44947,N_44500);
nand U45776 (N_45776,N_44132,N_44178);
or U45777 (N_45777,N_44110,N_44245);
or U45778 (N_45778,N_44320,N_44007);
and U45779 (N_45779,N_44757,N_44045);
and U45780 (N_45780,N_44582,N_44408);
nand U45781 (N_45781,N_44408,N_44972);
and U45782 (N_45782,N_44263,N_44823);
nor U45783 (N_45783,N_44507,N_44377);
and U45784 (N_45784,N_44433,N_44729);
nor U45785 (N_45785,N_44823,N_44551);
nor U45786 (N_45786,N_44370,N_44408);
or U45787 (N_45787,N_44198,N_44509);
nor U45788 (N_45788,N_44341,N_44909);
or U45789 (N_45789,N_44637,N_44866);
and U45790 (N_45790,N_44456,N_44021);
nand U45791 (N_45791,N_44990,N_44030);
nor U45792 (N_45792,N_44387,N_44315);
or U45793 (N_45793,N_44646,N_44576);
nand U45794 (N_45794,N_44817,N_44835);
xor U45795 (N_45795,N_44849,N_44460);
nand U45796 (N_45796,N_44530,N_44770);
nor U45797 (N_45797,N_44638,N_44226);
or U45798 (N_45798,N_44673,N_44106);
or U45799 (N_45799,N_44268,N_44693);
xnor U45800 (N_45800,N_44524,N_44802);
or U45801 (N_45801,N_44460,N_44425);
and U45802 (N_45802,N_44171,N_44124);
and U45803 (N_45803,N_44693,N_44770);
or U45804 (N_45804,N_44596,N_44753);
and U45805 (N_45805,N_44381,N_44728);
nand U45806 (N_45806,N_44219,N_44120);
nand U45807 (N_45807,N_44888,N_44542);
and U45808 (N_45808,N_44260,N_44618);
and U45809 (N_45809,N_44521,N_44913);
nor U45810 (N_45810,N_44032,N_44965);
or U45811 (N_45811,N_44434,N_44688);
nor U45812 (N_45812,N_44815,N_44621);
nand U45813 (N_45813,N_44588,N_44708);
xnor U45814 (N_45814,N_44749,N_44994);
or U45815 (N_45815,N_44025,N_44770);
nand U45816 (N_45816,N_44637,N_44753);
and U45817 (N_45817,N_44366,N_44936);
or U45818 (N_45818,N_44569,N_44155);
nand U45819 (N_45819,N_44557,N_44327);
xor U45820 (N_45820,N_44558,N_44538);
nor U45821 (N_45821,N_44888,N_44599);
xnor U45822 (N_45822,N_44759,N_44636);
and U45823 (N_45823,N_44036,N_44112);
or U45824 (N_45824,N_44418,N_44135);
nand U45825 (N_45825,N_44967,N_44052);
nand U45826 (N_45826,N_44219,N_44653);
nor U45827 (N_45827,N_44435,N_44331);
xor U45828 (N_45828,N_44776,N_44224);
nand U45829 (N_45829,N_44999,N_44171);
nand U45830 (N_45830,N_44453,N_44879);
and U45831 (N_45831,N_44928,N_44645);
nand U45832 (N_45832,N_44469,N_44053);
nor U45833 (N_45833,N_44338,N_44450);
nand U45834 (N_45834,N_44974,N_44839);
nand U45835 (N_45835,N_44772,N_44268);
and U45836 (N_45836,N_44426,N_44550);
nor U45837 (N_45837,N_44961,N_44208);
nor U45838 (N_45838,N_44126,N_44766);
nand U45839 (N_45839,N_44612,N_44291);
or U45840 (N_45840,N_44192,N_44455);
or U45841 (N_45841,N_44199,N_44126);
and U45842 (N_45842,N_44669,N_44547);
or U45843 (N_45843,N_44691,N_44514);
and U45844 (N_45844,N_44489,N_44767);
and U45845 (N_45845,N_44720,N_44118);
or U45846 (N_45846,N_44632,N_44051);
xor U45847 (N_45847,N_44760,N_44002);
and U45848 (N_45848,N_44439,N_44934);
nor U45849 (N_45849,N_44907,N_44208);
or U45850 (N_45850,N_44271,N_44689);
xnor U45851 (N_45851,N_44709,N_44437);
xor U45852 (N_45852,N_44805,N_44208);
or U45853 (N_45853,N_44711,N_44560);
xor U45854 (N_45854,N_44893,N_44484);
xnor U45855 (N_45855,N_44896,N_44039);
nand U45856 (N_45856,N_44130,N_44358);
and U45857 (N_45857,N_44480,N_44537);
and U45858 (N_45858,N_44235,N_44707);
or U45859 (N_45859,N_44763,N_44211);
and U45860 (N_45860,N_44629,N_44279);
nand U45861 (N_45861,N_44487,N_44825);
nand U45862 (N_45862,N_44093,N_44741);
nor U45863 (N_45863,N_44996,N_44048);
and U45864 (N_45864,N_44731,N_44968);
nor U45865 (N_45865,N_44533,N_44895);
nor U45866 (N_45866,N_44945,N_44857);
xor U45867 (N_45867,N_44844,N_44176);
nand U45868 (N_45868,N_44197,N_44523);
nand U45869 (N_45869,N_44089,N_44799);
xor U45870 (N_45870,N_44271,N_44649);
xnor U45871 (N_45871,N_44263,N_44034);
nor U45872 (N_45872,N_44931,N_44635);
xor U45873 (N_45873,N_44144,N_44205);
nor U45874 (N_45874,N_44642,N_44431);
nand U45875 (N_45875,N_44837,N_44118);
nand U45876 (N_45876,N_44351,N_44868);
and U45877 (N_45877,N_44244,N_44657);
and U45878 (N_45878,N_44795,N_44580);
nor U45879 (N_45879,N_44611,N_44593);
nor U45880 (N_45880,N_44296,N_44216);
nor U45881 (N_45881,N_44515,N_44051);
nor U45882 (N_45882,N_44720,N_44358);
or U45883 (N_45883,N_44655,N_44987);
xor U45884 (N_45884,N_44131,N_44003);
or U45885 (N_45885,N_44487,N_44155);
or U45886 (N_45886,N_44387,N_44694);
xnor U45887 (N_45887,N_44509,N_44237);
xor U45888 (N_45888,N_44547,N_44056);
nand U45889 (N_45889,N_44888,N_44894);
and U45890 (N_45890,N_44050,N_44199);
nand U45891 (N_45891,N_44591,N_44709);
xor U45892 (N_45892,N_44792,N_44201);
and U45893 (N_45893,N_44568,N_44796);
or U45894 (N_45894,N_44278,N_44888);
and U45895 (N_45895,N_44029,N_44193);
or U45896 (N_45896,N_44136,N_44962);
nand U45897 (N_45897,N_44561,N_44933);
nor U45898 (N_45898,N_44984,N_44085);
xor U45899 (N_45899,N_44396,N_44327);
and U45900 (N_45900,N_44516,N_44759);
or U45901 (N_45901,N_44645,N_44333);
xnor U45902 (N_45902,N_44141,N_44143);
or U45903 (N_45903,N_44968,N_44955);
or U45904 (N_45904,N_44947,N_44932);
xor U45905 (N_45905,N_44147,N_44266);
xnor U45906 (N_45906,N_44905,N_44919);
or U45907 (N_45907,N_44488,N_44081);
or U45908 (N_45908,N_44335,N_44011);
xnor U45909 (N_45909,N_44080,N_44362);
and U45910 (N_45910,N_44181,N_44349);
and U45911 (N_45911,N_44097,N_44861);
or U45912 (N_45912,N_44023,N_44116);
or U45913 (N_45913,N_44380,N_44445);
nand U45914 (N_45914,N_44086,N_44633);
or U45915 (N_45915,N_44480,N_44508);
nor U45916 (N_45916,N_44384,N_44248);
xnor U45917 (N_45917,N_44581,N_44540);
or U45918 (N_45918,N_44785,N_44248);
nand U45919 (N_45919,N_44776,N_44347);
nor U45920 (N_45920,N_44208,N_44465);
xor U45921 (N_45921,N_44225,N_44078);
nand U45922 (N_45922,N_44183,N_44268);
and U45923 (N_45923,N_44179,N_44477);
and U45924 (N_45924,N_44989,N_44775);
or U45925 (N_45925,N_44527,N_44515);
or U45926 (N_45926,N_44804,N_44572);
nand U45927 (N_45927,N_44261,N_44014);
nor U45928 (N_45928,N_44501,N_44084);
nand U45929 (N_45929,N_44944,N_44995);
and U45930 (N_45930,N_44993,N_44007);
nand U45931 (N_45931,N_44420,N_44917);
nand U45932 (N_45932,N_44976,N_44899);
xor U45933 (N_45933,N_44686,N_44900);
or U45934 (N_45934,N_44428,N_44007);
nand U45935 (N_45935,N_44376,N_44802);
or U45936 (N_45936,N_44296,N_44156);
xor U45937 (N_45937,N_44911,N_44458);
xnor U45938 (N_45938,N_44884,N_44119);
or U45939 (N_45939,N_44670,N_44380);
or U45940 (N_45940,N_44657,N_44297);
or U45941 (N_45941,N_44354,N_44003);
xor U45942 (N_45942,N_44234,N_44617);
nand U45943 (N_45943,N_44578,N_44290);
or U45944 (N_45944,N_44814,N_44317);
nor U45945 (N_45945,N_44289,N_44275);
nor U45946 (N_45946,N_44682,N_44851);
and U45947 (N_45947,N_44394,N_44244);
nand U45948 (N_45948,N_44807,N_44862);
xnor U45949 (N_45949,N_44653,N_44228);
xor U45950 (N_45950,N_44072,N_44246);
or U45951 (N_45951,N_44960,N_44987);
nand U45952 (N_45952,N_44357,N_44801);
nand U45953 (N_45953,N_44790,N_44378);
nor U45954 (N_45954,N_44921,N_44605);
nor U45955 (N_45955,N_44043,N_44326);
nor U45956 (N_45956,N_44808,N_44817);
and U45957 (N_45957,N_44001,N_44937);
and U45958 (N_45958,N_44881,N_44685);
and U45959 (N_45959,N_44186,N_44540);
and U45960 (N_45960,N_44240,N_44379);
and U45961 (N_45961,N_44365,N_44170);
and U45962 (N_45962,N_44865,N_44453);
or U45963 (N_45963,N_44740,N_44165);
nand U45964 (N_45964,N_44480,N_44370);
and U45965 (N_45965,N_44866,N_44613);
xor U45966 (N_45966,N_44882,N_44003);
or U45967 (N_45967,N_44723,N_44130);
or U45968 (N_45968,N_44043,N_44247);
nand U45969 (N_45969,N_44833,N_44783);
xor U45970 (N_45970,N_44967,N_44815);
nand U45971 (N_45971,N_44123,N_44715);
or U45972 (N_45972,N_44739,N_44711);
and U45973 (N_45973,N_44714,N_44226);
xnor U45974 (N_45974,N_44746,N_44088);
and U45975 (N_45975,N_44842,N_44897);
nand U45976 (N_45976,N_44250,N_44079);
xor U45977 (N_45977,N_44496,N_44537);
xor U45978 (N_45978,N_44704,N_44777);
xor U45979 (N_45979,N_44689,N_44962);
nand U45980 (N_45980,N_44667,N_44950);
nor U45981 (N_45981,N_44256,N_44469);
and U45982 (N_45982,N_44020,N_44441);
nor U45983 (N_45983,N_44935,N_44864);
or U45984 (N_45984,N_44804,N_44288);
xnor U45985 (N_45985,N_44448,N_44441);
and U45986 (N_45986,N_44455,N_44718);
xor U45987 (N_45987,N_44405,N_44705);
or U45988 (N_45988,N_44013,N_44861);
or U45989 (N_45989,N_44809,N_44558);
nor U45990 (N_45990,N_44093,N_44035);
and U45991 (N_45991,N_44230,N_44470);
nor U45992 (N_45992,N_44480,N_44083);
and U45993 (N_45993,N_44700,N_44538);
nand U45994 (N_45994,N_44112,N_44439);
and U45995 (N_45995,N_44246,N_44904);
xor U45996 (N_45996,N_44003,N_44524);
nor U45997 (N_45997,N_44636,N_44168);
and U45998 (N_45998,N_44831,N_44420);
nand U45999 (N_45999,N_44779,N_44240);
nor U46000 (N_46000,N_45174,N_45377);
or U46001 (N_46001,N_45934,N_45141);
nor U46002 (N_46002,N_45181,N_45721);
nor U46003 (N_46003,N_45283,N_45701);
or U46004 (N_46004,N_45384,N_45952);
and U46005 (N_46005,N_45186,N_45460);
nand U46006 (N_46006,N_45505,N_45179);
nand U46007 (N_46007,N_45447,N_45286);
nand U46008 (N_46008,N_45209,N_45289);
or U46009 (N_46009,N_45127,N_45909);
nand U46010 (N_46010,N_45243,N_45002);
and U46011 (N_46011,N_45651,N_45421);
and U46012 (N_46012,N_45249,N_45968);
or U46013 (N_46013,N_45821,N_45307);
xor U46014 (N_46014,N_45624,N_45938);
xor U46015 (N_46015,N_45622,N_45545);
nor U46016 (N_46016,N_45244,N_45414);
nor U46017 (N_46017,N_45389,N_45163);
or U46018 (N_46018,N_45479,N_45950);
or U46019 (N_46019,N_45071,N_45569);
nor U46020 (N_46020,N_45492,N_45866);
nor U46021 (N_46021,N_45014,N_45443);
nand U46022 (N_46022,N_45380,N_45501);
nand U46023 (N_46023,N_45874,N_45756);
nor U46024 (N_46024,N_45685,N_45812);
nand U46025 (N_46025,N_45082,N_45686);
xor U46026 (N_46026,N_45567,N_45769);
and U46027 (N_46027,N_45160,N_45195);
nand U46028 (N_46028,N_45172,N_45316);
and U46029 (N_46029,N_45425,N_45681);
or U46030 (N_46030,N_45099,N_45997);
xnor U46031 (N_46031,N_45493,N_45142);
nor U46032 (N_46032,N_45272,N_45930);
and U46033 (N_46033,N_45333,N_45649);
and U46034 (N_46034,N_45396,N_45003);
nand U46035 (N_46035,N_45969,N_45115);
xor U46036 (N_46036,N_45817,N_45836);
nor U46037 (N_46037,N_45096,N_45344);
nand U46038 (N_46038,N_45964,N_45843);
xor U46039 (N_46039,N_45779,N_45466);
and U46040 (N_46040,N_45093,N_45349);
nor U46041 (N_46041,N_45720,N_45089);
xor U46042 (N_46042,N_45111,N_45355);
xnor U46043 (N_46043,N_45457,N_45426);
or U46044 (N_46044,N_45700,N_45328);
or U46045 (N_46045,N_45925,N_45605);
nand U46046 (N_46046,N_45656,N_45102);
xnor U46047 (N_46047,N_45553,N_45269);
xor U46048 (N_46048,N_45016,N_45139);
or U46049 (N_46049,N_45473,N_45536);
nor U46050 (N_46050,N_45571,N_45413);
xnor U46051 (N_46051,N_45427,N_45156);
nand U46052 (N_46052,N_45816,N_45051);
nand U46053 (N_46053,N_45942,N_45653);
nor U46054 (N_46054,N_45595,N_45368);
and U46055 (N_46055,N_45372,N_45852);
or U46056 (N_46056,N_45664,N_45106);
or U46057 (N_46057,N_45130,N_45012);
nand U46058 (N_46058,N_45876,N_45728);
nor U46059 (N_46059,N_45445,N_45897);
or U46060 (N_46060,N_45116,N_45539);
xor U46061 (N_46061,N_45626,N_45914);
xnor U46062 (N_46062,N_45292,N_45066);
and U46063 (N_46063,N_45689,N_45528);
nor U46064 (N_46064,N_45207,N_45596);
or U46065 (N_46065,N_45642,N_45279);
or U46066 (N_46066,N_45036,N_45122);
and U46067 (N_46067,N_45798,N_45829);
xnor U46068 (N_46068,N_45235,N_45369);
and U46069 (N_46069,N_45119,N_45687);
or U46070 (N_46070,N_45494,N_45270);
xor U46071 (N_46071,N_45024,N_45191);
nor U46072 (N_46072,N_45205,N_45908);
nor U46073 (N_46073,N_45250,N_45778);
xnor U46074 (N_46074,N_45331,N_45029);
or U46075 (N_46075,N_45870,N_45586);
and U46076 (N_46076,N_45468,N_45076);
or U46077 (N_46077,N_45223,N_45497);
xnor U46078 (N_46078,N_45510,N_45159);
or U46079 (N_46079,N_45810,N_45788);
nor U46080 (N_46080,N_45251,N_45913);
xor U46081 (N_46081,N_45165,N_45170);
and U46082 (N_46082,N_45184,N_45435);
nor U46083 (N_46083,N_45827,N_45840);
nor U46084 (N_46084,N_45780,N_45933);
nand U46085 (N_46085,N_45234,N_45177);
nor U46086 (N_46086,N_45405,N_45782);
xor U46087 (N_46087,N_45903,N_45723);
or U46088 (N_46088,N_45302,N_45004);
xnor U46089 (N_46089,N_45169,N_45702);
nand U46090 (N_46090,N_45464,N_45027);
nor U46091 (N_46091,N_45814,N_45990);
nor U46092 (N_46092,N_45607,N_45297);
nor U46093 (N_46093,N_45200,N_45006);
nor U46094 (N_46094,N_45375,N_45485);
or U46095 (N_46095,N_45436,N_45247);
nand U46096 (N_46096,N_45703,N_45477);
or U46097 (N_46097,N_45916,N_45381);
nand U46098 (N_46098,N_45070,N_45192);
nor U46099 (N_46099,N_45188,N_45844);
xnor U46100 (N_46100,N_45920,N_45976);
nor U46101 (N_46101,N_45210,N_45786);
xor U46102 (N_46102,N_45740,N_45713);
or U46103 (N_46103,N_45676,N_45763);
nor U46104 (N_46104,N_45120,N_45290);
or U46105 (N_46105,N_45910,N_45345);
xnor U46106 (N_46106,N_45957,N_45047);
xnor U46107 (N_46107,N_45760,N_45404);
or U46108 (N_46108,N_45828,N_45987);
xor U46109 (N_46109,N_45078,N_45044);
and U46110 (N_46110,N_45892,N_45803);
and U46111 (N_46111,N_45341,N_45860);
nand U46112 (N_46112,N_45054,N_45893);
nand U46113 (N_46113,N_45011,N_45675);
or U46114 (N_46114,N_45409,N_45693);
and U46115 (N_46115,N_45100,N_45416);
nand U46116 (N_46116,N_45296,N_45264);
and U46117 (N_46117,N_45230,N_45848);
or U46118 (N_46118,N_45872,N_45972);
or U46119 (N_46119,N_45379,N_45879);
xnor U46120 (N_46120,N_45598,N_45294);
nand U46121 (N_46121,N_45726,N_45781);
nor U46122 (N_46122,N_45965,N_45901);
nand U46123 (N_46123,N_45877,N_45742);
nand U46124 (N_46124,N_45482,N_45562);
nand U46125 (N_46125,N_45696,N_45669);
or U46126 (N_46126,N_45880,N_45695);
nor U46127 (N_46127,N_45261,N_45513);
or U46128 (N_46128,N_45080,N_45481);
and U46129 (N_46129,N_45402,N_45772);
nand U46130 (N_46130,N_45144,N_45825);
nand U46131 (N_46131,N_45745,N_45017);
nand U46132 (N_46132,N_45537,N_45339);
nand U46133 (N_46133,N_45838,N_45912);
and U46134 (N_46134,N_45287,N_45523);
nand U46135 (N_46135,N_45180,N_45050);
or U46136 (N_46136,N_45796,N_45591);
or U46137 (N_46137,N_45735,N_45807);
nand U46138 (N_46138,N_45614,N_45835);
nor U46139 (N_46139,N_45398,N_45548);
nand U46140 (N_46140,N_45206,N_45657);
or U46141 (N_46141,N_45533,N_45441);
and U46142 (N_46142,N_45320,N_45574);
or U46143 (N_46143,N_45668,N_45940);
or U46144 (N_46144,N_45824,N_45581);
and U46145 (N_46145,N_45512,N_45855);
or U46146 (N_46146,N_45334,N_45609);
or U46147 (N_46147,N_45211,N_45588);
nor U46148 (N_46148,N_45258,N_45348);
or U46149 (N_46149,N_45376,N_45471);
xnor U46150 (N_46150,N_45061,N_45587);
nand U46151 (N_46151,N_45222,N_45224);
and U46152 (N_46152,N_45392,N_45145);
or U46153 (N_46153,N_45491,N_45883);
or U46154 (N_46154,N_45213,N_45431);
nand U46155 (N_46155,N_45672,N_45064);
nor U46156 (N_46156,N_45746,N_45280);
nand U46157 (N_46157,N_45982,N_45615);
xnor U46158 (N_46158,N_45551,N_45241);
xnor U46159 (N_46159,N_45303,N_45549);
xnor U46160 (N_46160,N_45087,N_45684);
and U46161 (N_46161,N_45500,N_45797);
xor U46162 (N_46162,N_45511,N_45691);
or U46163 (N_46163,N_45240,N_45789);
or U46164 (N_46164,N_45386,N_45488);
and U46165 (N_46165,N_45947,N_45366);
and U46166 (N_46166,N_45975,N_45639);
nor U46167 (N_46167,N_45801,N_45532);
xor U46168 (N_46168,N_45060,N_45709);
nor U46169 (N_46169,N_45863,N_45715);
xor U46170 (N_46170,N_45765,N_45845);
nand U46171 (N_46171,N_45319,N_45998);
and U46172 (N_46172,N_45086,N_45465);
nand U46173 (N_46173,N_45634,N_45531);
xnor U46174 (N_46174,N_45434,N_45295);
or U46175 (N_46175,N_45140,N_45198);
nand U46176 (N_46176,N_45476,N_45199);
or U46177 (N_46177,N_45365,N_45490);
and U46178 (N_46178,N_45022,N_45394);
and U46179 (N_46179,N_45853,N_45403);
nor U46180 (N_46180,N_45098,N_45800);
nand U46181 (N_46181,N_45682,N_45338);
nor U46182 (N_46182,N_45837,N_45677);
xor U46183 (N_46183,N_45045,N_45323);
nand U46184 (N_46184,N_45088,N_45919);
xnor U46185 (N_46185,N_45183,N_45229);
xnor U46186 (N_46186,N_45601,N_45805);
nand U46187 (N_46187,N_45226,N_45225);
xnor U46188 (N_46188,N_45636,N_45282);
and U46189 (N_46189,N_45541,N_45758);
nand U46190 (N_46190,N_45980,N_45887);
or U46191 (N_46191,N_45846,N_45025);
nand U46192 (N_46192,N_45711,N_45889);
or U46193 (N_46193,N_45967,N_45422);
nor U46194 (N_46194,N_45246,N_45655);
and U46195 (N_46195,N_45005,N_45019);
and U46196 (N_46196,N_45010,N_45278);
or U46197 (N_46197,N_45013,N_45898);
or U46198 (N_46198,N_45274,N_45550);
xor U46199 (N_46199,N_45714,N_45136);
nor U46200 (N_46200,N_45515,N_45298);
xor U46201 (N_46201,N_45630,N_45737);
xor U46202 (N_46202,N_45030,N_45260);
nand U46203 (N_46203,N_45208,N_45212);
xor U46204 (N_46204,N_45227,N_45754);
and U46205 (N_46205,N_45455,N_45881);
or U46206 (N_46206,N_45310,N_45809);
nand U46207 (N_46207,N_45775,N_45153);
and U46208 (N_46208,N_45750,N_45978);
or U46209 (N_46209,N_45231,N_45555);
nor U46210 (N_46210,N_45818,N_45839);
or U46211 (N_46211,N_45722,N_45654);
xnor U46212 (N_46212,N_45190,N_45018);
nor U46213 (N_46213,N_45128,N_45660);
xnor U46214 (N_46214,N_45032,N_45958);
nand U46215 (N_46215,N_45065,N_45802);
nand U46216 (N_46216,N_45167,N_45178);
nor U46217 (N_46217,N_45129,N_45804);
xor U46218 (N_46218,N_45830,N_45220);
and U46219 (N_46219,N_45641,N_45534);
nand U46220 (N_46220,N_45960,N_45945);
or U46221 (N_46221,N_45645,N_45203);
and U46222 (N_46222,N_45680,N_45164);
and U46223 (N_46223,N_45257,N_45033);
xnor U46224 (N_46224,N_45600,N_45411);
nor U46225 (N_46225,N_45196,N_45993);
xnor U46226 (N_46226,N_45939,N_45971);
and U46227 (N_46227,N_45834,N_45266);
and U46228 (N_46228,N_45718,N_45135);
xor U46229 (N_46229,N_45585,N_45273);
nand U46230 (N_46230,N_45351,N_45716);
nor U46231 (N_46231,N_45538,N_45977);
or U46232 (N_46232,N_45698,N_45520);
and U46233 (N_46233,N_45795,N_45517);
and U46234 (N_46234,N_45202,N_45518);
nor U46235 (N_46235,N_45604,N_45090);
and U46236 (N_46236,N_45899,N_45936);
and U46237 (N_46237,N_45276,N_45992);
nand U46238 (N_46238,N_45690,N_45059);
xor U46239 (N_46239,N_45643,N_45440);
and U46240 (N_46240,N_45000,N_45717);
or U46241 (N_46241,N_45900,N_45738);
nor U46242 (N_46242,N_45578,N_45193);
nor U46243 (N_46243,N_45955,N_45347);
xnor U46244 (N_46244,N_45524,N_45996);
or U46245 (N_46245,N_45766,N_45661);
nand U46246 (N_46246,N_45962,N_45057);
nand U46247 (N_46247,N_45566,N_45831);
nor U46248 (N_46248,N_45104,N_45579);
nor U46249 (N_46249,N_45388,N_45215);
and U46250 (N_46250,N_45813,N_45768);
nor U46251 (N_46251,N_45418,N_45390);
xnor U46252 (N_46252,N_45697,N_45154);
and U46253 (N_46253,N_45335,N_45616);
and U46254 (N_46254,N_45216,N_45420);
xnor U46255 (N_46255,N_45561,N_45640);
nor U46256 (N_46256,N_45478,N_45784);
or U46257 (N_46257,N_45509,N_45360);
or U46258 (N_46258,N_45162,N_45268);
xnor U46259 (N_46259,N_45646,N_45218);
nor U46260 (N_46260,N_45131,N_45073);
and U46261 (N_46261,N_45833,N_45168);
and U46262 (N_46262,N_45204,N_45451);
or U46263 (N_46263,N_45688,N_45439);
nand U46264 (N_46264,N_45028,N_45419);
or U46265 (N_46265,N_45707,N_45358);
and U46266 (N_46266,N_45725,N_45255);
nand U46267 (N_46267,N_45312,N_45037);
and U46268 (N_46268,N_45433,N_45068);
xor U46269 (N_46269,N_45951,N_45417);
and U46270 (N_46270,N_45484,N_45606);
nor U46271 (N_46271,N_45752,N_45808);
nand U46272 (N_46272,N_45741,N_45108);
or U46273 (N_46273,N_45387,N_45248);
xnor U46274 (N_46274,N_45461,N_45692);
and U46275 (N_46275,N_45429,N_45516);
xor U46276 (N_46276,N_45284,N_45861);
or U46277 (N_46277,N_45123,N_45792);
nor U46278 (N_46278,N_45446,N_45074);
and U46279 (N_46279,N_45385,N_45495);
xnor U46280 (N_46280,N_45905,N_45710);
and U46281 (N_46281,N_45974,N_45770);
xnor U46282 (N_46282,N_45767,N_45806);
or U46283 (N_46283,N_45041,N_45590);
nor U46284 (N_46284,N_45885,N_45592);
nand U46285 (N_46285,N_45790,N_45158);
nor U46286 (N_46286,N_45456,N_45869);
nand U46287 (N_46287,N_45083,N_45486);
nand U46288 (N_46288,N_45864,N_45105);
xor U46289 (N_46289,N_45932,N_45121);
xnor U46290 (N_46290,N_45391,N_45764);
and U46291 (N_46291,N_45113,N_45621);
nor U46292 (N_46292,N_45565,N_45175);
xnor U46293 (N_46293,N_45793,N_45753);
or U46294 (N_46294,N_45558,N_45020);
and U46295 (N_46295,N_45973,N_45034);
or U46296 (N_46296,N_45865,N_45890);
or U46297 (N_46297,N_45924,N_45705);
nand U46298 (N_46298,N_45617,N_45862);
xor U46299 (N_46299,N_45514,N_45126);
or U46300 (N_46300,N_45719,N_45777);
nor U46301 (N_46301,N_45091,N_45171);
nor U46302 (N_46302,N_45603,N_45929);
nand U46303 (N_46303,N_45543,N_45888);
or U46304 (N_46304,N_45743,N_45300);
nand U46305 (N_46305,N_45277,N_45330);
or U46306 (N_46306,N_45281,N_45927);
nand U46307 (N_46307,N_45730,N_45530);
and U46308 (N_46308,N_45739,N_45546);
and U46309 (N_46309,N_45859,N_45894);
nor U46310 (N_46310,N_45378,N_45291);
nand U46311 (N_46311,N_45773,N_45069);
or U46312 (N_46312,N_45125,N_45921);
nor U46313 (N_46313,N_45820,N_45428);
nand U46314 (N_46314,N_45991,N_45946);
nand U46315 (N_46315,N_45308,N_45503);
nor U46316 (N_46316,N_45635,N_45023);
or U46317 (N_46317,N_45662,N_45670);
xor U46318 (N_46318,N_45999,N_45611);
nor U46319 (N_46319,N_45309,N_45265);
xnor U46320 (N_46320,N_45540,N_45712);
xnor U46321 (N_46321,N_45573,N_45554);
or U46322 (N_46322,N_45529,N_45794);
and U46323 (N_46323,N_45917,N_45984);
nand U46324 (N_46324,N_45610,N_45103);
and U46325 (N_46325,N_45293,N_45733);
xnor U46326 (N_46326,N_45650,N_45665);
nand U46327 (N_46327,N_45467,N_45242);
nor U46328 (N_46328,N_45474,N_45233);
nand U46329 (N_46329,N_45432,N_45382);
or U46330 (N_46330,N_45631,N_45854);
or U46331 (N_46331,N_45744,N_45961);
or U46332 (N_46332,N_45480,N_45363);
nand U46333 (N_46333,N_45544,N_45079);
and U46334 (N_46334,N_45706,N_45075);
nand U46335 (N_46335,N_45393,N_45732);
nand U46336 (N_46336,N_45943,N_45849);
or U46337 (N_46337,N_45979,N_45150);
or U46338 (N_46338,N_45437,N_45954);
or U46339 (N_46339,N_45067,N_45847);
nor U46340 (N_46340,N_45340,N_45557);
nor U46341 (N_46341,N_45904,N_45949);
and U46342 (N_46342,N_45256,N_45462);
or U46343 (N_46343,N_45867,N_45499);
nand U46344 (N_46344,N_45875,N_45584);
nor U46345 (N_46345,N_45062,N_45931);
or U46346 (N_46346,N_45350,N_45217);
and U46347 (N_46347,N_45542,N_45053);
xnor U46348 (N_46348,N_45423,N_45058);
nor U46349 (N_46349,N_45252,N_45117);
nand U46350 (N_46350,N_45519,N_45771);
nor U46351 (N_46351,N_45408,N_45759);
nor U46352 (N_46352,N_45472,N_45629);
nand U46353 (N_46353,N_45995,N_45114);
or U46354 (N_46354,N_45666,N_45221);
and U46355 (N_46355,N_45001,N_45857);
xor U46356 (N_46356,N_45329,N_45507);
and U46357 (N_46357,N_45267,N_45245);
nand U46358 (N_46358,N_45325,N_45371);
nor U46359 (N_46359,N_45658,N_45774);
or U46360 (N_46360,N_45194,N_45459);
nor U46361 (N_46361,N_45487,N_45694);
or U46362 (N_46362,N_45956,N_45056);
nand U46363 (N_46363,N_45783,N_45356);
nand U46364 (N_46364,N_45747,N_45236);
nand U46365 (N_46365,N_45948,N_45580);
and U46366 (N_46366,N_45620,N_45757);
or U46367 (N_46367,N_45185,N_45253);
nand U46368 (N_46368,N_45346,N_45021);
nand U46369 (N_46369,N_45452,N_45438);
xnor U46370 (N_46370,N_45568,N_45966);
nor U46371 (N_46371,N_45151,N_45597);
xnor U46372 (N_46372,N_45077,N_45659);
and U46373 (N_46373,N_45370,N_45138);
nand U46374 (N_46374,N_45667,N_45444);
and U46375 (N_46375,N_45400,N_45674);
or U46376 (N_46376,N_45173,N_45575);
and U46377 (N_46377,N_45944,N_45623);
nor U46378 (N_46378,N_45547,N_45647);
or U46379 (N_46379,N_45124,N_45166);
and U46380 (N_46380,N_45084,N_45040);
and U46381 (N_46381,N_45092,N_45442);
nor U46382 (N_46382,N_45851,N_45787);
and U46383 (N_46383,N_45318,N_45981);
xor U46384 (N_46384,N_45594,N_45638);
or U46385 (N_46385,N_45357,N_45288);
nor U46386 (N_46386,N_45526,N_45858);
nand U46387 (N_46387,N_45353,N_45373);
and U46388 (N_46388,N_45989,N_45201);
or U46389 (N_46389,N_45699,N_45039);
nor U46390 (N_46390,N_45362,N_45301);
or U46391 (N_46391,N_45886,N_45147);
or U46392 (N_46392,N_45359,N_45095);
nor U46393 (N_46393,N_45475,N_45237);
and U46394 (N_46394,N_45755,N_45271);
and U46395 (N_46395,N_45628,N_45663);
and U46396 (N_46396,N_45959,N_45963);
xnor U46397 (N_46397,N_45454,N_45046);
or U46398 (N_46398,N_45397,N_45238);
nor U46399 (N_46399,N_45107,N_45727);
nor U46400 (N_46400,N_45315,N_45430);
nand U46401 (N_46401,N_45751,N_45826);
nor U46402 (N_46402,N_45923,N_45305);
nand U46403 (N_46403,N_45232,N_45842);
xor U46404 (N_46404,N_45583,N_45704);
xor U46405 (N_46405,N_45941,N_45327);
and U46406 (N_46406,N_45008,N_45915);
xnor U46407 (N_46407,N_45572,N_45593);
xnor U46408 (N_46408,N_45506,N_45508);
nor U46409 (N_46409,N_45907,N_45819);
or U46410 (N_46410,N_45239,N_45026);
or U46411 (N_46411,N_45407,N_45326);
and U46412 (N_46412,N_45577,N_45986);
or U46413 (N_46413,N_45453,N_45254);
nor U46414 (N_46414,N_45094,N_45731);
or U46415 (N_46415,N_45152,N_45724);
and U46416 (N_46416,N_45343,N_45134);
and U46417 (N_46417,N_45832,N_45354);
xnor U46418 (N_46418,N_45483,N_45321);
and U46419 (N_46419,N_45785,N_45361);
xor U46420 (N_46420,N_45791,N_45928);
nor U46421 (N_46421,N_45502,N_45560);
and U46422 (N_46422,N_45009,N_45926);
xnor U46423 (N_46423,N_45214,N_45148);
or U46424 (N_46424,N_45395,N_45157);
and U46425 (N_46425,N_45262,N_45504);
or U46426 (N_46426,N_45263,N_45182);
and U46427 (N_46427,N_45608,N_45463);
or U46428 (N_46428,N_45679,N_45856);
and U46429 (N_46429,N_45552,N_45161);
and U46430 (N_46430,N_45228,N_45884);
xnor U46431 (N_46431,N_45132,N_45342);
nand U46432 (N_46432,N_45850,N_45133);
or U46433 (N_46433,N_45563,N_45469);
nor U46434 (N_46434,N_45895,N_45306);
or U46435 (N_46435,N_45015,N_45776);
and U46436 (N_46436,N_45906,N_45424);
xor U46437 (N_46437,N_45868,N_45007);
nand U46438 (N_46438,N_45873,N_45085);
nand U46439 (N_46439,N_45599,N_45648);
nand U46440 (N_46440,N_45048,N_45891);
nand U46441 (N_46441,N_45613,N_45322);
and U46442 (N_46442,N_45644,N_45458);
and U46443 (N_46443,N_45337,N_45311);
and U46444 (N_46444,N_45527,N_45412);
nand U46445 (N_46445,N_45811,N_45734);
and U46446 (N_46446,N_45749,N_45364);
and U46447 (N_46447,N_45678,N_45799);
or U46448 (N_46448,N_45922,N_45304);
nor U46449 (N_46449,N_45761,N_45918);
xor U46450 (N_46450,N_45970,N_45822);
or U46451 (N_46451,N_45633,N_45612);
nor U46452 (N_46452,N_45521,N_45072);
nor U46453 (N_46453,N_45031,N_45299);
or U46454 (N_46454,N_45219,N_45602);
nand U46455 (N_46455,N_45823,N_45042);
xnor U46456 (N_46456,N_45189,N_45994);
xnor U46457 (N_46457,N_45937,N_45671);
and U46458 (N_46458,N_45275,N_45143);
and U46459 (N_46459,N_45582,N_45498);
and U46460 (N_46460,N_45559,N_45383);
nor U46461 (N_46461,N_45496,N_45197);
xor U46462 (N_46462,N_45259,N_45352);
or U46463 (N_46463,N_45564,N_45570);
nand U46464 (N_46464,N_45109,N_45762);
nor U46465 (N_46465,N_45415,N_45187);
nand U46466 (N_46466,N_45556,N_45576);
or U46467 (N_46467,N_45882,N_45406);
nor U46468 (N_46468,N_45841,N_45399);
and U46469 (N_46469,N_45324,N_45450);
nand U46470 (N_46470,N_45935,N_45055);
nor U46471 (N_46471,N_45625,N_45317);
or U46472 (N_46472,N_45522,N_45449);
nor U46473 (N_46473,N_45708,N_45049);
xor U46474 (N_46474,N_45652,N_45673);
or U46475 (N_46475,N_45902,N_45911);
nand U46476 (N_46476,N_45632,N_45637);
or U46477 (N_46477,N_45410,N_45367);
or U46478 (N_46478,N_45285,N_45101);
or U46479 (N_46479,N_45896,N_45043);
nand U46480 (N_46480,N_45149,N_45953);
xnor U46481 (N_46481,N_45332,N_45314);
nand U46482 (N_46482,N_45110,N_45118);
nor U46483 (N_46483,N_45097,N_45683);
nor U46484 (N_46484,N_45470,N_45815);
nor U46485 (N_46485,N_45146,N_45176);
and U46486 (N_46486,N_45589,N_45052);
or U46487 (N_46487,N_45983,N_45988);
xor U46488 (N_46488,N_45736,N_45535);
xor U46489 (N_46489,N_45878,N_45374);
nor U46490 (N_46490,N_45313,N_45448);
xor U46491 (N_46491,N_45038,N_45489);
nor U46492 (N_46492,N_45137,N_45112);
nor U46493 (N_46493,N_45155,N_45627);
or U46494 (N_46494,N_45729,N_45401);
nor U46495 (N_46495,N_45336,N_45748);
nand U46496 (N_46496,N_45035,N_45618);
nand U46497 (N_46497,N_45871,N_45619);
xor U46498 (N_46498,N_45985,N_45081);
nor U46499 (N_46499,N_45063,N_45525);
or U46500 (N_46500,N_45240,N_45371);
nand U46501 (N_46501,N_45156,N_45310);
and U46502 (N_46502,N_45724,N_45934);
nor U46503 (N_46503,N_45837,N_45070);
xnor U46504 (N_46504,N_45056,N_45823);
and U46505 (N_46505,N_45194,N_45053);
or U46506 (N_46506,N_45724,N_45682);
xnor U46507 (N_46507,N_45488,N_45531);
or U46508 (N_46508,N_45716,N_45051);
or U46509 (N_46509,N_45801,N_45450);
nand U46510 (N_46510,N_45412,N_45194);
or U46511 (N_46511,N_45217,N_45563);
or U46512 (N_46512,N_45966,N_45525);
nand U46513 (N_46513,N_45567,N_45495);
or U46514 (N_46514,N_45467,N_45855);
and U46515 (N_46515,N_45725,N_45959);
nand U46516 (N_46516,N_45094,N_45004);
nor U46517 (N_46517,N_45980,N_45766);
nor U46518 (N_46518,N_45174,N_45178);
or U46519 (N_46519,N_45003,N_45127);
and U46520 (N_46520,N_45936,N_45011);
nand U46521 (N_46521,N_45209,N_45315);
xor U46522 (N_46522,N_45950,N_45547);
nand U46523 (N_46523,N_45013,N_45234);
and U46524 (N_46524,N_45851,N_45566);
nor U46525 (N_46525,N_45383,N_45841);
or U46526 (N_46526,N_45239,N_45321);
nor U46527 (N_46527,N_45914,N_45261);
nor U46528 (N_46528,N_45735,N_45519);
nor U46529 (N_46529,N_45409,N_45424);
or U46530 (N_46530,N_45217,N_45890);
or U46531 (N_46531,N_45536,N_45282);
or U46532 (N_46532,N_45131,N_45404);
and U46533 (N_46533,N_45240,N_45937);
or U46534 (N_46534,N_45988,N_45944);
xor U46535 (N_46535,N_45618,N_45703);
or U46536 (N_46536,N_45318,N_45287);
or U46537 (N_46537,N_45686,N_45591);
xor U46538 (N_46538,N_45388,N_45216);
nand U46539 (N_46539,N_45430,N_45100);
xnor U46540 (N_46540,N_45344,N_45843);
nand U46541 (N_46541,N_45596,N_45999);
or U46542 (N_46542,N_45960,N_45207);
and U46543 (N_46543,N_45683,N_45421);
nor U46544 (N_46544,N_45503,N_45761);
nand U46545 (N_46545,N_45521,N_45401);
nor U46546 (N_46546,N_45133,N_45342);
xnor U46547 (N_46547,N_45579,N_45549);
and U46548 (N_46548,N_45108,N_45126);
nand U46549 (N_46549,N_45467,N_45900);
xnor U46550 (N_46550,N_45677,N_45009);
nand U46551 (N_46551,N_45563,N_45832);
nand U46552 (N_46552,N_45164,N_45081);
nor U46553 (N_46553,N_45610,N_45101);
and U46554 (N_46554,N_45520,N_45407);
nor U46555 (N_46555,N_45642,N_45784);
nor U46556 (N_46556,N_45382,N_45401);
or U46557 (N_46557,N_45424,N_45276);
nor U46558 (N_46558,N_45378,N_45790);
nor U46559 (N_46559,N_45106,N_45277);
and U46560 (N_46560,N_45362,N_45210);
nand U46561 (N_46561,N_45926,N_45218);
or U46562 (N_46562,N_45041,N_45585);
and U46563 (N_46563,N_45320,N_45575);
xnor U46564 (N_46564,N_45112,N_45201);
and U46565 (N_46565,N_45229,N_45894);
nand U46566 (N_46566,N_45406,N_45335);
or U46567 (N_46567,N_45236,N_45476);
xor U46568 (N_46568,N_45642,N_45043);
and U46569 (N_46569,N_45705,N_45214);
or U46570 (N_46570,N_45238,N_45482);
nand U46571 (N_46571,N_45155,N_45625);
xor U46572 (N_46572,N_45442,N_45836);
nor U46573 (N_46573,N_45106,N_45362);
xor U46574 (N_46574,N_45035,N_45823);
xor U46575 (N_46575,N_45895,N_45708);
and U46576 (N_46576,N_45294,N_45538);
and U46577 (N_46577,N_45679,N_45241);
or U46578 (N_46578,N_45859,N_45945);
nor U46579 (N_46579,N_45761,N_45754);
and U46580 (N_46580,N_45517,N_45927);
or U46581 (N_46581,N_45988,N_45764);
and U46582 (N_46582,N_45596,N_45845);
and U46583 (N_46583,N_45303,N_45046);
or U46584 (N_46584,N_45564,N_45013);
nand U46585 (N_46585,N_45722,N_45972);
nand U46586 (N_46586,N_45843,N_45246);
and U46587 (N_46587,N_45527,N_45192);
nor U46588 (N_46588,N_45434,N_45602);
nand U46589 (N_46589,N_45520,N_45197);
nor U46590 (N_46590,N_45753,N_45583);
or U46591 (N_46591,N_45597,N_45484);
xor U46592 (N_46592,N_45693,N_45173);
nor U46593 (N_46593,N_45344,N_45721);
or U46594 (N_46594,N_45147,N_45761);
nor U46595 (N_46595,N_45635,N_45177);
nor U46596 (N_46596,N_45415,N_45807);
and U46597 (N_46597,N_45148,N_45820);
and U46598 (N_46598,N_45999,N_45713);
xor U46599 (N_46599,N_45266,N_45281);
nor U46600 (N_46600,N_45664,N_45900);
nand U46601 (N_46601,N_45212,N_45304);
xnor U46602 (N_46602,N_45529,N_45511);
nand U46603 (N_46603,N_45822,N_45739);
or U46604 (N_46604,N_45152,N_45048);
nor U46605 (N_46605,N_45483,N_45263);
xnor U46606 (N_46606,N_45682,N_45526);
xnor U46607 (N_46607,N_45606,N_45316);
and U46608 (N_46608,N_45327,N_45709);
or U46609 (N_46609,N_45754,N_45935);
or U46610 (N_46610,N_45159,N_45939);
nand U46611 (N_46611,N_45232,N_45803);
and U46612 (N_46612,N_45254,N_45204);
or U46613 (N_46613,N_45833,N_45416);
nor U46614 (N_46614,N_45630,N_45691);
or U46615 (N_46615,N_45701,N_45633);
nor U46616 (N_46616,N_45294,N_45858);
or U46617 (N_46617,N_45154,N_45012);
or U46618 (N_46618,N_45680,N_45184);
or U46619 (N_46619,N_45599,N_45808);
nor U46620 (N_46620,N_45293,N_45634);
or U46621 (N_46621,N_45230,N_45415);
or U46622 (N_46622,N_45330,N_45662);
and U46623 (N_46623,N_45634,N_45408);
and U46624 (N_46624,N_45731,N_45092);
nand U46625 (N_46625,N_45112,N_45120);
xor U46626 (N_46626,N_45065,N_45631);
nand U46627 (N_46627,N_45989,N_45920);
xor U46628 (N_46628,N_45572,N_45053);
or U46629 (N_46629,N_45141,N_45128);
and U46630 (N_46630,N_45119,N_45987);
xnor U46631 (N_46631,N_45702,N_45270);
or U46632 (N_46632,N_45715,N_45896);
or U46633 (N_46633,N_45243,N_45494);
nand U46634 (N_46634,N_45622,N_45003);
and U46635 (N_46635,N_45552,N_45807);
xnor U46636 (N_46636,N_45845,N_45818);
or U46637 (N_46637,N_45204,N_45516);
nor U46638 (N_46638,N_45373,N_45328);
nand U46639 (N_46639,N_45467,N_45236);
nor U46640 (N_46640,N_45414,N_45394);
and U46641 (N_46641,N_45595,N_45448);
xnor U46642 (N_46642,N_45006,N_45928);
xor U46643 (N_46643,N_45245,N_45955);
nand U46644 (N_46644,N_45333,N_45243);
nand U46645 (N_46645,N_45434,N_45259);
or U46646 (N_46646,N_45852,N_45818);
xnor U46647 (N_46647,N_45506,N_45967);
and U46648 (N_46648,N_45350,N_45489);
nand U46649 (N_46649,N_45512,N_45394);
and U46650 (N_46650,N_45148,N_45387);
and U46651 (N_46651,N_45778,N_45796);
nand U46652 (N_46652,N_45212,N_45967);
xor U46653 (N_46653,N_45438,N_45378);
xnor U46654 (N_46654,N_45941,N_45093);
and U46655 (N_46655,N_45923,N_45042);
xor U46656 (N_46656,N_45321,N_45392);
nand U46657 (N_46657,N_45659,N_45939);
nand U46658 (N_46658,N_45664,N_45272);
nand U46659 (N_46659,N_45545,N_45392);
or U46660 (N_46660,N_45981,N_45645);
xor U46661 (N_46661,N_45658,N_45421);
or U46662 (N_46662,N_45563,N_45170);
nand U46663 (N_46663,N_45925,N_45439);
nor U46664 (N_46664,N_45636,N_45003);
xnor U46665 (N_46665,N_45993,N_45149);
and U46666 (N_46666,N_45742,N_45820);
nor U46667 (N_46667,N_45409,N_45817);
and U46668 (N_46668,N_45660,N_45530);
and U46669 (N_46669,N_45841,N_45798);
nor U46670 (N_46670,N_45378,N_45774);
nand U46671 (N_46671,N_45835,N_45264);
xnor U46672 (N_46672,N_45270,N_45669);
nor U46673 (N_46673,N_45321,N_45711);
nand U46674 (N_46674,N_45167,N_45060);
and U46675 (N_46675,N_45338,N_45097);
nor U46676 (N_46676,N_45405,N_45758);
and U46677 (N_46677,N_45869,N_45152);
or U46678 (N_46678,N_45273,N_45374);
xor U46679 (N_46679,N_45319,N_45672);
and U46680 (N_46680,N_45283,N_45051);
xor U46681 (N_46681,N_45678,N_45817);
xor U46682 (N_46682,N_45321,N_45983);
nor U46683 (N_46683,N_45991,N_45177);
or U46684 (N_46684,N_45214,N_45680);
and U46685 (N_46685,N_45710,N_45735);
nand U46686 (N_46686,N_45314,N_45947);
nor U46687 (N_46687,N_45664,N_45235);
nor U46688 (N_46688,N_45755,N_45310);
xnor U46689 (N_46689,N_45458,N_45928);
nand U46690 (N_46690,N_45744,N_45530);
and U46691 (N_46691,N_45019,N_45735);
xor U46692 (N_46692,N_45133,N_45972);
or U46693 (N_46693,N_45953,N_45983);
nand U46694 (N_46694,N_45793,N_45744);
xor U46695 (N_46695,N_45770,N_45246);
and U46696 (N_46696,N_45802,N_45103);
nor U46697 (N_46697,N_45393,N_45927);
and U46698 (N_46698,N_45217,N_45936);
xnor U46699 (N_46699,N_45131,N_45246);
xor U46700 (N_46700,N_45201,N_45756);
nor U46701 (N_46701,N_45211,N_45470);
nand U46702 (N_46702,N_45756,N_45530);
or U46703 (N_46703,N_45919,N_45308);
xor U46704 (N_46704,N_45168,N_45759);
xor U46705 (N_46705,N_45734,N_45549);
nand U46706 (N_46706,N_45498,N_45528);
or U46707 (N_46707,N_45204,N_45828);
or U46708 (N_46708,N_45352,N_45382);
nor U46709 (N_46709,N_45414,N_45326);
and U46710 (N_46710,N_45017,N_45854);
nand U46711 (N_46711,N_45726,N_45317);
nor U46712 (N_46712,N_45550,N_45637);
nand U46713 (N_46713,N_45004,N_45847);
and U46714 (N_46714,N_45859,N_45456);
nor U46715 (N_46715,N_45987,N_45712);
or U46716 (N_46716,N_45879,N_45517);
nand U46717 (N_46717,N_45633,N_45528);
nand U46718 (N_46718,N_45601,N_45174);
or U46719 (N_46719,N_45632,N_45371);
xnor U46720 (N_46720,N_45658,N_45198);
nand U46721 (N_46721,N_45341,N_45870);
or U46722 (N_46722,N_45899,N_45480);
nand U46723 (N_46723,N_45212,N_45378);
and U46724 (N_46724,N_45076,N_45498);
nand U46725 (N_46725,N_45959,N_45968);
xor U46726 (N_46726,N_45538,N_45025);
nand U46727 (N_46727,N_45742,N_45172);
xor U46728 (N_46728,N_45841,N_45990);
xor U46729 (N_46729,N_45726,N_45004);
nor U46730 (N_46730,N_45709,N_45577);
nor U46731 (N_46731,N_45137,N_45790);
nor U46732 (N_46732,N_45301,N_45646);
or U46733 (N_46733,N_45880,N_45740);
xnor U46734 (N_46734,N_45488,N_45460);
nand U46735 (N_46735,N_45999,N_45508);
xnor U46736 (N_46736,N_45831,N_45141);
and U46737 (N_46737,N_45295,N_45214);
or U46738 (N_46738,N_45276,N_45331);
or U46739 (N_46739,N_45274,N_45845);
nor U46740 (N_46740,N_45507,N_45137);
nand U46741 (N_46741,N_45811,N_45781);
nand U46742 (N_46742,N_45173,N_45497);
nand U46743 (N_46743,N_45379,N_45405);
nand U46744 (N_46744,N_45979,N_45295);
or U46745 (N_46745,N_45547,N_45513);
or U46746 (N_46746,N_45228,N_45865);
nor U46747 (N_46747,N_45790,N_45321);
and U46748 (N_46748,N_45109,N_45927);
or U46749 (N_46749,N_45879,N_45810);
nand U46750 (N_46750,N_45062,N_45662);
nand U46751 (N_46751,N_45692,N_45401);
xnor U46752 (N_46752,N_45305,N_45539);
or U46753 (N_46753,N_45255,N_45266);
and U46754 (N_46754,N_45918,N_45573);
or U46755 (N_46755,N_45226,N_45060);
nand U46756 (N_46756,N_45761,N_45769);
nand U46757 (N_46757,N_45684,N_45978);
nand U46758 (N_46758,N_45232,N_45515);
and U46759 (N_46759,N_45433,N_45602);
nand U46760 (N_46760,N_45654,N_45353);
xor U46761 (N_46761,N_45232,N_45469);
and U46762 (N_46762,N_45137,N_45281);
or U46763 (N_46763,N_45015,N_45748);
and U46764 (N_46764,N_45986,N_45390);
xnor U46765 (N_46765,N_45566,N_45134);
xnor U46766 (N_46766,N_45039,N_45915);
xor U46767 (N_46767,N_45999,N_45187);
or U46768 (N_46768,N_45117,N_45361);
and U46769 (N_46769,N_45585,N_45376);
and U46770 (N_46770,N_45890,N_45366);
nand U46771 (N_46771,N_45734,N_45403);
or U46772 (N_46772,N_45237,N_45083);
and U46773 (N_46773,N_45347,N_45711);
or U46774 (N_46774,N_45471,N_45342);
nand U46775 (N_46775,N_45723,N_45467);
xor U46776 (N_46776,N_45344,N_45578);
or U46777 (N_46777,N_45496,N_45559);
xor U46778 (N_46778,N_45898,N_45483);
or U46779 (N_46779,N_45413,N_45320);
nor U46780 (N_46780,N_45320,N_45846);
nand U46781 (N_46781,N_45885,N_45391);
and U46782 (N_46782,N_45719,N_45922);
xor U46783 (N_46783,N_45375,N_45645);
and U46784 (N_46784,N_45064,N_45826);
nand U46785 (N_46785,N_45905,N_45688);
xor U46786 (N_46786,N_45751,N_45687);
xor U46787 (N_46787,N_45931,N_45938);
nor U46788 (N_46788,N_45782,N_45843);
nor U46789 (N_46789,N_45568,N_45274);
nor U46790 (N_46790,N_45073,N_45915);
or U46791 (N_46791,N_45342,N_45900);
and U46792 (N_46792,N_45862,N_45535);
xnor U46793 (N_46793,N_45309,N_45662);
or U46794 (N_46794,N_45793,N_45315);
or U46795 (N_46795,N_45652,N_45995);
nand U46796 (N_46796,N_45973,N_45010);
or U46797 (N_46797,N_45510,N_45089);
and U46798 (N_46798,N_45544,N_45773);
nand U46799 (N_46799,N_45277,N_45237);
nand U46800 (N_46800,N_45949,N_45986);
nor U46801 (N_46801,N_45086,N_45724);
or U46802 (N_46802,N_45790,N_45007);
nor U46803 (N_46803,N_45251,N_45652);
or U46804 (N_46804,N_45487,N_45485);
and U46805 (N_46805,N_45430,N_45547);
or U46806 (N_46806,N_45497,N_45789);
and U46807 (N_46807,N_45864,N_45274);
xor U46808 (N_46808,N_45724,N_45323);
xnor U46809 (N_46809,N_45240,N_45646);
and U46810 (N_46810,N_45255,N_45969);
or U46811 (N_46811,N_45027,N_45887);
nor U46812 (N_46812,N_45085,N_45096);
or U46813 (N_46813,N_45385,N_45449);
nor U46814 (N_46814,N_45094,N_45363);
nor U46815 (N_46815,N_45858,N_45470);
nand U46816 (N_46816,N_45708,N_45248);
or U46817 (N_46817,N_45618,N_45473);
xor U46818 (N_46818,N_45622,N_45307);
nor U46819 (N_46819,N_45791,N_45638);
or U46820 (N_46820,N_45093,N_45542);
nor U46821 (N_46821,N_45527,N_45042);
xnor U46822 (N_46822,N_45576,N_45680);
or U46823 (N_46823,N_45433,N_45734);
and U46824 (N_46824,N_45241,N_45354);
nor U46825 (N_46825,N_45265,N_45032);
or U46826 (N_46826,N_45843,N_45721);
nor U46827 (N_46827,N_45892,N_45535);
xor U46828 (N_46828,N_45709,N_45541);
and U46829 (N_46829,N_45853,N_45065);
or U46830 (N_46830,N_45708,N_45692);
or U46831 (N_46831,N_45318,N_45782);
or U46832 (N_46832,N_45465,N_45686);
or U46833 (N_46833,N_45579,N_45046);
xor U46834 (N_46834,N_45858,N_45549);
and U46835 (N_46835,N_45757,N_45611);
nand U46836 (N_46836,N_45390,N_45559);
nor U46837 (N_46837,N_45259,N_45970);
nor U46838 (N_46838,N_45532,N_45230);
nor U46839 (N_46839,N_45223,N_45301);
nor U46840 (N_46840,N_45552,N_45933);
xnor U46841 (N_46841,N_45553,N_45200);
xnor U46842 (N_46842,N_45605,N_45163);
and U46843 (N_46843,N_45670,N_45789);
xnor U46844 (N_46844,N_45959,N_45435);
nor U46845 (N_46845,N_45921,N_45118);
nand U46846 (N_46846,N_45883,N_45555);
xnor U46847 (N_46847,N_45184,N_45289);
or U46848 (N_46848,N_45131,N_45248);
xnor U46849 (N_46849,N_45228,N_45006);
or U46850 (N_46850,N_45186,N_45846);
and U46851 (N_46851,N_45912,N_45096);
nor U46852 (N_46852,N_45511,N_45313);
or U46853 (N_46853,N_45252,N_45391);
or U46854 (N_46854,N_45451,N_45274);
nand U46855 (N_46855,N_45524,N_45476);
xnor U46856 (N_46856,N_45248,N_45180);
nand U46857 (N_46857,N_45286,N_45126);
nor U46858 (N_46858,N_45976,N_45836);
and U46859 (N_46859,N_45106,N_45263);
and U46860 (N_46860,N_45194,N_45260);
nand U46861 (N_46861,N_45917,N_45953);
or U46862 (N_46862,N_45154,N_45101);
and U46863 (N_46863,N_45175,N_45213);
nor U46864 (N_46864,N_45275,N_45558);
and U46865 (N_46865,N_45535,N_45241);
nand U46866 (N_46866,N_45744,N_45331);
nor U46867 (N_46867,N_45013,N_45695);
xnor U46868 (N_46868,N_45398,N_45934);
and U46869 (N_46869,N_45349,N_45938);
and U46870 (N_46870,N_45453,N_45845);
and U46871 (N_46871,N_45552,N_45748);
nor U46872 (N_46872,N_45407,N_45050);
nor U46873 (N_46873,N_45610,N_45133);
nand U46874 (N_46874,N_45619,N_45359);
nor U46875 (N_46875,N_45895,N_45360);
nor U46876 (N_46876,N_45512,N_45074);
xor U46877 (N_46877,N_45414,N_45737);
xnor U46878 (N_46878,N_45674,N_45023);
xor U46879 (N_46879,N_45661,N_45084);
xor U46880 (N_46880,N_45659,N_45656);
or U46881 (N_46881,N_45124,N_45659);
and U46882 (N_46882,N_45152,N_45431);
xnor U46883 (N_46883,N_45683,N_45248);
or U46884 (N_46884,N_45173,N_45374);
nand U46885 (N_46885,N_45803,N_45169);
xnor U46886 (N_46886,N_45716,N_45289);
nor U46887 (N_46887,N_45739,N_45795);
xor U46888 (N_46888,N_45144,N_45215);
or U46889 (N_46889,N_45070,N_45996);
or U46890 (N_46890,N_45494,N_45979);
and U46891 (N_46891,N_45309,N_45676);
or U46892 (N_46892,N_45504,N_45992);
nor U46893 (N_46893,N_45857,N_45479);
and U46894 (N_46894,N_45251,N_45601);
xnor U46895 (N_46895,N_45550,N_45991);
nand U46896 (N_46896,N_45500,N_45638);
nand U46897 (N_46897,N_45704,N_45271);
nor U46898 (N_46898,N_45048,N_45481);
xnor U46899 (N_46899,N_45029,N_45110);
nor U46900 (N_46900,N_45773,N_45534);
or U46901 (N_46901,N_45774,N_45922);
or U46902 (N_46902,N_45186,N_45670);
nor U46903 (N_46903,N_45839,N_45746);
nor U46904 (N_46904,N_45793,N_45542);
xnor U46905 (N_46905,N_45768,N_45700);
xnor U46906 (N_46906,N_45204,N_45968);
xnor U46907 (N_46907,N_45452,N_45944);
nor U46908 (N_46908,N_45359,N_45890);
xnor U46909 (N_46909,N_45594,N_45957);
nor U46910 (N_46910,N_45728,N_45674);
and U46911 (N_46911,N_45439,N_45099);
xor U46912 (N_46912,N_45505,N_45096);
nand U46913 (N_46913,N_45345,N_45189);
or U46914 (N_46914,N_45905,N_45754);
or U46915 (N_46915,N_45739,N_45828);
and U46916 (N_46916,N_45022,N_45675);
and U46917 (N_46917,N_45445,N_45666);
or U46918 (N_46918,N_45950,N_45328);
or U46919 (N_46919,N_45190,N_45779);
nor U46920 (N_46920,N_45341,N_45648);
nand U46921 (N_46921,N_45505,N_45172);
and U46922 (N_46922,N_45007,N_45397);
xor U46923 (N_46923,N_45132,N_45838);
nand U46924 (N_46924,N_45433,N_45406);
nand U46925 (N_46925,N_45859,N_45995);
nor U46926 (N_46926,N_45616,N_45609);
nand U46927 (N_46927,N_45479,N_45733);
xnor U46928 (N_46928,N_45659,N_45219);
nor U46929 (N_46929,N_45452,N_45510);
xnor U46930 (N_46930,N_45305,N_45641);
nor U46931 (N_46931,N_45399,N_45668);
xor U46932 (N_46932,N_45688,N_45767);
and U46933 (N_46933,N_45254,N_45933);
and U46934 (N_46934,N_45160,N_45253);
and U46935 (N_46935,N_45221,N_45479);
nor U46936 (N_46936,N_45842,N_45453);
and U46937 (N_46937,N_45794,N_45222);
nand U46938 (N_46938,N_45932,N_45370);
and U46939 (N_46939,N_45095,N_45672);
or U46940 (N_46940,N_45438,N_45832);
xor U46941 (N_46941,N_45701,N_45950);
xnor U46942 (N_46942,N_45229,N_45213);
and U46943 (N_46943,N_45553,N_45811);
or U46944 (N_46944,N_45803,N_45096);
nor U46945 (N_46945,N_45824,N_45784);
nor U46946 (N_46946,N_45881,N_45158);
nor U46947 (N_46947,N_45038,N_45059);
or U46948 (N_46948,N_45580,N_45783);
nor U46949 (N_46949,N_45094,N_45542);
or U46950 (N_46950,N_45838,N_45571);
nor U46951 (N_46951,N_45690,N_45646);
xor U46952 (N_46952,N_45644,N_45452);
nand U46953 (N_46953,N_45402,N_45066);
xnor U46954 (N_46954,N_45145,N_45652);
nand U46955 (N_46955,N_45559,N_45718);
nand U46956 (N_46956,N_45825,N_45531);
xor U46957 (N_46957,N_45943,N_45401);
and U46958 (N_46958,N_45601,N_45887);
nor U46959 (N_46959,N_45322,N_45342);
xor U46960 (N_46960,N_45750,N_45855);
nor U46961 (N_46961,N_45848,N_45246);
nor U46962 (N_46962,N_45570,N_45462);
nor U46963 (N_46963,N_45747,N_45686);
nand U46964 (N_46964,N_45209,N_45961);
and U46965 (N_46965,N_45015,N_45914);
nor U46966 (N_46966,N_45340,N_45022);
and U46967 (N_46967,N_45402,N_45821);
or U46968 (N_46968,N_45672,N_45426);
nand U46969 (N_46969,N_45048,N_45839);
nand U46970 (N_46970,N_45584,N_45865);
nor U46971 (N_46971,N_45736,N_45397);
nor U46972 (N_46972,N_45822,N_45362);
nor U46973 (N_46973,N_45355,N_45623);
or U46974 (N_46974,N_45539,N_45115);
or U46975 (N_46975,N_45503,N_45134);
xnor U46976 (N_46976,N_45066,N_45108);
or U46977 (N_46977,N_45807,N_45394);
xor U46978 (N_46978,N_45466,N_45241);
xor U46979 (N_46979,N_45972,N_45059);
nand U46980 (N_46980,N_45836,N_45016);
nand U46981 (N_46981,N_45288,N_45158);
or U46982 (N_46982,N_45599,N_45100);
nand U46983 (N_46983,N_45029,N_45336);
xnor U46984 (N_46984,N_45142,N_45520);
xnor U46985 (N_46985,N_45886,N_45233);
nand U46986 (N_46986,N_45858,N_45476);
nand U46987 (N_46987,N_45007,N_45162);
xor U46988 (N_46988,N_45618,N_45690);
nor U46989 (N_46989,N_45130,N_45905);
and U46990 (N_46990,N_45118,N_45914);
xor U46991 (N_46991,N_45965,N_45908);
nor U46992 (N_46992,N_45434,N_45093);
or U46993 (N_46993,N_45708,N_45208);
xor U46994 (N_46994,N_45363,N_45856);
and U46995 (N_46995,N_45382,N_45336);
xor U46996 (N_46996,N_45277,N_45168);
nand U46997 (N_46997,N_45794,N_45209);
nand U46998 (N_46998,N_45505,N_45461);
and U46999 (N_46999,N_45494,N_45371);
and U47000 (N_47000,N_46187,N_46208);
nand U47001 (N_47001,N_46936,N_46879);
nor U47002 (N_47002,N_46142,N_46821);
and U47003 (N_47003,N_46211,N_46532);
and U47004 (N_47004,N_46801,N_46100);
and U47005 (N_47005,N_46803,N_46109);
xor U47006 (N_47006,N_46155,N_46322);
and U47007 (N_47007,N_46463,N_46216);
and U47008 (N_47008,N_46627,N_46811);
nand U47009 (N_47009,N_46447,N_46711);
and U47010 (N_47010,N_46841,N_46396);
and U47011 (N_47011,N_46733,N_46658);
or U47012 (N_47012,N_46047,N_46415);
xor U47013 (N_47013,N_46413,N_46931);
and U47014 (N_47014,N_46700,N_46004);
or U47015 (N_47015,N_46701,N_46160);
nor U47016 (N_47016,N_46420,N_46778);
nand U47017 (N_47017,N_46351,N_46485);
xor U47018 (N_47018,N_46566,N_46753);
nand U47019 (N_47019,N_46853,N_46584);
nand U47020 (N_47020,N_46228,N_46596);
nand U47021 (N_47021,N_46417,N_46305);
xnor U47022 (N_47022,N_46430,N_46473);
and U47023 (N_47023,N_46054,N_46297);
and U47024 (N_47024,N_46095,N_46336);
and U47025 (N_47025,N_46661,N_46193);
and U47026 (N_47026,N_46314,N_46085);
or U47027 (N_47027,N_46338,N_46058);
nor U47028 (N_47028,N_46144,N_46895);
or U47029 (N_47029,N_46547,N_46401);
or U47030 (N_47030,N_46343,N_46275);
nor U47031 (N_47031,N_46785,N_46874);
nand U47032 (N_47032,N_46847,N_46183);
or U47033 (N_47033,N_46069,N_46747);
nor U47034 (N_47034,N_46556,N_46300);
nand U47035 (N_47035,N_46398,N_46744);
and U47036 (N_47036,N_46117,N_46453);
or U47037 (N_47037,N_46159,N_46974);
and U47038 (N_47038,N_46407,N_46018);
or U47039 (N_47039,N_46509,N_46716);
and U47040 (N_47040,N_46064,N_46775);
or U47041 (N_47041,N_46885,N_46713);
or U47042 (N_47042,N_46845,N_46145);
xor U47043 (N_47043,N_46198,N_46205);
nor U47044 (N_47044,N_46819,N_46151);
or U47045 (N_47045,N_46026,N_46599);
nor U47046 (N_47046,N_46023,N_46199);
xor U47047 (N_47047,N_46689,N_46461);
and U47048 (N_47048,N_46783,N_46993);
or U47049 (N_47049,N_46278,N_46587);
xor U47050 (N_47050,N_46104,N_46626);
nand U47051 (N_47051,N_46540,N_46549);
xnor U47052 (N_47052,N_46357,N_46638);
nand U47053 (N_47053,N_46210,N_46215);
and U47054 (N_47054,N_46075,N_46073);
nor U47055 (N_47055,N_46586,N_46515);
xnor U47056 (N_47056,N_46412,N_46537);
nand U47057 (N_47057,N_46260,N_46467);
and U47058 (N_47058,N_46489,N_46907);
or U47059 (N_47059,N_46954,N_46953);
nor U47060 (N_47060,N_46376,N_46423);
nor U47061 (N_47061,N_46720,N_46524);
or U47062 (N_47062,N_46288,N_46935);
or U47063 (N_47063,N_46868,N_46831);
nand U47064 (N_47064,N_46702,N_46866);
xnor U47065 (N_47065,N_46299,N_46225);
or U47066 (N_47066,N_46328,N_46286);
and U47067 (N_47067,N_46308,N_46139);
nand U47068 (N_47068,N_46408,N_46636);
xor U47069 (N_47069,N_46794,N_46083);
xnor U47070 (N_47070,N_46400,N_46873);
xnor U47071 (N_47071,N_46929,N_46967);
or U47072 (N_47072,N_46662,N_46884);
nor U47073 (N_47073,N_46670,N_46922);
nand U47074 (N_47074,N_46091,N_46544);
xor U47075 (N_47075,N_46686,N_46450);
nand U47076 (N_47076,N_46951,N_46072);
xor U47077 (N_47077,N_46536,N_46088);
and U47078 (N_47078,N_46007,N_46836);
nor U47079 (N_47079,N_46846,N_46692);
and U47080 (N_47080,N_46105,N_46699);
or U47081 (N_47081,N_46380,N_46855);
nor U47082 (N_47082,N_46800,N_46226);
and U47083 (N_47083,N_46588,N_46999);
xnor U47084 (N_47084,N_46383,N_46604);
or U47085 (N_47085,N_46416,N_46971);
or U47086 (N_47086,N_46878,N_46835);
xor U47087 (N_47087,N_46981,N_46452);
xor U47088 (N_47088,N_46984,N_46877);
nor U47089 (N_47089,N_46217,N_46833);
nand U47090 (N_47090,N_46046,N_46978);
or U47091 (N_47091,N_46983,N_46220);
nand U47092 (N_47092,N_46826,N_46212);
nand U47093 (N_47093,N_46313,N_46804);
nand U47094 (N_47094,N_46189,N_46221);
and U47095 (N_47095,N_46637,N_46528);
nand U47096 (N_47096,N_46272,N_46163);
nor U47097 (N_47097,N_46441,N_46323);
xor U47098 (N_47098,N_46522,N_46062);
nor U47099 (N_47099,N_46222,N_46332);
or U47100 (N_47100,N_46888,N_46042);
nor U47101 (N_47101,N_46548,N_46668);
and U47102 (N_47102,N_46592,N_46533);
xor U47103 (N_47103,N_46397,N_46937);
nor U47104 (N_47104,N_46737,N_46976);
and U47105 (N_47105,N_46863,N_46550);
nand U47106 (N_47106,N_46429,N_46606);
or U47107 (N_47107,N_46782,N_46455);
nand U47108 (N_47108,N_46965,N_46399);
or U47109 (N_47109,N_46697,N_46353);
nor U47110 (N_47110,N_46994,N_46280);
nand U47111 (N_47111,N_46200,N_46623);
nor U47112 (N_47112,N_46457,N_46178);
nand U47113 (N_47113,N_46108,N_46372);
xnor U47114 (N_47114,N_46789,N_46403);
and U47115 (N_47115,N_46518,N_46858);
and U47116 (N_47116,N_46945,N_46573);
or U47117 (N_47117,N_46112,N_46133);
xnor U47118 (N_47118,N_46092,N_46292);
and U47119 (N_47119,N_46291,N_46391);
and U47120 (N_47120,N_46389,N_46992);
or U47121 (N_47121,N_46458,N_46394);
nand U47122 (N_47122,N_46454,N_46277);
nand U47123 (N_47123,N_46614,N_46545);
nand U47124 (N_47124,N_46152,N_46107);
nor U47125 (N_47125,N_46237,N_46977);
or U47126 (N_47126,N_46456,N_46605);
or U47127 (N_47127,N_46156,N_46119);
and U47128 (N_47128,N_46704,N_46608);
nor U47129 (N_47129,N_46060,N_46952);
xnor U47130 (N_47130,N_46049,N_46194);
nor U47131 (N_47131,N_46908,N_46056);
nor U47132 (N_47132,N_46932,N_46395);
and U47133 (N_47133,N_46612,N_46552);
or U47134 (N_47134,N_46530,N_46666);
nand U47135 (N_47135,N_46121,N_46576);
nand U47136 (N_47136,N_46158,N_46138);
nand U47137 (N_47137,N_46184,N_46762);
nor U47138 (N_47138,N_46807,N_46961);
or U47139 (N_47139,N_46191,N_46683);
and U47140 (N_47140,N_46140,N_46887);
nand U47141 (N_47141,N_46779,N_46345);
or U47142 (N_47142,N_46563,N_46955);
nor U47143 (N_47143,N_46262,N_46926);
nand U47144 (N_47144,N_46525,N_46171);
xnor U47145 (N_47145,N_46862,N_46476);
or U47146 (N_47146,N_46712,N_46206);
and U47147 (N_47147,N_46244,N_46053);
or U47148 (N_47148,N_46165,N_46195);
or U47149 (N_47149,N_46368,N_46837);
or U47150 (N_47150,N_46769,N_46529);
nor U47151 (N_47151,N_46316,N_46864);
xnor U47152 (N_47152,N_46891,N_46341);
nor U47153 (N_47153,N_46102,N_46963);
nor U47154 (N_47154,N_46734,N_46125);
xor U47155 (N_47155,N_46721,N_46784);
or U47156 (N_47156,N_46861,N_46203);
and U47157 (N_47157,N_46498,N_46089);
nor U47158 (N_47158,N_46763,N_46619);
nor U47159 (N_47159,N_46911,N_46068);
or U47160 (N_47160,N_46507,N_46361);
nor U47161 (N_47161,N_46392,N_46465);
nand U47162 (N_47162,N_46362,N_46363);
xnor U47163 (N_47163,N_46204,N_46045);
nand U47164 (N_47164,N_46402,N_46066);
and U47165 (N_47165,N_46113,N_46366);
or U47166 (N_47166,N_46464,N_46688);
nand U47167 (N_47167,N_46828,N_46207);
nor U47168 (N_47168,N_46037,N_46186);
and U47169 (N_47169,N_46756,N_46387);
and U47170 (N_47170,N_46730,N_46311);
or U47171 (N_47171,N_46948,N_46590);
nand U47172 (N_47172,N_46657,N_46348);
nand U47173 (N_47173,N_46365,N_46038);
xnor U47174 (N_47174,N_46960,N_46093);
nor U47175 (N_47175,N_46153,N_46805);
nor U47176 (N_47176,N_46143,N_46468);
nor U47177 (N_47177,N_46051,N_46788);
nand U47178 (N_47178,N_46924,N_46164);
or U47179 (N_47179,N_46687,N_46249);
and U47180 (N_47180,N_46520,N_46806);
and U47181 (N_47181,N_46616,N_46504);
nand U47182 (N_47182,N_46912,N_46750);
nand U47183 (N_47183,N_46000,N_46296);
nor U47184 (N_47184,N_46337,N_46664);
and U47185 (N_47185,N_46268,N_46957);
nor U47186 (N_47186,N_46118,N_46621);
and U47187 (N_47187,N_46474,N_46684);
nand U47188 (N_47188,N_46531,N_46170);
nor U47189 (N_47189,N_46149,N_46674);
nand U47190 (N_47190,N_46869,N_46276);
xor U47191 (N_47191,N_46620,N_46982);
or U47192 (N_47192,N_46157,N_46640);
nor U47193 (N_47193,N_46479,N_46022);
nor U47194 (N_47194,N_46809,N_46724);
xnor U47195 (N_47195,N_46825,N_46695);
or U47196 (N_47196,N_46369,N_46190);
xor U47197 (N_47197,N_46493,N_46393);
xor U47198 (N_47198,N_46490,N_46168);
and U47199 (N_47199,N_46964,N_46405);
nor U47200 (N_47200,N_46135,N_46972);
nand U47201 (N_47201,N_46780,N_46443);
nor U47202 (N_47202,N_46943,N_46317);
xor U47203 (N_47203,N_46077,N_46834);
nand U47204 (N_47204,N_46609,N_46710);
nor U47205 (N_47205,N_46767,N_46654);
xnor U47206 (N_47206,N_46196,N_46364);
and U47207 (N_47207,N_46078,N_46039);
or U47208 (N_47208,N_46335,N_46015);
nor U47209 (N_47209,N_46557,N_46676);
nand U47210 (N_47210,N_46239,N_46421);
xor U47211 (N_47211,N_46057,N_46347);
xor U47212 (N_47212,N_46141,N_46264);
nand U47213 (N_47213,N_46944,N_46632);
or U47214 (N_47214,N_46927,N_46648);
or U47215 (N_47215,N_46790,N_46824);
nand U47216 (N_47216,N_46633,N_46578);
nand U47217 (N_47217,N_46367,N_46500);
nor U47218 (N_47218,N_46437,N_46802);
and U47219 (N_47219,N_46041,N_46079);
or U47220 (N_47220,N_46517,N_46466);
or U47221 (N_47221,N_46377,N_46772);
or U47222 (N_47222,N_46628,N_46975);
nand U47223 (N_47223,N_46917,N_46523);
xor U47224 (N_47224,N_46254,N_46630);
and U47225 (N_47225,N_46899,N_46958);
and U47226 (N_47226,N_46319,N_46705);
or U47227 (N_47227,N_46333,N_46012);
or U47228 (N_47228,N_46745,N_46581);
nor U47229 (N_47229,N_46428,N_46554);
nor U47230 (N_47230,N_46379,N_46867);
nand U47231 (N_47231,N_46792,N_46969);
nor U47232 (N_47232,N_46055,N_46898);
xor U47233 (N_47233,N_46514,N_46411);
and U47234 (N_47234,N_46404,N_46318);
nand U47235 (N_47235,N_46791,N_46127);
and U47236 (N_47236,N_46787,N_46257);
nor U47237 (N_47237,N_46099,N_46980);
and U47238 (N_47238,N_46950,N_46938);
xor U47239 (N_47239,N_46502,N_46355);
nor U47240 (N_47240,N_46034,N_46798);
xnor U47241 (N_47241,N_46488,N_46496);
and U47242 (N_47242,N_46080,N_46014);
xnor U47243 (N_47243,N_46499,N_46103);
or U47244 (N_47244,N_46624,N_46373);
nand U47245 (N_47245,N_46607,N_46562);
nand U47246 (N_47246,N_46303,N_46766);
nor U47247 (N_47247,N_46986,N_46253);
or U47248 (N_47248,N_46694,N_46346);
nor U47249 (N_47249,N_46832,N_46857);
or U47250 (N_47250,N_46973,N_46265);
nor U47251 (N_47251,N_46551,N_46358);
and U47252 (N_47252,N_46354,N_46860);
and U47253 (N_47253,N_46718,N_46988);
and U47254 (N_47254,N_46081,N_46647);
nor U47255 (N_47255,N_46914,N_46959);
nor U47256 (N_47256,N_46469,N_46659);
xor U47257 (N_47257,N_46167,N_46755);
nor U47258 (N_47258,N_46675,N_46166);
nor U47259 (N_47259,N_46344,N_46048);
nand U47260 (N_47260,N_46815,N_46896);
and U47261 (N_47261,N_46242,N_46998);
xnor U47262 (N_47262,N_46732,N_46933);
nor U47263 (N_47263,N_46555,N_46942);
nor U47264 (N_47264,N_46434,N_46735);
xor U47265 (N_47265,N_46374,N_46263);
nand U47266 (N_47266,N_46796,N_46880);
nand U47267 (N_47267,N_46459,N_46010);
or U47268 (N_47268,N_46610,N_46760);
nand U47269 (N_47269,N_46445,N_46375);
or U47270 (N_47270,N_46258,N_46480);
or U47271 (N_47271,N_46024,N_46897);
and U47272 (N_47272,N_46370,N_46229);
or U47273 (N_47273,N_46512,N_46040);
nor U47274 (N_47274,N_46234,N_46082);
nand U47275 (N_47275,N_46043,N_46582);
nand U47276 (N_47276,N_46731,N_46008);
nand U47277 (N_47277,N_46030,N_46589);
nand U47278 (N_47278,N_46134,N_46503);
or U47279 (N_47279,N_46970,N_46539);
xor U47280 (N_47280,N_46290,N_46989);
or U47281 (N_47281,N_46817,N_46174);
xor U47282 (N_47282,N_46180,N_46295);
nor U47283 (N_47283,N_46685,N_46385);
nor U47284 (N_47284,N_46651,N_46101);
and U47285 (N_47285,N_46340,N_46691);
nor U47286 (N_47286,N_46224,N_46070);
nand U47287 (N_47287,N_46865,N_46881);
or U47288 (N_47288,N_46765,N_46111);
xor U47289 (N_47289,N_46903,N_46820);
nor U47290 (N_47290,N_46513,N_46146);
nor U47291 (N_47291,N_46947,N_46137);
or U47292 (N_47292,N_46016,N_46324);
nor U47293 (N_47293,N_46919,N_46209);
nor U47294 (N_47294,N_46629,N_46067);
nand U47295 (N_47295,N_46904,N_46197);
xor U47296 (N_47296,N_46122,N_46505);
nand U47297 (N_47297,N_46682,N_46235);
nand U47298 (N_47298,N_46739,N_46631);
nor U47299 (N_47299,N_46245,N_46279);
and U47300 (N_47300,N_46856,N_46331);
nand U47301 (N_47301,N_46613,N_46427);
and U47302 (N_47302,N_46667,N_46492);
or U47303 (N_47303,N_46808,N_46444);
nand U47304 (N_47304,N_46130,N_46096);
nor U47305 (N_47305,N_46600,N_46294);
nand U47306 (N_47306,N_46131,N_46388);
or U47307 (N_47307,N_46129,N_46086);
xor U47308 (N_47308,N_46432,N_46915);
nand U47309 (N_47309,N_46598,N_46169);
nor U47310 (N_47310,N_46901,N_46939);
or U47311 (N_47311,N_46390,N_46192);
or U47312 (N_47312,N_46843,N_46565);
nor U47313 (N_47313,N_46923,N_46872);
and U47314 (N_47314,N_46987,N_46617);
nor U47315 (N_47315,N_46985,N_46406);
or U47316 (N_47316,N_46035,N_46890);
nor U47317 (N_47317,N_46672,N_46663);
or U47318 (N_47318,N_46946,N_46188);
and U47319 (N_47319,N_46273,N_46074);
nor U47320 (N_47320,N_46227,N_46644);
xor U47321 (N_47321,N_46535,N_46414);
or U47322 (N_47322,N_46997,N_46673);
and U47323 (N_47323,N_46776,N_46475);
or U47324 (N_47324,N_46564,N_46128);
and U47325 (N_47325,N_46321,N_46440);
xnor U47326 (N_47326,N_46851,N_46425);
or U47327 (N_47327,N_46813,N_46601);
or U47328 (N_47328,N_46840,N_46709);
nor U47329 (N_47329,N_46774,N_46910);
or U47330 (N_47330,N_46282,N_46717);
and U47331 (N_47331,N_46849,N_46893);
or U47332 (N_47332,N_46021,N_46930);
nor U47333 (N_47333,N_46449,N_46693);
nand U47334 (N_47334,N_46271,N_46219);
xor U47335 (N_47335,N_46526,N_46818);
and U47336 (N_47336,N_46838,N_46956);
nor U47337 (N_47337,N_46098,N_46017);
xor U47338 (N_47338,N_46516,N_46583);
nor U47339 (N_47339,N_46916,N_46669);
xnor U47340 (N_47340,N_46448,N_46678);
or U47341 (N_47341,N_46652,N_46602);
or U47342 (N_47342,N_46446,N_46266);
or U47343 (N_47343,N_46497,N_46593);
nor U47344 (N_47344,N_46003,N_46325);
nor U47345 (N_47345,N_46577,N_46307);
or U47346 (N_47346,N_46009,N_46698);
or U47347 (N_47347,N_46097,N_46251);
or U47348 (N_47348,N_46748,N_46470);
xor U47349 (N_47349,N_46132,N_46793);
nand U47350 (N_47350,N_46597,N_46646);
nor U47351 (N_47351,N_46360,N_46248);
or U47352 (N_47352,N_46768,N_46281);
and U47353 (N_47353,N_46736,N_46059);
and U47354 (N_47354,N_46491,N_46223);
nand U47355 (N_47355,N_46603,N_46542);
and U47356 (N_47356,N_46310,N_46287);
xor U47357 (N_47357,N_46622,N_46315);
nor U47358 (N_47358,N_46019,N_46025);
and U47359 (N_47359,N_46773,N_46810);
nand U47360 (N_47360,N_46011,N_46106);
and U47361 (N_47361,N_46690,N_46680);
and U47362 (N_47362,N_46241,N_46650);
nor U47363 (N_47363,N_46777,N_46634);
nand U47364 (N_47364,N_46063,N_46839);
nand U47365 (N_47365,N_46422,N_46339);
xnor U47366 (N_47366,N_46653,N_46738);
nor U47367 (N_47367,N_46848,N_46486);
xnor U47368 (N_47368,N_46386,N_46495);
or U47369 (N_47369,N_46087,N_46934);
xor U47370 (N_47370,N_46882,N_46641);
nor U47371 (N_47371,N_46746,N_46949);
nor U47372 (N_47372,N_46726,N_46725);
or U47373 (N_47373,N_46625,N_46381);
nor U47374 (N_47374,N_46574,N_46759);
nand U47375 (N_47375,N_46553,N_46797);
and U47376 (N_47376,N_46940,N_46708);
nand U47377 (N_47377,N_46202,N_46213);
or U47378 (N_47378,N_46786,N_46136);
nor U47379 (N_47379,N_46870,N_46615);
and U47380 (N_47380,N_46426,N_46635);
nand U47381 (N_47381,N_46905,N_46179);
nor U47382 (N_47382,N_46920,N_46844);
or U47383 (N_47383,N_46764,N_46006);
and U47384 (N_47384,N_46579,N_46722);
nor U47385 (N_47385,N_46883,N_46852);
xor U47386 (N_47386,N_46816,N_46494);
nor U47387 (N_47387,N_46028,N_46812);
and U47388 (N_47388,N_46771,N_46409);
xor U47389 (N_47389,N_46418,N_46232);
nand U47390 (N_47390,N_46289,N_46770);
nand U47391 (N_47391,N_46410,N_46116);
nor U47392 (N_47392,N_46875,N_46243);
nor U47393 (N_47393,N_46110,N_46740);
and U47394 (N_47394,N_46482,N_46681);
nand U47395 (N_47395,N_46928,N_46594);
and U47396 (N_47396,N_46230,N_46567);
xnor U47397 (N_47397,N_46558,N_46752);
and U47398 (N_47398,N_46591,N_46706);
or U47399 (N_47399,N_46501,N_46352);
xnor U47400 (N_47400,N_46126,N_46350);
or U47401 (N_47401,N_46246,N_46876);
nand U47402 (N_47402,N_46714,N_46534);
or U47403 (N_47403,N_46114,N_46124);
xnor U47404 (N_47404,N_46527,N_46029);
nor U47405 (N_47405,N_46487,N_46172);
xor U47406 (N_47406,N_46013,N_46032);
xor U47407 (N_47407,N_46538,N_46506);
xor U47408 (N_47408,N_46483,N_46642);
nor U47409 (N_47409,N_46656,N_46255);
or U47410 (N_47410,N_46546,N_46481);
nor U47411 (N_47411,N_46306,N_46541);
or U47412 (N_47412,N_46643,N_46442);
or U47413 (N_47413,N_46728,N_46719);
nand U47414 (N_47414,N_46309,N_46471);
nor U47415 (N_47415,N_46918,N_46148);
nand U47416 (N_47416,N_46559,N_46696);
or U47417 (N_47417,N_46349,N_46508);
or U47418 (N_47418,N_46120,N_46327);
and U47419 (N_47419,N_46001,N_46090);
or U47420 (N_47420,N_46052,N_46302);
or U47421 (N_47421,N_46886,N_46267);
nor U47422 (N_47422,N_46611,N_46757);
xor U47423 (N_47423,N_46384,N_46742);
xnor U47424 (N_47424,N_46889,N_46256);
nand U47425 (N_47425,N_46181,N_46749);
and U47426 (N_47426,N_46850,N_46568);
or U47427 (N_47427,N_46799,N_46094);
xor U47428 (N_47428,N_46218,N_46071);
and U47429 (N_47429,N_46065,N_46580);
and U47430 (N_47430,N_46161,N_46795);
xnor U47431 (N_47431,N_46044,N_46182);
nor U47432 (N_47432,N_46002,N_46084);
and U47433 (N_47433,N_46436,N_46312);
nand U47434 (N_47434,N_46284,N_46435);
nor U47435 (N_47435,N_46723,N_46259);
and U47436 (N_47436,N_46572,N_46511);
xor U47437 (N_47437,N_46460,N_46478);
xnor U47438 (N_47438,N_46283,N_46020);
nand U47439 (N_47439,N_46382,N_46031);
nor U47440 (N_47440,N_46741,N_46830);
and U47441 (N_47441,N_46510,N_46829);
nand U47442 (N_47442,N_46906,N_46236);
and U47443 (N_47443,N_46433,N_46177);
xor U47444 (N_47444,N_46703,N_46854);
xor U47445 (N_47445,N_46269,N_46660);
xnor U47446 (N_47446,N_46569,N_46274);
and U47447 (N_47447,N_46477,N_46781);
or U47448 (N_47448,N_46823,N_46729);
or U47449 (N_47449,N_46677,N_46909);
nor U47450 (N_47450,N_46595,N_46521);
xnor U47451 (N_47451,N_46050,N_46585);
nand U47452 (N_47452,N_46990,N_46727);
or U47453 (N_47453,N_46005,N_46329);
or U47454 (N_47454,N_46439,N_46560);
nor U47455 (N_47455,N_46293,N_46270);
xnor U47456 (N_47456,N_46162,N_46150);
nand U47457 (N_47457,N_46033,N_46438);
xor U47458 (N_47458,N_46173,N_46995);
or U47459 (N_47459,N_46231,N_46247);
and U47460 (N_47460,N_46892,N_46966);
or U47461 (N_47461,N_46941,N_46962);
and U47462 (N_47462,N_46175,N_46147);
nor U47463 (N_47463,N_46707,N_46240);
nand U47464 (N_47464,N_46827,N_46214);
xor U47465 (N_47465,N_46649,N_46671);
nor U47466 (N_47466,N_46996,N_46484);
and U47467 (N_47467,N_46356,N_46076);
or U47468 (N_47468,N_46334,N_46570);
nand U47469 (N_47469,N_46571,N_46061);
xnor U47470 (N_47470,N_46027,N_46645);
nand U47471 (N_47471,N_46419,N_46871);
nand U47472 (N_47472,N_46575,N_46304);
xor U47473 (N_47473,N_46359,N_46201);
or U47474 (N_47474,N_46639,N_46115);
xor U47475 (N_47475,N_46320,N_46814);
nor U47476 (N_47476,N_46462,N_46761);
nand U47477 (N_47477,N_46679,N_46472);
and U47478 (N_47478,N_46859,N_46715);
and U47479 (N_47479,N_46894,N_46751);
xnor U47480 (N_47480,N_46238,N_46233);
nor U47481 (N_47481,N_46123,N_46330);
xor U47482 (N_47482,N_46261,N_46991);
or U47483 (N_47483,N_46378,N_46301);
nor U47484 (N_47484,N_46655,N_46176);
nor U47485 (N_47485,N_46036,N_46342);
or U47486 (N_47486,N_46743,N_46902);
nand U47487 (N_47487,N_46154,N_46758);
nor U47488 (N_47488,N_46822,N_46968);
or U47489 (N_47489,N_46519,N_46451);
nor U47490 (N_47490,N_46185,N_46665);
nor U47491 (N_47491,N_46298,N_46913);
nand U47492 (N_47492,N_46842,N_46424);
nand U47493 (N_47493,N_46285,N_46431);
or U47494 (N_47494,N_46326,N_46561);
nor U47495 (N_47495,N_46754,N_46900);
or U47496 (N_47496,N_46252,N_46925);
xnor U47497 (N_47497,N_46543,N_46921);
or U47498 (N_47498,N_46250,N_46371);
xnor U47499 (N_47499,N_46979,N_46618);
or U47500 (N_47500,N_46070,N_46732);
nor U47501 (N_47501,N_46385,N_46632);
or U47502 (N_47502,N_46823,N_46957);
and U47503 (N_47503,N_46404,N_46525);
or U47504 (N_47504,N_46740,N_46813);
or U47505 (N_47505,N_46807,N_46619);
nand U47506 (N_47506,N_46561,N_46007);
xor U47507 (N_47507,N_46671,N_46064);
and U47508 (N_47508,N_46107,N_46243);
and U47509 (N_47509,N_46450,N_46589);
nor U47510 (N_47510,N_46268,N_46966);
nand U47511 (N_47511,N_46846,N_46546);
nand U47512 (N_47512,N_46742,N_46421);
nor U47513 (N_47513,N_46149,N_46377);
xnor U47514 (N_47514,N_46192,N_46143);
and U47515 (N_47515,N_46457,N_46331);
and U47516 (N_47516,N_46888,N_46083);
nor U47517 (N_47517,N_46060,N_46120);
xor U47518 (N_47518,N_46452,N_46534);
or U47519 (N_47519,N_46210,N_46468);
nor U47520 (N_47520,N_46610,N_46091);
nor U47521 (N_47521,N_46791,N_46819);
nor U47522 (N_47522,N_46501,N_46742);
nand U47523 (N_47523,N_46172,N_46088);
and U47524 (N_47524,N_46694,N_46120);
and U47525 (N_47525,N_46468,N_46765);
xnor U47526 (N_47526,N_46977,N_46474);
xnor U47527 (N_47527,N_46271,N_46774);
nand U47528 (N_47528,N_46726,N_46274);
xnor U47529 (N_47529,N_46394,N_46725);
or U47530 (N_47530,N_46275,N_46287);
xor U47531 (N_47531,N_46209,N_46671);
xor U47532 (N_47532,N_46290,N_46261);
or U47533 (N_47533,N_46494,N_46612);
xor U47534 (N_47534,N_46356,N_46032);
nand U47535 (N_47535,N_46569,N_46809);
nand U47536 (N_47536,N_46314,N_46191);
nor U47537 (N_47537,N_46081,N_46618);
nand U47538 (N_47538,N_46400,N_46709);
or U47539 (N_47539,N_46266,N_46087);
nand U47540 (N_47540,N_46863,N_46667);
and U47541 (N_47541,N_46839,N_46613);
nand U47542 (N_47542,N_46748,N_46150);
nand U47543 (N_47543,N_46381,N_46067);
or U47544 (N_47544,N_46692,N_46425);
and U47545 (N_47545,N_46424,N_46463);
nor U47546 (N_47546,N_46802,N_46596);
xnor U47547 (N_47547,N_46151,N_46941);
xnor U47548 (N_47548,N_46466,N_46275);
nor U47549 (N_47549,N_46736,N_46362);
xor U47550 (N_47550,N_46313,N_46686);
and U47551 (N_47551,N_46026,N_46296);
and U47552 (N_47552,N_46700,N_46629);
or U47553 (N_47553,N_46015,N_46158);
or U47554 (N_47554,N_46790,N_46674);
or U47555 (N_47555,N_46995,N_46659);
nor U47556 (N_47556,N_46626,N_46471);
xor U47557 (N_47557,N_46493,N_46009);
xnor U47558 (N_47558,N_46864,N_46116);
nand U47559 (N_47559,N_46764,N_46203);
nand U47560 (N_47560,N_46079,N_46040);
and U47561 (N_47561,N_46035,N_46775);
nor U47562 (N_47562,N_46253,N_46905);
and U47563 (N_47563,N_46825,N_46122);
or U47564 (N_47564,N_46779,N_46614);
or U47565 (N_47565,N_46741,N_46956);
nand U47566 (N_47566,N_46433,N_46941);
xnor U47567 (N_47567,N_46845,N_46468);
nor U47568 (N_47568,N_46378,N_46643);
xor U47569 (N_47569,N_46211,N_46967);
xnor U47570 (N_47570,N_46312,N_46018);
xor U47571 (N_47571,N_46959,N_46400);
xor U47572 (N_47572,N_46073,N_46365);
nor U47573 (N_47573,N_46764,N_46140);
nor U47574 (N_47574,N_46385,N_46378);
nor U47575 (N_47575,N_46004,N_46956);
nand U47576 (N_47576,N_46958,N_46714);
and U47577 (N_47577,N_46008,N_46713);
nor U47578 (N_47578,N_46212,N_46754);
nand U47579 (N_47579,N_46581,N_46460);
and U47580 (N_47580,N_46363,N_46775);
or U47581 (N_47581,N_46372,N_46973);
nor U47582 (N_47582,N_46098,N_46503);
and U47583 (N_47583,N_46505,N_46313);
or U47584 (N_47584,N_46704,N_46497);
nand U47585 (N_47585,N_46097,N_46824);
nand U47586 (N_47586,N_46106,N_46709);
nor U47587 (N_47587,N_46526,N_46006);
and U47588 (N_47588,N_46606,N_46623);
or U47589 (N_47589,N_46985,N_46088);
xnor U47590 (N_47590,N_46760,N_46453);
or U47591 (N_47591,N_46366,N_46461);
nor U47592 (N_47592,N_46652,N_46024);
xor U47593 (N_47593,N_46804,N_46819);
nor U47594 (N_47594,N_46079,N_46256);
nor U47595 (N_47595,N_46442,N_46137);
or U47596 (N_47596,N_46321,N_46661);
xnor U47597 (N_47597,N_46879,N_46595);
and U47598 (N_47598,N_46506,N_46182);
nand U47599 (N_47599,N_46919,N_46585);
xnor U47600 (N_47600,N_46279,N_46712);
or U47601 (N_47601,N_46454,N_46463);
xnor U47602 (N_47602,N_46602,N_46239);
or U47603 (N_47603,N_46519,N_46862);
or U47604 (N_47604,N_46520,N_46321);
or U47605 (N_47605,N_46379,N_46605);
nand U47606 (N_47606,N_46004,N_46220);
nor U47607 (N_47607,N_46192,N_46365);
and U47608 (N_47608,N_46745,N_46172);
and U47609 (N_47609,N_46676,N_46786);
xor U47610 (N_47610,N_46659,N_46207);
nand U47611 (N_47611,N_46884,N_46745);
nor U47612 (N_47612,N_46251,N_46394);
xor U47613 (N_47613,N_46053,N_46281);
nor U47614 (N_47614,N_46459,N_46235);
or U47615 (N_47615,N_46402,N_46122);
nor U47616 (N_47616,N_46957,N_46604);
or U47617 (N_47617,N_46742,N_46094);
nand U47618 (N_47618,N_46962,N_46102);
or U47619 (N_47619,N_46883,N_46164);
or U47620 (N_47620,N_46688,N_46257);
nor U47621 (N_47621,N_46329,N_46382);
xnor U47622 (N_47622,N_46909,N_46703);
xnor U47623 (N_47623,N_46505,N_46947);
nand U47624 (N_47624,N_46021,N_46680);
xnor U47625 (N_47625,N_46247,N_46782);
nand U47626 (N_47626,N_46551,N_46987);
nand U47627 (N_47627,N_46947,N_46295);
nand U47628 (N_47628,N_46385,N_46459);
xnor U47629 (N_47629,N_46690,N_46594);
nor U47630 (N_47630,N_46303,N_46003);
nand U47631 (N_47631,N_46775,N_46577);
and U47632 (N_47632,N_46996,N_46269);
nand U47633 (N_47633,N_46502,N_46081);
nand U47634 (N_47634,N_46393,N_46939);
or U47635 (N_47635,N_46929,N_46616);
or U47636 (N_47636,N_46464,N_46009);
nand U47637 (N_47637,N_46191,N_46611);
nand U47638 (N_47638,N_46716,N_46960);
nand U47639 (N_47639,N_46564,N_46119);
nand U47640 (N_47640,N_46855,N_46756);
or U47641 (N_47641,N_46794,N_46787);
and U47642 (N_47642,N_46721,N_46853);
xnor U47643 (N_47643,N_46323,N_46610);
or U47644 (N_47644,N_46955,N_46702);
or U47645 (N_47645,N_46849,N_46668);
and U47646 (N_47646,N_46915,N_46336);
nor U47647 (N_47647,N_46736,N_46376);
or U47648 (N_47648,N_46902,N_46825);
nor U47649 (N_47649,N_46395,N_46889);
nor U47650 (N_47650,N_46186,N_46764);
nand U47651 (N_47651,N_46942,N_46106);
nand U47652 (N_47652,N_46048,N_46898);
and U47653 (N_47653,N_46311,N_46946);
or U47654 (N_47654,N_46649,N_46689);
or U47655 (N_47655,N_46818,N_46828);
or U47656 (N_47656,N_46395,N_46453);
and U47657 (N_47657,N_46731,N_46948);
nor U47658 (N_47658,N_46116,N_46317);
nand U47659 (N_47659,N_46357,N_46626);
xor U47660 (N_47660,N_46126,N_46218);
nand U47661 (N_47661,N_46883,N_46866);
nand U47662 (N_47662,N_46717,N_46706);
nor U47663 (N_47663,N_46996,N_46052);
nand U47664 (N_47664,N_46200,N_46096);
nand U47665 (N_47665,N_46892,N_46634);
nor U47666 (N_47666,N_46534,N_46135);
and U47667 (N_47667,N_46711,N_46541);
xnor U47668 (N_47668,N_46659,N_46996);
and U47669 (N_47669,N_46590,N_46424);
or U47670 (N_47670,N_46851,N_46958);
xor U47671 (N_47671,N_46622,N_46317);
or U47672 (N_47672,N_46766,N_46966);
nor U47673 (N_47673,N_46783,N_46652);
nor U47674 (N_47674,N_46706,N_46675);
xor U47675 (N_47675,N_46865,N_46982);
or U47676 (N_47676,N_46959,N_46013);
or U47677 (N_47677,N_46696,N_46050);
or U47678 (N_47678,N_46764,N_46954);
nand U47679 (N_47679,N_46450,N_46534);
nor U47680 (N_47680,N_46283,N_46938);
and U47681 (N_47681,N_46985,N_46524);
xnor U47682 (N_47682,N_46642,N_46609);
and U47683 (N_47683,N_46257,N_46207);
xor U47684 (N_47684,N_46443,N_46510);
xor U47685 (N_47685,N_46850,N_46079);
xnor U47686 (N_47686,N_46920,N_46858);
or U47687 (N_47687,N_46945,N_46880);
xnor U47688 (N_47688,N_46859,N_46763);
nor U47689 (N_47689,N_46000,N_46428);
nor U47690 (N_47690,N_46850,N_46629);
and U47691 (N_47691,N_46519,N_46389);
xor U47692 (N_47692,N_46115,N_46454);
and U47693 (N_47693,N_46887,N_46937);
and U47694 (N_47694,N_46078,N_46415);
or U47695 (N_47695,N_46548,N_46155);
xnor U47696 (N_47696,N_46671,N_46699);
or U47697 (N_47697,N_46936,N_46998);
xor U47698 (N_47698,N_46751,N_46873);
and U47699 (N_47699,N_46557,N_46435);
and U47700 (N_47700,N_46216,N_46915);
nand U47701 (N_47701,N_46978,N_46073);
xnor U47702 (N_47702,N_46253,N_46616);
nor U47703 (N_47703,N_46316,N_46100);
or U47704 (N_47704,N_46266,N_46978);
xnor U47705 (N_47705,N_46876,N_46781);
xor U47706 (N_47706,N_46438,N_46595);
and U47707 (N_47707,N_46355,N_46330);
nand U47708 (N_47708,N_46333,N_46815);
nand U47709 (N_47709,N_46601,N_46296);
nand U47710 (N_47710,N_46931,N_46045);
nor U47711 (N_47711,N_46411,N_46010);
or U47712 (N_47712,N_46658,N_46199);
and U47713 (N_47713,N_46078,N_46904);
nand U47714 (N_47714,N_46823,N_46842);
nor U47715 (N_47715,N_46463,N_46288);
nand U47716 (N_47716,N_46995,N_46143);
nor U47717 (N_47717,N_46870,N_46792);
nand U47718 (N_47718,N_46837,N_46438);
nor U47719 (N_47719,N_46508,N_46950);
nor U47720 (N_47720,N_46355,N_46424);
nand U47721 (N_47721,N_46271,N_46595);
xnor U47722 (N_47722,N_46003,N_46129);
and U47723 (N_47723,N_46762,N_46729);
xnor U47724 (N_47724,N_46436,N_46224);
nand U47725 (N_47725,N_46541,N_46418);
nand U47726 (N_47726,N_46857,N_46063);
xor U47727 (N_47727,N_46800,N_46478);
xnor U47728 (N_47728,N_46119,N_46890);
or U47729 (N_47729,N_46796,N_46390);
nor U47730 (N_47730,N_46014,N_46016);
and U47731 (N_47731,N_46475,N_46701);
nor U47732 (N_47732,N_46603,N_46851);
or U47733 (N_47733,N_46629,N_46581);
nand U47734 (N_47734,N_46116,N_46227);
or U47735 (N_47735,N_46011,N_46238);
nor U47736 (N_47736,N_46816,N_46977);
nor U47737 (N_47737,N_46973,N_46665);
nand U47738 (N_47738,N_46650,N_46231);
or U47739 (N_47739,N_46097,N_46062);
nor U47740 (N_47740,N_46119,N_46843);
and U47741 (N_47741,N_46557,N_46768);
nand U47742 (N_47742,N_46064,N_46492);
nand U47743 (N_47743,N_46017,N_46983);
and U47744 (N_47744,N_46314,N_46662);
xnor U47745 (N_47745,N_46605,N_46022);
or U47746 (N_47746,N_46725,N_46443);
xor U47747 (N_47747,N_46507,N_46503);
or U47748 (N_47748,N_46456,N_46754);
or U47749 (N_47749,N_46487,N_46209);
nand U47750 (N_47750,N_46188,N_46807);
and U47751 (N_47751,N_46968,N_46358);
xnor U47752 (N_47752,N_46377,N_46590);
nor U47753 (N_47753,N_46051,N_46098);
and U47754 (N_47754,N_46370,N_46398);
nor U47755 (N_47755,N_46421,N_46356);
and U47756 (N_47756,N_46099,N_46865);
or U47757 (N_47757,N_46714,N_46618);
xor U47758 (N_47758,N_46803,N_46806);
xor U47759 (N_47759,N_46776,N_46361);
and U47760 (N_47760,N_46525,N_46280);
nor U47761 (N_47761,N_46424,N_46435);
nor U47762 (N_47762,N_46287,N_46143);
and U47763 (N_47763,N_46414,N_46112);
and U47764 (N_47764,N_46107,N_46141);
and U47765 (N_47765,N_46474,N_46533);
nor U47766 (N_47766,N_46285,N_46140);
xor U47767 (N_47767,N_46391,N_46232);
nor U47768 (N_47768,N_46639,N_46010);
or U47769 (N_47769,N_46031,N_46136);
nor U47770 (N_47770,N_46324,N_46110);
nor U47771 (N_47771,N_46323,N_46013);
or U47772 (N_47772,N_46810,N_46216);
xnor U47773 (N_47773,N_46588,N_46994);
nand U47774 (N_47774,N_46573,N_46466);
and U47775 (N_47775,N_46489,N_46810);
nand U47776 (N_47776,N_46898,N_46883);
and U47777 (N_47777,N_46859,N_46277);
and U47778 (N_47778,N_46500,N_46338);
or U47779 (N_47779,N_46729,N_46505);
nand U47780 (N_47780,N_46964,N_46214);
nand U47781 (N_47781,N_46023,N_46007);
and U47782 (N_47782,N_46573,N_46545);
nor U47783 (N_47783,N_46368,N_46883);
or U47784 (N_47784,N_46035,N_46791);
or U47785 (N_47785,N_46645,N_46940);
xor U47786 (N_47786,N_46607,N_46980);
or U47787 (N_47787,N_46826,N_46649);
and U47788 (N_47788,N_46499,N_46799);
and U47789 (N_47789,N_46942,N_46548);
xnor U47790 (N_47790,N_46718,N_46007);
nor U47791 (N_47791,N_46160,N_46222);
xor U47792 (N_47792,N_46366,N_46888);
xor U47793 (N_47793,N_46768,N_46669);
nor U47794 (N_47794,N_46912,N_46367);
nand U47795 (N_47795,N_46086,N_46666);
or U47796 (N_47796,N_46712,N_46343);
xnor U47797 (N_47797,N_46624,N_46062);
or U47798 (N_47798,N_46135,N_46077);
and U47799 (N_47799,N_46257,N_46553);
xnor U47800 (N_47800,N_46223,N_46559);
xor U47801 (N_47801,N_46064,N_46046);
and U47802 (N_47802,N_46852,N_46567);
nand U47803 (N_47803,N_46783,N_46171);
and U47804 (N_47804,N_46132,N_46177);
or U47805 (N_47805,N_46194,N_46593);
and U47806 (N_47806,N_46948,N_46823);
xor U47807 (N_47807,N_46457,N_46292);
nor U47808 (N_47808,N_46886,N_46429);
or U47809 (N_47809,N_46925,N_46895);
and U47810 (N_47810,N_46041,N_46163);
xor U47811 (N_47811,N_46031,N_46809);
nand U47812 (N_47812,N_46866,N_46963);
nand U47813 (N_47813,N_46960,N_46033);
and U47814 (N_47814,N_46463,N_46571);
and U47815 (N_47815,N_46843,N_46709);
nand U47816 (N_47816,N_46745,N_46452);
and U47817 (N_47817,N_46098,N_46497);
xnor U47818 (N_47818,N_46362,N_46319);
and U47819 (N_47819,N_46673,N_46940);
nor U47820 (N_47820,N_46160,N_46850);
or U47821 (N_47821,N_46582,N_46489);
nand U47822 (N_47822,N_46125,N_46603);
nor U47823 (N_47823,N_46488,N_46793);
or U47824 (N_47824,N_46332,N_46790);
and U47825 (N_47825,N_46640,N_46793);
xor U47826 (N_47826,N_46454,N_46774);
nand U47827 (N_47827,N_46412,N_46442);
nor U47828 (N_47828,N_46968,N_46423);
and U47829 (N_47829,N_46745,N_46421);
xnor U47830 (N_47830,N_46578,N_46708);
xor U47831 (N_47831,N_46792,N_46550);
or U47832 (N_47832,N_46921,N_46413);
nor U47833 (N_47833,N_46593,N_46576);
nor U47834 (N_47834,N_46034,N_46094);
nor U47835 (N_47835,N_46798,N_46553);
or U47836 (N_47836,N_46076,N_46644);
or U47837 (N_47837,N_46285,N_46758);
nand U47838 (N_47838,N_46987,N_46591);
nor U47839 (N_47839,N_46017,N_46139);
nor U47840 (N_47840,N_46516,N_46473);
and U47841 (N_47841,N_46489,N_46001);
xor U47842 (N_47842,N_46833,N_46752);
and U47843 (N_47843,N_46122,N_46837);
or U47844 (N_47844,N_46252,N_46751);
and U47845 (N_47845,N_46004,N_46099);
nor U47846 (N_47846,N_46262,N_46575);
xor U47847 (N_47847,N_46044,N_46512);
nor U47848 (N_47848,N_46191,N_46095);
nor U47849 (N_47849,N_46005,N_46278);
nor U47850 (N_47850,N_46614,N_46964);
xor U47851 (N_47851,N_46385,N_46062);
xnor U47852 (N_47852,N_46781,N_46906);
and U47853 (N_47853,N_46405,N_46559);
xor U47854 (N_47854,N_46612,N_46081);
and U47855 (N_47855,N_46659,N_46572);
and U47856 (N_47856,N_46310,N_46352);
xor U47857 (N_47857,N_46968,N_46901);
nand U47858 (N_47858,N_46249,N_46483);
and U47859 (N_47859,N_46851,N_46823);
nor U47860 (N_47860,N_46318,N_46873);
nor U47861 (N_47861,N_46752,N_46614);
or U47862 (N_47862,N_46176,N_46895);
nor U47863 (N_47863,N_46193,N_46688);
xnor U47864 (N_47864,N_46791,N_46829);
and U47865 (N_47865,N_46409,N_46490);
or U47866 (N_47866,N_46256,N_46725);
or U47867 (N_47867,N_46232,N_46022);
or U47868 (N_47868,N_46090,N_46050);
xnor U47869 (N_47869,N_46033,N_46305);
nor U47870 (N_47870,N_46474,N_46416);
or U47871 (N_47871,N_46180,N_46199);
and U47872 (N_47872,N_46990,N_46386);
and U47873 (N_47873,N_46169,N_46529);
and U47874 (N_47874,N_46132,N_46644);
xnor U47875 (N_47875,N_46578,N_46658);
and U47876 (N_47876,N_46399,N_46154);
xor U47877 (N_47877,N_46375,N_46057);
nor U47878 (N_47878,N_46119,N_46644);
xor U47879 (N_47879,N_46430,N_46410);
and U47880 (N_47880,N_46273,N_46331);
or U47881 (N_47881,N_46694,N_46582);
nor U47882 (N_47882,N_46416,N_46229);
or U47883 (N_47883,N_46695,N_46315);
xor U47884 (N_47884,N_46590,N_46704);
nand U47885 (N_47885,N_46826,N_46627);
nor U47886 (N_47886,N_46881,N_46367);
and U47887 (N_47887,N_46549,N_46418);
xnor U47888 (N_47888,N_46953,N_46689);
or U47889 (N_47889,N_46846,N_46076);
nand U47890 (N_47890,N_46004,N_46690);
nor U47891 (N_47891,N_46874,N_46963);
nand U47892 (N_47892,N_46171,N_46296);
and U47893 (N_47893,N_46525,N_46161);
or U47894 (N_47894,N_46604,N_46715);
xnor U47895 (N_47895,N_46954,N_46582);
and U47896 (N_47896,N_46257,N_46458);
and U47897 (N_47897,N_46090,N_46003);
nor U47898 (N_47898,N_46129,N_46333);
nor U47899 (N_47899,N_46493,N_46189);
and U47900 (N_47900,N_46733,N_46942);
xor U47901 (N_47901,N_46267,N_46538);
or U47902 (N_47902,N_46038,N_46796);
nand U47903 (N_47903,N_46392,N_46546);
or U47904 (N_47904,N_46796,N_46502);
nand U47905 (N_47905,N_46428,N_46318);
xnor U47906 (N_47906,N_46681,N_46025);
or U47907 (N_47907,N_46876,N_46394);
or U47908 (N_47908,N_46630,N_46237);
nand U47909 (N_47909,N_46944,N_46107);
nor U47910 (N_47910,N_46281,N_46724);
nor U47911 (N_47911,N_46600,N_46353);
and U47912 (N_47912,N_46595,N_46479);
nor U47913 (N_47913,N_46793,N_46231);
nand U47914 (N_47914,N_46620,N_46230);
and U47915 (N_47915,N_46373,N_46174);
and U47916 (N_47916,N_46421,N_46179);
xor U47917 (N_47917,N_46848,N_46373);
and U47918 (N_47918,N_46682,N_46325);
or U47919 (N_47919,N_46819,N_46729);
nor U47920 (N_47920,N_46759,N_46567);
or U47921 (N_47921,N_46905,N_46444);
or U47922 (N_47922,N_46105,N_46790);
xnor U47923 (N_47923,N_46531,N_46154);
xnor U47924 (N_47924,N_46122,N_46797);
nand U47925 (N_47925,N_46908,N_46317);
nand U47926 (N_47926,N_46350,N_46468);
and U47927 (N_47927,N_46177,N_46116);
or U47928 (N_47928,N_46586,N_46710);
or U47929 (N_47929,N_46883,N_46767);
and U47930 (N_47930,N_46673,N_46434);
nor U47931 (N_47931,N_46728,N_46375);
nor U47932 (N_47932,N_46844,N_46832);
nand U47933 (N_47933,N_46971,N_46672);
and U47934 (N_47934,N_46268,N_46724);
nor U47935 (N_47935,N_46671,N_46564);
or U47936 (N_47936,N_46026,N_46866);
nand U47937 (N_47937,N_46689,N_46009);
or U47938 (N_47938,N_46862,N_46162);
nor U47939 (N_47939,N_46580,N_46756);
xnor U47940 (N_47940,N_46248,N_46286);
or U47941 (N_47941,N_46086,N_46034);
nand U47942 (N_47942,N_46215,N_46714);
and U47943 (N_47943,N_46534,N_46658);
or U47944 (N_47944,N_46990,N_46857);
nor U47945 (N_47945,N_46690,N_46057);
nor U47946 (N_47946,N_46826,N_46390);
and U47947 (N_47947,N_46366,N_46889);
xnor U47948 (N_47948,N_46011,N_46523);
and U47949 (N_47949,N_46383,N_46695);
nand U47950 (N_47950,N_46163,N_46726);
nor U47951 (N_47951,N_46689,N_46228);
nor U47952 (N_47952,N_46036,N_46010);
nor U47953 (N_47953,N_46663,N_46693);
xor U47954 (N_47954,N_46901,N_46540);
nor U47955 (N_47955,N_46729,N_46685);
and U47956 (N_47956,N_46115,N_46450);
or U47957 (N_47957,N_46680,N_46173);
nand U47958 (N_47958,N_46448,N_46153);
and U47959 (N_47959,N_46494,N_46442);
xnor U47960 (N_47960,N_46903,N_46813);
xnor U47961 (N_47961,N_46021,N_46647);
and U47962 (N_47962,N_46354,N_46788);
and U47963 (N_47963,N_46333,N_46192);
nor U47964 (N_47964,N_46987,N_46214);
and U47965 (N_47965,N_46621,N_46952);
xnor U47966 (N_47966,N_46247,N_46585);
xnor U47967 (N_47967,N_46247,N_46429);
xnor U47968 (N_47968,N_46706,N_46598);
nand U47969 (N_47969,N_46307,N_46966);
xor U47970 (N_47970,N_46247,N_46826);
xor U47971 (N_47971,N_46850,N_46169);
nor U47972 (N_47972,N_46522,N_46277);
nand U47973 (N_47973,N_46978,N_46946);
nand U47974 (N_47974,N_46268,N_46581);
and U47975 (N_47975,N_46818,N_46325);
nor U47976 (N_47976,N_46907,N_46626);
or U47977 (N_47977,N_46650,N_46376);
and U47978 (N_47978,N_46463,N_46874);
nor U47979 (N_47979,N_46330,N_46001);
xor U47980 (N_47980,N_46658,N_46257);
or U47981 (N_47981,N_46014,N_46609);
and U47982 (N_47982,N_46246,N_46565);
nand U47983 (N_47983,N_46089,N_46768);
and U47984 (N_47984,N_46116,N_46871);
nor U47985 (N_47985,N_46820,N_46361);
xor U47986 (N_47986,N_46240,N_46829);
or U47987 (N_47987,N_46226,N_46639);
and U47988 (N_47988,N_46393,N_46271);
nand U47989 (N_47989,N_46612,N_46434);
xnor U47990 (N_47990,N_46290,N_46620);
and U47991 (N_47991,N_46905,N_46310);
nand U47992 (N_47992,N_46259,N_46956);
and U47993 (N_47993,N_46673,N_46288);
and U47994 (N_47994,N_46482,N_46303);
or U47995 (N_47995,N_46940,N_46999);
and U47996 (N_47996,N_46291,N_46413);
or U47997 (N_47997,N_46910,N_46870);
nor U47998 (N_47998,N_46629,N_46050);
and U47999 (N_47999,N_46638,N_46325);
or U48000 (N_48000,N_47610,N_47219);
nand U48001 (N_48001,N_47568,N_47869);
and U48002 (N_48002,N_47136,N_47073);
and U48003 (N_48003,N_47200,N_47825);
nand U48004 (N_48004,N_47277,N_47202);
nand U48005 (N_48005,N_47244,N_47261);
nor U48006 (N_48006,N_47583,N_47086);
xnor U48007 (N_48007,N_47749,N_47538);
or U48008 (N_48008,N_47924,N_47569);
or U48009 (N_48009,N_47993,N_47632);
and U48010 (N_48010,N_47486,N_47352);
or U48011 (N_48011,N_47496,N_47917);
nor U48012 (N_48012,N_47243,N_47897);
or U48013 (N_48013,N_47540,N_47753);
xnor U48014 (N_48014,N_47468,N_47638);
xor U48015 (N_48015,N_47589,N_47393);
and U48016 (N_48016,N_47672,N_47595);
nor U48017 (N_48017,N_47420,N_47249);
nand U48018 (N_48018,N_47682,N_47828);
nand U48019 (N_48019,N_47535,N_47091);
nand U48020 (N_48020,N_47108,N_47305);
nor U48021 (N_48021,N_47203,N_47157);
xor U48022 (N_48022,N_47930,N_47520);
and U48023 (N_48023,N_47892,N_47973);
nand U48024 (N_48024,N_47054,N_47752);
nor U48025 (N_48025,N_47623,N_47692);
xor U48026 (N_48026,N_47737,N_47185);
nor U48027 (N_48027,N_47548,N_47374);
or U48028 (N_48028,N_47600,N_47436);
and U48029 (N_48029,N_47193,N_47693);
xnor U48030 (N_48030,N_47636,N_47717);
or U48031 (N_48031,N_47452,N_47571);
xor U48032 (N_48032,N_47195,N_47780);
nand U48033 (N_48033,N_47818,N_47796);
and U48034 (N_48034,N_47552,N_47017);
or U48035 (N_48035,N_47167,N_47088);
nor U48036 (N_48036,N_47918,N_47143);
xor U48037 (N_48037,N_47804,N_47162);
nand U48038 (N_48038,N_47702,N_47123);
and U48039 (N_48039,N_47547,N_47497);
nor U48040 (N_48040,N_47968,N_47529);
nor U48041 (N_48041,N_47264,N_47508);
or U48042 (N_48042,N_47052,N_47239);
or U48043 (N_48043,N_47362,N_47634);
and U48044 (N_48044,N_47401,N_47430);
or U48045 (N_48045,N_47906,N_47232);
nand U48046 (N_48046,N_47210,N_47332);
and U48047 (N_48047,N_47138,N_47706);
nor U48048 (N_48048,N_47487,N_47810);
xnor U48049 (N_48049,N_47093,N_47466);
nor U48050 (N_48050,N_47795,N_47546);
nor U48051 (N_48051,N_47381,N_47281);
and U48052 (N_48052,N_47592,N_47330);
nand U48053 (N_48053,N_47894,N_47373);
nand U48054 (N_48054,N_47423,N_47683);
xnor U48055 (N_48055,N_47863,N_47907);
nand U48056 (N_48056,N_47932,N_47619);
or U48057 (N_48057,N_47778,N_47492);
nand U48058 (N_48058,N_47675,N_47343);
nand U48059 (N_48059,N_47442,N_47990);
or U48060 (N_48060,N_47910,N_47635);
xnor U48061 (N_48061,N_47615,N_47340);
or U48062 (N_48062,N_47586,N_47833);
xnor U48063 (N_48063,N_47758,N_47633);
or U48064 (N_48064,N_47901,N_47186);
nand U48065 (N_48065,N_47426,N_47333);
xor U48066 (N_48066,N_47037,N_47139);
and U48067 (N_48067,N_47156,N_47253);
xor U48068 (N_48068,N_47987,N_47198);
xor U48069 (N_48069,N_47409,N_47325);
or U48070 (N_48070,N_47671,N_47835);
nor U48071 (N_48071,N_47178,N_47904);
and U48072 (N_48072,N_47214,N_47027);
or U48073 (N_48073,N_47188,N_47970);
xnor U48074 (N_48074,N_47781,N_47356);
or U48075 (N_48075,N_47351,N_47687);
or U48076 (N_48076,N_47981,N_47129);
xnor U48077 (N_48077,N_47019,N_47344);
nor U48078 (N_48078,N_47455,N_47992);
and U48079 (N_48079,N_47991,N_47609);
nand U48080 (N_48080,N_47493,N_47388);
or U48081 (N_48081,N_47861,N_47296);
nor U48082 (N_48082,N_47120,N_47695);
and U48083 (N_48083,N_47740,N_47895);
xor U48084 (N_48084,N_47310,N_47912);
and U48085 (N_48085,N_47231,N_47848);
or U48086 (N_48086,N_47130,N_47885);
xnor U48087 (N_48087,N_47680,N_47590);
nand U48088 (N_48088,N_47501,N_47889);
and U48089 (N_48089,N_47255,N_47179);
or U48090 (N_48090,N_47223,N_47342);
nand U48091 (N_48091,N_47950,N_47553);
nand U48092 (N_48092,N_47629,N_47103);
or U48093 (N_48093,N_47639,N_47582);
nor U48094 (N_48094,N_47371,N_47471);
or U48095 (N_48095,N_47331,N_47982);
nor U48096 (N_48096,N_47016,N_47560);
or U48097 (N_48097,N_47036,N_47840);
or U48098 (N_48098,N_47997,N_47826);
nand U48099 (N_48099,N_47247,N_47656);
nand U48100 (N_48100,N_47542,N_47563);
nor U48101 (N_48101,N_47106,N_47837);
or U48102 (N_48102,N_47743,N_47564);
xnor U48103 (N_48103,N_47598,N_47943);
nand U48104 (N_48104,N_47725,N_47699);
or U48105 (N_48105,N_47944,N_47849);
nand U48106 (N_48106,N_47134,N_47380);
or U48107 (N_48107,N_47655,N_47700);
nor U48108 (N_48108,N_47248,N_47797);
nor U48109 (N_48109,N_47360,N_47843);
or U48110 (N_48110,N_47511,N_47483);
xor U48111 (N_48111,N_47128,N_47385);
and U48112 (N_48112,N_47858,N_47477);
and U48113 (N_48113,N_47321,N_47659);
xor U48114 (N_48114,N_47710,N_47882);
xor U48115 (N_48115,N_47958,N_47928);
and U48116 (N_48116,N_47116,N_47408);
nor U48117 (N_48117,N_47578,N_47631);
or U48118 (N_48118,N_47080,N_47624);
nand U48119 (N_48119,N_47131,N_47983);
and U48120 (N_48120,N_47888,N_47320);
nand U48121 (N_48121,N_47067,N_47199);
xor U48122 (N_48122,N_47323,N_47505);
xnor U48123 (N_48123,N_47896,N_47579);
nor U48124 (N_48124,N_47570,N_47478);
nor U48125 (N_48125,N_47645,N_47312);
or U48126 (N_48126,N_47031,N_47163);
nor U48127 (N_48127,N_47857,N_47878);
nand U48128 (N_48128,N_47046,N_47847);
xnor U48129 (N_48129,N_47284,N_47921);
nand U48130 (N_48130,N_47757,N_47257);
or U48131 (N_48131,N_47591,N_47033);
nand U48132 (N_48132,N_47694,N_47276);
or U48133 (N_48133,N_47577,N_47761);
or U48134 (N_48134,N_47502,N_47809);
and U48135 (N_48135,N_47141,N_47403);
or U48136 (N_48136,N_47751,N_47491);
nor U48137 (N_48137,N_47147,N_47812);
nand U48138 (N_48138,N_47098,N_47567);
nor U48139 (N_48139,N_47750,N_47020);
nand U48140 (N_48140,N_47875,N_47597);
nand U48141 (N_48141,N_47585,N_47337);
nor U48142 (N_48142,N_47053,N_47267);
xnor U48143 (N_48143,N_47929,N_47291);
or U48144 (N_48144,N_47476,N_47329);
or U48145 (N_48145,N_47024,N_47125);
or U48146 (N_48146,N_47457,N_47306);
and U48147 (N_48147,N_47318,N_47169);
xnor U48148 (N_48148,N_47148,N_47177);
xor U48149 (N_48149,N_47738,N_47599);
nor U48150 (N_48150,N_47470,N_47839);
nor U48151 (N_48151,N_47820,N_47015);
nor U48152 (N_48152,N_47841,N_47448);
nand U48153 (N_48153,N_47786,N_47940);
nand U48154 (N_48154,N_47007,N_47165);
and U48155 (N_48155,N_47049,N_47714);
or U48156 (N_48156,N_47627,N_47949);
nand U48157 (N_48157,N_47899,N_47545);
xnor U48158 (N_48158,N_47925,N_47686);
nand U48159 (N_48159,N_47967,N_47241);
and U48160 (N_48160,N_47137,N_47115);
nor U48161 (N_48161,N_47431,N_47341);
and U48162 (N_48162,N_47022,N_47372);
and U48163 (N_48163,N_47399,N_47217);
or U48164 (N_48164,N_47759,N_47461);
or U48165 (N_48165,N_47962,N_47608);
or U48166 (N_48166,N_47669,N_47530);
or U48167 (N_48167,N_47250,N_47090);
nand U48168 (N_48168,N_47954,N_47268);
nand U48169 (N_48169,N_47065,N_47258);
nor U48170 (N_48170,N_47395,N_47868);
nand U48171 (N_48171,N_47969,N_47621);
or U48172 (N_48172,N_47440,N_47755);
xnor U48173 (N_48173,N_47390,N_47679);
or U48174 (N_48174,N_47112,N_47988);
nor U48175 (N_48175,N_47166,N_47913);
xnor U48176 (N_48176,N_47298,N_47605);
or U48177 (N_48177,N_47415,N_47503);
xnor U48178 (N_48178,N_47941,N_47014);
xor U48179 (N_48179,N_47495,N_47911);
nor U48180 (N_48180,N_47230,N_47300);
and U48181 (N_48181,N_47664,N_47557);
or U48182 (N_48182,N_47023,N_47043);
and U48183 (N_48183,N_47445,N_47561);
nor U48184 (N_48184,N_47152,N_47056);
nor U48185 (N_48185,N_47234,N_47428);
and U48186 (N_48186,N_47102,N_47213);
and U48187 (N_48187,N_47489,N_47688);
xnor U48188 (N_48188,N_47512,N_47978);
nand U48189 (N_48189,N_47051,N_47095);
and U48190 (N_48190,N_47174,N_47462);
and U48191 (N_48191,N_47574,N_47382);
nor U48192 (N_48192,N_47637,N_47190);
and U48193 (N_48193,N_47070,N_47101);
xor U48194 (N_48194,N_47003,N_47760);
or U48195 (N_48195,N_47813,N_47201);
and U48196 (N_48196,N_47773,N_47209);
nand U48197 (N_48197,N_47718,N_47047);
or U48198 (N_48198,N_47111,N_47283);
nor U48199 (N_48199,N_47834,N_47221);
and U48200 (N_48200,N_47957,N_47293);
or U48201 (N_48201,N_47425,N_47229);
and U48202 (N_48202,N_47458,N_47235);
nand U48203 (N_48203,N_47935,N_47322);
nor U48204 (N_48204,N_47916,N_47660);
nor U48205 (N_48205,N_47326,N_47554);
xnor U48206 (N_48206,N_47391,N_47886);
or U48207 (N_48207,N_47075,N_47058);
nand U48208 (N_48208,N_47346,N_47711);
or U48209 (N_48209,N_47048,N_47816);
xnor U48210 (N_48210,N_47593,N_47551);
xor U48211 (N_48211,N_47729,N_47062);
and U48212 (N_48212,N_47533,N_47010);
xnor U48213 (N_48213,N_47044,N_47411);
or U48214 (N_48214,N_47526,N_47110);
nand U48215 (N_48215,N_47085,N_47994);
and U48216 (N_48216,N_47197,N_47744);
nand U48217 (N_48217,N_47063,N_47794);
or U48218 (N_48218,N_47069,N_47713);
or U48219 (N_48219,N_47354,N_47450);
nor U48220 (N_48220,N_47865,N_47846);
and U48221 (N_48221,N_47588,N_47626);
nor U48222 (N_48222,N_47731,N_47733);
or U48223 (N_48223,N_47364,N_47734);
or U48224 (N_48224,N_47665,N_47275);
or U48225 (N_48225,N_47406,N_47011);
xnor U48226 (N_48226,N_47777,N_47290);
xor U48227 (N_48227,N_47790,N_47289);
or U48228 (N_48228,N_47338,N_47034);
nand U48229 (N_48229,N_47164,N_47715);
or U48230 (N_48230,N_47870,N_47437);
xnor U48231 (N_48231,N_47353,N_47055);
and U48232 (N_48232,N_47959,N_47802);
nor U48233 (N_48233,N_47674,N_47328);
nor U48234 (N_48234,N_47377,N_47575);
nand U48235 (N_48235,N_47704,N_47871);
nor U48236 (N_48236,N_47923,N_47741);
nand U48237 (N_48237,N_47192,N_47412);
nor U48238 (N_48238,N_47498,N_47182);
or U48239 (N_48239,N_47936,N_47601);
xnor U48240 (N_48240,N_47914,N_47453);
nor U48241 (N_48241,N_47117,N_47228);
nor U48242 (N_48242,N_47596,N_47386);
xor U48243 (N_48243,N_47927,N_47237);
nor U48244 (N_48244,N_47236,N_47287);
nand U48245 (N_48245,N_47720,N_47850);
and U48246 (N_48246,N_47295,N_47971);
xor U48247 (N_48247,N_47685,N_47534);
or U48248 (N_48248,N_47989,N_47335);
nor U48249 (N_48249,N_47006,N_47181);
nor U48250 (N_48250,N_47821,N_47113);
nand U48251 (N_48251,N_47414,N_47159);
xnor U48252 (N_48252,N_47464,N_47506);
nand U48253 (N_48253,N_47819,N_47856);
nor U48254 (N_48254,N_47874,N_47648);
or U48255 (N_48255,N_47025,N_47806);
nor U48256 (N_48256,N_47183,N_47173);
and U48257 (N_48257,N_47404,N_47867);
xor U48258 (N_48258,N_47726,N_47272);
or U48259 (N_48259,N_47807,N_47145);
nand U48260 (N_48260,N_47479,N_47836);
nor U48261 (N_48261,N_47972,N_47303);
nand U48262 (N_48262,N_47771,N_47697);
nand U48263 (N_48263,N_47233,N_47643);
and U48264 (N_48264,N_47050,N_47407);
and U48265 (N_48265,N_47334,N_47422);
nor U48266 (N_48266,N_47500,N_47032);
and U48267 (N_48267,N_47747,N_47038);
or U48268 (N_48268,N_47532,N_47937);
xnor U48269 (N_48269,N_47363,N_47082);
xnor U48270 (N_48270,N_47614,N_47456);
nand U48271 (N_48271,N_47227,N_47948);
or U48272 (N_48272,N_47375,N_47555);
and U48273 (N_48273,N_47424,N_47860);
nand U48274 (N_48274,N_47772,N_47449);
nor U48275 (N_48275,N_47616,N_47663);
and U48276 (N_48276,N_47522,N_47286);
nor U48277 (N_48277,N_47387,N_47876);
xor U48278 (N_48278,N_47525,N_47719);
xnor U48279 (N_48279,N_47122,N_47142);
or U48280 (N_48280,N_47104,N_47297);
nand U48281 (N_48281,N_47081,N_47893);
or U48282 (N_48282,N_47844,N_47218);
nand U48283 (N_48283,N_47961,N_47008);
xnor U48284 (N_48284,N_47770,N_47435);
nand U48285 (N_48285,N_47434,N_47676);
and U48286 (N_48286,N_47060,N_47240);
nand U48287 (N_48287,N_47144,N_47026);
xnor U48288 (N_48288,N_47212,N_47984);
and U48289 (N_48289,N_47698,N_47767);
or U48290 (N_48290,N_47207,N_47028);
xor U48291 (N_48291,N_47262,N_47963);
xnor U48292 (N_48292,N_47775,N_47280);
and U48293 (N_48293,N_47225,N_47955);
nor U48294 (N_48294,N_47985,N_47299);
nor U48295 (N_48295,N_47365,N_47433);
and U48296 (N_48296,N_47580,N_47266);
and U48297 (N_48297,N_47979,N_47446);
xnor U48298 (N_48298,N_47667,N_47204);
nor U48299 (N_48299,N_47915,N_47762);
xor U48300 (N_48300,N_47238,N_47576);
and U48301 (N_48301,N_47400,N_47716);
nand U48302 (N_48302,N_47278,N_47691);
xor U48303 (N_48303,N_47180,N_47150);
nand U48304 (N_48304,N_47739,N_47622);
or U48305 (N_48305,N_47071,N_47319);
nand U48306 (N_48306,N_47891,N_47079);
xnor U48307 (N_48307,N_47603,N_47832);
nand U48308 (N_48308,N_47784,N_47805);
xnor U48309 (N_48309,N_47438,N_47559);
xor U48310 (N_48310,N_47735,N_47304);
xnor U48311 (N_48311,N_47763,N_47900);
nand U48312 (N_48312,N_47402,N_47273);
nor U48313 (N_48313,N_47184,N_47824);
xor U48314 (N_48314,N_47594,N_47154);
nor U48315 (N_48315,N_47644,N_47421);
nand U48316 (N_48316,N_47996,N_47474);
nor U48317 (N_48317,N_47254,N_47662);
and U48318 (N_48318,N_47160,N_47000);
nor U48319 (N_48319,N_47654,N_47158);
nand U48320 (N_48320,N_47830,N_47612);
nor U48321 (N_48321,N_47708,N_47469);
nor U48322 (N_48322,N_47168,N_47852);
xnor U48323 (N_48323,N_47851,N_47723);
nor U48324 (N_48324,N_47339,N_47109);
xor U48325 (N_48325,N_47539,N_47822);
nor U48326 (N_48326,N_47271,N_47001);
xnor U48327 (N_48327,N_47013,N_47368);
and U48328 (N_48328,N_47441,N_47947);
or U48329 (N_48329,N_47705,N_47021);
or U48330 (N_48330,N_47384,N_47730);
xor U48331 (N_48331,N_47389,N_47317);
nand U48332 (N_48332,N_47514,N_47454);
or U48333 (N_48333,N_47220,N_47998);
nand U48334 (N_48334,N_47721,N_47587);
nand U48335 (N_48335,N_47413,N_47211);
nor U48336 (N_48336,N_47114,N_47269);
and U48337 (N_48337,N_47460,N_47712);
nor U48338 (N_48338,N_47661,N_47061);
xor U48339 (N_48339,N_47484,N_47611);
and U48340 (N_48340,N_47367,N_47282);
nor U48341 (N_48341,N_47313,N_47245);
nor U48342 (N_48342,N_47827,N_47172);
and U48343 (N_48343,N_47242,N_47155);
or U48344 (N_48344,N_47581,N_47879);
xnor U48345 (N_48345,N_47709,N_47494);
xor U48346 (N_48346,N_47764,N_47541);
or U48347 (N_48347,N_47938,N_47926);
and U48348 (N_48348,N_47976,N_47419);
xor U48349 (N_48349,N_47531,N_47765);
nand U48350 (N_48350,N_47292,N_47416);
or U48351 (N_48351,N_47964,N_47519);
xnor U48352 (N_48352,N_47149,N_47064);
nor U48353 (N_48353,N_47222,N_47931);
nand U48354 (N_48354,N_47118,N_47724);
or U48355 (N_48355,N_47756,N_47315);
and U48356 (N_48356,N_47902,N_47722);
nand U48357 (N_48357,N_47398,N_47518);
xnor U48358 (N_48358,N_47057,N_47628);
xnor U48359 (N_48359,N_47550,N_47378);
xor U48360 (N_48360,N_47584,N_47690);
nor U48361 (N_48361,N_47041,N_47383);
and U48362 (N_48362,N_47919,N_47279);
or U48363 (N_48363,N_47429,N_47647);
or U48364 (N_48364,N_47042,N_47853);
xor U48365 (N_48365,N_47653,N_47808);
xor U48366 (N_48366,N_47370,N_47396);
xor U48367 (N_48367,N_47405,N_47171);
or U48368 (N_48368,N_47397,N_47087);
or U48369 (N_48369,N_47696,N_47092);
nor U48370 (N_48370,N_47030,N_47175);
xnor U48371 (N_48371,N_47394,N_47153);
xnor U48372 (N_48372,N_47543,N_47838);
nor U48373 (N_48373,N_47132,N_47005);
xor U48374 (N_48374,N_47606,N_47135);
nor U48375 (N_48375,N_47376,N_47074);
nand U48376 (N_48376,N_47681,N_47473);
or U48377 (N_48377,N_47146,N_47189);
and U48378 (N_48378,N_47521,N_47727);
and U48379 (N_48379,N_47814,N_47572);
and U48380 (N_48380,N_47226,N_47977);
xor U48381 (N_48381,N_47004,N_47732);
xnor U48382 (N_48382,N_47309,N_47613);
xnor U48383 (N_48383,N_47078,N_47980);
nor U48384 (N_48384,N_47651,N_47094);
nor U48385 (N_48385,N_47418,N_47782);
xnor U48386 (N_48386,N_47256,N_47191);
and U48387 (N_48387,N_47270,N_47754);
and U48388 (N_48388,N_47842,N_47045);
nor U48389 (N_48389,N_47946,N_47307);
nor U48390 (N_48390,N_47345,N_47068);
or U48391 (N_48391,N_47083,N_47864);
nand U48392 (N_48392,N_47536,N_47507);
nor U48393 (N_48393,N_47668,N_47862);
nand U48394 (N_48394,N_47537,N_47785);
xnor U48395 (N_48395,N_47766,N_47815);
and U48396 (N_48396,N_47800,N_47974);
or U48397 (N_48397,N_47811,N_47866);
or U48398 (N_48398,N_47650,N_47649);
xor U48399 (N_48399,N_47347,N_47658);
nand U48400 (N_48400,N_47607,N_47742);
nor U48401 (N_48401,N_47793,N_47076);
or U48402 (N_48402,N_47707,N_47516);
xnor U48403 (N_48403,N_47194,N_47642);
nor U48404 (N_48404,N_47039,N_47481);
xor U48405 (N_48405,N_47829,N_47205);
and U48406 (N_48406,N_47909,N_47084);
and U48407 (N_48407,N_47922,N_47573);
or U48408 (N_48408,N_47410,N_47187);
and U48409 (N_48409,N_47002,N_47602);
nand U48410 (N_48410,N_47107,N_47736);
or U48411 (N_48411,N_47485,N_47096);
and U48412 (N_48412,N_47965,N_47465);
nand U48413 (N_48413,N_47678,N_47975);
nor U48414 (N_48414,N_47285,N_47504);
and U48415 (N_48415,N_47792,N_47327);
xnor U48416 (N_48416,N_47788,N_47951);
xor U48417 (N_48417,N_47472,N_47939);
or U48418 (N_48418,N_47884,N_47488);
nor U48419 (N_48419,N_47224,N_47369);
xor U48420 (N_48420,N_47350,N_47215);
xnor U48421 (N_48421,N_47314,N_47854);
xor U48422 (N_48422,N_47952,N_47288);
nor U48423 (N_48423,N_47170,N_47934);
nor U48424 (N_48424,N_47728,N_47887);
nand U48425 (N_48425,N_47995,N_47549);
xor U48426 (N_48426,N_47956,N_47881);
and U48427 (N_48427,N_47779,N_47432);
or U48428 (N_48428,N_47510,N_47089);
or U48429 (N_48429,N_47480,N_47641);
nor U48430 (N_48430,N_47515,N_47029);
and U48431 (N_48431,N_47776,N_47873);
nor U48432 (N_48432,N_47294,N_47960);
nor U48433 (N_48433,N_47748,N_47625);
and U48434 (N_48434,N_47012,N_47801);
nand U48435 (N_48435,N_47124,N_47140);
nor U48436 (N_48436,N_47348,N_47308);
or U48437 (N_48437,N_47392,N_47905);
nand U48438 (N_48438,N_47791,N_47746);
nor U48439 (N_48439,N_47877,N_47872);
nor U48440 (N_48440,N_47439,N_47259);
nand U48441 (N_48441,N_47336,N_47427);
nor U48442 (N_48442,N_47798,N_47459);
or U48443 (N_48443,N_47127,N_47880);
nand U48444 (N_48444,N_47783,N_47523);
xor U48445 (N_48445,N_47077,N_47883);
nand U48446 (N_48446,N_47366,N_47524);
or U48447 (N_48447,N_47774,N_47357);
or U48448 (N_48448,N_47684,N_47799);
or U48449 (N_48449,N_47509,N_47196);
nor U48450 (N_48450,N_47040,N_47789);
xor U48451 (N_48451,N_47490,N_47126);
xor U48452 (N_48452,N_47677,N_47652);
nor U48453 (N_48453,N_47562,N_47817);
nand U48454 (N_48454,N_47513,N_47035);
nor U48455 (N_48455,N_47845,N_47358);
or U48456 (N_48456,N_47208,N_47920);
or U48457 (N_48457,N_47604,N_47059);
and U48458 (N_48458,N_47265,N_47666);
and U48459 (N_48459,N_47018,N_47640);
or U48460 (N_48460,N_47066,N_47855);
and U48461 (N_48461,N_47246,N_47119);
or U48462 (N_48462,N_47646,N_47349);
xor U48463 (N_48463,N_47617,N_47703);
nand U48464 (N_48464,N_47673,N_47769);
nor U48465 (N_48465,N_47121,N_47966);
nand U48466 (N_48466,N_47903,N_47986);
and U48467 (N_48467,N_47176,N_47528);
nor U48468 (N_48468,N_47745,N_47463);
nand U48469 (N_48469,N_47565,N_47898);
xnor U48470 (N_48470,N_47527,N_47803);
or U48471 (N_48471,N_47274,N_47072);
xnor U48472 (N_48472,N_47206,N_47657);
and U48473 (N_48473,N_47620,N_47482);
xnor U48474 (N_48474,N_47451,N_47859);
and U48475 (N_48475,N_47324,N_47544);
nand U48476 (N_48476,N_47999,N_47133);
xnor U48477 (N_48477,N_47099,N_47105);
xor U48478 (N_48478,N_47252,N_47701);
xnor U48479 (N_48479,N_47499,N_47689);
and U48480 (N_48480,N_47823,N_47953);
and U48481 (N_48481,N_47942,N_47100);
xor U48482 (N_48482,N_47444,N_47216);
or U48483 (N_48483,N_47443,N_47890);
or U48484 (N_48484,N_47302,N_47359);
nand U48485 (N_48485,N_47566,N_47768);
nand U48486 (N_48486,N_47558,N_47475);
or U48487 (N_48487,N_47361,N_47009);
nor U48488 (N_48488,N_47630,N_47556);
or U48489 (N_48489,N_47161,N_47263);
nor U48490 (N_48490,N_47908,N_47517);
nand U48491 (N_48491,N_47311,N_47379);
or U48492 (N_48492,N_47301,N_47670);
nor U48493 (N_48493,N_47933,N_47467);
or U48494 (N_48494,N_47316,N_47355);
and U48495 (N_48495,N_47260,N_47831);
nor U48496 (N_48496,N_47151,N_47945);
or U48497 (N_48497,N_47787,N_47447);
xnor U48498 (N_48498,N_47251,N_47417);
nand U48499 (N_48499,N_47618,N_47097);
xnor U48500 (N_48500,N_47593,N_47217);
nand U48501 (N_48501,N_47309,N_47870);
nor U48502 (N_48502,N_47998,N_47467);
and U48503 (N_48503,N_47305,N_47971);
xnor U48504 (N_48504,N_47877,N_47805);
or U48505 (N_48505,N_47510,N_47032);
or U48506 (N_48506,N_47860,N_47015);
nand U48507 (N_48507,N_47182,N_47747);
and U48508 (N_48508,N_47544,N_47727);
and U48509 (N_48509,N_47080,N_47948);
or U48510 (N_48510,N_47252,N_47414);
and U48511 (N_48511,N_47219,N_47921);
nor U48512 (N_48512,N_47790,N_47771);
nand U48513 (N_48513,N_47404,N_47633);
and U48514 (N_48514,N_47357,N_47754);
and U48515 (N_48515,N_47233,N_47349);
nor U48516 (N_48516,N_47182,N_47948);
xnor U48517 (N_48517,N_47435,N_47083);
nor U48518 (N_48518,N_47968,N_47560);
nand U48519 (N_48519,N_47334,N_47701);
nand U48520 (N_48520,N_47882,N_47494);
xor U48521 (N_48521,N_47802,N_47088);
and U48522 (N_48522,N_47039,N_47042);
nand U48523 (N_48523,N_47435,N_47499);
nor U48524 (N_48524,N_47993,N_47205);
xnor U48525 (N_48525,N_47538,N_47988);
and U48526 (N_48526,N_47415,N_47232);
or U48527 (N_48527,N_47264,N_47835);
and U48528 (N_48528,N_47690,N_47026);
and U48529 (N_48529,N_47685,N_47460);
nand U48530 (N_48530,N_47349,N_47712);
nand U48531 (N_48531,N_47086,N_47016);
or U48532 (N_48532,N_47902,N_47030);
and U48533 (N_48533,N_47885,N_47785);
and U48534 (N_48534,N_47605,N_47337);
and U48535 (N_48535,N_47231,N_47708);
and U48536 (N_48536,N_47631,N_47222);
or U48537 (N_48537,N_47236,N_47188);
xor U48538 (N_48538,N_47538,N_47585);
xor U48539 (N_48539,N_47639,N_47032);
and U48540 (N_48540,N_47321,N_47763);
or U48541 (N_48541,N_47708,N_47346);
nand U48542 (N_48542,N_47132,N_47271);
and U48543 (N_48543,N_47822,N_47630);
or U48544 (N_48544,N_47047,N_47352);
and U48545 (N_48545,N_47777,N_47619);
and U48546 (N_48546,N_47539,N_47548);
and U48547 (N_48547,N_47821,N_47608);
and U48548 (N_48548,N_47553,N_47588);
and U48549 (N_48549,N_47883,N_47457);
and U48550 (N_48550,N_47091,N_47163);
and U48551 (N_48551,N_47685,N_47594);
xor U48552 (N_48552,N_47276,N_47700);
nor U48553 (N_48553,N_47000,N_47661);
nand U48554 (N_48554,N_47602,N_47817);
or U48555 (N_48555,N_47056,N_47322);
or U48556 (N_48556,N_47150,N_47038);
nor U48557 (N_48557,N_47508,N_47047);
or U48558 (N_48558,N_47012,N_47655);
nor U48559 (N_48559,N_47499,N_47172);
nand U48560 (N_48560,N_47945,N_47249);
xnor U48561 (N_48561,N_47484,N_47739);
xnor U48562 (N_48562,N_47800,N_47746);
xnor U48563 (N_48563,N_47422,N_47800);
nand U48564 (N_48564,N_47758,N_47508);
xnor U48565 (N_48565,N_47228,N_47693);
nand U48566 (N_48566,N_47242,N_47753);
nand U48567 (N_48567,N_47663,N_47539);
and U48568 (N_48568,N_47902,N_47383);
nand U48569 (N_48569,N_47810,N_47578);
or U48570 (N_48570,N_47368,N_47917);
and U48571 (N_48571,N_47456,N_47075);
nand U48572 (N_48572,N_47497,N_47009);
or U48573 (N_48573,N_47752,N_47853);
nand U48574 (N_48574,N_47185,N_47889);
or U48575 (N_48575,N_47768,N_47798);
xor U48576 (N_48576,N_47437,N_47162);
and U48577 (N_48577,N_47074,N_47362);
xnor U48578 (N_48578,N_47275,N_47132);
xor U48579 (N_48579,N_47202,N_47436);
nand U48580 (N_48580,N_47704,N_47754);
nand U48581 (N_48581,N_47212,N_47547);
nand U48582 (N_48582,N_47794,N_47684);
or U48583 (N_48583,N_47946,N_47243);
and U48584 (N_48584,N_47431,N_47619);
nand U48585 (N_48585,N_47364,N_47708);
nor U48586 (N_48586,N_47558,N_47845);
nor U48587 (N_48587,N_47976,N_47288);
and U48588 (N_48588,N_47851,N_47306);
nor U48589 (N_48589,N_47850,N_47893);
nand U48590 (N_48590,N_47399,N_47481);
xnor U48591 (N_48591,N_47218,N_47517);
nor U48592 (N_48592,N_47998,N_47924);
xnor U48593 (N_48593,N_47644,N_47677);
nand U48594 (N_48594,N_47775,N_47010);
xnor U48595 (N_48595,N_47998,N_47562);
nor U48596 (N_48596,N_47809,N_47564);
nor U48597 (N_48597,N_47529,N_47917);
nand U48598 (N_48598,N_47389,N_47522);
nand U48599 (N_48599,N_47238,N_47667);
or U48600 (N_48600,N_47434,N_47019);
or U48601 (N_48601,N_47594,N_47119);
xnor U48602 (N_48602,N_47113,N_47747);
and U48603 (N_48603,N_47616,N_47287);
and U48604 (N_48604,N_47345,N_47240);
nor U48605 (N_48605,N_47178,N_47221);
xor U48606 (N_48606,N_47672,N_47593);
or U48607 (N_48607,N_47189,N_47805);
or U48608 (N_48608,N_47648,N_47572);
xor U48609 (N_48609,N_47336,N_47465);
xnor U48610 (N_48610,N_47213,N_47782);
nand U48611 (N_48611,N_47946,N_47494);
nand U48612 (N_48612,N_47479,N_47832);
nand U48613 (N_48613,N_47751,N_47968);
nor U48614 (N_48614,N_47260,N_47346);
nand U48615 (N_48615,N_47863,N_47613);
nand U48616 (N_48616,N_47640,N_47088);
and U48617 (N_48617,N_47034,N_47718);
or U48618 (N_48618,N_47795,N_47626);
or U48619 (N_48619,N_47367,N_47181);
nor U48620 (N_48620,N_47203,N_47720);
nand U48621 (N_48621,N_47499,N_47356);
nand U48622 (N_48622,N_47016,N_47774);
or U48623 (N_48623,N_47783,N_47850);
and U48624 (N_48624,N_47520,N_47286);
and U48625 (N_48625,N_47960,N_47390);
or U48626 (N_48626,N_47897,N_47661);
nor U48627 (N_48627,N_47123,N_47080);
and U48628 (N_48628,N_47172,N_47123);
and U48629 (N_48629,N_47874,N_47969);
nand U48630 (N_48630,N_47104,N_47025);
or U48631 (N_48631,N_47467,N_47808);
or U48632 (N_48632,N_47338,N_47421);
nand U48633 (N_48633,N_47809,N_47726);
nand U48634 (N_48634,N_47659,N_47879);
or U48635 (N_48635,N_47567,N_47661);
or U48636 (N_48636,N_47689,N_47783);
and U48637 (N_48637,N_47870,N_47050);
and U48638 (N_48638,N_47386,N_47066);
xor U48639 (N_48639,N_47111,N_47607);
or U48640 (N_48640,N_47931,N_47101);
nor U48641 (N_48641,N_47288,N_47881);
nor U48642 (N_48642,N_47937,N_47864);
xnor U48643 (N_48643,N_47039,N_47866);
nor U48644 (N_48644,N_47647,N_47847);
nand U48645 (N_48645,N_47556,N_47564);
xnor U48646 (N_48646,N_47374,N_47963);
and U48647 (N_48647,N_47954,N_47048);
nor U48648 (N_48648,N_47403,N_47188);
xor U48649 (N_48649,N_47134,N_47238);
and U48650 (N_48650,N_47124,N_47930);
nor U48651 (N_48651,N_47455,N_47466);
xnor U48652 (N_48652,N_47499,N_47745);
nor U48653 (N_48653,N_47958,N_47727);
xor U48654 (N_48654,N_47467,N_47041);
or U48655 (N_48655,N_47456,N_47194);
nor U48656 (N_48656,N_47172,N_47956);
nand U48657 (N_48657,N_47607,N_47996);
nand U48658 (N_48658,N_47789,N_47632);
and U48659 (N_48659,N_47739,N_47205);
nand U48660 (N_48660,N_47146,N_47903);
nand U48661 (N_48661,N_47061,N_47336);
nor U48662 (N_48662,N_47784,N_47361);
xnor U48663 (N_48663,N_47370,N_47419);
or U48664 (N_48664,N_47945,N_47881);
nor U48665 (N_48665,N_47405,N_47245);
and U48666 (N_48666,N_47982,N_47094);
and U48667 (N_48667,N_47516,N_47697);
xor U48668 (N_48668,N_47480,N_47091);
or U48669 (N_48669,N_47271,N_47649);
or U48670 (N_48670,N_47558,N_47727);
xor U48671 (N_48671,N_47306,N_47738);
nor U48672 (N_48672,N_47304,N_47734);
nand U48673 (N_48673,N_47755,N_47133);
and U48674 (N_48674,N_47837,N_47756);
and U48675 (N_48675,N_47776,N_47767);
and U48676 (N_48676,N_47325,N_47454);
and U48677 (N_48677,N_47292,N_47250);
nand U48678 (N_48678,N_47006,N_47195);
or U48679 (N_48679,N_47606,N_47685);
or U48680 (N_48680,N_47131,N_47292);
nand U48681 (N_48681,N_47121,N_47139);
or U48682 (N_48682,N_47441,N_47054);
xor U48683 (N_48683,N_47281,N_47647);
or U48684 (N_48684,N_47121,N_47249);
nand U48685 (N_48685,N_47996,N_47948);
nor U48686 (N_48686,N_47600,N_47903);
xnor U48687 (N_48687,N_47585,N_47341);
nor U48688 (N_48688,N_47915,N_47155);
xnor U48689 (N_48689,N_47860,N_47007);
nor U48690 (N_48690,N_47904,N_47790);
or U48691 (N_48691,N_47782,N_47134);
and U48692 (N_48692,N_47311,N_47449);
nand U48693 (N_48693,N_47527,N_47658);
nand U48694 (N_48694,N_47402,N_47411);
or U48695 (N_48695,N_47852,N_47510);
nand U48696 (N_48696,N_47073,N_47077);
and U48697 (N_48697,N_47667,N_47684);
xnor U48698 (N_48698,N_47408,N_47879);
xor U48699 (N_48699,N_47442,N_47720);
xnor U48700 (N_48700,N_47288,N_47146);
nand U48701 (N_48701,N_47827,N_47469);
xor U48702 (N_48702,N_47507,N_47422);
and U48703 (N_48703,N_47944,N_47951);
nor U48704 (N_48704,N_47990,N_47225);
and U48705 (N_48705,N_47301,N_47110);
nor U48706 (N_48706,N_47650,N_47195);
and U48707 (N_48707,N_47876,N_47022);
and U48708 (N_48708,N_47545,N_47384);
nor U48709 (N_48709,N_47853,N_47077);
or U48710 (N_48710,N_47959,N_47108);
or U48711 (N_48711,N_47698,N_47571);
nand U48712 (N_48712,N_47067,N_47670);
xnor U48713 (N_48713,N_47004,N_47586);
nor U48714 (N_48714,N_47309,N_47499);
or U48715 (N_48715,N_47882,N_47040);
and U48716 (N_48716,N_47694,N_47435);
nand U48717 (N_48717,N_47220,N_47654);
nand U48718 (N_48718,N_47638,N_47957);
or U48719 (N_48719,N_47347,N_47083);
nor U48720 (N_48720,N_47732,N_47344);
or U48721 (N_48721,N_47486,N_47697);
and U48722 (N_48722,N_47323,N_47116);
xnor U48723 (N_48723,N_47344,N_47493);
nor U48724 (N_48724,N_47872,N_47403);
and U48725 (N_48725,N_47491,N_47799);
nand U48726 (N_48726,N_47975,N_47023);
xor U48727 (N_48727,N_47773,N_47894);
nand U48728 (N_48728,N_47942,N_47869);
xor U48729 (N_48729,N_47158,N_47251);
nor U48730 (N_48730,N_47196,N_47043);
nor U48731 (N_48731,N_47668,N_47923);
and U48732 (N_48732,N_47825,N_47206);
or U48733 (N_48733,N_47632,N_47752);
and U48734 (N_48734,N_47042,N_47949);
nor U48735 (N_48735,N_47251,N_47157);
nand U48736 (N_48736,N_47096,N_47472);
or U48737 (N_48737,N_47783,N_47759);
and U48738 (N_48738,N_47248,N_47190);
xnor U48739 (N_48739,N_47094,N_47025);
or U48740 (N_48740,N_47705,N_47079);
nor U48741 (N_48741,N_47305,N_47348);
or U48742 (N_48742,N_47026,N_47587);
or U48743 (N_48743,N_47773,N_47914);
xnor U48744 (N_48744,N_47159,N_47617);
and U48745 (N_48745,N_47308,N_47156);
and U48746 (N_48746,N_47345,N_47381);
nand U48747 (N_48747,N_47522,N_47929);
xnor U48748 (N_48748,N_47936,N_47494);
xor U48749 (N_48749,N_47155,N_47490);
or U48750 (N_48750,N_47671,N_47555);
and U48751 (N_48751,N_47742,N_47076);
xnor U48752 (N_48752,N_47009,N_47743);
and U48753 (N_48753,N_47024,N_47673);
or U48754 (N_48754,N_47000,N_47799);
nor U48755 (N_48755,N_47736,N_47256);
xnor U48756 (N_48756,N_47736,N_47368);
nor U48757 (N_48757,N_47910,N_47130);
or U48758 (N_48758,N_47837,N_47164);
and U48759 (N_48759,N_47189,N_47412);
or U48760 (N_48760,N_47797,N_47871);
and U48761 (N_48761,N_47692,N_47943);
and U48762 (N_48762,N_47586,N_47201);
nor U48763 (N_48763,N_47649,N_47837);
or U48764 (N_48764,N_47022,N_47033);
nand U48765 (N_48765,N_47643,N_47326);
xor U48766 (N_48766,N_47784,N_47558);
and U48767 (N_48767,N_47109,N_47272);
nor U48768 (N_48768,N_47364,N_47405);
or U48769 (N_48769,N_47811,N_47455);
and U48770 (N_48770,N_47843,N_47416);
nor U48771 (N_48771,N_47567,N_47020);
and U48772 (N_48772,N_47728,N_47213);
or U48773 (N_48773,N_47283,N_47780);
nand U48774 (N_48774,N_47868,N_47077);
nand U48775 (N_48775,N_47126,N_47936);
and U48776 (N_48776,N_47727,N_47001);
nand U48777 (N_48777,N_47436,N_47649);
or U48778 (N_48778,N_47092,N_47872);
nand U48779 (N_48779,N_47538,N_47033);
xnor U48780 (N_48780,N_47153,N_47281);
xnor U48781 (N_48781,N_47627,N_47970);
and U48782 (N_48782,N_47785,N_47894);
nand U48783 (N_48783,N_47423,N_47111);
nand U48784 (N_48784,N_47089,N_47585);
or U48785 (N_48785,N_47937,N_47463);
or U48786 (N_48786,N_47192,N_47721);
xor U48787 (N_48787,N_47524,N_47165);
and U48788 (N_48788,N_47050,N_47770);
and U48789 (N_48789,N_47955,N_47966);
nor U48790 (N_48790,N_47736,N_47543);
xnor U48791 (N_48791,N_47163,N_47464);
xor U48792 (N_48792,N_47517,N_47366);
and U48793 (N_48793,N_47014,N_47348);
xor U48794 (N_48794,N_47422,N_47637);
and U48795 (N_48795,N_47072,N_47686);
nand U48796 (N_48796,N_47003,N_47969);
xnor U48797 (N_48797,N_47169,N_47552);
or U48798 (N_48798,N_47676,N_47982);
xnor U48799 (N_48799,N_47067,N_47900);
or U48800 (N_48800,N_47003,N_47197);
nor U48801 (N_48801,N_47656,N_47018);
nand U48802 (N_48802,N_47841,N_47875);
xor U48803 (N_48803,N_47064,N_47567);
xnor U48804 (N_48804,N_47868,N_47894);
nor U48805 (N_48805,N_47016,N_47534);
and U48806 (N_48806,N_47368,N_47546);
or U48807 (N_48807,N_47140,N_47752);
and U48808 (N_48808,N_47996,N_47306);
or U48809 (N_48809,N_47509,N_47317);
nor U48810 (N_48810,N_47398,N_47662);
xor U48811 (N_48811,N_47359,N_47260);
and U48812 (N_48812,N_47927,N_47577);
nor U48813 (N_48813,N_47510,N_47750);
nand U48814 (N_48814,N_47095,N_47339);
or U48815 (N_48815,N_47553,N_47027);
and U48816 (N_48816,N_47155,N_47889);
or U48817 (N_48817,N_47445,N_47018);
nor U48818 (N_48818,N_47816,N_47821);
and U48819 (N_48819,N_47445,N_47363);
xor U48820 (N_48820,N_47228,N_47198);
or U48821 (N_48821,N_47798,N_47491);
nor U48822 (N_48822,N_47145,N_47095);
and U48823 (N_48823,N_47926,N_47249);
xor U48824 (N_48824,N_47980,N_47979);
or U48825 (N_48825,N_47553,N_47475);
xor U48826 (N_48826,N_47122,N_47267);
nor U48827 (N_48827,N_47863,N_47869);
or U48828 (N_48828,N_47555,N_47789);
nor U48829 (N_48829,N_47680,N_47838);
and U48830 (N_48830,N_47026,N_47029);
nor U48831 (N_48831,N_47019,N_47608);
xor U48832 (N_48832,N_47407,N_47245);
xnor U48833 (N_48833,N_47779,N_47528);
and U48834 (N_48834,N_47199,N_47394);
or U48835 (N_48835,N_47908,N_47144);
nand U48836 (N_48836,N_47454,N_47301);
and U48837 (N_48837,N_47670,N_47807);
nor U48838 (N_48838,N_47322,N_47848);
nand U48839 (N_48839,N_47587,N_47604);
nand U48840 (N_48840,N_47199,N_47493);
nand U48841 (N_48841,N_47312,N_47253);
or U48842 (N_48842,N_47136,N_47447);
nor U48843 (N_48843,N_47184,N_47532);
or U48844 (N_48844,N_47126,N_47772);
or U48845 (N_48845,N_47599,N_47189);
and U48846 (N_48846,N_47259,N_47441);
or U48847 (N_48847,N_47766,N_47143);
nor U48848 (N_48848,N_47328,N_47485);
and U48849 (N_48849,N_47754,N_47538);
nor U48850 (N_48850,N_47199,N_47530);
and U48851 (N_48851,N_47475,N_47063);
xnor U48852 (N_48852,N_47821,N_47941);
xnor U48853 (N_48853,N_47385,N_47535);
nor U48854 (N_48854,N_47072,N_47906);
nand U48855 (N_48855,N_47063,N_47734);
nor U48856 (N_48856,N_47855,N_47917);
nand U48857 (N_48857,N_47683,N_47809);
and U48858 (N_48858,N_47262,N_47142);
and U48859 (N_48859,N_47575,N_47522);
or U48860 (N_48860,N_47505,N_47592);
nand U48861 (N_48861,N_47362,N_47386);
nand U48862 (N_48862,N_47395,N_47806);
xor U48863 (N_48863,N_47149,N_47086);
xnor U48864 (N_48864,N_47738,N_47845);
xnor U48865 (N_48865,N_47838,N_47748);
xnor U48866 (N_48866,N_47613,N_47096);
and U48867 (N_48867,N_47008,N_47912);
xor U48868 (N_48868,N_47575,N_47631);
nand U48869 (N_48869,N_47512,N_47831);
and U48870 (N_48870,N_47654,N_47243);
and U48871 (N_48871,N_47514,N_47559);
nand U48872 (N_48872,N_47785,N_47185);
and U48873 (N_48873,N_47290,N_47486);
and U48874 (N_48874,N_47305,N_47285);
xor U48875 (N_48875,N_47920,N_47641);
or U48876 (N_48876,N_47310,N_47847);
nand U48877 (N_48877,N_47068,N_47975);
xor U48878 (N_48878,N_47916,N_47778);
xnor U48879 (N_48879,N_47787,N_47812);
nor U48880 (N_48880,N_47519,N_47793);
and U48881 (N_48881,N_47831,N_47284);
nand U48882 (N_48882,N_47952,N_47012);
and U48883 (N_48883,N_47843,N_47780);
xnor U48884 (N_48884,N_47865,N_47025);
nand U48885 (N_48885,N_47032,N_47146);
and U48886 (N_48886,N_47965,N_47273);
and U48887 (N_48887,N_47471,N_47349);
or U48888 (N_48888,N_47074,N_47947);
nor U48889 (N_48889,N_47321,N_47758);
xnor U48890 (N_48890,N_47018,N_47938);
and U48891 (N_48891,N_47449,N_47883);
and U48892 (N_48892,N_47312,N_47846);
nor U48893 (N_48893,N_47020,N_47639);
nor U48894 (N_48894,N_47286,N_47646);
nor U48895 (N_48895,N_47416,N_47817);
xor U48896 (N_48896,N_47087,N_47554);
and U48897 (N_48897,N_47365,N_47279);
or U48898 (N_48898,N_47968,N_47957);
or U48899 (N_48899,N_47153,N_47441);
and U48900 (N_48900,N_47938,N_47302);
nor U48901 (N_48901,N_47557,N_47821);
or U48902 (N_48902,N_47389,N_47346);
nand U48903 (N_48903,N_47508,N_47516);
or U48904 (N_48904,N_47995,N_47174);
xor U48905 (N_48905,N_47911,N_47416);
xnor U48906 (N_48906,N_47749,N_47931);
xnor U48907 (N_48907,N_47751,N_47041);
nand U48908 (N_48908,N_47928,N_47426);
nor U48909 (N_48909,N_47581,N_47360);
and U48910 (N_48910,N_47923,N_47239);
nand U48911 (N_48911,N_47616,N_47926);
nand U48912 (N_48912,N_47041,N_47546);
or U48913 (N_48913,N_47779,N_47247);
xor U48914 (N_48914,N_47646,N_47272);
and U48915 (N_48915,N_47008,N_47790);
nand U48916 (N_48916,N_47133,N_47792);
nor U48917 (N_48917,N_47003,N_47728);
xor U48918 (N_48918,N_47486,N_47359);
nor U48919 (N_48919,N_47228,N_47687);
xnor U48920 (N_48920,N_47754,N_47168);
nor U48921 (N_48921,N_47562,N_47640);
nand U48922 (N_48922,N_47220,N_47646);
and U48923 (N_48923,N_47707,N_47965);
xnor U48924 (N_48924,N_47896,N_47688);
nor U48925 (N_48925,N_47225,N_47454);
and U48926 (N_48926,N_47744,N_47485);
and U48927 (N_48927,N_47070,N_47529);
or U48928 (N_48928,N_47856,N_47224);
xor U48929 (N_48929,N_47878,N_47578);
or U48930 (N_48930,N_47559,N_47104);
and U48931 (N_48931,N_47118,N_47734);
nor U48932 (N_48932,N_47684,N_47470);
xnor U48933 (N_48933,N_47515,N_47948);
nor U48934 (N_48934,N_47885,N_47831);
nor U48935 (N_48935,N_47439,N_47378);
or U48936 (N_48936,N_47902,N_47768);
nand U48937 (N_48937,N_47412,N_47565);
and U48938 (N_48938,N_47984,N_47306);
xnor U48939 (N_48939,N_47299,N_47716);
or U48940 (N_48940,N_47876,N_47880);
and U48941 (N_48941,N_47889,N_47275);
or U48942 (N_48942,N_47961,N_47236);
or U48943 (N_48943,N_47802,N_47415);
nand U48944 (N_48944,N_47588,N_47135);
or U48945 (N_48945,N_47127,N_47934);
nand U48946 (N_48946,N_47852,N_47554);
nand U48947 (N_48947,N_47464,N_47109);
nand U48948 (N_48948,N_47383,N_47382);
or U48949 (N_48949,N_47646,N_47545);
or U48950 (N_48950,N_47407,N_47185);
nand U48951 (N_48951,N_47281,N_47869);
or U48952 (N_48952,N_47578,N_47665);
xor U48953 (N_48953,N_47298,N_47774);
nand U48954 (N_48954,N_47920,N_47127);
or U48955 (N_48955,N_47627,N_47535);
nand U48956 (N_48956,N_47003,N_47311);
xnor U48957 (N_48957,N_47605,N_47892);
nor U48958 (N_48958,N_47226,N_47110);
and U48959 (N_48959,N_47419,N_47197);
xor U48960 (N_48960,N_47534,N_47261);
nor U48961 (N_48961,N_47437,N_47390);
xnor U48962 (N_48962,N_47297,N_47672);
nor U48963 (N_48963,N_47900,N_47324);
nor U48964 (N_48964,N_47799,N_47760);
xnor U48965 (N_48965,N_47512,N_47515);
xor U48966 (N_48966,N_47150,N_47752);
xnor U48967 (N_48967,N_47340,N_47290);
nor U48968 (N_48968,N_47194,N_47684);
xnor U48969 (N_48969,N_47802,N_47869);
xor U48970 (N_48970,N_47151,N_47622);
nor U48971 (N_48971,N_47674,N_47563);
xor U48972 (N_48972,N_47636,N_47395);
nor U48973 (N_48973,N_47666,N_47299);
xnor U48974 (N_48974,N_47398,N_47746);
or U48975 (N_48975,N_47083,N_47876);
xor U48976 (N_48976,N_47890,N_47281);
xnor U48977 (N_48977,N_47674,N_47299);
or U48978 (N_48978,N_47784,N_47131);
nand U48979 (N_48979,N_47567,N_47627);
nor U48980 (N_48980,N_47956,N_47214);
nand U48981 (N_48981,N_47867,N_47749);
xnor U48982 (N_48982,N_47862,N_47242);
nand U48983 (N_48983,N_47611,N_47247);
nand U48984 (N_48984,N_47214,N_47655);
xor U48985 (N_48985,N_47706,N_47755);
nand U48986 (N_48986,N_47538,N_47454);
nor U48987 (N_48987,N_47720,N_47331);
nor U48988 (N_48988,N_47431,N_47340);
or U48989 (N_48989,N_47264,N_47187);
or U48990 (N_48990,N_47000,N_47794);
or U48991 (N_48991,N_47310,N_47889);
nand U48992 (N_48992,N_47530,N_47610);
nand U48993 (N_48993,N_47889,N_47896);
xor U48994 (N_48994,N_47056,N_47300);
and U48995 (N_48995,N_47702,N_47238);
nand U48996 (N_48996,N_47714,N_47890);
nand U48997 (N_48997,N_47103,N_47314);
xnor U48998 (N_48998,N_47536,N_47561);
and U48999 (N_48999,N_47484,N_47780);
nor U49000 (N_49000,N_48614,N_48992);
nor U49001 (N_49001,N_48321,N_48786);
and U49002 (N_49002,N_48456,N_48060);
xor U49003 (N_49003,N_48235,N_48026);
and U49004 (N_49004,N_48656,N_48336);
or U49005 (N_49005,N_48081,N_48800);
nor U49006 (N_49006,N_48188,N_48035);
nor U49007 (N_49007,N_48548,N_48449);
nor U49008 (N_49008,N_48770,N_48885);
and U49009 (N_49009,N_48911,N_48636);
nor U49010 (N_49010,N_48093,N_48458);
or U49011 (N_49011,N_48995,N_48806);
and U49012 (N_49012,N_48605,N_48005);
or U49013 (N_49013,N_48750,N_48086);
nand U49014 (N_49014,N_48138,N_48370);
nand U49015 (N_49015,N_48867,N_48454);
nor U49016 (N_49016,N_48464,N_48246);
xnor U49017 (N_49017,N_48483,N_48008);
nand U49018 (N_49018,N_48597,N_48587);
nand U49019 (N_49019,N_48242,N_48499);
and U49020 (N_49020,N_48355,N_48725);
or U49021 (N_49021,N_48652,N_48999);
and U49022 (N_49022,N_48453,N_48259);
and U49023 (N_49023,N_48072,N_48882);
or U49024 (N_49024,N_48645,N_48788);
xor U49025 (N_49025,N_48304,N_48599);
nand U49026 (N_49026,N_48669,N_48533);
xor U49027 (N_49027,N_48479,N_48367);
nand U49028 (N_49028,N_48576,N_48433);
and U49029 (N_49029,N_48823,N_48975);
or U49030 (N_49030,N_48022,N_48088);
and U49031 (N_49031,N_48435,N_48870);
or U49032 (N_49032,N_48303,N_48831);
or U49033 (N_49033,N_48696,N_48878);
nor U49034 (N_49034,N_48708,N_48327);
and U49035 (N_49035,N_48879,N_48043);
or U49036 (N_49036,N_48232,N_48863);
nor U49037 (N_49037,N_48318,N_48324);
and U49038 (N_49038,N_48263,N_48399);
nor U49039 (N_49039,N_48796,N_48205);
or U49040 (N_49040,N_48736,N_48952);
xnor U49041 (N_49041,N_48991,N_48312);
nand U49042 (N_49042,N_48465,N_48100);
and U49043 (N_49043,N_48906,N_48646);
nor U49044 (N_49044,N_48233,N_48032);
nor U49045 (N_49045,N_48843,N_48401);
and U49046 (N_49046,N_48753,N_48168);
nand U49047 (N_49047,N_48943,N_48210);
nor U49048 (N_49048,N_48441,N_48761);
nand U49049 (N_49049,N_48888,N_48459);
nor U49050 (N_49050,N_48281,N_48398);
and U49051 (N_49051,N_48683,N_48670);
or U49052 (N_49052,N_48294,N_48524);
xor U49053 (N_49053,N_48891,N_48311);
xor U49054 (N_49054,N_48490,N_48865);
nand U49055 (N_49055,N_48536,N_48221);
nor U49056 (N_49056,N_48258,N_48358);
nor U49057 (N_49057,N_48171,N_48353);
xnor U49058 (N_49058,N_48837,N_48586);
and U49059 (N_49059,N_48684,N_48756);
xnor U49060 (N_49060,N_48222,N_48296);
nor U49061 (N_49061,N_48512,N_48182);
or U49062 (N_49062,N_48762,N_48780);
nor U49063 (N_49063,N_48859,N_48640);
and U49064 (N_49064,N_48821,N_48105);
or U49065 (N_49065,N_48930,N_48570);
nand U49066 (N_49066,N_48767,N_48234);
or U49067 (N_49067,N_48572,N_48905);
or U49068 (N_49068,N_48307,N_48286);
or U49069 (N_49069,N_48076,N_48065);
and U49070 (N_49070,N_48320,N_48824);
nand U49071 (N_49071,N_48298,N_48694);
or U49072 (N_49072,N_48771,N_48365);
or U49073 (N_49073,N_48066,N_48342);
xnor U49074 (N_49074,N_48501,N_48302);
nand U49075 (N_49075,N_48054,N_48247);
and U49076 (N_49076,N_48810,N_48002);
nand U49077 (N_49077,N_48630,N_48067);
nor U49078 (N_49078,N_48229,N_48804);
nor U49079 (N_49079,N_48983,N_48580);
and U49080 (N_49080,N_48404,N_48956);
nor U49081 (N_49081,N_48244,N_48153);
nand U49082 (N_49082,N_48047,N_48164);
or U49083 (N_49083,N_48732,N_48634);
nor U49084 (N_49084,N_48175,N_48275);
or U49085 (N_49085,N_48900,N_48903);
nand U49086 (N_49086,N_48299,N_48016);
xor U49087 (N_49087,N_48291,N_48883);
and U49088 (N_49088,N_48469,N_48498);
or U49089 (N_49089,N_48369,N_48792);
or U49090 (N_49090,N_48739,N_48612);
or U49091 (N_49091,N_48775,N_48840);
and U49092 (N_49092,N_48755,N_48161);
xnor U49093 (N_49093,N_48591,N_48363);
xnor U49094 (N_49094,N_48288,N_48011);
nand U49095 (N_49095,N_48797,N_48256);
and U49096 (N_49096,N_48720,N_48149);
nand U49097 (N_49097,N_48808,N_48935);
xor U49098 (N_49098,N_48013,N_48420);
xor U49099 (N_49099,N_48946,N_48389);
or U49100 (N_49100,N_48410,N_48970);
nor U49101 (N_49101,N_48908,N_48923);
nor U49102 (N_49102,N_48575,N_48354);
or U49103 (N_49103,N_48230,N_48451);
xor U49104 (N_49104,N_48960,N_48414);
xor U49105 (N_49105,N_48892,N_48812);
and U49106 (N_49106,N_48754,N_48904);
and U49107 (N_49107,N_48541,N_48637);
and U49108 (N_49108,N_48620,N_48196);
and U49109 (N_49109,N_48283,N_48961);
or U49110 (N_49110,N_48818,N_48078);
or U49111 (N_49111,N_48660,N_48390);
or U49112 (N_49112,N_48200,N_48562);
nand U49113 (N_49113,N_48914,N_48212);
and U49114 (N_49114,N_48145,N_48962);
nand U49115 (N_49115,N_48163,N_48317);
and U49116 (N_49116,N_48589,N_48098);
nor U49117 (N_49117,N_48293,N_48107);
nor U49118 (N_49118,N_48610,N_48740);
nor U49119 (N_49119,N_48554,N_48368);
nand U49120 (N_49120,N_48503,N_48994);
xor U49121 (N_49121,N_48531,N_48866);
nor U49122 (N_49122,N_48735,N_48239);
or U49123 (N_49123,N_48111,N_48176);
and U49124 (N_49124,N_48073,N_48071);
xor U49125 (N_49125,N_48019,N_48186);
nor U49126 (N_49126,N_48722,N_48147);
nand U49127 (N_49127,N_48329,N_48347);
nor U49128 (N_49128,N_48091,N_48516);
nor U49129 (N_49129,N_48919,N_48829);
xnor U49130 (N_49130,N_48384,N_48687);
nor U49131 (N_49131,N_48967,N_48551);
and U49132 (N_49132,N_48190,N_48521);
nand U49133 (N_49133,N_48253,N_48462);
xnor U49134 (N_49134,N_48036,N_48228);
or U49135 (N_49135,N_48189,N_48468);
xor U49136 (N_49136,N_48314,N_48836);
nor U49137 (N_49137,N_48833,N_48596);
or U49138 (N_49138,N_48477,N_48124);
and U49139 (N_49139,N_48731,N_48243);
xnor U49140 (N_49140,N_48933,N_48674);
and U49141 (N_49141,N_48197,N_48592);
nand U49142 (N_49142,N_48033,N_48951);
or U49143 (N_49143,N_48573,N_48350);
nand U49144 (N_49144,N_48495,N_48707);
nor U49145 (N_49145,N_48622,N_48759);
xor U49146 (N_49146,N_48403,N_48858);
or U49147 (N_49147,N_48340,N_48260);
xnor U49148 (N_49148,N_48719,N_48856);
nand U49149 (N_49149,N_48909,N_48565);
or U49150 (N_49150,N_48344,N_48009);
or U49151 (N_49151,N_48306,N_48313);
xor U49152 (N_49152,N_48621,N_48703);
or U49153 (N_49153,N_48953,N_48538);
nor U49154 (N_49154,N_48902,N_48884);
or U49155 (N_49155,N_48828,N_48448);
nand U49156 (N_49156,N_48997,N_48006);
and U49157 (N_49157,N_48623,N_48550);
xnor U49158 (N_49158,N_48931,N_48120);
and U49159 (N_49159,N_48766,N_48848);
or U49160 (N_49160,N_48986,N_48174);
xnor U49161 (N_49161,N_48184,N_48845);
or U49162 (N_49162,N_48126,N_48747);
xnor U49163 (N_49163,N_48038,N_48532);
xnor U49164 (N_49164,N_48134,N_48880);
or U49165 (N_49165,N_48711,N_48505);
or U49166 (N_49166,N_48555,N_48582);
nand U49167 (N_49167,N_48603,N_48106);
nand U49168 (N_49168,N_48852,N_48549);
nand U49169 (N_49169,N_48560,N_48136);
nand U49170 (N_49170,N_48236,N_48042);
nor U49171 (N_49171,N_48334,N_48791);
xor U49172 (N_49172,N_48665,N_48201);
xnor U49173 (N_49173,N_48942,N_48092);
and U49174 (N_49174,N_48130,N_48869);
nand U49175 (N_49175,N_48509,N_48271);
or U49176 (N_49176,N_48095,N_48478);
or U49177 (N_49177,N_48827,N_48346);
nand U49178 (N_49178,N_48380,N_48333);
nand U49179 (N_49179,N_48728,N_48693);
nor U49180 (N_49180,N_48300,N_48557);
and U49181 (N_49181,N_48172,N_48981);
xor U49182 (N_49182,N_48868,N_48938);
nor U49183 (N_49183,N_48309,N_48604);
xnor U49184 (N_49184,N_48180,N_48624);
and U49185 (N_49185,N_48497,N_48724);
and U49186 (N_49186,N_48280,N_48393);
nand U49187 (N_49187,N_48328,N_48613);
or U49188 (N_49188,N_48262,N_48772);
and U49189 (N_49189,N_48543,N_48682);
and U49190 (N_49190,N_48816,N_48673);
nor U49191 (N_49191,N_48199,N_48917);
xor U49192 (N_49192,N_48830,N_48746);
xor U49193 (N_49193,N_48413,N_48422);
xnor U49194 (N_49194,N_48697,N_48437);
or U49195 (N_49195,N_48101,N_48455);
xor U49196 (N_49196,N_48366,N_48698);
and U49197 (N_49197,N_48940,N_48305);
or U49198 (N_49198,N_48431,N_48204);
or U49199 (N_49199,N_48726,N_48547);
or U49200 (N_49200,N_48945,N_48899);
or U49201 (N_49201,N_48208,N_48650);
nand U49202 (N_49202,N_48504,N_48659);
xnor U49203 (N_49203,N_48950,N_48397);
or U49204 (N_49204,N_48491,N_48926);
or U49205 (N_49205,N_48779,N_48826);
or U49206 (N_49206,N_48820,N_48556);
nand U49207 (N_49207,N_48450,N_48948);
nand U49208 (N_49208,N_48096,N_48715);
nor U49209 (N_49209,N_48117,N_48502);
and U49210 (N_49210,N_48987,N_48461);
and U49211 (N_49211,N_48089,N_48338);
and U49212 (N_49212,N_48023,N_48255);
or U49213 (N_49213,N_48721,N_48000);
nor U49214 (N_49214,N_48520,N_48424);
and U49215 (N_49215,N_48638,N_48661);
nand U49216 (N_49216,N_48297,N_48225);
or U49217 (N_49217,N_48781,N_48064);
or U49218 (N_49218,N_48341,N_48679);
and U49219 (N_49219,N_48423,N_48574);
or U49220 (N_49220,N_48738,N_48608);
nor U49221 (N_49221,N_48663,N_48177);
or U49222 (N_49222,N_48457,N_48654);
nand U49223 (N_49223,N_48672,N_48323);
and U49224 (N_49224,N_48484,N_48851);
and U49225 (N_49225,N_48568,N_48626);
nor U49226 (N_49226,N_48331,N_48277);
and U49227 (N_49227,N_48332,N_48052);
nor U49228 (N_49228,N_48114,N_48954);
and U49229 (N_49229,N_48802,N_48156);
xnor U49230 (N_49230,N_48889,N_48787);
nor U49231 (N_49231,N_48021,N_48525);
or U49232 (N_49232,N_48061,N_48944);
nor U49233 (N_49233,N_48896,N_48068);
nand U49234 (N_49234,N_48815,N_48492);
xor U49235 (N_49235,N_48727,N_48170);
or U49236 (N_49236,N_48211,N_48743);
and U49237 (N_49237,N_48741,N_48158);
nand U49238 (N_49238,N_48700,N_48295);
nor U49239 (N_49239,N_48110,N_48920);
xor U49240 (N_49240,N_48062,N_48044);
xor U49241 (N_49241,N_48439,N_48601);
nor U49242 (N_49242,N_48801,N_48213);
xor U49243 (N_49243,N_48097,N_48482);
and U49244 (N_49244,N_48860,N_48475);
and U49245 (N_49245,N_48769,N_48075);
xor U49246 (N_49246,N_48119,N_48958);
or U49247 (N_49247,N_48701,N_48123);
nor U49248 (N_49248,N_48966,N_48515);
xnor U49249 (N_49249,N_48273,N_48730);
nor U49250 (N_49250,N_48357,N_48713);
nor U49251 (N_49251,N_48877,N_48973);
xor U49252 (N_49252,N_48248,N_48361);
nand U49253 (N_49253,N_48705,N_48631);
nand U49254 (N_49254,N_48427,N_48977);
xor U49255 (N_49255,N_48990,N_48471);
xor U49256 (N_49256,N_48018,N_48817);
or U49257 (N_49257,N_48090,N_48402);
nor U49258 (N_49258,N_48157,N_48343);
xor U49259 (N_49259,N_48546,N_48267);
and U49260 (N_49260,N_48734,N_48718);
xor U49261 (N_49261,N_48014,N_48162);
nor U49262 (N_49262,N_48165,N_48207);
and U49263 (N_49263,N_48785,N_48028);
nor U49264 (N_49264,N_48675,N_48443);
nand U49265 (N_49265,N_48602,N_48894);
nand U49266 (N_49266,N_48566,N_48777);
and U49267 (N_49267,N_48773,N_48488);
nand U49268 (N_49268,N_48195,N_48396);
and U49269 (N_49269,N_48627,N_48362);
nor U49270 (N_49270,N_48425,N_48031);
and U49271 (N_49271,N_48989,N_48657);
xor U49272 (N_49272,N_48308,N_48760);
xor U49273 (N_49273,N_48445,N_48223);
nor U49274 (N_49274,N_48326,N_48594);
nor U49275 (N_49275,N_48392,N_48379);
or U49276 (N_49276,N_48901,N_48409);
nand U49277 (N_49277,N_48473,N_48274);
or U49278 (N_49278,N_48978,N_48415);
xor U49279 (N_49279,N_48063,N_48662);
nor U49280 (N_49280,N_48191,N_48964);
and U49281 (N_49281,N_48202,N_48615);
nand U49282 (N_49282,N_48751,N_48446);
nand U49283 (N_49283,N_48629,N_48535);
xnor U49284 (N_49284,N_48783,N_48144);
or U49285 (N_49285,N_48434,N_48272);
nor U49286 (N_49286,N_48486,N_48692);
nand U49287 (N_49287,N_48215,N_48737);
xnor U49288 (N_49288,N_48558,N_48511);
nor U49289 (N_49289,N_48041,N_48789);
and U49290 (N_49290,N_48963,N_48050);
or U49291 (N_49291,N_48857,N_48135);
or U49292 (N_49292,N_48844,N_48676);
or U49293 (N_49293,N_48527,N_48809);
nand U49294 (N_49294,N_48481,N_48220);
and U49295 (N_49295,N_48351,N_48412);
xor U49296 (N_49296,N_48742,N_48400);
or U49297 (N_49297,N_48160,N_48982);
xnor U49298 (N_49298,N_48744,N_48416);
nand U49299 (N_49299,N_48421,N_48411);
and U49300 (N_49300,N_48643,N_48752);
nor U49301 (N_49301,N_48537,N_48348);
and U49302 (N_49302,N_48394,N_48984);
nand U49303 (N_49303,N_48265,N_48927);
or U49304 (N_49304,N_48763,N_48758);
and U49305 (N_49305,N_48284,N_48876);
and U49306 (N_49306,N_48915,N_48778);
xnor U49307 (N_49307,N_48112,N_48765);
or U49308 (N_49308,N_48632,N_48364);
nor U49309 (N_49309,N_48048,N_48579);
or U49310 (N_49310,N_48678,N_48001);
and U49311 (N_49311,N_48748,N_48198);
and U49312 (N_49312,N_48764,N_48282);
xnor U49313 (N_49313,N_48939,N_48360);
nand U49314 (N_49314,N_48137,N_48007);
or U49315 (N_49315,N_48386,N_48955);
nor U49316 (N_49316,N_48179,N_48807);
nand U49317 (N_49317,N_48356,N_48417);
and U49318 (N_49318,N_48897,N_48118);
or U49319 (N_49319,N_48226,N_48528);
or U49320 (N_49320,N_48635,N_48745);
or U49321 (N_49321,N_48552,N_48214);
nor U49322 (N_49322,N_48872,N_48373);
nor U49323 (N_49323,N_48934,N_48178);
nand U49324 (N_49324,N_48998,N_48887);
and U49325 (N_49325,N_48059,N_48034);
xor U49326 (N_49326,N_48968,N_48664);
xnor U49327 (N_49327,N_48907,N_48474);
and U49328 (N_49328,N_48493,N_48058);
nor U49329 (N_49329,N_48561,N_48181);
or U49330 (N_49330,N_48056,N_48979);
nand U49331 (N_49331,N_48835,N_48849);
and U49332 (N_49332,N_48671,N_48173);
and U49333 (N_49333,N_48714,N_48642);
and U49334 (N_49334,N_48667,N_48330);
xnor U49335 (N_49335,N_48681,N_48290);
and U49336 (N_49336,N_48301,N_48463);
and U49337 (N_49337,N_48127,N_48980);
nand U49338 (N_49338,N_48030,N_48749);
nor U49339 (N_49339,N_48709,N_48686);
and U49340 (N_49340,N_48680,N_48717);
and U49341 (N_49341,N_48012,N_48405);
xnor U49342 (N_49342,N_48972,N_48542);
nand U49343 (N_49343,N_48315,N_48187);
nor U49344 (N_49344,N_48559,N_48893);
nor U49345 (N_49345,N_48245,N_48025);
or U49346 (N_49346,N_48834,N_48500);
nand U49347 (N_49347,N_48432,N_48774);
nand U49348 (N_49348,N_48850,N_48151);
nand U49349 (N_49349,N_48139,N_48924);
nor U49350 (N_49350,N_48037,N_48069);
xor U49351 (N_49351,N_48974,N_48494);
nor U49352 (N_49352,N_48252,N_48436);
xnor U49353 (N_49353,N_48371,N_48116);
or U49354 (N_49354,N_48508,N_48154);
or U49355 (N_49355,N_48733,N_48419);
nor U49356 (N_49356,N_48082,N_48203);
xnor U49357 (N_49357,N_48159,N_48814);
nor U49358 (N_49358,N_48768,N_48985);
or U49359 (N_49359,N_48625,N_48480);
and U49360 (N_49360,N_48466,N_48653);
xnor U49361 (N_49361,N_48581,N_48699);
or U49362 (N_49362,N_48140,N_48046);
nand U49363 (N_49363,N_48529,N_48024);
nand U49364 (N_49364,N_48237,N_48925);
xor U49365 (N_49365,N_48442,N_48563);
nor U49366 (N_49366,N_48606,N_48352);
xnor U49367 (N_49367,N_48251,N_48706);
xor U49368 (N_49368,N_48375,N_48916);
or U49369 (N_49369,N_48143,N_48969);
or U49370 (N_49370,N_48257,N_48131);
and U49371 (N_49371,N_48152,N_48838);
xnor U49372 (N_49372,N_48704,N_48633);
nor U49373 (N_49373,N_48649,N_48583);
and U49374 (N_49374,N_48619,N_48285);
and U49375 (N_49375,N_48003,N_48438);
xor U49376 (N_49376,N_48910,N_48051);
nor U49377 (N_49377,N_48617,N_48359);
and U49378 (N_49378,N_48276,N_48799);
or U49379 (N_49379,N_48485,N_48841);
nand U49380 (N_49380,N_48349,N_48099);
and U49381 (N_49381,N_48846,N_48150);
and U49382 (N_49382,N_48460,N_48094);
nand U49383 (N_49383,N_48618,N_48847);
xor U49384 (N_49384,N_48010,N_48132);
and U49385 (N_49385,N_48122,N_48685);
xnor U49386 (N_49386,N_48567,N_48489);
nor U49387 (N_49387,N_48142,N_48996);
nor U49388 (N_49388,N_48240,N_48936);
xor U49389 (N_49389,N_48655,N_48447);
nor U49390 (N_49390,N_48217,N_48264);
xnor U49391 (N_49391,N_48790,N_48155);
or U49392 (N_49392,N_48861,N_48584);
or U49393 (N_49393,N_48224,N_48569);
and U49394 (N_49394,N_48383,N_48795);
nor U49395 (N_49395,N_48947,N_48971);
and U49396 (N_49396,N_48855,N_48496);
and U49397 (N_49397,N_48571,N_48476);
and U49398 (N_49398,N_48219,N_48206);
nor U49399 (N_49399,N_48873,N_48539);
and U49400 (N_49400,N_48027,N_48084);
or U49401 (N_49401,N_48015,N_48270);
nor U49402 (N_49402,N_48322,N_48598);
and U49403 (N_49403,N_48085,N_48381);
xor U49404 (N_49404,N_48929,N_48169);
nand U49405 (N_49405,N_48049,N_48695);
nand U49406 (N_49406,N_48238,N_48522);
xor U49407 (N_49407,N_48129,N_48874);
and U49408 (N_49408,N_48641,N_48510);
or U49409 (N_49409,N_48125,N_48912);
or U49410 (N_49410,N_48784,N_48020);
xor U49411 (N_49411,N_48487,N_48639);
and U49412 (N_49412,N_48854,N_48523);
nand U49413 (N_49413,N_48842,N_48600);
nand U49414 (N_49414,N_48374,N_48553);
nand U49415 (N_49415,N_48167,N_48070);
xnor U49416 (N_49416,N_48794,N_48941);
or U49417 (N_49417,N_48287,N_48585);
and U49418 (N_49418,N_48871,N_48121);
xnor U49419 (N_49419,N_48976,N_48757);
or U49420 (N_49420,N_48577,N_48029);
and U49421 (N_49421,N_48932,N_48530);
nand U49422 (N_49422,N_48517,N_48688);
xnor U49423 (N_49423,N_48077,N_48337);
and U49424 (N_49424,N_48444,N_48004);
xor U49425 (N_49425,N_48544,N_48702);
or U49426 (N_49426,N_48113,N_48039);
or U49427 (N_49427,N_48918,N_48241);
or U49428 (N_49428,N_48729,N_48227);
nor U49429 (N_49429,N_48185,N_48853);
nor U49430 (N_49430,N_48166,N_48319);
nand U49431 (N_49431,N_48382,N_48616);
or U49432 (N_49432,N_48339,N_48593);
and U49433 (N_49433,N_48055,N_48895);
and U49434 (N_49434,N_48578,N_48250);
and U49435 (N_49435,N_48839,N_48921);
xor U49436 (N_49436,N_48254,N_48644);
nand U49437 (N_49437,N_48666,N_48148);
nand U49438 (N_49438,N_48040,N_48832);
and U49439 (N_49439,N_48193,N_48782);
or U49440 (N_49440,N_48928,N_48723);
or U49441 (N_49441,N_48875,N_48988);
nand U49442 (N_49442,N_48133,N_48430);
or U49443 (N_49443,N_48278,N_48428);
xor U49444 (N_49444,N_48526,N_48218);
xnor U49445 (N_49445,N_48507,N_48949);
and U49446 (N_49446,N_48231,N_48289);
nor U49447 (N_49447,N_48564,N_48376);
xor U49448 (N_49448,N_48937,N_48609);
xnor U49449 (N_49449,N_48691,N_48922);
xor U49450 (N_49450,N_48518,N_48103);
nor U49451 (N_49451,N_48388,N_48045);
or U49452 (N_49452,N_48426,N_48325);
and U49453 (N_49453,N_48391,N_48053);
or U49454 (N_49454,N_48017,N_48607);
and U49455 (N_49455,N_48590,N_48534);
xor U49456 (N_49456,N_48648,N_48372);
and U49457 (N_49457,N_48080,N_48811);
nand U49458 (N_49458,N_48776,N_48345);
xnor U49459 (N_49459,N_48519,N_48825);
nor U49460 (N_49460,N_48104,N_48881);
nand U49461 (N_49461,N_48886,N_48712);
nand U49462 (N_49462,N_48993,N_48588);
nand U49463 (N_49463,N_48965,N_48819);
nand U49464 (N_49464,N_48385,N_48377);
nand U49465 (N_49465,N_48269,N_48141);
or U49466 (N_49466,N_48710,N_48079);
nand U49467 (N_49467,N_48467,N_48611);
and U49468 (N_49468,N_48109,N_48470);
nand U49469 (N_49469,N_48418,N_48115);
or U49470 (N_49470,N_48913,N_48249);
nand U49471 (N_49471,N_48658,N_48890);
nor U49472 (N_49472,N_48862,N_48266);
nand U49473 (N_49473,N_48472,N_48102);
nand U49474 (N_49474,N_48651,N_48074);
and U49475 (N_49475,N_48803,N_48395);
nand U49476 (N_49476,N_48595,N_48440);
or U49477 (N_49477,N_48387,N_48677);
and U49478 (N_49478,N_48864,N_48083);
nand U49479 (N_49479,N_48128,N_48647);
nor U49480 (N_49480,N_48216,N_48514);
or U49481 (N_49481,N_48429,N_48057);
xor U49482 (N_49482,N_48959,N_48813);
xnor U49483 (N_49483,N_48668,N_48316);
nor U49484 (N_49484,N_48805,N_48628);
or U49485 (N_49485,N_48292,N_48716);
nor U49486 (N_49486,N_48268,N_48310);
nor U49487 (N_49487,N_48108,N_48378);
nor U49488 (N_49488,N_48087,N_48406);
or U49489 (N_49489,N_48540,N_48545);
or U49490 (N_49490,N_48335,N_48194);
nand U49491 (N_49491,N_48798,N_48822);
or U49492 (N_49492,N_48898,N_48793);
xor U49493 (N_49493,N_48506,N_48690);
and U49494 (N_49494,N_48452,N_48146);
nor U49495 (N_49495,N_48209,N_48183);
or U49496 (N_49496,N_48957,N_48407);
or U49497 (N_49497,N_48408,N_48513);
and U49498 (N_49498,N_48689,N_48279);
and U49499 (N_49499,N_48261,N_48192);
and U49500 (N_49500,N_48062,N_48924);
and U49501 (N_49501,N_48071,N_48768);
nand U49502 (N_49502,N_48570,N_48102);
and U49503 (N_49503,N_48642,N_48545);
or U49504 (N_49504,N_48645,N_48270);
xnor U49505 (N_49505,N_48124,N_48630);
or U49506 (N_49506,N_48333,N_48994);
xor U49507 (N_49507,N_48836,N_48204);
and U49508 (N_49508,N_48950,N_48925);
or U49509 (N_49509,N_48070,N_48340);
nand U49510 (N_49510,N_48585,N_48314);
xnor U49511 (N_49511,N_48894,N_48809);
nand U49512 (N_49512,N_48329,N_48003);
and U49513 (N_49513,N_48449,N_48028);
nand U49514 (N_49514,N_48568,N_48523);
or U49515 (N_49515,N_48041,N_48617);
or U49516 (N_49516,N_48818,N_48222);
nor U49517 (N_49517,N_48401,N_48914);
nand U49518 (N_49518,N_48348,N_48874);
or U49519 (N_49519,N_48346,N_48180);
and U49520 (N_49520,N_48845,N_48454);
nand U49521 (N_49521,N_48398,N_48606);
xor U49522 (N_49522,N_48635,N_48442);
or U49523 (N_49523,N_48452,N_48347);
nand U49524 (N_49524,N_48291,N_48625);
and U49525 (N_49525,N_48281,N_48433);
and U49526 (N_49526,N_48861,N_48233);
xor U49527 (N_49527,N_48853,N_48661);
nand U49528 (N_49528,N_48078,N_48400);
and U49529 (N_49529,N_48384,N_48618);
nor U49530 (N_49530,N_48440,N_48768);
xnor U49531 (N_49531,N_48836,N_48020);
nor U49532 (N_49532,N_48061,N_48702);
xnor U49533 (N_49533,N_48447,N_48560);
and U49534 (N_49534,N_48183,N_48972);
and U49535 (N_49535,N_48533,N_48614);
nor U49536 (N_49536,N_48899,N_48568);
nor U49537 (N_49537,N_48701,N_48554);
nand U49538 (N_49538,N_48581,N_48765);
xnor U49539 (N_49539,N_48976,N_48846);
or U49540 (N_49540,N_48351,N_48222);
or U49541 (N_49541,N_48481,N_48506);
or U49542 (N_49542,N_48169,N_48185);
nand U49543 (N_49543,N_48799,N_48015);
nor U49544 (N_49544,N_48504,N_48620);
xnor U49545 (N_49545,N_48667,N_48061);
nand U49546 (N_49546,N_48780,N_48884);
and U49547 (N_49547,N_48239,N_48434);
and U49548 (N_49548,N_48422,N_48477);
nand U49549 (N_49549,N_48366,N_48425);
or U49550 (N_49550,N_48781,N_48955);
and U49551 (N_49551,N_48324,N_48848);
or U49552 (N_49552,N_48516,N_48731);
nand U49553 (N_49553,N_48975,N_48965);
or U49554 (N_49554,N_48762,N_48435);
nand U49555 (N_49555,N_48157,N_48951);
nor U49556 (N_49556,N_48343,N_48701);
xnor U49557 (N_49557,N_48796,N_48192);
nand U49558 (N_49558,N_48438,N_48948);
nand U49559 (N_49559,N_48798,N_48152);
xnor U49560 (N_49560,N_48268,N_48609);
nor U49561 (N_49561,N_48609,N_48584);
xor U49562 (N_49562,N_48098,N_48824);
or U49563 (N_49563,N_48244,N_48877);
nor U49564 (N_49564,N_48967,N_48140);
nand U49565 (N_49565,N_48417,N_48712);
nor U49566 (N_49566,N_48776,N_48977);
and U49567 (N_49567,N_48128,N_48482);
nor U49568 (N_49568,N_48481,N_48671);
nand U49569 (N_49569,N_48324,N_48777);
nor U49570 (N_49570,N_48952,N_48218);
nor U49571 (N_49571,N_48496,N_48122);
or U49572 (N_49572,N_48505,N_48426);
nand U49573 (N_49573,N_48317,N_48786);
and U49574 (N_49574,N_48538,N_48693);
or U49575 (N_49575,N_48099,N_48404);
nor U49576 (N_49576,N_48101,N_48200);
nor U49577 (N_49577,N_48404,N_48130);
nor U49578 (N_49578,N_48125,N_48119);
nand U49579 (N_49579,N_48529,N_48179);
or U49580 (N_49580,N_48839,N_48498);
xnor U49581 (N_49581,N_48148,N_48123);
nand U49582 (N_49582,N_48412,N_48225);
and U49583 (N_49583,N_48407,N_48990);
or U49584 (N_49584,N_48770,N_48431);
xnor U49585 (N_49585,N_48923,N_48173);
nand U49586 (N_49586,N_48868,N_48408);
nand U49587 (N_49587,N_48046,N_48420);
and U49588 (N_49588,N_48314,N_48780);
xnor U49589 (N_49589,N_48242,N_48280);
nand U49590 (N_49590,N_48443,N_48458);
or U49591 (N_49591,N_48009,N_48458);
or U49592 (N_49592,N_48002,N_48984);
or U49593 (N_49593,N_48308,N_48404);
nor U49594 (N_49594,N_48511,N_48830);
and U49595 (N_49595,N_48158,N_48014);
nor U49596 (N_49596,N_48429,N_48807);
or U49597 (N_49597,N_48094,N_48600);
and U49598 (N_49598,N_48583,N_48846);
nand U49599 (N_49599,N_48731,N_48296);
xnor U49600 (N_49600,N_48996,N_48026);
nor U49601 (N_49601,N_48293,N_48159);
or U49602 (N_49602,N_48923,N_48986);
nor U49603 (N_49603,N_48501,N_48137);
and U49604 (N_49604,N_48664,N_48673);
nand U49605 (N_49605,N_48029,N_48252);
nor U49606 (N_49606,N_48848,N_48349);
xnor U49607 (N_49607,N_48533,N_48905);
and U49608 (N_49608,N_48455,N_48331);
or U49609 (N_49609,N_48196,N_48504);
nand U49610 (N_49610,N_48264,N_48841);
and U49611 (N_49611,N_48793,N_48137);
and U49612 (N_49612,N_48410,N_48255);
and U49613 (N_49613,N_48964,N_48204);
nand U49614 (N_49614,N_48464,N_48349);
xnor U49615 (N_49615,N_48801,N_48582);
nand U49616 (N_49616,N_48358,N_48187);
or U49617 (N_49617,N_48635,N_48140);
or U49618 (N_49618,N_48734,N_48926);
or U49619 (N_49619,N_48410,N_48452);
or U49620 (N_49620,N_48156,N_48998);
xor U49621 (N_49621,N_48974,N_48945);
and U49622 (N_49622,N_48956,N_48700);
or U49623 (N_49623,N_48038,N_48980);
xor U49624 (N_49624,N_48722,N_48645);
nor U49625 (N_49625,N_48768,N_48875);
nor U49626 (N_49626,N_48895,N_48321);
nand U49627 (N_49627,N_48890,N_48517);
nor U49628 (N_49628,N_48532,N_48984);
nor U49629 (N_49629,N_48909,N_48175);
nand U49630 (N_49630,N_48742,N_48970);
nand U49631 (N_49631,N_48616,N_48535);
and U49632 (N_49632,N_48139,N_48849);
xor U49633 (N_49633,N_48698,N_48812);
nor U49634 (N_49634,N_48577,N_48230);
nor U49635 (N_49635,N_48306,N_48648);
and U49636 (N_49636,N_48341,N_48707);
xnor U49637 (N_49637,N_48033,N_48051);
or U49638 (N_49638,N_48788,N_48310);
xnor U49639 (N_49639,N_48133,N_48387);
nand U49640 (N_49640,N_48633,N_48362);
or U49641 (N_49641,N_48194,N_48236);
xnor U49642 (N_49642,N_48878,N_48660);
nor U49643 (N_49643,N_48351,N_48902);
nor U49644 (N_49644,N_48848,N_48171);
or U49645 (N_49645,N_48369,N_48281);
xnor U49646 (N_49646,N_48259,N_48690);
nor U49647 (N_49647,N_48456,N_48584);
or U49648 (N_49648,N_48462,N_48931);
xor U49649 (N_49649,N_48919,N_48895);
xnor U49650 (N_49650,N_48600,N_48390);
nand U49651 (N_49651,N_48857,N_48479);
or U49652 (N_49652,N_48168,N_48047);
and U49653 (N_49653,N_48454,N_48748);
xor U49654 (N_49654,N_48681,N_48908);
nand U49655 (N_49655,N_48042,N_48492);
and U49656 (N_49656,N_48597,N_48640);
xor U49657 (N_49657,N_48651,N_48944);
and U49658 (N_49658,N_48007,N_48669);
or U49659 (N_49659,N_48688,N_48728);
or U49660 (N_49660,N_48142,N_48602);
and U49661 (N_49661,N_48646,N_48607);
and U49662 (N_49662,N_48124,N_48548);
or U49663 (N_49663,N_48887,N_48068);
and U49664 (N_49664,N_48893,N_48932);
xnor U49665 (N_49665,N_48394,N_48108);
and U49666 (N_49666,N_48292,N_48071);
nor U49667 (N_49667,N_48970,N_48518);
nand U49668 (N_49668,N_48111,N_48050);
xnor U49669 (N_49669,N_48389,N_48097);
and U49670 (N_49670,N_48896,N_48462);
or U49671 (N_49671,N_48151,N_48923);
xor U49672 (N_49672,N_48108,N_48202);
xnor U49673 (N_49673,N_48025,N_48199);
xnor U49674 (N_49674,N_48959,N_48406);
nor U49675 (N_49675,N_48955,N_48553);
nor U49676 (N_49676,N_48538,N_48393);
nor U49677 (N_49677,N_48981,N_48083);
and U49678 (N_49678,N_48057,N_48436);
nand U49679 (N_49679,N_48975,N_48709);
nand U49680 (N_49680,N_48104,N_48168);
nor U49681 (N_49681,N_48454,N_48210);
xnor U49682 (N_49682,N_48311,N_48948);
nand U49683 (N_49683,N_48451,N_48970);
nand U49684 (N_49684,N_48893,N_48521);
xor U49685 (N_49685,N_48115,N_48962);
nor U49686 (N_49686,N_48083,N_48576);
or U49687 (N_49687,N_48590,N_48346);
or U49688 (N_49688,N_48587,N_48096);
nand U49689 (N_49689,N_48209,N_48220);
xnor U49690 (N_49690,N_48811,N_48178);
nand U49691 (N_49691,N_48084,N_48267);
nor U49692 (N_49692,N_48503,N_48745);
nand U49693 (N_49693,N_48426,N_48417);
xnor U49694 (N_49694,N_48888,N_48223);
nor U49695 (N_49695,N_48467,N_48664);
or U49696 (N_49696,N_48266,N_48404);
xnor U49697 (N_49697,N_48551,N_48039);
nand U49698 (N_49698,N_48230,N_48963);
and U49699 (N_49699,N_48405,N_48345);
or U49700 (N_49700,N_48284,N_48450);
nor U49701 (N_49701,N_48509,N_48560);
and U49702 (N_49702,N_48167,N_48671);
nand U49703 (N_49703,N_48292,N_48068);
or U49704 (N_49704,N_48403,N_48987);
nand U49705 (N_49705,N_48257,N_48340);
xnor U49706 (N_49706,N_48296,N_48522);
nor U49707 (N_49707,N_48815,N_48551);
xnor U49708 (N_49708,N_48987,N_48712);
nor U49709 (N_49709,N_48773,N_48709);
nor U49710 (N_49710,N_48088,N_48283);
and U49711 (N_49711,N_48243,N_48701);
xnor U49712 (N_49712,N_48965,N_48779);
xnor U49713 (N_49713,N_48984,N_48079);
or U49714 (N_49714,N_48503,N_48112);
nor U49715 (N_49715,N_48611,N_48909);
nor U49716 (N_49716,N_48392,N_48664);
nor U49717 (N_49717,N_48770,N_48335);
and U49718 (N_49718,N_48137,N_48233);
and U49719 (N_49719,N_48554,N_48715);
nor U49720 (N_49720,N_48479,N_48972);
nand U49721 (N_49721,N_48287,N_48300);
or U49722 (N_49722,N_48278,N_48300);
xnor U49723 (N_49723,N_48588,N_48188);
and U49724 (N_49724,N_48142,N_48915);
or U49725 (N_49725,N_48412,N_48931);
nor U49726 (N_49726,N_48854,N_48157);
nand U49727 (N_49727,N_48033,N_48216);
nand U49728 (N_49728,N_48737,N_48411);
or U49729 (N_49729,N_48132,N_48805);
nand U49730 (N_49730,N_48212,N_48830);
or U49731 (N_49731,N_48788,N_48711);
xor U49732 (N_49732,N_48431,N_48332);
or U49733 (N_49733,N_48251,N_48130);
nand U49734 (N_49734,N_48545,N_48733);
and U49735 (N_49735,N_48418,N_48178);
nand U49736 (N_49736,N_48340,N_48358);
and U49737 (N_49737,N_48212,N_48441);
xor U49738 (N_49738,N_48947,N_48965);
xnor U49739 (N_49739,N_48562,N_48466);
and U49740 (N_49740,N_48656,N_48434);
or U49741 (N_49741,N_48529,N_48394);
or U49742 (N_49742,N_48467,N_48484);
and U49743 (N_49743,N_48085,N_48178);
xor U49744 (N_49744,N_48876,N_48666);
nor U49745 (N_49745,N_48941,N_48457);
and U49746 (N_49746,N_48981,N_48998);
nor U49747 (N_49747,N_48684,N_48555);
nand U49748 (N_49748,N_48983,N_48889);
nor U49749 (N_49749,N_48926,N_48084);
or U49750 (N_49750,N_48780,N_48232);
and U49751 (N_49751,N_48830,N_48843);
and U49752 (N_49752,N_48216,N_48336);
nor U49753 (N_49753,N_48777,N_48528);
nand U49754 (N_49754,N_48692,N_48747);
nand U49755 (N_49755,N_48383,N_48431);
xnor U49756 (N_49756,N_48687,N_48550);
xnor U49757 (N_49757,N_48778,N_48530);
nor U49758 (N_49758,N_48078,N_48846);
or U49759 (N_49759,N_48890,N_48957);
and U49760 (N_49760,N_48216,N_48023);
nand U49761 (N_49761,N_48544,N_48646);
nor U49762 (N_49762,N_48040,N_48397);
xnor U49763 (N_49763,N_48522,N_48211);
nand U49764 (N_49764,N_48912,N_48548);
xor U49765 (N_49765,N_48502,N_48563);
nor U49766 (N_49766,N_48568,N_48701);
or U49767 (N_49767,N_48319,N_48516);
nand U49768 (N_49768,N_48794,N_48335);
nor U49769 (N_49769,N_48711,N_48631);
xor U49770 (N_49770,N_48651,N_48277);
xnor U49771 (N_49771,N_48536,N_48553);
nor U49772 (N_49772,N_48888,N_48057);
xor U49773 (N_49773,N_48715,N_48217);
nor U49774 (N_49774,N_48966,N_48005);
nand U49775 (N_49775,N_48045,N_48264);
nand U49776 (N_49776,N_48143,N_48052);
or U49777 (N_49777,N_48783,N_48252);
nand U49778 (N_49778,N_48450,N_48203);
or U49779 (N_49779,N_48985,N_48264);
nand U49780 (N_49780,N_48310,N_48363);
xnor U49781 (N_49781,N_48864,N_48056);
or U49782 (N_49782,N_48923,N_48175);
nand U49783 (N_49783,N_48673,N_48428);
nand U49784 (N_49784,N_48377,N_48499);
nor U49785 (N_49785,N_48787,N_48617);
xor U49786 (N_49786,N_48380,N_48198);
or U49787 (N_49787,N_48126,N_48972);
or U49788 (N_49788,N_48867,N_48446);
nor U49789 (N_49789,N_48236,N_48996);
xor U49790 (N_49790,N_48249,N_48360);
or U49791 (N_49791,N_48286,N_48099);
nor U49792 (N_49792,N_48774,N_48214);
or U49793 (N_49793,N_48522,N_48074);
nand U49794 (N_49794,N_48515,N_48638);
nor U49795 (N_49795,N_48275,N_48240);
xnor U49796 (N_49796,N_48226,N_48533);
xor U49797 (N_49797,N_48290,N_48842);
nand U49798 (N_49798,N_48331,N_48113);
or U49799 (N_49799,N_48811,N_48050);
and U49800 (N_49800,N_48874,N_48044);
and U49801 (N_49801,N_48561,N_48477);
and U49802 (N_49802,N_48796,N_48062);
nand U49803 (N_49803,N_48093,N_48911);
or U49804 (N_49804,N_48457,N_48722);
and U49805 (N_49805,N_48541,N_48180);
or U49806 (N_49806,N_48750,N_48522);
nand U49807 (N_49807,N_48719,N_48819);
or U49808 (N_49808,N_48771,N_48882);
nor U49809 (N_49809,N_48458,N_48340);
nor U49810 (N_49810,N_48185,N_48492);
nor U49811 (N_49811,N_48887,N_48326);
nor U49812 (N_49812,N_48215,N_48055);
and U49813 (N_49813,N_48340,N_48743);
and U49814 (N_49814,N_48502,N_48115);
xnor U49815 (N_49815,N_48329,N_48236);
or U49816 (N_49816,N_48933,N_48618);
or U49817 (N_49817,N_48852,N_48603);
nor U49818 (N_49818,N_48318,N_48026);
nand U49819 (N_49819,N_48830,N_48588);
and U49820 (N_49820,N_48267,N_48624);
or U49821 (N_49821,N_48608,N_48328);
xnor U49822 (N_49822,N_48871,N_48325);
nand U49823 (N_49823,N_48259,N_48838);
or U49824 (N_49824,N_48721,N_48783);
xor U49825 (N_49825,N_48207,N_48367);
nand U49826 (N_49826,N_48517,N_48431);
or U49827 (N_49827,N_48859,N_48038);
xnor U49828 (N_49828,N_48728,N_48310);
nand U49829 (N_49829,N_48446,N_48960);
xnor U49830 (N_49830,N_48774,N_48656);
xor U49831 (N_49831,N_48321,N_48673);
xnor U49832 (N_49832,N_48473,N_48160);
or U49833 (N_49833,N_48410,N_48634);
nand U49834 (N_49834,N_48979,N_48453);
and U49835 (N_49835,N_48992,N_48474);
or U49836 (N_49836,N_48135,N_48299);
nor U49837 (N_49837,N_48927,N_48371);
and U49838 (N_49838,N_48244,N_48931);
and U49839 (N_49839,N_48696,N_48727);
xnor U49840 (N_49840,N_48924,N_48477);
and U49841 (N_49841,N_48210,N_48662);
xor U49842 (N_49842,N_48466,N_48252);
nor U49843 (N_49843,N_48021,N_48337);
or U49844 (N_49844,N_48572,N_48438);
or U49845 (N_49845,N_48790,N_48793);
nand U49846 (N_49846,N_48988,N_48267);
nand U49847 (N_49847,N_48142,N_48882);
and U49848 (N_49848,N_48575,N_48469);
xnor U49849 (N_49849,N_48326,N_48106);
xnor U49850 (N_49850,N_48811,N_48396);
nor U49851 (N_49851,N_48910,N_48101);
nand U49852 (N_49852,N_48046,N_48862);
nor U49853 (N_49853,N_48693,N_48501);
nand U49854 (N_49854,N_48058,N_48189);
nand U49855 (N_49855,N_48041,N_48047);
nand U49856 (N_49856,N_48896,N_48275);
nor U49857 (N_49857,N_48215,N_48192);
xor U49858 (N_49858,N_48044,N_48438);
nor U49859 (N_49859,N_48847,N_48556);
nand U49860 (N_49860,N_48765,N_48539);
xnor U49861 (N_49861,N_48971,N_48433);
nand U49862 (N_49862,N_48867,N_48483);
or U49863 (N_49863,N_48854,N_48534);
nand U49864 (N_49864,N_48245,N_48741);
xor U49865 (N_49865,N_48613,N_48677);
xor U49866 (N_49866,N_48006,N_48964);
and U49867 (N_49867,N_48488,N_48272);
or U49868 (N_49868,N_48625,N_48844);
nor U49869 (N_49869,N_48881,N_48225);
or U49870 (N_49870,N_48759,N_48816);
xnor U49871 (N_49871,N_48519,N_48009);
and U49872 (N_49872,N_48730,N_48999);
nor U49873 (N_49873,N_48712,N_48025);
nor U49874 (N_49874,N_48452,N_48719);
xor U49875 (N_49875,N_48967,N_48278);
nand U49876 (N_49876,N_48810,N_48454);
xor U49877 (N_49877,N_48812,N_48899);
xor U49878 (N_49878,N_48550,N_48841);
and U49879 (N_49879,N_48074,N_48138);
xor U49880 (N_49880,N_48839,N_48550);
xor U49881 (N_49881,N_48099,N_48448);
nor U49882 (N_49882,N_48348,N_48119);
or U49883 (N_49883,N_48236,N_48244);
and U49884 (N_49884,N_48892,N_48912);
nand U49885 (N_49885,N_48512,N_48207);
xnor U49886 (N_49886,N_48640,N_48156);
and U49887 (N_49887,N_48401,N_48822);
nand U49888 (N_49888,N_48129,N_48304);
nor U49889 (N_49889,N_48320,N_48202);
xor U49890 (N_49890,N_48741,N_48305);
xor U49891 (N_49891,N_48933,N_48676);
xor U49892 (N_49892,N_48623,N_48254);
nand U49893 (N_49893,N_48308,N_48621);
and U49894 (N_49894,N_48697,N_48627);
xor U49895 (N_49895,N_48808,N_48183);
xnor U49896 (N_49896,N_48626,N_48992);
nor U49897 (N_49897,N_48843,N_48709);
nand U49898 (N_49898,N_48428,N_48821);
nand U49899 (N_49899,N_48553,N_48099);
and U49900 (N_49900,N_48976,N_48811);
and U49901 (N_49901,N_48418,N_48846);
nor U49902 (N_49902,N_48337,N_48956);
nor U49903 (N_49903,N_48630,N_48599);
or U49904 (N_49904,N_48318,N_48968);
or U49905 (N_49905,N_48653,N_48301);
xnor U49906 (N_49906,N_48227,N_48845);
xor U49907 (N_49907,N_48808,N_48087);
xor U49908 (N_49908,N_48816,N_48397);
and U49909 (N_49909,N_48038,N_48462);
or U49910 (N_49910,N_48642,N_48256);
or U49911 (N_49911,N_48132,N_48709);
nor U49912 (N_49912,N_48252,N_48048);
nand U49913 (N_49913,N_48666,N_48538);
xor U49914 (N_49914,N_48251,N_48186);
and U49915 (N_49915,N_48088,N_48200);
nand U49916 (N_49916,N_48811,N_48002);
xnor U49917 (N_49917,N_48840,N_48769);
nand U49918 (N_49918,N_48154,N_48991);
and U49919 (N_49919,N_48283,N_48559);
nor U49920 (N_49920,N_48575,N_48915);
nor U49921 (N_49921,N_48985,N_48949);
nor U49922 (N_49922,N_48209,N_48770);
nand U49923 (N_49923,N_48772,N_48900);
xor U49924 (N_49924,N_48269,N_48018);
xnor U49925 (N_49925,N_48394,N_48262);
or U49926 (N_49926,N_48077,N_48191);
nor U49927 (N_49927,N_48338,N_48305);
nand U49928 (N_49928,N_48572,N_48953);
nor U49929 (N_49929,N_48893,N_48605);
and U49930 (N_49930,N_48941,N_48857);
nand U49931 (N_49931,N_48582,N_48044);
and U49932 (N_49932,N_48386,N_48008);
nor U49933 (N_49933,N_48125,N_48549);
xnor U49934 (N_49934,N_48868,N_48675);
and U49935 (N_49935,N_48035,N_48063);
and U49936 (N_49936,N_48550,N_48866);
nand U49937 (N_49937,N_48937,N_48395);
nor U49938 (N_49938,N_48633,N_48714);
and U49939 (N_49939,N_48575,N_48403);
nand U49940 (N_49940,N_48814,N_48855);
and U49941 (N_49941,N_48526,N_48514);
and U49942 (N_49942,N_48116,N_48581);
or U49943 (N_49943,N_48330,N_48720);
nand U49944 (N_49944,N_48477,N_48672);
xnor U49945 (N_49945,N_48723,N_48845);
nand U49946 (N_49946,N_48212,N_48187);
xor U49947 (N_49947,N_48775,N_48265);
nand U49948 (N_49948,N_48211,N_48259);
nor U49949 (N_49949,N_48147,N_48527);
or U49950 (N_49950,N_48043,N_48146);
and U49951 (N_49951,N_48427,N_48370);
and U49952 (N_49952,N_48675,N_48260);
and U49953 (N_49953,N_48092,N_48088);
nand U49954 (N_49954,N_48440,N_48919);
nand U49955 (N_49955,N_48679,N_48277);
xor U49956 (N_49956,N_48979,N_48514);
and U49957 (N_49957,N_48574,N_48551);
and U49958 (N_49958,N_48210,N_48095);
nand U49959 (N_49959,N_48734,N_48597);
and U49960 (N_49960,N_48375,N_48790);
and U49961 (N_49961,N_48263,N_48144);
nor U49962 (N_49962,N_48715,N_48066);
or U49963 (N_49963,N_48799,N_48136);
and U49964 (N_49964,N_48978,N_48663);
nand U49965 (N_49965,N_48067,N_48993);
nor U49966 (N_49966,N_48970,N_48260);
nand U49967 (N_49967,N_48429,N_48372);
xnor U49968 (N_49968,N_48435,N_48734);
nor U49969 (N_49969,N_48235,N_48681);
nand U49970 (N_49970,N_48769,N_48603);
or U49971 (N_49971,N_48464,N_48147);
nand U49972 (N_49972,N_48801,N_48766);
nand U49973 (N_49973,N_48605,N_48111);
and U49974 (N_49974,N_48721,N_48121);
nand U49975 (N_49975,N_48352,N_48976);
nand U49976 (N_49976,N_48001,N_48647);
or U49977 (N_49977,N_48955,N_48628);
nor U49978 (N_49978,N_48366,N_48939);
xnor U49979 (N_49979,N_48460,N_48081);
nor U49980 (N_49980,N_48362,N_48809);
nor U49981 (N_49981,N_48106,N_48573);
xnor U49982 (N_49982,N_48982,N_48244);
nor U49983 (N_49983,N_48608,N_48645);
or U49984 (N_49984,N_48407,N_48167);
nor U49985 (N_49985,N_48245,N_48339);
xor U49986 (N_49986,N_48431,N_48259);
and U49987 (N_49987,N_48109,N_48783);
xnor U49988 (N_49988,N_48898,N_48112);
or U49989 (N_49989,N_48896,N_48316);
nand U49990 (N_49990,N_48727,N_48777);
xor U49991 (N_49991,N_48015,N_48577);
xor U49992 (N_49992,N_48314,N_48620);
xnor U49993 (N_49993,N_48233,N_48707);
nor U49994 (N_49994,N_48136,N_48686);
nand U49995 (N_49995,N_48536,N_48483);
nor U49996 (N_49996,N_48548,N_48586);
or U49997 (N_49997,N_48929,N_48768);
nand U49998 (N_49998,N_48145,N_48059);
and U49999 (N_49999,N_48854,N_48019);
xor UO_0 (O_0,N_49219,N_49972);
nor UO_1 (O_1,N_49160,N_49203);
or UO_2 (O_2,N_49380,N_49879);
nand UO_3 (O_3,N_49782,N_49664);
xnor UO_4 (O_4,N_49937,N_49572);
xnor UO_5 (O_5,N_49147,N_49079);
or UO_6 (O_6,N_49653,N_49104);
and UO_7 (O_7,N_49202,N_49614);
and UO_8 (O_8,N_49932,N_49454);
and UO_9 (O_9,N_49019,N_49018);
and UO_10 (O_10,N_49978,N_49119);
nor UO_11 (O_11,N_49707,N_49961);
and UO_12 (O_12,N_49680,N_49379);
nand UO_13 (O_13,N_49074,N_49523);
nor UO_14 (O_14,N_49519,N_49336);
or UO_15 (O_15,N_49657,N_49716);
nor UO_16 (O_16,N_49512,N_49719);
nand UO_17 (O_17,N_49113,N_49303);
nor UO_18 (O_18,N_49890,N_49128);
xor UO_19 (O_19,N_49212,N_49730);
and UO_20 (O_20,N_49810,N_49675);
or UO_21 (O_21,N_49737,N_49451);
and UO_22 (O_22,N_49267,N_49249);
or UO_23 (O_23,N_49643,N_49211);
nand UO_24 (O_24,N_49992,N_49189);
and UO_25 (O_25,N_49618,N_49943);
xnor UO_26 (O_26,N_49724,N_49229);
or UO_27 (O_27,N_49656,N_49067);
and UO_28 (O_28,N_49773,N_49838);
xnor UO_29 (O_29,N_49770,N_49860);
nor UO_30 (O_30,N_49504,N_49445);
or UO_31 (O_31,N_49644,N_49630);
xor UO_32 (O_32,N_49489,N_49156);
nand UO_33 (O_33,N_49853,N_49260);
nor UO_34 (O_34,N_49026,N_49514);
nand UO_35 (O_35,N_49101,N_49279);
xor UO_36 (O_36,N_49377,N_49503);
nand UO_37 (O_37,N_49208,N_49049);
nor UO_38 (O_38,N_49486,N_49422);
and UO_39 (O_39,N_49850,N_49798);
xnor UO_40 (O_40,N_49530,N_49914);
nand UO_41 (O_41,N_49066,N_49428);
nor UO_42 (O_42,N_49100,N_49287);
or UO_43 (O_43,N_49632,N_49949);
nor UO_44 (O_44,N_49294,N_49887);
and UO_45 (O_45,N_49224,N_49785);
or UO_46 (O_46,N_49615,N_49579);
nand UO_47 (O_47,N_49401,N_49641);
or UO_48 (O_48,N_49369,N_49538);
and UO_49 (O_49,N_49700,N_49966);
and UO_50 (O_50,N_49330,N_49452);
xor UO_51 (O_51,N_49291,N_49064);
or UO_52 (O_52,N_49031,N_49884);
nor UO_53 (O_53,N_49243,N_49767);
and UO_54 (O_54,N_49662,N_49776);
and UO_55 (O_55,N_49911,N_49044);
and UO_56 (O_56,N_49419,N_49829);
nor UO_57 (O_57,N_49324,N_49755);
or UO_58 (O_58,N_49546,N_49576);
or UO_59 (O_59,N_49191,N_49574);
nor UO_60 (O_60,N_49054,N_49387);
or UO_61 (O_61,N_49868,N_49094);
and UO_62 (O_62,N_49397,N_49305);
nor UO_63 (O_63,N_49723,N_49935);
xnor UO_64 (O_64,N_49593,N_49692);
or UO_65 (O_65,N_49312,N_49315);
xor UO_66 (O_66,N_49455,N_49591);
nand UO_67 (O_67,N_49928,N_49245);
or UO_68 (O_68,N_49023,N_49652);
and UO_69 (O_69,N_49485,N_49424);
xor UO_70 (O_70,N_49908,N_49597);
nand UO_71 (O_71,N_49133,N_49871);
or UO_72 (O_72,N_49665,N_49624);
nand UO_73 (O_73,N_49216,N_49363);
xor UO_74 (O_74,N_49490,N_49043);
and UO_75 (O_75,N_49543,N_49919);
and UO_76 (O_76,N_49778,N_49011);
or UO_77 (O_77,N_49434,N_49750);
nor UO_78 (O_78,N_49760,N_49950);
xor UO_79 (O_79,N_49289,N_49258);
and UO_80 (O_80,N_49600,N_49703);
and UO_81 (O_81,N_49851,N_49320);
or UO_82 (O_82,N_49276,N_49870);
xor UO_83 (O_83,N_49561,N_49448);
nand UO_84 (O_84,N_49999,N_49277);
or UO_85 (O_85,N_49759,N_49227);
nor UO_86 (O_86,N_49002,N_49126);
nor UO_87 (O_87,N_49529,N_49974);
nand UO_88 (O_88,N_49599,N_49836);
xnor UO_89 (O_89,N_49635,N_49352);
or UO_90 (O_90,N_49651,N_49459);
nor UO_91 (O_91,N_49481,N_49153);
nand UO_92 (O_92,N_49115,N_49034);
and UO_93 (O_93,N_49441,N_49461);
nand UO_94 (O_94,N_49112,N_49959);
or UO_95 (O_95,N_49150,N_49117);
nand UO_96 (O_96,N_49030,N_49149);
xnor UO_97 (O_97,N_49779,N_49982);
nand UO_98 (O_98,N_49958,N_49247);
nor UO_99 (O_99,N_49582,N_49334);
and UO_100 (O_100,N_49364,N_49796);
xor UO_101 (O_101,N_49876,N_49041);
and UO_102 (O_102,N_49864,N_49414);
xor UO_103 (O_103,N_49823,N_49148);
nand UO_104 (O_104,N_49934,N_49040);
and UO_105 (O_105,N_49076,N_49408);
xnor UO_106 (O_106,N_49244,N_49904);
xor UO_107 (O_107,N_49403,N_49511);
xor UO_108 (O_108,N_49936,N_49924);
nor UO_109 (O_109,N_49262,N_49215);
nand UO_110 (O_110,N_49736,N_49610);
xor UO_111 (O_111,N_49298,N_49728);
nand UO_112 (O_112,N_49433,N_49797);
and UO_113 (O_113,N_49533,N_49087);
and UO_114 (O_114,N_49883,N_49028);
xnor UO_115 (O_115,N_49078,N_49346);
nor UO_116 (O_116,N_49717,N_49713);
or UO_117 (O_117,N_49619,N_49192);
and UO_118 (O_118,N_49920,N_49093);
nand UO_119 (O_119,N_49359,N_49035);
xnor UO_120 (O_120,N_49912,N_49948);
nand UO_121 (O_121,N_49270,N_49856);
nor UO_122 (O_122,N_49390,N_49991);
xor UO_123 (O_123,N_49726,N_49005);
and UO_124 (O_124,N_49556,N_49129);
nand UO_125 (O_125,N_49568,N_49118);
xnor UO_126 (O_126,N_49575,N_49131);
or UO_127 (O_127,N_49465,N_49627);
and UO_128 (O_128,N_49300,N_49472);
and UO_129 (O_129,N_49400,N_49348);
nand UO_130 (O_130,N_49855,N_49373);
nor UO_131 (O_131,N_49721,N_49701);
xor UO_132 (O_132,N_49432,N_49648);
nand UO_133 (O_133,N_49695,N_49881);
or UO_134 (O_134,N_49009,N_49402);
and UO_135 (O_135,N_49092,N_49822);
and UO_136 (O_136,N_49449,N_49038);
nand UO_137 (O_137,N_49050,N_49492);
or UO_138 (O_138,N_49913,N_49204);
nor UO_139 (O_139,N_49872,N_49562);
nand UO_140 (O_140,N_49537,N_49356);
nand UO_141 (O_141,N_49319,N_49273);
and UO_142 (O_142,N_49174,N_49399);
or UO_143 (O_143,N_49800,N_49226);
and UO_144 (O_144,N_49214,N_49105);
nor UO_145 (O_145,N_49583,N_49354);
and UO_146 (O_146,N_49989,N_49184);
nand UO_147 (O_147,N_49740,N_49951);
or UO_148 (O_148,N_49253,N_49768);
xor UO_149 (O_149,N_49199,N_49251);
nand UO_150 (O_150,N_49467,N_49283);
nand UO_151 (O_151,N_49114,N_49110);
or UO_152 (O_152,N_49848,N_49998);
nor UO_153 (O_153,N_49570,N_49086);
nand UO_154 (O_154,N_49844,N_49517);
nor UO_155 (O_155,N_49068,N_49965);
or UO_156 (O_156,N_49888,N_49731);
nand UO_157 (O_157,N_49024,N_49132);
nor UO_158 (O_158,N_49483,N_49636);
and UO_159 (O_159,N_49197,N_49569);
or UO_160 (O_160,N_49698,N_49140);
nand UO_161 (O_161,N_49438,N_49560);
nand UO_162 (O_162,N_49477,N_49621);
or UO_163 (O_163,N_49286,N_49167);
or UO_164 (O_164,N_49613,N_49764);
and UO_165 (O_165,N_49163,N_49654);
nor UO_166 (O_166,N_49393,N_49825);
nand UO_167 (O_167,N_49317,N_49460);
nand UO_168 (O_168,N_49012,N_49734);
xor UO_169 (O_169,N_49803,N_49802);
nor UO_170 (O_170,N_49997,N_49281);
xnor UO_171 (O_171,N_49754,N_49183);
or UO_172 (O_172,N_49967,N_49268);
and UO_173 (O_173,N_49077,N_49344);
nand UO_174 (O_174,N_49788,N_49687);
or UO_175 (O_175,N_49793,N_49275);
nor UO_176 (O_176,N_49584,N_49639);
xor UO_177 (O_177,N_49993,N_49097);
xor UO_178 (O_178,N_49440,N_49103);
nor UO_179 (O_179,N_49370,N_49099);
and UO_180 (O_180,N_49240,N_49263);
or UO_181 (O_181,N_49906,N_49386);
nor UO_182 (O_182,N_49338,N_49187);
nor UO_183 (O_183,N_49743,N_49238);
or UO_184 (O_184,N_49052,N_49121);
xnor UO_185 (O_185,N_49349,N_49955);
xnor UO_186 (O_186,N_49302,N_49784);
and UO_187 (O_187,N_49055,N_49427);
and UO_188 (O_188,N_49689,N_49587);
xor UO_189 (O_189,N_49415,N_49106);
or UO_190 (O_190,N_49237,N_49827);
nand UO_191 (O_191,N_49350,N_49495);
and UO_192 (O_192,N_49033,N_49491);
nor UO_193 (O_193,N_49817,N_49531);
or UO_194 (O_194,N_49882,N_49235);
nor UO_195 (O_195,N_49196,N_49616);
or UO_196 (O_196,N_49674,N_49606);
or UO_197 (O_197,N_49013,N_49479);
nand UO_198 (O_198,N_49910,N_49786);
nor UO_199 (O_199,N_49371,N_49201);
or UO_200 (O_200,N_49308,N_49520);
and UO_201 (O_201,N_49650,N_49663);
or UO_202 (O_202,N_49304,N_49590);
or UO_203 (O_203,N_49357,N_49378);
nand UO_204 (O_204,N_49930,N_49791);
xor UO_205 (O_205,N_49200,N_49471);
xnor UO_206 (O_206,N_49775,N_49682);
and UO_207 (O_207,N_49343,N_49466);
or UO_208 (O_208,N_49130,N_49946);
xor UO_209 (O_209,N_49231,N_49765);
nor UO_210 (O_210,N_49640,N_49804);
and UO_211 (O_211,N_49248,N_49814);
or UO_212 (O_212,N_49282,N_49548);
nor UO_213 (O_213,N_49411,N_49994);
or UO_214 (O_214,N_49795,N_49554);
and UO_215 (O_215,N_49525,N_49162);
nand UO_216 (O_216,N_49852,N_49507);
nor UO_217 (O_217,N_49960,N_49892);
or UO_218 (O_218,N_49952,N_49666);
nor UO_219 (O_219,N_49351,N_49956);
and UO_220 (O_220,N_49181,N_49145);
or UO_221 (O_221,N_49790,N_49072);
and UO_222 (O_222,N_49685,N_49720);
nor UO_223 (O_223,N_49637,N_49116);
or UO_224 (O_224,N_49984,N_49893);
nor UO_225 (O_225,N_49981,N_49292);
nor UO_226 (O_226,N_49439,N_49316);
nor UO_227 (O_227,N_49323,N_49135);
nand UO_228 (O_228,N_49484,N_49749);
and UO_229 (O_229,N_49176,N_49604);
or UO_230 (O_230,N_49339,N_49392);
xnor UO_231 (O_231,N_49396,N_49372);
and UO_232 (O_232,N_49845,N_49333);
or UO_233 (O_233,N_49430,N_49239);
nor UO_234 (O_234,N_49022,N_49830);
and UO_235 (O_235,N_49787,N_49633);
nand UO_236 (O_236,N_49272,N_49847);
nor UO_237 (O_237,N_49464,N_49611);
nand UO_238 (O_238,N_49712,N_49036);
nor UO_239 (O_239,N_49123,N_49975);
and UO_240 (O_240,N_49220,N_49082);
nor UO_241 (O_241,N_49686,N_49746);
nand UO_242 (O_242,N_49745,N_49898);
nor UO_243 (O_243,N_49539,N_49681);
nor UO_244 (O_244,N_49059,N_49668);
xnor UO_245 (O_245,N_49091,N_49168);
nand UO_246 (O_246,N_49544,N_49917);
nor UO_247 (O_247,N_49058,N_49524);
nand UO_248 (O_248,N_49173,N_49406);
nor UO_249 (O_249,N_49290,N_49969);
xnor UO_250 (O_250,N_49098,N_49274);
and UO_251 (O_251,N_49667,N_49842);
nor UO_252 (O_252,N_49833,N_49269);
and UO_253 (O_253,N_49706,N_49837);
or UO_254 (O_254,N_49062,N_49185);
and UO_255 (O_255,N_49622,N_49704);
xor UO_256 (O_256,N_49549,N_49580);
nand UO_257 (O_257,N_49766,N_49360);
xnor UO_258 (O_258,N_49510,N_49337);
or UO_259 (O_259,N_49482,N_49285);
nor UO_260 (O_260,N_49178,N_49927);
nor UO_261 (O_261,N_49468,N_49809);
and UO_262 (O_262,N_49816,N_49096);
nor UO_263 (O_263,N_49006,N_49980);
nor UO_264 (O_264,N_49107,N_49264);
and UO_265 (O_265,N_49714,N_49391);
nor UO_266 (O_266,N_49996,N_49697);
nor UO_267 (O_267,N_49436,N_49340);
nor UO_268 (O_268,N_49863,N_49221);
xnor UO_269 (O_269,N_49088,N_49299);
nor UO_270 (O_270,N_49532,N_49954);
nor UO_271 (O_271,N_49988,N_49756);
xnor UO_272 (O_272,N_49874,N_49541);
nand UO_273 (O_273,N_49688,N_49313);
nand UO_274 (O_274,N_49679,N_49909);
and UO_275 (O_275,N_49938,N_49362);
nand UO_276 (O_276,N_49535,N_49581);
and UO_277 (O_277,N_49421,N_49170);
xor UO_278 (O_278,N_49306,N_49550);
xor UO_279 (O_279,N_49004,N_49854);
or UO_280 (O_280,N_49151,N_49210);
xnor UO_281 (O_281,N_49839,N_49374);
or UO_282 (O_282,N_49715,N_49841);
and UO_283 (O_283,N_49138,N_49916);
nor UO_284 (O_284,N_49236,N_49931);
and UO_285 (O_285,N_49065,N_49442);
and UO_286 (O_286,N_49186,N_49806);
and UO_287 (O_287,N_49326,N_49241);
nand UO_288 (O_288,N_49522,N_49301);
or UO_289 (O_289,N_49047,N_49940);
xnor UO_290 (O_290,N_49891,N_49557);
nand UO_291 (O_291,N_49894,N_49683);
nor UO_292 (O_292,N_49709,N_49412);
nand UO_293 (O_293,N_49783,N_49869);
nor UO_294 (O_294,N_49901,N_49771);
xor UO_295 (O_295,N_49029,N_49458);
and UO_296 (O_296,N_49003,N_49693);
and UO_297 (O_297,N_49069,N_49670);
and UO_298 (O_298,N_49862,N_49090);
xnor UO_299 (O_299,N_49473,N_49015);
nor UO_300 (O_300,N_49521,N_49496);
xnor UO_301 (O_301,N_49843,N_49398);
or UO_302 (O_302,N_49218,N_49016);
nor UO_303 (O_303,N_49699,N_49645);
xnor UO_304 (O_304,N_49875,N_49188);
nand UO_305 (O_305,N_49945,N_49332);
nor UO_306 (O_306,N_49589,N_49696);
xnor UO_307 (O_307,N_49345,N_49375);
and UO_308 (O_308,N_49195,N_49500);
and UO_309 (O_309,N_49045,N_49708);
or UO_310 (O_310,N_49620,N_49807);
and UO_311 (O_311,N_49388,N_49903);
nand UO_312 (O_312,N_49564,N_49758);
xnor UO_313 (O_313,N_49381,N_49608);
or UO_314 (O_314,N_49027,N_49502);
nor UO_315 (O_315,N_49772,N_49646);
or UO_316 (O_316,N_49939,N_49676);
xor UO_317 (O_317,N_49612,N_49444);
nand UO_318 (O_318,N_49056,N_49628);
xnor UO_319 (O_319,N_49410,N_49143);
xnor UO_320 (O_320,N_49799,N_49694);
xor UO_321 (O_321,N_49254,N_49983);
or UO_322 (O_322,N_49563,N_49233);
xnor UO_323 (O_323,N_49310,N_49813);
xnor UO_324 (O_324,N_49915,N_49747);
and UO_325 (O_325,N_49124,N_49476);
nor UO_326 (O_326,N_49677,N_49329);
xnor UO_327 (O_327,N_49607,N_49897);
xor UO_328 (O_328,N_49480,N_49820);
xor UO_329 (O_329,N_49494,N_49518);
xor UO_330 (O_330,N_49508,N_49858);
xnor UO_331 (O_331,N_49205,N_49780);
or UO_332 (O_332,N_49182,N_49443);
nand UO_333 (O_333,N_49265,N_49985);
nor UO_334 (O_334,N_49416,N_49953);
and UO_335 (O_335,N_49293,N_49230);
nand UO_336 (O_336,N_49136,N_49769);
and UO_337 (O_337,N_49857,N_49849);
nand UO_338 (O_338,N_49487,N_49061);
nor UO_339 (O_339,N_49762,N_49976);
or UO_340 (O_340,N_49598,N_49774);
and UO_341 (O_341,N_49322,N_49342);
or UO_342 (O_342,N_49944,N_49020);
xor UO_343 (O_343,N_49710,N_49559);
nor UO_344 (O_344,N_49672,N_49886);
nor UO_345 (O_345,N_49417,N_49603);
and UO_346 (O_346,N_49111,N_49658);
and UO_347 (O_347,N_49609,N_49327);
nand UO_348 (O_348,N_49134,N_49592);
nand UO_349 (O_349,N_49634,N_49499);
nor UO_350 (O_350,N_49588,N_49425);
or UO_351 (O_351,N_49970,N_49341);
or UO_352 (O_352,N_49384,N_49781);
nand UO_353 (O_353,N_49190,N_49542);
nand UO_354 (O_354,N_49659,N_49311);
or UO_355 (O_355,N_49741,N_49832);
and UO_356 (O_356,N_49246,N_49353);
or UO_357 (O_357,N_49513,N_49962);
and UO_358 (O_358,N_49109,N_49545);
or UO_359 (O_359,N_49083,N_49252);
nor UO_360 (O_360,N_49361,N_49926);
xor UO_361 (O_361,N_49552,N_49501);
or UO_362 (O_362,N_49206,N_49266);
nand UO_363 (O_363,N_49623,N_49021);
and UO_364 (O_364,N_49039,N_49761);
nand UO_365 (O_365,N_49821,N_49727);
xor UO_366 (O_366,N_49081,N_49159);
and UO_367 (O_367,N_49540,N_49566);
nand UO_368 (O_368,N_49318,N_49777);
or UO_369 (O_369,N_49866,N_49335);
nor UO_370 (O_370,N_49325,N_49684);
or UO_371 (O_371,N_49179,N_49296);
nand UO_372 (O_372,N_49042,N_49601);
nor UO_373 (O_373,N_49395,N_49987);
or UO_374 (O_374,N_49046,N_49942);
xor UO_375 (O_375,N_49722,N_49394);
xor UO_376 (O_376,N_49376,N_49933);
nor UO_377 (O_377,N_49437,N_49923);
and UO_378 (O_378,N_49578,N_49702);
and UO_379 (O_379,N_49194,N_49127);
or UO_380 (O_380,N_49405,N_49895);
xor UO_381 (O_381,N_49649,N_49158);
or UO_382 (O_382,N_49475,N_49732);
or UO_383 (O_383,N_49748,N_49057);
nand UO_384 (O_384,N_49493,N_49735);
nand UO_385 (O_385,N_49558,N_49474);
xor UO_386 (O_386,N_49155,N_49014);
and UO_387 (O_387,N_49596,N_49261);
or UO_388 (O_388,N_49037,N_49831);
nand UO_389 (O_389,N_49000,N_49918);
nand UO_390 (O_390,N_49661,N_49407);
xnor UO_391 (O_391,N_49551,N_49565);
nor UO_392 (O_392,N_49125,N_49102);
xnor UO_393 (O_393,N_49811,N_49161);
or UO_394 (O_394,N_49690,N_49420);
nand UO_395 (O_395,N_49986,N_49008);
or UO_396 (O_396,N_49409,N_49073);
xnor UO_397 (O_397,N_49385,N_49122);
and UO_398 (O_398,N_49217,N_49642);
xnor UO_399 (O_399,N_49164,N_49457);
or UO_400 (O_400,N_49509,N_49053);
or UO_401 (O_401,N_49141,N_49120);
nand UO_402 (O_402,N_49142,N_49669);
nand UO_403 (O_403,N_49171,N_49228);
xor UO_404 (O_404,N_49367,N_49154);
nand UO_405 (O_405,N_49095,N_49840);
xor UO_406 (O_406,N_49812,N_49577);
nand UO_407 (O_407,N_49172,N_49922);
and UO_408 (O_408,N_49470,N_49469);
nand UO_409 (O_409,N_49085,N_49070);
or UO_410 (O_410,N_49973,N_49536);
nand UO_411 (O_411,N_49250,N_49413);
nand UO_412 (O_412,N_49166,N_49242);
nor UO_413 (O_413,N_49571,N_49025);
nor UO_414 (O_414,N_49157,N_49358);
or UO_415 (O_415,N_49859,N_49647);
or UO_416 (O_416,N_49744,N_49144);
nand UO_417 (O_417,N_49789,N_49383);
xnor UO_418 (O_418,N_49080,N_49175);
and UO_419 (O_419,N_49404,N_49515);
or UO_420 (O_420,N_49365,N_49828);
nor UO_421 (O_421,N_49453,N_49655);
nor UO_422 (O_422,N_49213,N_49929);
nand UO_423 (O_423,N_49921,N_49617);
or UO_424 (O_424,N_49705,N_49673);
and UO_425 (O_425,N_49995,N_49625);
or UO_426 (O_426,N_49818,N_49051);
nor UO_427 (O_427,N_49739,N_49007);
or UO_428 (O_428,N_49389,N_49060);
or UO_429 (O_429,N_49314,N_49139);
and UO_430 (O_430,N_49729,N_49063);
xor UO_431 (O_431,N_49947,N_49152);
and UO_432 (O_432,N_49382,N_49516);
nand UO_433 (O_433,N_49177,N_49885);
nand UO_434 (O_434,N_49462,N_49463);
nor UO_435 (O_435,N_49718,N_49447);
xnor UO_436 (O_436,N_49017,N_49256);
nand UO_437 (O_437,N_49567,N_49826);
and UO_438 (O_438,N_49108,N_49257);
or UO_439 (O_439,N_49819,N_49595);
or UO_440 (O_440,N_49137,N_49878);
nand UO_441 (O_441,N_49278,N_49280);
or UO_442 (O_442,N_49497,N_49259);
xor UO_443 (O_443,N_49309,N_49288);
or UO_444 (O_444,N_49331,N_49255);
or UO_445 (O_445,N_49146,N_49071);
nor UO_446 (O_446,N_49297,N_49763);
and UO_447 (O_447,N_49971,N_49963);
nand UO_448 (O_448,N_49547,N_49602);
xor UO_449 (O_449,N_49001,N_49232);
or UO_450 (O_450,N_49307,N_49977);
and UO_451 (O_451,N_49691,N_49629);
and UO_452 (O_452,N_49880,N_49805);
nand UO_453 (O_453,N_49671,N_49834);
and UO_454 (O_454,N_49222,N_49907);
nand UO_455 (O_455,N_49586,N_49355);
nand UO_456 (O_456,N_49861,N_49808);
nand UO_457 (O_457,N_49794,N_49426);
nor UO_458 (O_458,N_49867,N_49506);
and UO_459 (O_459,N_49638,N_49631);
nand UO_460 (O_460,N_49865,N_49225);
nor UO_461 (O_461,N_49979,N_49498);
nor UO_462 (O_462,N_49824,N_49792);
nor UO_463 (O_463,N_49207,N_49169);
and UO_464 (O_464,N_49450,N_49964);
xor UO_465 (O_465,N_49368,N_49815);
xnor UO_466 (O_466,N_49347,N_49478);
or UO_467 (O_467,N_49873,N_49446);
or UO_468 (O_468,N_49527,N_49526);
and UO_469 (O_469,N_49431,N_49678);
or UO_470 (O_470,N_49321,N_49534);
or UO_471 (O_471,N_49553,N_49010);
nor UO_472 (O_472,N_49084,N_49835);
and UO_473 (O_473,N_49505,N_49198);
nor UO_474 (O_474,N_49456,N_49846);
nand UO_475 (O_475,N_49896,N_49733);
nor UO_476 (O_476,N_49905,N_49752);
nand UO_477 (O_477,N_49271,N_49234);
nor UO_478 (O_478,N_49573,N_49957);
or UO_479 (O_479,N_49742,N_49165);
xor UO_480 (O_480,N_49990,N_49626);
nor UO_481 (O_481,N_49295,N_49209);
or UO_482 (O_482,N_49180,N_49418);
xnor UO_483 (O_483,N_49284,N_49594);
nand UO_484 (O_484,N_49555,N_49941);
xnor UO_485 (O_485,N_49032,N_49757);
and UO_486 (O_486,N_49075,N_49738);
or UO_487 (O_487,N_49925,N_49193);
nor UO_488 (O_488,N_49968,N_49751);
or UO_489 (O_489,N_49889,N_49605);
or UO_490 (O_490,N_49725,N_49899);
or UO_491 (O_491,N_49435,N_49423);
or UO_492 (O_492,N_49528,N_49753);
nand UO_493 (O_493,N_49711,N_49048);
or UO_494 (O_494,N_49801,N_49366);
xnor UO_495 (O_495,N_49660,N_49877);
or UO_496 (O_496,N_49585,N_49488);
or UO_497 (O_497,N_49089,N_49223);
and UO_498 (O_498,N_49902,N_49328);
and UO_499 (O_499,N_49900,N_49429);
or UO_500 (O_500,N_49128,N_49168);
or UO_501 (O_501,N_49450,N_49730);
or UO_502 (O_502,N_49427,N_49942);
or UO_503 (O_503,N_49431,N_49436);
or UO_504 (O_504,N_49982,N_49091);
and UO_505 (O_505,N_49432,N_49675);
xor UO_506 (O_506,N_49253,N_49955);
or UO_507 (O_507,N_49424,N_49374);
or UO_508 (O_508,N_49764,N_49263);
nand UO_509 (O_509,N_49405,N_49420);
or UO_510 (O_510,N_49168,N_49010);
and UO_511 (O_511,N_49524,N_49734);
nand UO_512 (O_512,N_49088,N_49086);
nor UO_513 (O_513,N_49833,N_49466);
and UO_514 (O_514,N_49885,N_49322);
and UO_515 (O_515,N_49242,N_49246);
nor UO_516 (O_516,N_49625,N_49437);
nand UO_517 (O_517,N_49861,N_49362);
xor UO_518 (O_518,N_49667,N_49073);
or UO_519 (O_519,N_49458,N_49920);
and UO_520 (O_520,N_49967,N_49698);
xnor UO_521 (O_521,N_49175,N_49520);
or UO_522 (O_522,N_49549,N_49907);
nand UO_523 (O_523,N_49009,N_49549);
nor UO_524 (O_524,N_49134,N_49849);
or UO_525 (O_525,N_49797,N_49611);
nor UO_526 (O_526,N_49613,N_49109);
or UO_527 (O_527,N_49403,N_49555);
nand UO_528 (O_528,N_49849,N_49119);
nor UO_529 (O_529,N_49229,N_49438);
xor UO_530 (O_530,N_49681,N_49101);
nor UO_531 (O_531,N_49730,N_49968);
nand UO_532 (O_532,N_49843,N_49112);
or UO_533 (O_533,N_49253,N_49268);
nor UO_534 (O_534,N_49744,N_49805);
xor UO_535 (O_535,N_49939,N_49977);
or UO_536 (O_536,N_49582,N_49163);
and UO_537 (O_537,N_49634,N_49755);
xnor UO_538 (O_538,N_49494,N_49637);
or UO_539 (O_539,N_49160,N_49737);
or UO_540 (O_540,N_49835,N_49312);
nor UO_541 (O_541,N_49725,N_49918);
nand UO_542 (O_542,N_49231,N_49125);
nor UO_543 (O_543,N_49272,N_49868);
nand UO_544 (O_544,N_49927,N_49210);
nor UO_545 (O_545,N_49057,N_49975);
and UO_546 (O_546,N_49881,N_49353);
xor UO_547 (O_547,N_49564,N_49275);
nand UO_548 (O_548,N_49359,N_49421);
and UO_549 (O_549,N_49426,N_49418);
and UO_550 (O_550,N_49793,N_49516);
nand UO_551 (O_551,N_49450,N_49099);
or UO_552 (O_552,N_49200,N_49532);
and UO_553 (O_553,N_49832,N_49243);
and UO_554 (O_554,N_49765,N_49876);
nor UO_555 (O_555,N_49443,N_49162);
nor UO_556 (O_556,N_49766,N_49504);
nand UO_557 (O_557,N_49199,N_49329);
and UO_558 (O_558,N_49441,N_49687);
or UO_559 (O_559,N_49970,N_49220);
or UO_560 (O_560,N_49860,N_49933);
nor UO_561 (O_561,N_49096,N_49942);
nor UO_562 (O_562,N_49317,N_49195);
or UO_563 (O_563,N_49699,N_49288);
nand UO_564 (O_564,N_49597,N_49921);
and UO_565 (O_565,N_49057,N_49924);
nor UO_566 (O_566,N_49790,N_49378);
nand UO_567 (O_567,N_49050,N_49938);
and UO_568 (O_568,N_49706,N_49811);
or UO_569 (O_569,N_49455,N_49900);
nor UO_570 (O_570,N_49326,N_49396);
nor UO_571 (O_571,N_49399,N_49564);
or UO_572 (O_572,N_49724,N_49620);
nor UO_573 (O_573,N_49450,N_49001);
nand UO_574 (O_574,N_49673,N_49297);
xor UO_575 (O_575,N_49532,N_49334);
or UO_576 (O_576,N_49339,N_49958);
nand UO_577 (O_577,N_49588,N_49744);
nor UO_578 (O_578,N_49125,N_49605);
or UO_579 (O_579,N_49548,N_49352);
nor UO_580 (O_580,N_49734,N_49257);
or UO_581 (O_581,N_49622,N_49053);
nor UO_582 (O_582,N_49357,N_49849);
nand UO_583 (O_583,N_49276,N_49469);
nor UO_584 (O_584,N_49522,N_49749);
nand UO_585 (O_585,N_49008,N_49874);
nand UO_586 (O_586,N_49125,N_49796);
xor UO_587 (O_587,N_49878,N_49731);
xor UO_588 (O_588,N_49640,N_49544);
xnor UO_589 (O_589,N_49403,N_49491);
nand UO_590 (O_590,N_49511,N_49204);
nor UO_591 (O_591,N_49867,N_49815);
nor UO_592 (O_592,N_49836,N_49123);
nand UO_593 (O_593,N_49619,N_49079);
or UO_594 (O_594,N_49827,N_49717);
nand UO_595 (O_595,N_49507,N_49619);
nor UO_596 (O_596,N_49611,N_49807);
and UO_597 (O_597,N_49860,N_49144);
xor UO_598 (O_598,N_49080,N_49307);
nand UO_599 (O_599,N_49255,N_49253);
nor UO_600 (O_600,N_49093,N_49266);
nand UO_601 (O_601,N_49194,N_49506);
xor UO_602 (O_602,N_49638,N_49673);
or UO_603 (O_603,N_49024,N_49079);
xnor UO_604 (O_604,N_49153,N_49650);
nor UO_605 (O_605,N_49220,N_49874);
xor UO_606 (O_606,N_49983,N_49678);
nor UO_607 (O_607,N_49373,N_49899);
and UO_608 (O_608,N_49026,N_49846);
and UO_609 (O_609,N_49640,N_49512);
nand UO_610 (O_610,N_49445,N_49883);
nand UO_611 (O_611,N_49177,N_49620);
nand UO_612 (O_612,N_49642,N_49236);
or UO_613 (O_613,N_49301,N_49777);
and UO_614 (O_614,N_49020,N_49934);
nor UO_615 (O_615,N_49299,N_49633);
nor UO_616 (O_616,N_49884,N_49024);
nand UO_617 (O_617,N_49192,N_49111);
xnor UO_618 (O_618,N_49584,N_49342);
and UO_619 (O_619,N_49304,N_49878);
nand UO_620 (O_620,N_49409,N_49871);
or UO_621 (O_621,N_49762,N_49559);
nand UO_622 (O_622,N_49354,N_49534);
and UO_623 (O_623,N_49723,N_49783);
and UO_624 (O_624,N_49146,N_49943);
or UO_625 (O_625,N_49857,N_49760);
nand UO_626 (O_626,N_49840,N_49749);
nand UO_627 (O_627,N_49780,N_49009);
nand UO_628 (O_628,N_49906,N_49379);
and UO_629 (O_629,N_49423,N_49191);
and UO_630 (O_630,N_49781,N_49120);
nor UO_631 (O_631,N_49796,N_49582);
or UO_632 (O_632,N_49049,N_49064);
and UO_633 (O_633,N_49576,N_49754);
nand UO_634 (O_634,N_49786,N_49693);
xor UO_635 (O_635,N_49111,N_49355);
nor UO_636 (O_636,N_49353,N_49278);
xor UO_637 (O_637,N_49114,N_49880);
nor UO_638 (O_638,N_49834,N_49397);
nand UO_639 (O_639,N_49978,N_49387);
or UO_640 (O_640,N_49506,N_49200);
and UO_641 (O_641,N_49243,N_49725);
and UO_642 (O_642,N_49684,N_49864);
xor UO_643 (O_643,N_49989,N_49122);
xnor UO_644 (O_644,N_49332,N_49360);
and UO_645 (O_645,N_49615,N_49526);
nand UO_646 (O_646,N_49512,N_49405);
nand UO_647 (O_647,N_49090,N_49483);
nor UO_648 (O_648,N_49576,N_49273);
or UO_649 (O_649,N_49642,N_49203);
xnor UO_650 (O_650,N_49908,N_49914);
and UO_651 (O_651,N_49548,N_49564);
nand UO_652 (O_652,N_49197,N_49306);
xor UO_653 (O_653,N_49276,N_49928);
nor UO_654 (O_654,N_49953,N_49441);
or UO_655 (O_655,N_49575,N_49386);
or UO_656 (O_656,N_49623,N_49343);
nand UO_657 (O_657,N_49592,N_49206);
xor UO_658 (O_658,N_49563,N_49467);
or UO_659 (O_659,N_49063,N_49417);
or UO_660 (O_660,N_49533,N_49304);
nor UO_661 (O_661,N_49580,N_49313);
and UO_662 (O_662,N_49831,N_49415);
xnor UO_663 (O_663,N_49060,N_49089);
or UO_664 (O_664,N_49527,N_49760);
nor UO_665 (O_665,N_49380,N_49381);
xnor UO_666 (O_666,N_49171,N_49397);
and UO_667 (O_667,N_49043,N_49584);
nor UO_668 (O_668,N_49835,N_49948);
xor UO_669 (O_669,N_49664,N_49396);
or UO_670 (O_670,N_49095,N_49724);
and UO_671 (O_671,N_49123,N_49278);
xnor UO_672 (O_672,N_49541,N_49425);
xor UO_673 (O_673,N_49321,N_49545);
or UO_674 (O_674,N_49562,N_49008);
xnor UO_675 (O_675,N_49249,N_49831);
xor UO_676 (O_676,N_49309,N_49544);
and UO_677 (O_677,N_49749,N_49131);
nor UO_678 (O_678,N_49553,N_49714);
nor UO_679 (O_679,N_49623,N_49863);
nor UO_680 (O_680,N_49429,N_49009);
or UO_681 (O_681,N_49203,N_49721);
and UO_682 (O_682,N_49811,N_49483);
nand UO_683 (O_683,N_49314,N_49605);
nand UO_684 (O_684,N_49533,N_49004);
nor UO_685 (O_685,N_49315,N_49624);
nand UO_686 (O_686,N_49051,N_49000);
nor UO_687 (O_687,N_49430,N_49092);
xor UO_688 (O_688,N_49150,N_49714);
xnor UO_689 (O_689,N_49339,N_49628);
xor UO_690 (O_690,N_49029,N_49841);
nor UO_691 (O_691,N_49124,N_49644);
nand UO_692 (O_692,N_49051,N_49695);
and UO_693 (O_693,N_49996,N_49541);
nor UO_694 (O_694,N_49716,N_49747);
nor UO_695 (O_695,N_49616,N_49662);
nor UO_696 (O_696,N_49359,N_49495);
and UO_697 (O_697,N_49723,N_49289);
and UO_698 (O_698,N_49229,N_49883);
nand UO_699 (O_699,N_49264,N_49345);
or UO_700 (O_700,N_49636,N_49463);
or UO_701 (O_701,N_49089,N_49518);
or UO_702 (O_702,N_49104,N_49735);
and UO_703 (O_703,N_49362,N_49623);
or UO_704 (O_704,N_49910,N_49124);
xor UO_705 (O_705,N_49886,N_49932);
nand UO_706 (O_706,N_49987,N_49537);
nor UO_707 (O_707,N_49724,N_49430);
or UO_708 (O_708,N_49690,N_49469);
xor UO_709 (O_709,N_49775,N_49108);
xor UO_710 (O_710,N_49128,N_49321);
or UO_711 (O_711,N_49970,N_49823);
or UO_712 (O_712,N_49275,N_49545);
xor UO_713 (O_713,N_49797,N_49750);
or UO_714 (O_714,N_49247,N_49375);
nor UO_715 (O_715,N_49105,N_49191);
or UO_716 (O_716,N_49090,N_49234);
nor UO_717 (O_717,N_49948,N_49714);
and UO_718 (O_718,N_49426,N_49268);
nand UO_719 (O_719,N_49130,N_49456);
and UO_720 (O_720,N_49051,N_49692);
nand UO_721 (O_721,N_49415,N_49077);
or UO_722 (O_722,N_49569,N_49201);
nor UO_723 (O_723,N_49264,N_49814);
xnor UO_724 (O_724,N_49275,N_49696);
xor UO_725 (O_725,N_49702,N_49670);
or UO_726 (O_726,N_49427,N_49948);
or UO_727 (O_727,N_49799,N_49520);
or UO_728 (O_728,N_49461,N_49053);
xnor UO_729 (O_729,N_49160,N_49654);
or UO_730 (O_730,N_49396,N_49506);
xor UO_731 (O_731,N_49832,N_49103);
nand UO_732 (O_732,N_49748,N_49555);
nand UO_733 (O_733,N_49391,N_49437);
nand UO_734 (O_734,N_49078,N_49837);
or UO_735 (O_735,N_49733,N_49109);
nand UO_736 (O_736,N_49589,N_49543);
and UO_737 (O_737,N_49650,N_49917);
xor UO_738 (O_738,N_49409,N_49200);
xor UO_739 (O_739,N_49798,N_49103);
or UO_740 (O_740,N_49450,N_49146);
and UO_741 (O_741,N_49709,N_49878);
and UO_742 (O_742,N_49248,N_49222);
or UO_743 (O_743,N_49605,N_49347);
and UO_744 (O_744,N_49699,N_49723);
xor UO_745 (O_745,N_49163,N_49523);
and UO_746 (O_746,N_49599,N_49111);
nand UO_747 (O_747,N_49458,N_49250);
nor UO_748 (O_748,N_49645,N_49745);
nor UO_749 (O_749,N_49935,N_49043);
and UO_750 (O_750,N_49029,N_49862);
nand UO_751 (O_751,N_49585,N_49480);
nor UO_752 (O_752,N_49231,N_49001);
nand UO_753 (O_753,N_49486,N_49907);
and UO_754 (O_754,N_49309,N_49294);
nor UO_755 (O_755,N_49643,N_49809);
nor UO_756 (O_756,N_49839,N_49913);
or UO_757 (O_757,N_49134,N_49987);
or UO_758 (O_758,N_49086,N_49178);
or UO_759 (O_759,N_49565,N_49842);
and UO_760 (O_760,N_49361,N_49800);
xor UO_761 (O_761,N_49229,N_49730);
nand UO_762 (O_762,N_49320,N_49567);
or UO_763 (O_763,N_49687,N_49458);
or UO_764 (O_764,N_49174,N_49661);
nand UO_765 (O_765,N_49513,N_49426);
or UO_766 (O_766,N_49337,N_49944);
or UO_767 (O_767,N_49955,N_49639);
nand UO_768 (O_768,N_49399,N_49092);
xor UO_769 (O_769,N_49373,N_49737);
or UO_770 (O_770,N_49632,N_49316);
or UO_771 (O_771,N_49612,N_49558);
and UO_772 (O_772,N_49539,N_49678);
xor UO_773 (O_773,N_49296,N_49709);
or UO_774 (O_774,N_49123,N_49372);
and UO_775 (O_775,N_49379,N_49131);
xor UO_776 (O_776,N_49148,N_49399);
and UO_777 (O_777,N_49525,N_49286);
or UO_778 (O_778,N_49030,N_49676);
and UO_779 (O_779,N_49609,N_49847);
xnor UO_780 (O_780,N_49225,N_49449);
and UO_781 (O_781,N_49106,N_49292);
xor UO_782 (O_782,N_49012,N_49897);
or UO_783 (O_783,N_49448,N_49061);
nand UO_784 (O_784,N_49015,N_49197);
nor UO_785 (O_785,N_49221,N_49878);
nor UO_786 (O_786,N_49148,N_49075);
and UO_787 (O_787,N_49185,N_49292);
nand UO_788 (O_788,N_49936,N_49220);
or UO_789 (O_789,N_49720,N_49747);
or UO_790 (O_790,N_49779,N_49740);
nor UO_791 (O_791,N_49794,N_49648);
nand UO_792 (O_792,N_49159,N_49905);
nand UO_793 (O_793,N_49628,N_49843);
nand UO_794 (O_794,N_49583,N_49947);
nor UO_795 (O_795,N_49701,N_49889);
and UO_796 (O_796,N_49915,N_49556);
xnor UO_797 (O_797,N_49408,N_49984);
xor UO_798 (O_798,N_49441,N_49657);
nor UO_799 (O_799,N_49605,N_49111);
or UO_800 (O_800,N_49762,N_49412);
xor UO_801 (O_801,N_49352,N_49538);
or UO_802 (O_802,N_49788,N_49833);
xnor UO_803 (O_803,N_49296,N_49551);
nand UO_804 (O_804,N_49376,N_49055);
nand UO_805 (O_805,N_49213,N_49666);
and UO_806 (O_806,N_49283,N_49903);
nor UO_807 (O_807,N_49727,N_49800);
xnor UO_808 (O_808,N_49289,N_49453);
or UO_809 (O_809,N_49160,N_49168);
and UO_810 (O_810,N_49395,N_49075);
or UO_811 (O_811,N_49738,N_49246);
and UO_812 (O_812,N_49025,N_49736);
or UO_813 (O_813,N_49027,N_49706);
xor UO_814 (O_814,N_49160,N_49632);
and UO_815 (O_815,N_49598,N_49299);
nor UO_816 (O_816,N_49486,N_49901);
or UO_817 (O_817,N_49900,N_49542);
or UO_818 (O_818,N_49975,N_49879);
xnor UO_819 (O_819,N_49171,N_49099);
nand UO_820 (O_820,N_49681,N_49083);
or UO_821 (O_821,N_49999,N_49258);
or UO_822 (O_822,N_49694,N_49767);
nor UO_823 (O_823,N_49310,N_49951);
and UO_824 (O_824,N_49540,N_49811);
or UO_825 (O_825,N_49504,N_49454);
nand UO_826 (O_826,N_49535,N_49988);
or UO_827 (O_827,N_49943,N_49428);
or UO_828 (O_828,N_49213,N_49164);
and UO_829 (O_829,N_49077,N_49218);
nor UO_830 (O_830,N_49212,N_49387);
xor UO_831 (O_831,N_49295,N_49134);
xor UO_832 (O_832,N_49652,N_49956);
and UO_833 (O_833,N_49887,N_49250);
and UO_834 (O_834,N_49590,N_49607);
nand UO_835 (O_835,N_49497,N_49793);
nand UO_836 (O_836,N_49360,N_49847);
and UO_837 (O_837,N_49222,N_49708);
nor UO_838 (O_838,N_49621,N_49935);
nor UO_839 (O_839,N_49455,N_49674);
xor UO_840 (O_840,N_49574,N_49007);
nand UO_841 (O_841,N_49331,N_49128);
nand UO_842 (O_842,N_49939,N_49603);
or UO_843 (O_843,N_49724,N_49090);
and UO_844 (O_844,N_49952,N_49860);
and UO_845 (O_845,N_49107,N_49524);
nor UO_846 (O_846,N_49885,N_49231);
or UO_847 (O_847,N_49442,N_49512);
nand UO_848 (O_848,N_49002,N_49338);
nand UO_849 (O_849,N_49912,N_49962);
and UO_850 (O_850,N_49215,N_49457);
or UO_851 (O_851,N_49187,N_49242);
nand UO_852 (O_852,N_49581,N_49923);
and UO_853 (O_853,N_49951,N_49033);
and UO_854 (O_854,N_49178,N_49400);
and UO_855 (O_855,N_49813,N_49449);
xor UO_856 (O_856,N_49921,N_49258);
and UO_857 (O_857,N_49337,N_49113);
nand UO_858 (O_858,N_49204,N_49715);
and UO_859 (O_859,N_49238,N_49702);
nor UO_860 (O_860,N_49290,N_49990);
xor UO_861 (O_861,N_49191,N_49098);
and UO_862 (O_862,N_49730,N_49493);
or UO_863 (O_863,N_49498,N_49561);
or UO_864 (O_864,N_49598,N_49561);
nand UO_865 (O_865,N_49920,N_49621);
xnor UO_866 (O_866,N_49168,N_49772);
nor UO_867 (O_867,N_49698,N_49736);
or UO_868 (O_868,N_49305,N_49364);
nor UO_869 (O_869,N_49985,N_49085);
and UO_870 (O_870,N_49056,N_49850);
or UO_871 (O_871,N_49177,N_49831);
and UO_872 (O_872,N_49770,N_49432);
nand UO_873 (O_873,N_49388,N_49230);
xnor UO_874 (O_874,N_49888,N_49210);
or UO_875 (O_875,N_49531,N_49801);
and UO_876 (O_876,N_49676,N_49719);
xnor UO_877 (O_877,N_49733,N_49197);
and UO_878 (O_878,N_49649,N_49990);
or UO_879 (O_879,N_49408,N_49450);
and UO_880 (O_880,N_49645,N_49555);
nor UO_881 (O_881,N_49799,N_49215);
or UO_882 (O_882,N_49936,N_49064);
nand UO_883 (O_883,N_49196,N_49401);
and UO_884 (O_884,N_49245,N_49191);
xor UO_885 (O_885,N_49763,N_49224);
xor UO_886 (O_886,N_49033,N_49263);
nand UO_887 (O_887,N_49950,N_49707);
or UO_888 (O_888,N_49862,N_49120);
nand UO_889 (O_889,N_49555,N_49743);
and UO_890 (O_890,N_49231,N_49482);
nor UO_891 (O_891,N_49983,N_49969);
nand UO_892 (O_892,N_49107,N_49379);
nand UO_893 (O_893,N_49641,N_49771);
and UO_894 (O_894,N_49421,N_49600);
nor UO_895 (O_895,N_49118,N_49269);
nand UO_896 (O_896,N_49471,N_49431);
nand UO_897 (O_897,N_49055,N_49925);
nor UO_898 (O_898,N_49526,N_49764);
and UO_899 (O_899,N_49259,N_49525);
and UO_900 (O_900,N_49859,N_49128);
nor UO_901 (O_901,N_49400,N_49608);
or UO_902 (O_902,N_49043,N_49581);
nor UO_903 (O_903,N_49174,N_49158);
xor UO_904 (O_904,N_49929,N_49356);
nand UO_905 (O_905,N_49859,N_49578);
nand UO_906 (O_906,N_49002,N_49341);
or UO_907 (O_907,N_49006,N_49022);
or UO_908 (O_908,N_49848,N_49857);
or UO_909 (O_909,N_49393,N_49283);
nor UO_910 (O_910,N_49166,N_49516);
or UO_911 (O_911,N_49290,N_49368);
or UO_912 (O_912,N_49730,N_49540);
xnor UO_913 (O_913,N_49876,N_49136);
xnor UO_914 (O_914,N_49957,N_49398);
and UO_915 (O_915,N_49392,N_49645);
and UO_916 (O_916,N_49975,N_49482);
nor UO_917 (O_917,N_49856,N_49994);
and UO_918 (O_918,N_49457,N_49046);
or UO_919 (O_919,N_49384,N_49099);
nor UO_920 (O_920,N_49356,N_49646);
nor UO_921 (O_921,N_49346,N_49422);
nor UO_922 (O_922,N_49248,N_49287);
and UO_923 (O_923,N_49731,N_49171);
and UO_924 (O_924,N_49997,N_49569);
and UO_925 (O_925,N_49702,N_49106);
nor UO_926 (O_926,N_49906,N_49991);
and UO_927 (O_927,N_49955,N_49789);
nor UO_928 (O_928,N_49526,N_49433);
xnor UO_929 (O_929,N_49516,N_49623);
and UO_930 (O_930,N_49451,N_49986);
nor UO_931 (O_931,N_49465,N_49236);
or UO_932 (O_932,N_49795,N_49868);
nand UO_933 (O_933,N_49659,N_49837);
nor UO_934 (O_934,N_49221,N_49809);
or UO_935 (O_935,N_49111,N_49031);
xor UO_936 (O_936,N_49243,N_49507);
xor UO_937 (O_937,N_49066,N_49104);
and UO_938 (O_938,N_49254,N_49372);
nand UO_939 (O_939,N_49908,N_49804);
nand UO_940 (O_940,N_49778,N_49308);
nand UO_941 (O_941,N_49359,N_49494);
or UO_942 (O_942,N_49225,N_49437);
nor UO_943 (O_943,N_49777,N_49312);
or UO_944 (O_944,N_49738,N_49805);
nor UO_945 (O_945,N_49439,N_49385);
and UO_946 (O_946,N_49596,N_49056);
nor UO_947 (O_947,N_49522,N_49172);
and UO_948 (O_948,N_49757,N_49030);
or UO_949 (O_949,N_49261,N_49416);
nand UO_950 (O_950,N_49464,N_49873);
and UO_951 (O_951,N_49193,N_49858);
nor UO_952 (O_952,N_49685,N_49775);
nor UO_953 (O_953,N_49816,N_49936);
xor UO_954 (O_954,N_49400,N_49055);
nor UO_955 (O_955,N_49961,N_49970);
nor UO_956 (O_956,N_49041,N_49013);
xor UO_957 (O_957,N_49910,N_49282);
and UO_958 (O_958,N_49643,N_49857);
and UO_959 (O_959,N_49967,N_49800);
nand UO_960 (O_960,N_49571,N_49731);
nand UO_961 (O_961,N_49958,N_49865);
xnor UO_962 (O_962,N_49928,N_49442);
xor UO_963 (O_963,N_49483,N_49898);
or UO_964 (O_964,N_49781,N_49678);
xor UO_965 (O_965,N_49483,N_49985);
nor UO_966 (O_966,N_49857,N_49171);
nand UO_967 (O_967,N_49064,N_49671);
nand UO_968 (O_968,N_49074,N_49481);
xor UO_969 (O_969,N_49703,N_49814);
xor UO_970 (O_970,N_49819,N_49115);
and UO_971 (O_971,N_49941,N_49559);
nor UO_972 (O_972,N_49850,N_49531);
nand UO_973 (O_973,N_49664,N_49740);
and UO_974 (O_974,N_49164,N_49809);
nand UO_975 (O_975,N_49067,N_49219);
xnor UO_976 (O_976,N_49701,N_49217);
nand UO_977 (O_977,N_49048,N_49084);
and UO_978 (O_978,N_49640,N_49718);
nand UO_979 (O_979,N_49699,N_49956);
nor UO_980 (O_980,N_49789,N_49538);
and UO_981 (O_981,N_49086,N_49564);
xnor UO_982 (O_982,N_49926,N_49145);
xnor UO_983 (O_983,N_49183,N_49996);
xnor UO_984 (O_984,N_49800,N_49021);
or UO_985 (O_985,N_49393,N_49338);
nor UO_986 (O_986,N_49375,N_49272);
nor UO_987 (O_987,N_49873,N_49266);
or UO_988 (O_988,N_49023,N_49511);
nor UO_989 (O_989,N_49776,N_49109);
nand UO_990 (O_990,N_49644,N_49089);
or UO_991 (O_991,N_49541,N_49895);
nor UO_992 (O_992,N_49178,N_49871);
or UO_993 (O_993,N_49018,N_49823);
nor UO_994 (O_994,N_49657,N_49356);
nand UO_995 (O_995,N_49362,N_49952);
and UO_996 (O_996,N_49012,N_49249);
xnor UO_997 (O_997,N_49982,N_49634);
xor UO_998 (O_998,N_49139,N_49208);
nor UO_999 (O_999,N_49399,N_49047);
or UO_1000 (O_1000,N_49193,N_49170);
and UO_1001 (O_1001,N_49487,N_49489);
and UO_1002 (O_1002,N_49636,N_49831);
or UO_1003 (O_1003,N_49069,N_49293);
and UO_1004 (O_1004,N_49226,N_49805);
nor UO_1005 (O_1005,N_49183,N_49024);
nand UO_1006 (O_1006,N_49942,N_49575);
and UO_1007 (O_1007,N_49654,N_49676);
xor UO_1008 (O_1008,N_49429,N_49882);
nand UO_1009 (O_1009,N_49431,N_49011);
or UO_1010 (O_1010,N_49739,N_49979);
nor UO_1011 (O_1011,N_49277,N_49216);
or UO_1012 (O_1012,N_49021,N_49554);
nand UO_1013 (O_1013,N_49203,N_49447);
nand UO_1014 (O_1014,N_49004,N_49334);
nor UO_1015 (O_1015,N_49739,N_49501);
nor UO_1016 (O_1016,N_49659,N_49461);
and UO_1017 (O_1017,N_49086,N_49082);
nor UO_1018 (O_1018,N_49174,N_49220);
or UO_1019 (O_1019,N_49981,N_49803);
and UO_1020 (O_1020,N_49233,N_49772);
or UO_1021 (O_1021,N_49229,N_49743);
or UO_1022 (O_1022,N_49788,N_49630);
and UO_1023 (O_1023,N_49092,N_49801);
or UO_1024 (O_1024,N_49487,N_49671);
nor UO_1025 (O_1025,N_49417,N_49655);
or UO_1026 (O_1026,N_49665,N_49943);
nand UO_1027 (O_1027,N_49907,N_49541);
and UO_1028 (O_1028,N_49239,N_49506);
xor UO_1029 (O_1029,N_49871,N_49564);
xor UO_1030 (O_1030,N_49671,N_49825);
and UO_1031 (O_1031,N_49159,N_49046);
and UO_1032 (O_1032,N_49291,N_49071);
xor UO_1033 (O_1033,N_49292,N_49174);
and UO_1034 (O_1034,N_49845,N_49521);
or UO_1035 (O_1035,N_49021,N_49388);
or UO_1036 (O_1036,N_49850,N_49260);
and UO_1037 (O_1037,N_49648,N_49720);
nand UO_1038 (O_1038,N_49404,N_49903);
and UO_1039 (O_1039,N_49050,N_49127);
or UO_1040 (O_1040,N_49853,N_49703);
or UO_1041 (O_1041,N_49278,N_49460);
nand UO_1042 (O_1042,N_49134,N_49613);
or UO_1043 (O_1043,N_49062,N_49060);
and UO_1044 (O_1044,N_49002,N_49829);
or UO_1045 (O_1045,N_49939,N_49132);
nand UO_1046 (O_1046,N_49606,N_49147);
nand UO_1047 (O_1047,N_49771,N_49097);
nand UO_1048 (O_1048,N_49241,N_49792);
nand UO_1049 (O_1049,N_49149,N_49915);
nand UO_1050 (O_1050,N_49310,N_49509);
or UO_1051 (O_1051,N_49203,N_49347);
and UO_1052 (O_1052,N_49145,N_49411);
xnor UO_1053 (O_1053,N_49296,N_49661);
or UO_1054 (O_1054,N_49270,N_49857);
nor UO_1055 (O_1055,N_49583,N_49612);
xnor UO_1056 (O_1056,N_49357,N_49020);
nand UO_1057 (O_1057,N_49859,N_49976);
xnor UO_1058 (O_1058,N_49777,N_49235);
nand UO_1059 (O_1059,N_49058,N_49326);
and UO_1060 (O_1060,N_49553,N_49864);
xnor UO_1061 (O_1061,N_49647,N_49089);
or UO_1062 (O_1062,N_49613,N_49097);
nand UO_1063 (O_1063,N_49141,N_49210);
and UO_1064 (O_1064,N_49072,N_49069);
nand UO_1065 (O_1065,N_49788,N_49155);
or UO_1066 (O_1066,N_49913,N_49200);
and UO_1067 (O_1067,N_49621,N_49016);
nand UO_1068 (O_1068,N_49259,N_49462);
nor UO_1069 (O_1069,N_49013,N_49191);
nand UO_1070 (O_1070,N_49795,N_49840);
nand UO_1071 (O_1071,N_49555,N_49031);
xor UO_1072 (O_1072,N_49569,N_49328);
or UO_1073 (O_1073,N_49684,N_49617);
or UO_1074 (O_1074,N_49330,N_49394);
xnor UO_1075 (O_1075,N_49203,N_49908);
or UO_1076 (O_1076,N_49160,N_49790);
nor UO_1077 (O_1077,N_49183,N_49046);
and UO_1078 (O_1078,N_49893,N_49834);
and UO_1079 (O_1079,N_49371,N_49400);
xnor UO_1080 (O_1080,N_49595,N_49329);
and UO_1081 (O_1081,N_49189,N_49666);
or UO_1082 (O_1082,N_49318,N_49426);
nor UO_1083 (O_1083,N_49494,N_49005);
xor UO_1084 (O_1084,N_49246,N_49352);
nand UO_1085 (O_1085,N_49086,N_49612);
nor UO_1086 (O_1086,N_49580,N_49865);
nor UO_1087 (O_1087,N_49510,N_49300);
nor UO_1088 (O_1088,N_49144,N_49639);
nor UO_1089 (O_1089,N_49477,N_49467);
or UO_1090 (O_1090,N_49205,N_49427);
nor UO_1091 (O_1091,N_49557,N_49860);
nand UO_1092 (O_1092,N_49351,N_49888);
xor UO_1093 (O_1093,N_49083,N_49910);
nand UO_1094 (O_1094,N_49440,N_49126);
nor UO_1095 (O_1095,N_49637,N_49172);
xor UO_1096 (O_1096,N_49063,N_49513);
xnor UO_1097 (O_1097,N_49588,N_49656);
nand UO_1098 (O_1098,N_49659,N_49247);
xor UO_1099 (O_1099,N_49786,N_49394);
nand UO_1100 (O_1100,N_49814,N_49391);
nor UO_1101 (O_1101,N_49413,N_49264);
nand UO_1102 (O_1102,N_49202,N_49841);
xnor UO_1103 (O_1103,N_49654,N_49968);
and UO_1104 (O_1104,N_49498,N_49495);
and UO_1105 (O_1105,N_49052,N_49161);
or UO_1106 (O_1106,N_49714,N_49378);
xnor UO_1107 (O_1107,N_49398,N_49095);
and UO_1108 (O_1108,N_49814,N_49754);
nand UO_1109 (O_1109,N_49063,N_49272);
nor UO_1110 (O_1110,N_49070,N_49461);
nand UO_1111 (O_1111,N_49189,N_49080);
nand UO_1112 (O_1112,N_49577,N_49861);
nor UO_1113 (O_1113,N_49938,N_49574);
and UO_1114 (O_1114,N_49364,N_49096);
nor UO_1115 (O_1115,N_49020,N_49780);
nor UO_1116 (O_1116,N_49144,N_49260);
and UO_1117 (O_1117,N_49650,N_49665);
nor UO_1118 (O_1118,N_49339,N_49754);
xnor UO_1119 (O_1119,N_49688,N_49553);
nor UO_1120 (O_1120,N_49366,N_49311);
nor UO_1121 (O_1121,N_49657,N_49699);
nand UO_1122 (O_1122,N_49135,N_49156);
xnor UO_1123 (O_1123,N_49988,N_49971);
nand UO_1124 (O_1124,N_49282,N_49010);
and UO_1125 (O_1125,N_49880,N_49623);
xor UO_1126 (O_1126,N_49209,N_49764);
nor UO_1127 (O_1127,N_49182,N_49352);
xnor UO_1128 (O_1128,N_49855,N_49388);
nor UO_1129 (O_1129,N_49364,N_49139);
xor UO_1130 (O_1130,N_49343,N_49770);
or UO_1131 (O_1131,N_49216,N_49997);
and UO_1132 (O_1132,N_49301,N_49045);
nor UO_1133 (O_1133,N_49362,N_49490);
or UO_1134 (O_1134,N_49873,N_49792);
nand UO_1135 (O_1135,N_49816,N_49314);
nor UO_1136 (O_1136,N_49089,N_49173);
nand UO_1137 (O_1137,N_49129,N_49370);
or UO_1138 (O_1138,N_49800,N_49169);
and UO_1139 (O_1139,N_49464,N_49953);
xnor UO_1140 (O_1140,N_49345,N_49917);
nand UO_1141 (O_1141,N_49131,N_49378);
nand UO_1142 (O_1142,N_49960,N_49312);
and UO_1143 (O_1143,N_49210,N_49439);
nor UO_1144 (O_1144,N_49032,N_49920);
nand UO_1145 (O_1145,N_49759,N_49325);
nor UO_1146 (O_1146,N_49529,N_49932);
nor UO_1147 (O_1147,N_49926,N_49020);
nand UO_1148 (O_1148,N_49481,N_49913);
and UO_1149 (O_1149,N_49711,N_49219);
nor UO_1150 (O_1150,N_49168,N_49012);
or UO_1151 (O_1151,N_49780,N_49916);
nand UO_1152 (O_1152,N_49740,N_49299);
or UO_1153 (O_1153,N_49700,N_49722);
nor UO_1154 (O_1154,N_49937,N_49303);
nand UO_1155 (O_1155,N_49937,N_49979);
and UO_1156 (O_1156,N_49983,N_49258);
nor UO_1157 (O_1157,N_49315,N_49111);
xnor UO_1158 (O_1158,N_49819,N_49333);
or UO_1159 (O_1159,N_49587,N_49183);
xnor UO_1160 (O_1160,N_49617,N_49901);
nor UO_1161 (O_1161,N_49768,N_49817);
nor UO_1162 (O_1162,N_49091,N_49993);
nor UO_1163 (O_1163,N_49586,N_49059);
xor UO_1164 (O_1164,N_49722,N_49377);
and UO_1165 (O_1165,N_49157,N_49869);
or UO_1166 (O_1166,N_49175,N_49984);
xor UO_1167 (O_1167,N_49174,N_49025);
nand UO_1168 (O_1168,N_49797,N_49516);
xnor UO_1169 (O_1169,N_49028,N_49178);
or UO_1170 (O_1170,N_49961,N_49131);
and UO_1171 (O_1171,N_49048,N_49420);
nor UO_1172 (O_1172,N_49850,N_49171);
and UO_1173 (O_1173,N_49650,N_49349);
xor UO_1174 (O_1174,N_49178,N_49370);
and UO_1175 (O_1175,N_49460,N_49056);
nand UO_1176 (O_1176,N_49413,N_49762);
nor UO_1177 (O_1177,N_49237,N_49238);
nand UO_1178 (O_1178,N_49818,N_49614);
xnor UO_1179 (O_1179,N_49249,N_49143);
nand UO_1180 (O_1180,N_49508,N_49115);
nor UO_1181 (O_1181,N_49739,N_49152);
nor UO_1182 (O_1182,N_49423,N_49646);
nor UO_1183 (O_1183,N_49651,N_49888);
or UO_1184 (O_1184,N_49342,N_49047);
nand UO_1185 (O_1185,N_49255,N_49744);
nor UO_1186 (O_1186,N_49289,N_49469);
or UO_1187 (O_1187,N_49281,N_49301);
and UO_1188 (O_1188,N_49167,N_49625);
nand UO_1189 (O_1189,N_49121,N_49977);
xor UO_1190 (O_1190,N_49228,N_49349);
xor UO_1191 (O_1191,N_49411,N_49225);
and UO_1192 (O_1192,N_49414,N_49171);
nor UO_1193 (O_1193,N_49923,N_49419);
nand UO_1194 (O_1194,N_49681,N_49547);
and UO_1195 (O_1195,N_49035,N_49033);
xor UO_1196 (O_1196,N_49915,N_49159);
xnor UO_1197 (O_1197,N_49743,N_49808);
and UO_1198 (O_1198,N_49062,N_49239);
nand UO_1199 (O_1199,N_49237,N_49234);
or UO_1200 (O_1200,N_49882,N_49957);
or UO_1201 (O_1201,N_49088,N_49583);
nand UO_1202 (O_1202,N_49501,N_49284);
nand UO_1203 (O_1203,N_49393,N_49022);
xnor UO_1204 (O_1204,N_49170,N_49998);
or UO_1205 (O_1205,N_49907,N_49699);
or UO_1206 (O_1206,N_49177,N_49333);
and UO_1207 (O_1207,N_49349,N_49365);
nand UO_1208 (O_1208,N_49636,N_49747);
and UO_1209 (O_1209,N_49880,N_49961);
nor UO_1210 (O_1210,N_49129,N_49135);
and UO_1211 (O_1211,N_49127,N_49263);
or UO_1212 (O_1212,N_49846,N_49704);
or UO_1213 (O_1213,N_49763,N_49418);
xor UO_1214 (O_1214,N_49557,N_49892);
or UO_1215 (O_1215,N_49278,N_49566);
and UO_1216 (O_1216,N_49709,N_49693);
nor UO_1217 (O_1217,N_49170,N_49601);
nand UO_1218 (O_1218,N_49268,N_49923);
nor UO_1219 (O_1219,N_49761,N_49100);
xnor UO_1220 (O_1220,N_49814,N_49424);
nand UO_1221 (O_1221,N_49065,N_49370);
nand UO_1222 (O_1222,N_49317,N_49214);
xor UO_1223 (O_1223,N_49068,N_49117);
nor UO_1224 (O_1224,N_49438,N_49443);
nand UO_1225 (O_1225,N_49401,N_49436);
nand UO_1226 (O_1226,N_49495,N_49775);
and UO_1227 (O_1227,N_49328,N_49378);
or UO_1228 (O_1228,N_49082,N_49818);
nand UO_1229 (O_1229,N_49138,N_49796);
and UO_1230 (O_1230,N_49410,N_49358);
xor UO_1231 (O_1231,N_49546,N_49860);
xnor UO_1232 (O_1232,N_49098,N_49998);
xnor UO_1233 (O_1233,N_49831,N_49423);
or UO_1234 (O_1234,N_49722,N_49708);
nand UO_1235 (O_1235,N_49844,N_49202);
xnor UO_1236 (O_1236,N_49595,N_49237);
and UO_1237 (O_1237,N_49214,N_49292);
and UO_1238 (O_1238,N_49663,N_49331);
nor UO_1239 (O_1239,N_49375,N_49393);
or UO_1240 (O_1240,N_49173,N_49376);
and UO_1241 (O_1241,N_49479,N_49464);
nand UO_1242 (O_1242,N_49513,N_49079);
nor UO_1243 (O_1243,N_49895,N_49176);
nor UO_1244 (O_1244,N_49497,N_49656);
or UO_1245 (O_1245,N_49457,N_49910);
and UO_1246 (O_1246,N_49046,N_49507);
nand UO_1247 (O_1247,N_49652,N_49261);
and UO_1248 (O_1248,N_49094,N_49345);
nor UO_1249 (O_1249,N_49906,N_49683);
or UO_1250 (O_1250,N_49275,N_49668);
and UO_1251 (O_1251,N_49482,N_49594);
xnor UO_1252 (O_1252,N_49156,N_49942);
or UO_1253 (O_1253,N_49631,N_49426);
nand UO_1254 (O_1254,N_49088,N_49441);
nand UO_1255 (O_1255,N_49390,N_49864);
nand UO_1256 (O_1256,N_49461,N_49674);
and UO_1257 (O_1257,N_49246,N_49711);
or UO_1258 (O_1258,N_49590,N_49818);
or UO_1259 (O_1259,N_49330,N_49475);
xor UO_1260 (O_1260,N_49583,N_49630);
and UO_1261 (O_1261,N_49023,N_49194);
nand UO_1262 (O_1262,N_49164,N_49284);
and UO_1263 (O_1263,N_49182,N_49642);
nor UO_1264 (O_1264,N_49861,N_49605);
and UO_1265 (O_1265,N_49124,N_49701);
nor UO_1266 (O_1266,N_49069,N_49709);
or UO_1267 (O_1267,N_49452,N_49862);
and UO_1268 (O_1268,N_49814,N_49024);
nor UO_1269 (O_1269,N_49697,N_49006);
xnor UO_1270 (O_1270,N_49645,N_49230);
xor UO_1271 (O_1271,N_49961,N_49492);
nand UO_1272 (O_1272,N_49277,N_49119);
and UO_1273 (O_1273,N_49916,N_49429);
nor UO_1274 (O_1274,N_49377,N_49224);
and UO_1275 (O_1275,N_49658,N_49775);
or UO_1276 (O_1276,N_49665,N_49280);
or UO_1277 (O_1277,N_49946,N_49462);
or UO_1278 (O_1278,N_49155,N_49026);
or UO_1279 (O_1279,N_49347,N_49262);
xnor UO_1280 (O_1280,N_49557,N_49035);
and UO_1281 (O_1281,N_49272,N_49139);
and UO_1282 (O_1282,N_49956,N_49992);
and UO_1283 (O_1283,N_49195,N_49567);
or UO_1284 (O_1284,N_49809,N_49906);
and UO_1285 (O_1285,N_49256,N_49791);
and UO_1286 (O_1286,N_49763,N_49589);
and UO_1287 (O_1287,N_49163,N_49164);
nor UO_1288 (O_1288,N_49944,N_49418);
or UO_1289 (O_1289,N_49873,N_49584);
nor UO_1290 (O_1290,N_49899,N_49204);
nor UO_1291 (O_1291,N_49232,N_49184);
or UO_1292 (O_1292,N_49382,N_49906);
nor UO_1293 (O_1293,N_49047,N_49703);
xnor UO_1294 (O_1294,N_49052,N_49532);
and UO_1295 (O_1295,N_49463,N_49094);
nor UO_1296 (O_1296,N_49419,N_49938);
and UO_1297 (O_1297,N_49529,N_49628);
xnor UO_1298 (O_1298,N_49982,N_49449);
nand UO_1299 (O_1299,N_49358,N_49711);
nor UO_1300 (O_1300,N_49610,N_49630);
nand UO_1301 (O_1301,N_49585,N_49475);
or UO_1302 (O_1302,N_49274,N_49574);
and UO_1303 (O_1303,N_49812,N_49874);
nor UO_1304 (O_1304,N_49684,N_49715);
nor UO_1305 (O_1305,N_49929,N_49741);
xnor UO_1306 (O_1306,N_49654,N_49396);
xor UO_1307 (O_1307,N_49830,N_49411);
nor UO_1308 (O_1308,N_49660,N_49760);
or UO_1309 (O_1309,N_49040,N_49619);
nand UO_1310 (O_1310,N_49257,N_49519);
or UO_1311 (O_1311,N_49550,N_49277);
or UO_1312 (O_1312,N_49982,N_49509);
xnor UO_1313 (O_1313,N_49341,N_49312);
nor UO_1314 (O_1314,N_49351,N_49341);
xor UO_1315 (O_1315,N_49304,N_49815);
and UO_1316 (O_1316,N_49827,N_49640);
or UO_1317 (O_1317,N_49234,N_49229);
or UO_1318 (O_1318,N_49197,N_49889);
and UO_1319 (O_1319,N_49717,N_49913);
nor UO_1320 (O_1320,N_49935,N_49472);
nand UO_1321 (O_1321,N_49850,N_49819);
and UO_1322 (O_1322,N_49862,N_49326);
xnor UO_1323 (O_1323,N_49811,N_49178);
nor UO_1324 (O_1324,N_49516,N_49250);
or UO_1325 (O_1325,N_49287,N_49566);
xor UO_1326 (O_1326,N_49032,N_49185);
or UO_1327 (O_1327,N_49260,N_49614);
nand UO_1328 (O_1328,N_49685,N_49047);
and UO_1329 (O_1329,N_49341,N_49335);
nor UO_1330 (O_1330,N_49486,N_49293);
and UO_1331 (O_1331,N_49978,N_49795);
nor UO_1332 (O_1332,N_49668,N_49140);
and UO_1333 (O_1333,N_49463,N_49156);
and UO_1334 (O_1334,N_49264,N_49036);
xnor UO_1335 (O_1335,N_49434,N_49756);
and UO_1336 (O_1336,N_49545,N_49148);
and UO_1337 (O_1337,N_49547,N_49577);
or UO_1338 (O_1338,N_49970,N_49240);
nand UO_1339 (O_1339,N_49343,N_49414);
nor UO_1340 (O_1340,N_49005,N_49169);
and UO_1341 (O_1341,N_49022,N_49175);
nand UO_1342 (O_1342,N_49181,N_49025);
and UO_1343 (O_1343,N_49213,N_49015);
nor UO_1344 (O_1344,N_49625,N_49715);
xnor UO_1345 (O_1345,N_49558,N_49573);
nor UO_1346 (O_1346,N_49047,N_49930);
xnor UO_1347 (O_1347,N_49108,N_49252);
xnor UO_1348 (O_1348,N_49839,N_49773);
or UO_1349 (O_1349,N_49285,N_49068);
xnor UO_1350 (O_1350,N_49509,N_49631);
nor UO_1351 (O_1351,N_49418,N_49295);
xor UO_1352 (O_1352,N_49443,N_49245);
or UO_1353 (O_1353,N_49742,N_49472);
xor UO_1354 (O_1354,N_49138,N_49995);
and UO_1355 (O_1355,N_49987,N_49097);
nor UO_1356 (O_1356,N_49858,N_49270);
nor UO_1357 (O_1357,N_49862,N_49502);
or UO_1358 (O_1358,N_49622,N_49886);
xnor UO_1359 (O_1359,N_49196,N_49362);
and UO_1360 (O_1360,N_49988,N_49891);
nor UO_1361 (O_1361,N_49197,N_49036);
xor UO_1362 (O_1362,N_49914,N_49449);
or UO_1363 (O_1363,N_49589,N_49580);
xor UO_1364 (O_1364,N_49348,N_49375);
nor UO_1365 (O_1365,N_49810,N_49598);
nor UO_1366 (O_1366,N_49642,N_49233);
and UO_1367 (O_1367,N_49581,N_49538);
and UO_1368 (O_1368,N_49774,N_49884);
and UO_1369 (O_1369,N_49669,N_49371);
or UO_1370 (O_1370,N_49010,N_49369);
or UO_1371 (O_1371,N_49220,N_49544);
nor UO_1372 (O_1372,N_49312,N_49099);
nand UO_1373 (O_1373,N_49875,N_49572);
nor UO_1374 (O_1374,N_49550,N_49982);
xnor UO_1375 (O_1375,N_49647,N_49865);
and UO_1376 (O_1376,N_49711,N_49191);
nand UO_1377 (O_1377,N_49700,N_49164);
xor UO_1378 (O_1378,N_49081,N_49810);
nor UO_1379 (O_1379,N_49082,N_49772);
and UO_1380 (O_1380,N_49416,N_49135);
nor UO_1381 (O_1381,N_49013,N_49635);
xor UO_1382 (O_1382,N_49444,N_49057);
or UO_1383 (O_1383,N_49820,N_49880);
xnor UO_1384 (O_1384,N_49184,N_49593);
xnor UO_1385 (O_1385,N_49967,N_49619);
and UO_1386 (O_1386,N_49758,N_49272);
or UO_1387 (O_1387,N_49670,N_49261);
nand UO_1388 (O_1388,N_49637,N_49205);
nand UO_1389 (O_1389,N_49300,N_49257);
and UO_1390 (O_1390,N_49181,N_49663);
or UO_1391 (O_1391,N_49806,N_49166);
and UO_1392 (O_1392,N_49010,N_49316);
nand UO_1393 (O_1393,N_49048,N_49816);
nand UO_1394 (O_1394,N_49788,N_49514);
xnor UO_1395 (O_1395,N_49876,N_49594);
nor UO_1396 (O_1396,N_49238,N_49025);
nand UO_1397 (O_1397,N_49653,N_49138);
or UO_1398 (O_1398,N_49219,N_49221);
nor UO_1399 (O_1399,N_49996,N_49124);
or UO_1400 (O_1400,N_49719,N_49198);
or UO_1401 (O_1401,N_49003,N_49160);
or UO_1402 (O_1402,N_49973,N_49046);
nand UO_1403 (O_1403,N_49757,N_49860);
xnor UO_1404 (O_1404,N_49180,N_49312);
and UO_1405 (O_1405,N_49529,N_49108);
nor UO_1406 (O_1406,N_49914,N_49984);
nor UO_1407 (O_1407,N_49621,N_49134);
nand UO_1408 (O_1408,N_49600,N_49920);
and UO_1409 (O_1409,N_49466,N_49812);
and UO_1410 (O_1410,N_49805,N_49951);
and UO_1411 (O_1411,N_49768,N_49108);
and UO_1412 (O_1412,N_49314,N_49456);
xor UO_1413 (O_1413,N_49320,N_49558);
nand UO_1414 (O_1414,N_49955,N_49256);
xor UO_1415 (O_1415,N_49725,N_49889);
or UO_1416 (O_1416,N_49291,N_49019);
or UO_1417 (O_1417,N_49944,N_49171);
or UO_1418 (O_1418,N_49882,N_49981);
and UO_1419 (O_1419,N_49380,N_49990);
xnor UO_1420 (O_1420,N_49258,N_49697);
and UO_1421 (O_1421,N_49502,N_49056);
and UO_1422 (O_1422,N_49666,N_49771);
xnor UO_1423 (O_1423,N_49765,N_49697);
nor UO_1424 (O_1424,N_49383,N_49462);
or UO_1425 (O_1425,N_49174,N_49614);
or UO_1426 (O_1426,N_49853,N_49368);
xor UO_1427 (O_1427,N_49571,N_49256);
and UO_1428 (O_1428,N_49047,N_49452);
xnor UO_1429 (O_1429,N_49480,N_49730);
nor UO_1430 (O_1430,N_49318,N_49554);
nor UO_1431 (O_1431,N_49353,N_49920);
or UO_1432 (O_1432,N_49285,N_49433);
or UO_1433 (O_1433,N_49502,N_49462);
nor UO_1434 (O_1434,N_49758,N_49728);
nand UO_1435 (O_1435,N_49488,N_49537);
or UO_1436 (O_1436,N_49564,N_49286);
nor UO_1437 (O_1437,N_49809,N_49561);
nor UO_1438 (O_1438,N_49877,N_49641);
nor UO_1439 (O_1439,N_49842,N_49849);
or UO_1440 (O_1440,N_49167,N_49441);
and UO_1441 (O_1441,N_49666,N_49069);
or UO_1442 (O_1442,N_49136,N_49068);
xor UO_1443 (O_1443,N_49600,N_49856);
and UO_1444 (O_1444,N_49398,N_49631);
nand UO_1445 (O_1445,N_49740,N_49146);
xnor UO_1446 (O_1446,N_49401,N_49500);
nor UO_1447 (O_1447,N_49185,N_49714);
or UO_1448 (O_1448,N_49480,N_49613);
xnor UO_1449 (O_1449,N_49315,N_49005);
or UO_1450 (O_1450,N_49982,N_49824);
xnor UO_1451 (O_1451,N_49483,N_49482);
nand UO_1452 (O_1452,N_49015,N_49415);
or UO_1453 (O_1453,N_49191,N_49348);
xnor UO_1454 (O_1454,N_49616,N_49716);
xor UO_1455 (O_1455,N_49250,N_49109);
nor UO_1456 (O_1456,N_49729,N_49218);
nor UO_1457 (O_1457,N_49816,N_49648);
or UO_1458 (O_1458,N_49215,N_49205);
nor UO_1459 (O_1459,N_49546,N_49179);
nand UO_1460 (O_1460,N_49468,N_49426);
xor UO_1461 (O_1461,N_49538,N_49619);
nor UO_1462 (O_1462,N_49500,N_49793);
nor UO_1463 (O_1463,N_49471,N_49856);
nand UO_1464 (O_1464,N_49125,N_49571);
and UO_1465 (O_1465,N_49435,N_49974);
and UO_1466 (O_1466,N_49927,N_49698);
and UO_1467 (O_1467,N_49864,N_49944);
or UO_1468 (O_1468,N_49480,N_49870);
or UO_1469 (O_1469,N_49373,N_49441);
nor UO_1470 (O_1470,N_49060,N_49138);
and UO_1471 (O_1471,N_49386,N_49838);
or UO_1472 (O_1472,N_49103,N_49255);
or UO_1473 (O_1473,N_49982,N_49904);
nand UO_1474 (O_1474,N_49483,N_49513);
and UO_1475 (O_1475,N_49316,N_49394);
and UO_1476 (O_1476,N_49811,N_49845);
or UO_1477 (O_1477,N_49322,N_49160);
or UO_1478 (O_1478,N_49146,N_49947);
nor UO_1479 (O_1479,N_49698,N_49310);
nor UO_1480 (O_1480,N_49803,N_49836);
or UO_1481 (O_1481,N_49668,N_49636);
xnor UO_1482 (O_1482,N_49108,N_49869);
xnor UO_1483 (O_1483,N_49373,N_49105);
nand UO_1484 (O_1484,N_49176,N_49548);
nor UO_1485 (O_1485,N_49082,N_49692);
nand UO_1486 (O_1486,N_49639,N_49234);
or UO_1487 (O_1487,N_49114,N_49120);
nand UO_1488 (O_1488,N_49949,N_49211);
and UO_1489 (O_1489,N_49680,N_49694);
nand UO_1490 (O_1490,N_49954,N_49783);
or UO_1491 (O_1491,N_49474,N_49890);
xnor UO_1492 (O_1492,N_49400,N_49799);
nand UO_1493 (O_1493,N_49502,N_49464);
and UO_1494 (O_1494,N_49789,N_49422);
nand UO_1495 (O_1495,N_49999,N_49895);
nor UO_1496 (O_1496,N_49852,N_49288);
xnor UO_1497 (O_1497,N_49737,N_49212);
nand UO_1498 (O_1498,N_49830,N_49959);
nor UO_1499 (O_1499,N_49325,N_49400);
xnor UO_1500 (O_1500,N_49458,N_49412);
or UO_1501 (O_1501,N_49243,N_49462);
nor UO_1502 (O_1502,N_49961,N_49677);
or UO_1503 (O_1503,N_49795,N_49743);
nor UO_1504 (O_1504,N_49245,N_49600);
and UO_1505 (O_1505,N_49691,N_49554);
xor UO_1506 (O_1506,N_49639,N_49996);
or UO_1507 (O_1507,N_49189,N_49706);
or UO_1508 (O_1508,N_49629,N_49376);
xnor UO_1509 (O_1509,N_49988,N_49043);
nor UO_1510 (O_1510,N_49673,N_49825);
xnor UO_1511 (O_1511,N_49697,N_49085);
and UO_1512 (O_1512,N_49831,N_49330);
nand UO_1513 (O_1513,N_49885,N_49491);
nand UO_1514 (O_1514,N_49371,N_49429);
xnor UO_1515 (O_1515,N_49667,N_49305);
nor UO_1516 (O_1516,N_49855,N_49674);
or UO_1517 (O_1517,N_49686,N_49479);
nand UO_1518 (O_1518,N_49513,N_49864);
xor UO_1519 (O_1519,N_49610,N_49135);
and UO_1520 (O_1520,N_49917,N_49941);
or UO_1521 (O_1521,N_49639,N_49853);
or UO_1522 (O_1522,N_49487,N_49966);
and UO_1523 (O_1523,N_49138,N_49580);
xnor UO_1524 (O_1524,N_49876,N_49978);
nor UO_1525 (O_1525,N_49521,N_49950);
nor UO_1526 (O_1526,N_49053,N_49813);
xor UO_1527 (O_1527,N_49405,N_49720);
and UO_1528 (O_1528,N_49440,N_49222);
or UO_1529 (O_1529,N_49875,N_49457);
and UO_1530 (O_1530,N_49158,N_49494);
nand UO_1531 (O_1531,N_49228,N_49090);
nand UO_1532 (O_1532,N_49592,N_49596);
nor UO_1533 (O_1533,N_49991,N_49715);
and UO_1534 (O_1534,N_49422,N_49156);
nand UO_1535 (O_1535,N_49609,N_49498);
nor UO_1536 (O_1536,N_49037,N_49401);
nor UO_1537 (O_1537,N_49762,N_49923);
or UO_1538 (O_1538,N_49092,N_49935);
nand UO_1539 (O_1539,N_49071,N_49729);
and UO_1540 (O_1540,N_49358,N_49454);
xnor UO_1541 (O_1541,N_49328,N_49668);
nand UO_1542 (O_1542,N_49878,N_49662);
and UO_1543 (O_1543,N_49473,N_49365);
nor UO_1544 (O_1544,N_49203,N_49044);
nor UO_1545 (O_1545,N_49488,N_49415);
nand UO_1546 (O_1546,N_49545,N_49160);
xor UO_1547 (O_1547,N_49483,N_49970);
nand UO_1548 (O_1548,N_49650,N_49342);
xnor UO_1549 (O_1549,N_49776,N_49550);
nor UO_1550 (O_1550,N_49488,N_49908);
nand UO_1551 (O_1551,N_49673,N_49141);
or UO_1552 (O_1552,N_49132,N_49281);
xnor UO_1553 (O_1553,N_49567,N_49521);
nand UO_1554 (O_1554,N_49305,N_49343);
and UO_1555 (O_1555,N_49382,N_49782);
xnor UO_1556 (O_1556,N_49774,N_49173);
or UO_1557 (O_1557,N_49600,N_49432);
and UO_1558 (O_1558,N_49172,N_49817);
xor UO_1559 (O_1559,N_49000,N_49937);
xor UO_1560 (O_1560,N_49579,N_49503);
or UO_1561 (O_1561,N_49991,N_49496);
nor UO_1562 (O_1562,N_49851,N_49865);
or UO_1563 (O_1563,N_49262,N_49856);
xnor UO_1564 (O_1564,N_49426,N_49903);
xor UO_1565 (O_1565,N_49141,N_49503);
or UO_1566 (O_1566,N_49568,N_49365);
and UO_1567 (O_1567,N_49574,N_49648);
or UO_1568 (O_1568,N_49173,N_49760);
nand UO_1569 (O_1569,N_49266,N_49955);
or UO_1570 (O_1570,N_49424,N_49620);
xnor UO_1571 (O_1571,N_49877,N_49821);
or UO_1572 (O_1572,N_49861,N_49584);
nor UO_1573 (O_1573,N_49392,N_49968);
and UO_1574 (O_1574,N_49834,N_49837);
or UO_1575 (O_1575,N_49134,N_49674);
nand UO_1576 (O_1576,N_49604,N_49675);
nand UO_1577 (O_1577,N_49484,N_49550);
nor UO_1578 (O_1578,N_49330,N_49459);
xnor UO_1579 (O_1579,N_49422,N_49544);
and UO_1580 (O_1580,N_49945,N_49129);
nor UO_1581 (O_1581,N_49131,N_49930);
or UO_1582 (O_1582,N_49395,N_49873);
or UO_1583 (O_1583,N_49356,N_49089);
nand UO_1584 (O_1584,N_49456,N_49521);
or UO_1585 (O_1585,N_49185,N_49132);
nand UO_1586 (O_1586,N_49982,N_49765);
nand UO_1587 (O_1587,N_49131,N_49491);
or UO_1588 (O_1588,N_49507,N_49442);
xnor UO_1589 (O_1589,N_49332,N_49093);
xnor UO_1590 (O_1590,N_49583,N_49292);
nor UO_1591 (O_1591,N_49210,N_49379);
xor UO_1592 (O_1592,N_49690,N_49048);
nor UO_1593 (O_1593,N_49833,N_49605);
nand UO_1594 (O_1594,N_49677,N_49003);
and UO_1595 (O_1595,N_49735,N_49503);
or UO_1596 (O_1596,N_49175,N_49827);
xor UO_1597 (O_1597,N_49222,N_49850);
xnor UO_1598 (O_1598,N_49607,N_49017);
nand UO_1599 (O_1599,N_49896,N_49670);
nand UO_1600 (O_1600,N_49627,N_49309);
nand UO_1601 (O_1601,N_49683,N_49508);
nor UO_1602 (O_1602,N_49055,N_49256);
nor UO_1603 (O_1603,N_49426,N_49082);
and UO_1604 (O_1604,N_49073,N_49499);
and UO_1605 (O_1605,N_49815,N_49704);
or UO_1606 (O_1606,N_49087,N_49606);
xor UO_1607 (O_1607,N_49615,N_49468);
or UO_1608 (O_1608,N_49064,N_49577);
xor UO_1609 (O_1609,N_49006,N_49515);
xnor UO_1610 (O_1610,N_49035,N_49473);
nand UO_1611 (O_1611,N_49339,N_49687);
or UO_1612 (O_1612,N_49908,N_49402);
nor UO_1613 (O_1613,N_49726,N_49104);
or UO_1614 (O_1614,N_49310,N_49561);
nand UO_1615 (O_1615,N_49694,N_49908);
nand UO_1616 (O_1616,N_49205,N_49066);
nor UO_1617 (O_1617,N_49881,N_49874);
and UO_1618 (O_1618,N_49162,N_49773);
nand UO_1619 (O_1619,N_49209,N_49330);
and UO_1620 (O_1620,N_49865,N_49181);
xnor UO_1621 (O_1621,N_49040,N_49893);
xnor UO_1622 (O_1622,N_49407,N_49120);
nor UO_1623 (O_1623,N_49098,N_49568);
or UO_1624 (O_1624,N_49970,N_49102);
nand UO_1625 (O_1625,N_49236,N_49734);
xnor UO_1626 (O_1626,N_49421,N_49688);
or UO_1627 (O_1627,N_49607,N_49953);
and UO_1628 (O_1628,N_49267,N_49885);
xor UO_1629 (O_1629,N_49657,N_49933);
nor UO_1630 (O_1630,N_49703,N_49291);
nand UO_1631 (O_1631,N_49541,N_49222);
and UO_1632 (O_1632,N_49863,N_49101);
nor UO_1633 (O_1633,N_49285,N_49451);
and UO_1634 (O_1634,N_49718,N_49476);
and UO_1635 (O_1635,N_49820,N_49669);
xor UO_1636 (O_1636,N_49782,N_49155);
nor UO_1637 (O_1637,N_49454,N_49609);
nor UO_1638 (O_1638,N_49670,N_49586);
nor UO_1639 (O_1639,N_49170,N_49143);
or UO_1640 (O_1640,N_49842,N_49656);
and UO_1641 (O_1641,N_49231,N_49053);
xnor UO_1642 (O_1642,N_49317,N_49814);
xnor UO_1643 (O_1643,N_49832,N_49381);
or UO_1644 (O_1644,N_49319,N_49628);
or UO_1645 (O_1645,N_49240,N_49158);
and UO_1646 (O_1646,N_49964,N_49363);
nor UO_1647 (O_1647,N_49364,N_49538);
xor UO_1648 (O_1648,N_49501,N_49425);
xor UO_1649 (O_1649,N_49273,N_49103);
and UO_1650 (O_1650,N_49156,N_49994);
xor UO_1651 (O_1651,N_49156,N_49334);
nand UO_1652 (O_1652,N_49109,N_49540);
or UO_1653 (O_1653,N_49059,N_49781);
xnor UO_1654 (O_1654,N_49530,N_49025);
nand UO_1655 (O_1655,N_49792,N_49427);
nand UO_1656 (O_1656,N_49018,N_49027);
xnor UO_1657 (O_1657,N_49908,N_49910);
xor UO_1658 (O_1658,N_49627,N_49110);
nand UO_1659 (O_1659,N_49721,N_49972);
nand UO_1660 (O_1660,N_49655,N_49477);
and UO_1661 (O_1661,N_49239,N_49594);
nor UO_1662 (O_1662,N_49073,N_49754);
xor UO_1663 (O_1663,N_49659,N_49025);
and UO_1664 (O_1664,N_49634,N_49611);
or UO_1665 (O_1665,N_49460,N_49982);
and UO_1666 (O_1666,N_49522,N_49774);
nand UO_1667 (O_1667,N_49473,N_49087);
nand UO_1668 (O_1668,N_49850,N_49320);
and UO_1669 (O_1669,N_49216,N_49085);
xor UO_1670 (O_1670,N_49468,N_49539);
and UO_1671 (O_1671,N_49705,N_49361);
nor UO_1672 (O_1672,N_49003,N_49138);
and UO_1673 (O_1673,N_49143,N_49493);
or UO_1674 (O_1674,N_49607,N_49470);
nand UO_1675 (O_1675,N_49182,N_49196);
and UO_1676 (O_1676,N_49658,N_49799);
nor UO_1677 (O_1677,N_49505,N_49151);
nor UO_1678 (O_1678,N_49981,N_49917);
xnor UO_1679 (O_1679,N_49328,N_49600);
nor UO_1680 (O_1680,N_49851,N_49716);
or UO_1681 (O_1681,N_49037,N_49259);
nand UO_1682 (O_1682,N_49770,N_49053);
or UO_1683 (O_1683,N_49752,N_49442);
nand UO_1684 (O_1684,N_49583,N_49664);
and UO_1685 (O_1685,N_49721,N_49405);
nor UO_1686 (O_1686,N_49816,N_49027);
xor UO_1687 (O_1687,N_49835,N_49569);
and UO_1688 (O_1688,N_49876,N_49859);
nand UO_1689 (O_1689,N_49264,N_49553);
or UO_1690 (O_1690,N_49808,N_49476);
and UO_1691 (O_1691,N_49069,N_49292);
or UO_1692 (O_1692,N_49873,N_49998);
nor UO_1693 (O_1693,N_49873,N_49922);
or UO_1694 (O_1694,N_49911,N_49380);
and UO_1695 (O_1695,N_49657,N_49643);
nor UO_1696 (O_1696,N_49828,N_49026);
and UO_1697 (O_1697,N_49293,N_49136);
and UO_1698 (O_1698,N_49379,N_49331);
nor UO_1699 (O_1699,N_49806,N_49256);
and UO_1700 (O_1700,N_49491,N_49081);
nor UO_1701 (O_1701,N_49990,N_49097);
nor UO_1702 (O_1702,N_49589,N_49514);
nand UO_1703 (O_1703,N_49993,N_49792);
xnor UO_1704 (O_1704,N_49697,N_49810);
nand UO_1705 (O_1705,N_49920,N_49862);
nand UO_1706 (O_1706,N_49750,N_49408);
and UO_1707 (O_1707,N_49634,N_49915);
xor UO_1708 (O_1708,N_49585,N_49950);
nand UO_1709 (O_1709,N_49794,N_49725);
nand UO_1710 (O_1710,N_49928,N_49400);
or UO_1711 (O_1711,N_49077,N_49477);
nand UO_1712 (O_1712,N_49375,N_49650);
and UO_1713 (O_1713,N_49695,N_49327);
nor UO_1714 (O_1714,N_49354,N_49529);
or UO_1715 (O_1715,N_49052,N_49860);
and UO_1716 (O_1716,N_49063,N_49187);
nor UO_1717 (O_1717,N_49020,N_49791);
and UO_1718 (O_1718,N_49342,N_49522);
or UO_1719 (O_1719,N_49091,N_49894);
nand UO_1720 (O_1720,N_49632,N_49106);
and UO_1721 (O_1721,N_49391,N_49344);
nor UO_1722 (O_1722,N_49816,N_49078);
or UO_1723 (O_1723,N_49479,N_49155);
nor UO_1724 (O_1724,N_49593,N_49158);
nor UO_1725 (O_1725,N_49596,N_49074);
nand UO_1726 (O_1726,N_49244,N_49329);
nor UO_1727 (O_1727,N_49571,N_49224);
or UO_1728 (O_1728,N_49220,N_49159);
nand UO_1729 (O_1729,N_49562,N_49595);
xor UO_1730 (O_1730,N_49754,N_49819);
or UO_1731 (O_1731,N_49875,N_49654);
or UO_1732 (O_1732,N_49136,N_49106);
nor UO_1733 (O_1733,N_49507,N_49106);
xnor UO_1734 (O_1734,N_49155,N_49827);
and UO_1735 (O_1735,N_49661,N_49597);
and UO_1736 (O_1736,N_49314,N_49262);
xor UO_1737 (O_1737,N_49107,N_49764);
and UO_1738 (O_1738,N_49653,N_49807);
nor UO_1739 (O_1739,N_49134,N_49876);
nor UO_1740 (O_1740,N_49801,N_49038);
nor UO_1741 (O_1741,N_49258,N_49107);
nor UO_1742 (O_1742,N_49984,N_49123);
nand UO_1743 (O_1743,N_49623,N_49713);
xnor UO_1744 (O_1744,N_49360,N_49859);
or UO_1745 (O_1745,N_49204,N_49196);
and UO_1746 (O_1746,N_49371,N_49045);
xnor UO_1747 (O_1747,N_49040,N_49611);
nor UO_1748 (O_1748,N_49659,N_49865);
or UO_1749 (O_1749,N_49042,N_49986);
and UO_1750 (O_1750,N_49123,N_49839);
xnor UO_1751 (O_1751,N_49179,N_49005);
nor UO_1752 (O_1752,N_49439,N_49273);
xor UO_1753 (O_1753,N_49854,N_49383);
or UO_1754 (O_1754,N_49594,N_49124);
xor UO_1755 (O_1755,N_49658,N_49474);
nand UO_1756 (O_1756,N_49699,N_49032);
or UO_1757 (O_1757,N_49655,N_49554);
nor UO_1758 (O_1758,N_49353,N_49256);
and UO_1759 (O_1759,N_49075,N_49951);
xnor UO_1760 (O_1760,N_49281,N_49289);
xnor UO_1761 (O_1761,N_49633,N_49499);
nand UO_1762 (O_1762,N_49428,N_49539);
nand UO_1763 (O_1763,N_49497,N_49539);
nand UO_1764 (O_1764,N_49799,N_49284);
or UO_1765 (O_1765,N_49362,N_49880);
or UO_1766 (O_1766,N_49058,N_49120);
nand UO_1767 (O_1767,N_49882,N_49738);
and UO_1768 (O_1768,N_49655,N_49080);
xor UO_1769 (O_1769,N_49185,N_49979);
xor UO_1770 (O_1770,N_49151,N_49945);
nand UO_1771 (O_1771,N_49636,N_49248);
nor UO_1772 (O_1772,N_49850,N_49027);
and UO_1773 (O_1773,N_49179,N_49031);
and UO_1774 (O_1774,N_49829,N_49781);
xor UO_1775 (O_1775,N_49832,N_49575);
xor UO_1776 (O_1776,N_49312,N_49871);
and UO_1777 (O_1777,N_49509,N_49565);
or UO_1778 (O_1778,N_49539,N_49189);
xnor UO_1779 (O_1779,N_49180,N_49967);
nor UO_1780 (O_1780,N_49041,N_49207);
xnor UO_1781 (O_1781,N_49333,N_49656);
nand UO_1782 (O_1782,N_49458,N_49204);
xnor UO_1783 (O_1783,N_49245,N_49888);
nand UO_1784 (O_1784,N_49727,N_49561);
and UO_1785 (O_1785,N_49944,N_49899);
and UO_1786 (O_1786,N_49687,N_49016);
xor UO_1787 (O_1787,N_49931,N_49450);
or UO_1788 (O_1788,N_49733,N_49755);
nand UO_1789 (O_1789,N_49969,N_49770);
xor UO_1790 (O_1790,N_49737,N_49557);
or UO_1791 (O_1791,N_49185,N_49417);
xor UO_1792 (O_1792,N_49630,N_49481);
nand UO_1793 (O_1793,N_49407,N_49900);
nor UO_1794 (O_1794,N_49836,N_49496);
nor UO_1795 (O_1795,N_49855,N_49697);
xnor UO_1796 (O_1796,N_49969,N_49142);
nor UO_1797 (O_1797,N_49725,N_49160);
xor UO_1798 (O_1798,N_49798,N_49635);
xnor UO_1799 (O_1799,N_49332,N_49284);
and UO_1800 (O_1800,N_49869,N_49704);
xor UO_1801 (O_1801,N_49693,N_49828);
and UO_1802 (O_1802,N_49853,N_49234);
xnor UO_1803 (O_1803,N_49069,N_49585);
or UO_1804 (O_1804,N_49545,N_49848);
and UO_1805 (O_1805,N_49461,N_49348);
and UO_1806 (O_1806,N_49876,N_49165);
nand UO_1807 (O_1807,N_49888,N_49864);
nor UO_1808 (O_1808,N_49078,N_49508);
and UO_1809 (O_1809,N_49610,N_49400);
or UO_1810 (O_1810,N_49273,N_49128);
nand UO_1811 (O_1811,N_49435,N_49748);
and UO_1812 (O_1812,N_49892,N_49248);
nand UO_1813 (O_1813,N_49072,N_49066);
and UO_1814 (O_1814,N_49216,N_49914);
nand UO_1815 (O_1815,N_49468,N_49776);
and UO_1816 (O_1816,N_49820,N_49418);
nor UO_1817 (O_1817,N_49244,N_49130);
or UO_1818 (O_1818,N_49547,N_49536);
or UO_1819 (O_1819,N_49940,N_49970);
xor UO_1820 (O_1820,N_49821,N_49297);
nor UO_1821 (O_1821,N_49314,N_49564);
and UO_1822 (O_1822,N_49029,N_49638);
or UO_1823 (O_1823,N_49388,N_49255);
nand UO_1824 (O_1824,N_49681,N_49795);
nand UO_1825 (O_1825,N_49573,N_49969);
xnor UO_1826 (O_1826,N_49423,N_49269);
nor UO_1827 (O_1827,N_49499,N_49252);
nor UO_1828 (O_1828,N_49580,N_49474);
and UO_1829 (O_1829,N_49225,N_49492);
xor UO_1830 (O_1830,N_49867,N_49916);
xor UO_1831 (O_1831,N_49667,N_49231);
or UO_1832 (O_1832,N_49034,N_49221);
xnor UO_1833 (O_1833,N_49633,N_49885);
or UO_1834 (O_1834,N_49971,N_49321);
or UO_1835 (O_1835,N_49680,N_49901);
xor UO_1836 (O_1836,N_49537,N_49479);
and UO_1837 (O_1837,N_49697,N_49787);
nor UO_1838 (O_1838,N_49849,N_49605);
nand UO_1839 (O_1839,N_49789,N_49892);
nand UO_1840 (O_1840,N_49912,N_49671);
xor UO_1841 (O_1841,N_49818,N_49226);
xor UO_1842 (O_1842,N_49702,N_49262);
nor UO_1843 (O_1843,N_49436,N_49148);
nor UO_1844 (O_1844,N_49934,N_49168);
nand UO_1845 (O_1845,N_49541,N_49712);
nor UO_1846 (O_1846,N_49230,N_49950);
nand UO_1847 (O_1847,N_49887,N_49619);
nand UO_1848 (O_1848,N_49246,N_49652);
or UO_1849 (O_1849,N_49403,N_49618);
or UO_1850 (O_1850,N_49697,N_49156);
or UO_1851 (O_1851,N_49935,N_49924);
or UO_1852 (O_1852,N_49829,N_49302);
nand UO_1853 (O_1853,N_49881,N_49434);
and UO_1854 (O_1854,N_49451,N_49796);
and UO_1855 (O_1855,N_49112,N_49835);
and UO_1856 (O_1856,N_49312,N_49203);
and UO_1857 (O_1857,N_49756,N_49891);
or UO_1858 (O_1858,N_49360,N_49651);
or UO_1859 (O_1859,N_49135,N_49175);
xor UO_1860 (O_1860,N_49632,N_49310);
nor UO_1861 (O_1861,N_49084,N_49460);
xnor UO_1862 (O_1862,N_49210,N_49322);
or UO_1863 (O_1863,N_49320,N_49948);
and UO_1864 (O_1864,N_49367,N_49580);
nor UO_1865 (O_1865,N_49765,N_49449);
nor UO_1866 (O_1866,N_49610,N_49914);
and UO_1867 (O_1867,N_49243,N_49465);
nor UO_1868 (O_1868,N_49059,N_49706);
and UO_1869 (O_1869,N_49150,N_49474);
nand UO_1870 (O_1870,N_49228,N_49876);
nand UO_1871 (O_1871,N_49237,N_49969);
xnor UO_1872 (O_1872,N_49959,N_49241);
nor UO_1873 (O_1873,N_49403,N_49662);
and UO_1874 (O_1874,N_49374,N_49622);
nand UO_1875 (O_1875,N_49876,N_49925);
and UO_1876 (O_1876,N_49005,N_49698);
and UO_1877 (O_1877,N_49549,N_49782);
nand UO_1878 (O_1878,N_49407,N_49879);
and UO_1879 (O_1879,N_49299,N_49092);
nand UO_1880 (O_1880,N_49384,N_49385);
or UO_1881 (O_1881,N_49868,N_49308);
xor UO_1882 (O_1882,N_49347,N_49044);
xor UO_1883 (O_1883,N_49243,N_49436);
and UO_1884 (O_1884,N_49149,N_49069);
nor UO_1885 (O_1885,N_49791,N_49680);
nand UO_1886 (O_1886,N_49032,N_49151);
xor UO_1887 (O_1887,N_49672,N_49654);
or UO_1888 (O_1888,N_49555,N_49084);
or UO_1889 (O_1889,N_49946,N_49196);
or UO_1890 (O_1890,N_49557,N_49863);
and UO_1891 (O_1891,N_49820,N_49359);
and UO_1892 (O_1892,N_49850,N_49595);
nor UO_1893 (O_1893,N_49166,N_49460);
or UO_1894 (O_1894,N_49472,N_49692);
nand UO_1895 (O_1895,N_49587,N_49806);
nor UO_1896 (O_1896,N_49595,N_49903);
nand UO_1897 (O_1897,N_49603,N_49182);
xnor UO_1898 (O_1898,N_49458,N_49949);
nand UO_1899 (O_1899,N_49051,N_49835);
or UO_1900 (O_1900,N_49447,N_49345);
nand UO_1901 (O_1901,N_49011,N_49841);
nand UO_1902 (O_1902,N_49463,N_49307);
and UO_1903 (O_1903,N_49297,N_49042);
and UO_1904 (O_1904,N_49260,N_49658);
xor UO_1905 (O_1905,N_49437,N_49558);
and UO_1906 (O_1906,N_49784,N_49592);
xnor UO_1907 (O_1907,N_49244,N_49983);
xor UO_1908 (O_1908,N_49547,N_49885);
nand UO_1909 (O_1909,N_49128,N_49469);
or UO_1910 (O_1910,N_49909,N_49484);
nand UO_1911 (O_1911,N_49274,N_49977);
xnor UO_1912 (O_1912,N_49217,N_49866);
nor UO_1913 (O_1913,N_49567,N_49302);
nand UO_1914 (O_1914,N_49932,N_49281);
and UO_1915 (O_1915,N_49942,N_49879);
nand UO_1916 (O_1916,N_49616,N_49999);
xor UO_1917 (O_1917,N_49500,N_49595);
and UO_1918 (O_1918,N_49042,N_49599);
and UO_1919 (O_1919,N_49468,N_49521);
nand UO_1920 (O_1920,N_49602,N_49565);
nand UO_1921 (O_1921,N_49380,N_49971);
nand UO_1922 (O_1922,N_49092,N_49467);
nor UO_1923 (O_1923,N_49992,N_49319);
nand UO_1924 (O_1924,N_49808,N_49078);
xor UO_1925 (O_1925,N_49441,N_49707);
xor UO_1926 (O_1926,N_49313,N_49491);
or UO_1927 (O_1927,N_49037,N_49822);
nand UO_1928 (O_1928,N_49361,N_49992);
or UO_1929 (O_1929,N_49920,N_49199);
nand UO_1930 (O_1930,N_49969,N_49111);
xor UO_1931 (O_1931,N_49269,N_49304);
nand UO_1932 (O_1932,N_49063,N_49962);
or UO_1933 (O_1933,N_49281,N_49456);
nor UO_1934 (O_1934,N_49026,N_49741);
or UO_1935 (O_1935,N_49013,N_49414);
or UO_1936 (O_1936,N_49656,N_49081);
nand UO_1937 (O_1937,N_49681,N_49981);
nand UO_1938 (O_1938,N_49081,N_49867);
and UO_1939 (O_1939,N_49065,N_49624);
xor UO_1940 (O_1940,N_49849,N_49571);
xor UO_1941 (O_1941,N_49623,N_49548);
and UO_1942 (O_1942,N_49212,N_49882);
nand UO_1943 (O_1943,N_49141,N_49945);
or UO_1944 (O_1944,N_49960,N_49427);
and UO_1945 (O_1945,N_49523,N_49034);
or UO_1946 (O_1946,N_49299,N_49002);
nand UO_1947 (O_1947,N_49213,N_49055);
nand UO_1948 (O_1948,N_49245,N_49300);
and UO_1949 (O_1949,N_49217,N_49504);
nor UO_1950 (O_1950,N_49401,N_49116);
nor UO_1951 (O_1951,N_49729,N_49508);
xnor UO_1952 (O_1952,N_49684,N_49506);
and UO_1953 (O_1953,N_49364,N_49426);
or UO_1954 (O_1954,N_49474,N_49567);
nor UO_1955 (O_1955,N_49076,N_49470);
nor UO_1956 (O_1956,N_49689,N_49983);
nor UO_1957 (O_1957,N_49045,N_49794);
xor UO_1958 (O_1958,N_49468,N_49579);
and UO_1959 (O_1959,N_49766,N_49339);
nor UO_1960 (O_1960,N_49588,N_49475);
nand UO_1961 (O_1961,N_49659,N_49103);
nand UO_1962 (O_1962,N_49254,N_49305);
nor UO_1963 (O_1963,N_49586,N_49540);
xnor UO_1964 (O_1964,N_49624,N_49101);
nor UO_1965 (O_1965,N_49996,N_49344);
or UO_1966 (O_1966,N_49214,N_49202);
and UO_1967 (O_1967,N_49449,N_49219);
nand UO_1968 (O_1968,N_49306,N_49369);
and UO_1969 (O_1969,N_49206,N_49880);
or UO_1970 (O_1970,N_49803,N_49284);
or UO_1971 (O_1971,N_49713,N_49317);
or UO_1972 (O_1972,N_49767,N_49335);
nand UO_1973 (O_1973,N_49552,N_49556);
nand UO_1974 (O_1974,N_49377,N_49353);
and UO_1975 (O_1975,N_49996,N_49994);
or UO_1976 (O_1976,N_49967,N_49144);
or UO_1977 (O_1977,N_49325,N_49983);
and UO_1978 (O_1978,N_49136,N_49389);
or UO_1979 (O_1979,N_49601,N_49954);
xor UO_1980 (O_1980,N_49470,N_49752);
nor UO_1981 (O_1981,N_49593,N_49929);
and UO_1982 (O_1982,N_49985,N_49668);
xor UO_1983 (O_1983,N_49033,N_49649);
nor UO_1984 (O_1984,N_49394,N_49168);
nand UO_1985 (O_1985,N_49589,N_49979);
xor UO_1986 (O_1986,N_49935,N_49570);
and UO_1987 (O_1987,N_49100,N_49904);
and UO_1988 (O_1988,N_49354,N_49078);
and UO_1989 (O_1989,N_49810,N_49906);
nor UO_1990 (O_1990,N_49466,N_49420);
nand UO_1991 (O_1991,N_49060,N_49522);
or UO_1992 (O_1992,N_49792,N_49965);
and UO_1993 (O_1993,N_49401,N_49336);
nor UO_1994 (O_1994,N_49962,N_49795);
nand UO_1995 (O_1995,N_49775,N_49449);
and UO_1996 (O_1996,N_49558,N_49457);
and UO_1997 (O_1997,N_49696,N_49870);
nor UO_1998 (O_1998,N_49838,N_49080);
nor UO_1999 (O_1999,N_49019,N_49570);
or UO_2000 (O_2000,N_49206,N_49515);
and UO_2001 (O_2001,N_49586,N_49228);
or UO_2002 (O_2002,N_49105,N_49882);
or UO_2003 (O_2003,N_49956,N_49299);
xnor UO_2004 (O_2004,N_49276,N_49347);
or UO_2005 (O_2005,N_49956,N_49540);
and UO_2006 (O_2006,N_49710,N_49009);
and UO_2007 (O_2007,N_49895,N_49084);
nand UO_2008 (O_2008,N_49484,N_49986);
nand UO_2009 (O_2009,N_49960,N_49067);
and UO_2010 (O_2010,N_49716,N_49357);
or UO_2011 (O_2011,N_49095,N_49509);
or UO_2012 (O_2012,N_49582,N_49471);
nand UO_2013 (O_2013,N_49233,N_49146);
and UO_2014 (O_2014,N_49428,N_49766);
and UO_2015 (O_2015,N_49920,N_49094);
nand UO_2016 (O_2016,N_49229,N_49964);
and UO_2017 (O_2017,N_49059,N_49785);
and UO_2018 (O_2018,N_49454,N_49258);
and UO_2019 (O_2019,N_49196,N_49612);
nor UO_2020 (O_2020,N_49406,N_49270);
and UO_2021 (O_2021,N_49821,N_49784);
or UO_2022 (O_2022,N_49278,N_49416);
nor UO_2023 (O_2023,N_49218,N_49280);
nand UO_2024 (O_2024,N_49004,N_49859);
or UO_2025 (O_2025,N_49696,N_49562);
xnor UO_2026 (O_2026,N_49346,N_49310);
nand UO_2027 (O_2027,N_49713,N_49142);
and UO_2028 (O_2028,N_49408,N_49834);
nor UO_2029 (O_2029,N_49602,N_49866);
and UO_2030 (O_2030,N_49934,N_49758);
xnor UO_2031 (O_2031,N_49591,N_49742);
and UO_2032 (O_2032,N_49083,N_49245);
nand UO_2033 (O_2033,N_49540,N_49213);
nand UO_2034 (O_2034,N_49506,N_49032);
xor UO_2035 (O_2035,N_49700,N_49239);
nand UO_2036 (O_2036,N_49273,N_49227);
xor UO_2037 (O_2037,N_49547,N_49311);
nor UO_2038 (O_2038,N_49810,N_49163);
and UO_2039 (O_2039,N_49831,N_49329);
xor UO_2040 (O_2040,N_49444,N_49552);
and UO_2041 (O_2041,N_49939,N_49502);
or UO_2042 (O_2042,N_49974,N_49387);
xnor UO_2043 (O_2043,N_49653,N_49295);
nand UO_2044 (O_2044,N_49479,N_49229);
or UO_2045 (O_2045,N_49726,N_49849);
nor UO_2046 (O_2046,N_49940,N_49208);
xor UO_2047 (O_2047,N_49382,N_49779);
and UO_2048 (O_2048,N_49091,N_49298);
and UO_2049 (O_2049,N_49578,N_49343);
nand UO_2050 (O_2050,N_49224,N_49686);
nor UO_2051 (O_2051,N_49612,N_49794);
nor UO_2052 (O_2052,N_49735,N_49730);
nor UO_2053 (O_2053,N_49932,N_49075);
or UO_2054 (O_2054,N_49498,N_49135);
nand UO_2055 (O_2055,N_49791,N_49199);
xor UO_2056 (O_2056,N_49248,N_49909);
or UO_2057 (O_2057,N_49395,N_49866);
nor UO_2058 (O_2058,N_49617,N_49969);
or UO_2059 (O_2059,N_49264,N_49932);
or UO_2060 (O_2060,N_49983,N_49851);
xnor UO_2061 (O_2061,N_49371,N_49227);
xnor UO_2062 (O_2062,N_49771,N_49850);
xnor UO_2063 (O_2063,N_49153,N_49047);
or UO_2064 (O_2064,N_49987,N_49379);
nor UO_2065 (O_2065,N_49379,N_49596);
xor UO_2066 (O_2066,N_49033,N_49512);
xnor UO_2067 (O_2067,N_49076,N_49014);
and UO_2068 (O_2068,N_49720,N_49483);
xor UO_2069 (O_2069,N_49290,N_49017);
and UO_2070 (O_2070,N_49463,N_49879);
or UO_2071 (O_2071,N_49324,N_49167);
or UO_2072 (O_2072,N_49809,N_49908);
nor UO_2073 (O_2073,N_49291,N_49812);
and UO_2074 (O_2074,N_49012,N_49365);
or UO_2075 (O_2075,N_49613,N_49374);
or UO_2076 (O_2076,N_49754,N_49972);
or UO_2077 (O_2077,N_49914,N_49303);
xnor UO_2078 (O_2078,N_49141,N_49772);
xnor UO_2079 (O_2079,N_49185,N_49240);
and UO_2080 (O_2080,N_49708,N_49680);
or UO_2081 (O_2081,N_49796,N_49971);
xor UO_2082 (O_2082,N_49184,N_49529);
nor UO_2083 (O_2083,N_49904,N_49095);
or UO_2084 (O_2084,N_49321,N_49247);
xor UO_2085 (O_2085,N_49911,N_49844);
nor UO_2086 (O_2086,N_49944,N_49765);
and UO_2087 (O_2087,N_49272,N_49693);
nor UO_2088 (O_2088,N_49755,N_49764);
or UO_2089 (O_2089,N_49779,N_49712);
or UO_2090 (O_2090,N_49235,N_49657);
or UO_2091 (O_2091,N_49522,N_49413);
nor UO_2092 (O_2092,N_49955,N_49736);
nand UO_2093 (O_2093,N_49314,N_49036);
or UO_2094 (O_2094,N_49502,N_49183);
or UO_2095 (O_2095,N_49658,N_49809);
nor UO_2096 (O_2096,N_49721,N_49702);
and UO_2097 (O_2097,N_49719,N_49923);
nand UO_2098 (O_2098,N_49911,N_49155);
and UO_2099 (O_2099,N_49905,N_49187);
xor UO_2100 (O_2100,N_49245,N_49583);
or UO_2101 (O_2101,N_49079,N_49402);
and UO_2102 (O_2102,N_49813,N_49031);
xnor UO_2103 (O_2103,N_49475,N_49008);
or UO_2104 (O_2104,N_49744,N_49698);
nand UO_2105 (O_2105,N_49646,N_49026);
and UO_2106 (O_2106,N_49311,N_49488);
or UO_2107 (O_2107,N_49973,N_49528);
or UO_2108 (O_2108,N_49110,N_49644);
and UO_2109 (O_2109,N_49936,N_49933);
nor UO_2110 (O_2110,N_49476,N_49911);
xor UO_2111 (O_2111,N_49897,N_49419);
xor UO_2112 (O_2112,N_49309,N_49630);
or UO_2113 (O_2113,N_49152,N_49842);
nand UO_2114 (O_2114,N_49195,N_49219);
nand UO_2115 (O_2115,N_49702,N_49788);
and UO_2116 (O_2116,N_49552,N_49419);
or UO_2117 (O_2117,N_49790,N_49470);
xor UO_2118 (O_2118,N_49413,N_49374);
and UO_2119 (O_2119,N_49616,N_49049);
xor UO_2120 (O_2120,N_49742,N_49794);
xor UO_2121 (O_2121,N_49342,N_49950);
xnor UO_2122 (O_2122,N_49427,N_49133);
or UO_2123 (O_2123,N_49221,N_49728);
or UO_2124 (O_2124,N_49321,N_49288);
nor UO_2125 (O_2125,N_49923,N_49651);
and UO_2126 (O_2126,N_49492,N_49887);
or UO_2127 (O_2127,N_49978,N_49505);
xnor UO_2128 (O_2128,N_49976,N_49645);
xnor UO_2129 (O_2129,N_49657,N_49391);
xnor UO_2130 (O_2130,N_49344,N_49869);
xnor UO_2131 (O_2131,N_49379,N_49077);
or UO_2132 (O_2132,N_49151,N_49953);
or UO_2133 (O_2133,N_49653,N_49333);
xnor UO_2134 (O_2134,N_49686,N_49135);
or UO_2135 (O_2135,N_49855,N_49745);
or UO_2136 (O_2136,N_49118,N_49750);
nor UO_2137 (O_2137,N_49611,N_49670);
and UO_2138 (O_2138,N_49878,N_49702);
xor UO_2139 (O_2139,N_49288,N_49934);
xnor UO_2140 (O_2140,N_49169,N_49431);
xnor UO_2141 (O_2141,N_49001,N_49929);
and UO_2142 (O_2142,N_49594,N_49464);
xnor UO_2143 (O_2143,N_49780,N_49728);
and UO_2144 (O_2144,N_49891,N_49334);
nand UO_2145 (O_2145,N_49084,N_49967);
xor UO_2146 (O_2146,N_49942,N_49587);
xnor UO_2147 (O_2147,N_49646,N_49374);
or UO_2148 (O_2148,N_49114,N_49012);
or UO_2149 (O_2149,N_49564,N_49144);
and UO_2150 (O_2150,N_49497,N_49484);
or UO_2151 (O_2151,N_49971,N_49225);
and UO_2152 (O_2152,N_49664,N_49682);
nand UO_2153 (O_2153,N_49093,N_49925);
nor UO_2154 (O_2154,N_49390,N_49093);
nand UO_2155 (O_2155,N_49297,N_49278);
nor UO_2156 (O_2156,N_49544,N_49274);
nand UO_2157 (O_2157,N_49923,N_49975);
and UO_2158 (O_2158,N_49443,N_49708);
and UO_2159 (O_2159,N_49034,N_49623);
nor UO_2160 (O_2160,N_49409,N_49652);
xor UO_2161 (O_2161,N_49498,N_49375);
nor UO_2162 (O_2162,N_49267,N_49617);
xor UO_2163 (O_2163,N_49190,N_49128);
nor UO_2164 (O_2164,N_49624,N_49639);
xnor UO_2165 (O_2165,N_49234,N_49067);
and UO_2166 (O_2166,N_49824,N_49643);
nor UO_2167 (O_2167,N_49440,N_49027);
or UO_2168 (O_2168,N_49605,N_49543);
or UO_2169 (O_2169,N_49707,N_49812);
nand UO_2170 (O_2170,N_49775,N_49188);
nor UO_2171 (O_2171,N_49271,N_49018);
or UO_2172 (O_2172,N_49553,N_49508);
xor UO_2173 (O_2173,N_49121,N_49125);
or UO_2174 (O_2174,N_49239,N_49922);
xnor UO_2175 (O_2175,N_49576,N_49246);
xor UO_2176 (O_2176,N_49067,N_49245);
nand UO_2177 (O_2177,N_49082,N_49929);
nor UO_2178 (O_2178,N_49683,N_49070);
xor UO_2179 (O_2179,N_49300,N_49919);
or UO_2180 (O_2180,N_49761,N_49328);
and UO_2181 (O_2181,N_49138,N_49497);
nor UO_2182 (O_2182,N_49876,N_49329);
nand UO_2183 (O_2183,N_49987,N_49451);
xor UO_2184 (O_2184,N_49325,N_49288);
and UO_2185 (O_2185,N_49087,N_49241);
xor UO_2186 (O_2186,N_49034,N_49176);
or UO_2187 (O_2187,N_49224,N_49288);
nor UO_2188 (O_2188,N_49920,N_49301);
xor UO_2189 (O_2189,N_49354,N_49080);
nor UO_2190 (O_2190,N_49850,N_49302);
nand UO_2191 (O_2191,N_49338,N_49201);
nor UO_2192 (O_2192,N_49493,N_49363);
and UO_2193 (O_2193,N_49800,N_49538);
and UO_2194 (O_2194,N_49209,N_49662);
or UO_2195 (O_2195,N_49158,N_49609);
nor UO_2196 (O_2196,N_49748,N_49364);
or UO_2197 (O_2197,N_49548,N_49126);
nor UO_2198 (O_2198,N_49275,N_49437);
xnor UO_2199 (O_2199,N_49038,N_49635);
xor UO_2200 (O_2200,N_49247,N_49461);
xor UO_2201 (O_2201,N_49856,N_49913);
nor UO_2202 (O_2202,N_49922,N_49002);
or UO_2203 (O_2203,N_49745,N_49616);
or UO_2204 (O_2204,N_49938,N_49395);
nand UO_2205 (O_2205,N_49076,N_49279);
nor UO_2206 (O_2206,N_49289,N_49176);
or UO_2207 (O_2207,N_49295,N_49315);
or UO_2208 (O_2208,N_49553,N_49903);
or UO_2209 (O_2209,N_49801,N_49100);
nand UO_2210 (O_2210,N_49398,N_49616);
nand UO_2211 (O_2211,N_49197,N_49520);
nor UO_2212 (O_2212,N_49502,N_49224);
xnor UO_2213 (O_2213,N_49957,N_49020);
xor UO_2214 (O_2214,N_49888,N_49690);
nor UO_2215 (O_2215,N_49804,N_49999);
nand UO_2216 (O_2216,N_49199,N_49060);
nand UO_2217 (O_2217,N_49763,N_49784);
nand UO_2218 (O_2218,N_49160,N_49883);
and UO_2219 (O_2219,N_49775,N_49809);
xnor UO_2220 (O_2220,N_49855,N_49413);
or UO_2221 (O_2221,N_49451,N_49950);
nor UO_2222 (O_2222,N_49074,N_49601);
nand UO_2223 (O_2223,N_49477,N_49110);
or UO_2224 (O_2224,N_49959,N_49410);
nand UO_2225 (O_2225,N_49415,N_49177);
nor UO_2226 (O_2226,N_49026,N_49942);
or UO_2227 (O_2227,N_49116,N_49097);
nor UO_2228 (O_2228,N_49325,N_49801);
nand UO_2229 (O_2229,N_49008,N_49207);
and UO_2230 (O_2230,N_49558,N_49492);
nand UO_2231 (O_2231,N_49377,N_49616);
or UO_2232 (O_2232,N_49467,N_49287);
and UO_2233 (O_2233,N_49864,N_49214);
and UO_2234 (O_2234,N_49592,N_49301);
nand UO_2235 (O_2235,N_49229,N_49230);
xor UO_2236 (O_2236,N_49274,N_49332);
xnor UO_2237 (O_2237,N_49267,N_49558);
and UO_2238 (O_2238,N_49982,N_49256);
nor UO_2239 (O_2239,N_49494,N_49768);
or UO_2240 (O_2240,N_49193,N_49247);
and UO_2241 (O_2241,N_49439,N_49629);
xor UO_2242 (O_2242,N_49503,N_49482);
and UO_2243 (O_2243,N_49276,N_49352);
or UO_2244 (O_2244,N_49948,N_49382);
nand UO_2245 (O_2245,N_49630,N_49812);
and UO_2246 (O_2246,N_49799,N_49263);
nor UO_2247 (O_2247,N_49164,N_49670);
nor UO_2248 (O_2248,N_49533,N_49320);
or UO_2249 (O_2249,N_49303,N_49860);
and UO_2250 (O_2250,N_49944,N_49112);
nor UO_2251 (O_2251,N_49560,N_49974);
xnor UO_2252 (O_2252,N_49913,N_49277);
nor UO_2253 (O_2253,N_49682,N_49429);
nand UO_2254 (O_2254,N_49708,N_49725);
xor UO_2255 (O_2255,N_49404,N_49320);
or UO_2256 (O_2256,N_49212,N_49424);
nand UO_2257 (O_2257,N_49644,N_49408);
nor UO_2258 (O_2258,N_49642,N_49479);
nor UO_2259 (O_2259,N_49500,N_49211);
nor UO_2260 (O_2260,N_49184,N_49969);
nor UO_2261 (O_2261,N_49123,N_49302);
nor UO_2262 (O_2262,N_49974,N_49002);
xor UO_2263 (O_2263,N_49553,N_49452);
nor UO_2264 (O_2264,N_49926,N_49546);
nor UO_2265 (O_2265,N_49438,N_49412);
nand UO_2266 (O_2266,N_49998,N_49365);
or UO_2267 (O_2267,N_49311,N_49373);
or UO_2268 (O_2268,N_49171,N_49679);
nor UO_2269 (O_2269,N_49493,N_49342);
and UO_2270 (O_2270,N_49681,N_49265);
nand UO_2271 (O_2271,N_49809,N_49459);
and UO_2272 (O_2272,N_49109,N_49888);
xnor UO_2273 (O_2273,N_49413,N_49608);
nand UO_2274 (O_2274,N_49038,N_49542);
and UO_2275 (O_2275,N_49737,N_49402);
or UO_2276 (O_2276,N_49885,N_49746);
and UO_2277 (O_2277,N_49176,N_49763);
xnor UO_2278 (O_2278,N_49483,N_49102);
nor UO_2279 (O_2279,N_49762,N_49455);
and UO_2280 (O_2280,N_49584,N_49778);
nor UO_2281 (O_2281,N_49228,N_49748);
or UO_2282 (O_2282,N_49860,N_49917);
and UO_2283 (O_2283,N_49213,N_49150);
nand UO_2284 (O_2284,N_49494,N_49003);
xor UO_2285 (O_2285,N_49081,N_49495);
nand UO_2286 (O_2286,N_49984,N_49060);
nor UO_2287 (O_2287,N_49020,N_49849);
xor UO_2288 (O_2288,N_49852,N_49267);
nor UO_2289 (O_2289,N_49775,N_49807);
nor UO_2290 (O_2290,N_49236,N_49409);
nand UO_2291 (O_2291,N_49439,N_49130);
and UO_2292 (O_2292,N_49306,N_49673);
xor UO_2293 (O_2293,N_49592,N_49044);
and UO_2294 (O_2294,N_49994,N_49732);
xor UO_2295 (O_2295,N_49739,N_49605);
nor UO_2296 (O_2296,N_49645,N_49383);
nand UO_2297 (O_2297,N_49942,N_49817);
nor UO_2298 (O_2298,N_49657,N_49727);
xnor UO_2299 (O_2299,N_49194,N_49881);
and UO_2300 (O_2300,N_49645,N_49439);
nand UO_2301 (O_2301,N_49195,N_49375);
nor UO_2302 (O_2302,N_49373,N_49050);
xor UO_2303 (O_2303,N_49401,N_49549);
and UO_2304 (O_2304,N_49466,N_49825);
or UO_2305 (O_2305,N_49316,N_49795);
or UO_2306 (O_2306,N_49443,N_49621);
or UO_2307 (O_2307,N_49421,N_49823);
and UO_2308 (O_2308,N_49710,N_49033);
or UO_2309 (O_2309,N_49769,N_49968);
nor UO_2310 (O_2310,N_49331,N_49042);
and UO_2311 (O_2311,N_49270,N_49540);
nor UO_2312 (O_2312,N_49970,N_49213);
and UO_2313 (O_2313,N_49998,N_49947);
or UO_2314 (O_2314,N_49429,N_49132);
and UO_2315 (O_2315,N_49891,N_49122);
xnor UO_2316 (O_2316,N_49965,N_49731);
xor UO_2317 (O_2317,N_49397,N_49375);
or UO_2318 (O_2318,N_49151,N_49395);
and UO_2319 (O_2319,N_49630,N_49338);
and UO_2320 (O_2320,N_49645,N_49809);
and UO_2321 (O_2321,N_49360,N_49689);
xor UO_2322 (O_2322,N_49616,N_49434);
nand UO_2323 (O_2323,N_49568,N_49271);
nor UO_2324 (O_2324,N_49103,N_49540);
or UO_2325 (O_2325,N_49969,N_49372);
or UO_2326 (O_2326,N_49489,N_49435);
and UO_2327 (O_2327,N_49429,N_49231);
nor UO_2328 (O_2328,N_49081,N_49576);
or UO_2329 (O_2329,N_49620,N_49474);
or UO_2330 (O_2330,N_49160,N_49836);
xor UO_2331 (O_2331,N_49213,N_49679);
or UO_2332 (O_2332,N_49328,N_49919);
xnor UO_2333 (O_2333,N_49357,N_49210);
xnor UO_2334 (O_2334,N_49396,N_49789);
and UO_2335 (O_2335,N_49842,N_49799);
nand UO_2336 (O_2336,N_49460,N_49176);
nand UO_2337 (O_2337,N_49127,N_49914);
and UO_2338 (O_2338,N_49002,N_49228);
or UO_2339 (O_2339,N_49724,N_49844);
nor UO_2340 (O_2340,N_49841,N_49788);
and UO_2341 (O_2341,N_49721,N_49820);
xor UO_2342 (O_2342,N_49726,N_49749);
and UO_2343 (O_2343,N_49873,N_49257);
or UO_2344 (O_2344,N_49654,N_49986);
nand UO_2345 (O_2345,N_49560,N_49561);
nor UO_2346 (O_2346,N_49992,N_49009);
xnor UO_2347 (O_2347,N_49156,N_49167);
nor UO_2348 (O_2348,N_49942,N_49635);
or UO_2349 (O_2349,N_49319,N_49811);
or UO_2350 (O_2350,N_49944,N_49767);
xor UO_2351 (O_2351,N_49772,N_49600);
nand UO_2352 (O_2352,N_49330,N_49045);
nand UO_2353 (O_2353,N_49447,N_49990);
or UO_2354 (O_2354,N_49002,N_49668);
xor UO_2355 (O_2355,N_49853,N_49263);
nor UO_2356 (O_2356,N_49923,N_49184);
nor UO_2357 (O_2357,N_49917,N_49316);
nor UO_2358 (O_2358,N_49266,N_49423);
or UO_2359 (O_2359,N_49346,N_49055);
nor UO_2360 (O_2360,N_49090,N_49852);
xnor UO_2361 (O_2361,N_49823,N_49573);
or UO_2362 (O_2362,N_49197,N_49404);
nor UO_2363 (O_2363,N_49599,N_49070);
nor UO_2364 (O_2364,N_49419,N_49282);
nand UO_2365 (O_2365,N_49662,N_49615);
xor UO_2366 (O_2366,N_49560,N_49661);
or UO_2367 (O_2367,N_49907,N_49807);
and UO_2368 (O_2368,N_49036,N_49225);
nand UO_2369 (O_2369,N_49905,N_49098);
and UO_2370 (O_2370,N_49070,N_49118);
or UO_2371 (O_2371,N_49154,N_49348);
nor UO_2372 (O_2372,N_49639,N_49473);
xnor UO_2373 (O_2373,N_49920,N_49978);
nor UO_2374 (O_2374,N_49776,N_49412);
or UO_2375 (O_2375,N_49219,N_49317);
nand UO_2376 (O_2376,N_49200,N_49814);
and UO_2377 (O_2377,N_49415,N_49834);
nand UO_2378 (O_2378,N_49678,N_49551);
nor UO_2379 (O_2379,N_49296,N_49333);
or UO_2380 (O_2380,N_49494,N_49305);
xnor UO_2381 (O_2381,N_49466,N_49285);
nand UO_2382 (O_2382,N_49428,N_49523);
nand UO_2383 (O_2383,N_49206,N_49853);
xor UO_2384 (O_2384,N_49995,N_49016);
xor UO_2385 (O_2385,N_49667,N_49097);
nand UO_2386 (O_2386,N_49555,N_49489);
nor UO_2387 (O_2387,N_49451,N_49761);
xor UO_2388 (O_2388,N_49448,N_49343);
xor UO_2389 (O_2389,N_49412,N_49892);
xor UO_2390 (O_2390,N_49362,N_49223);
nor UO_2391 (O_2391,N_49230,N_49797);
and UO_2392 (O_2392,N_49233,N_49767);
or UO_2393 (O_2393,N_49380,N_49092);
xnor UO_2394 (O_2394,N_49117,N_49662);
and UO_2395 (O_2395,N_49824,N_49622);
and UO_2396 (O_2396,N_49036,N_49660);
nor UO_2397 (O_2397,N_49695,N_49715);
nor UO_2398 (O_2398,N_49208,N_49636);
and UO_2399 (O_2399,N_49488,N_49501);
nor UO_2400 (O_2400,N_49387,N_49168);
nor UO_2401 (O_2401,N_49697,N_49801);
nand UO_2402 (O_2402,N_49198,N_49346);
and UO_2403 (O_2403,N_49195,N_49415);
or UO_2404 (O_2404,N_49483,N_49282);
nand UO_2405 (O_2405,N_49488,N_49944);
or UO_2406 (O_2406,N_49056,N_49813);
xnor UO_2407 (O_2407,N_49653,N_49302);
or UO_2408 (O_2408,N_49336,N_49853);
and UO_2409 (O_2409,N_49586,N_49337);
or UO_2410 (O_2410,N_49038,N_49869);
nor UO_2411 (O_2411,N_49624,N_49786);
xor UO_2412 (O_2412,N_49014,N_49166);
or UO_2413 (O_2413,N_49472,N_49436);
nor UO_2414 (O_2414,N_49994,N_49695);
nand UO_2415 (O_2415,N_49563,N_49052);
xor UO_2416 (O_2416,N_49621,N_49955);
xnor UO_2417 (O_2417,N_49460,N_49426);
xnor UO_2418 (O_2418,N_49423,N_49906);
or UO_2419 (O_2419,N_49286,N_49380);
nor UO_2420 (O_2420,N_49937,N_49938);
and UO_2421 (O_2421,N_49367,N_49801);
nor UO_2422 (O_2422,N_49530,N_49177);
xnor UO_2423 (O_2423,N_49194,N_49936);
or UO_2424 (O_2424,N_49800,N_49460);
nor UO_2425 (O_2425,N_49613,N_49581);
or UO_2426 (O_2426,N_49098,N_49606);
xor UO_2427 (O_2427,N_49745,N_49683);
nor UO_2428 (O_2428,N_49077,N_49286);
nor UO_2429 (O_2429,N_49432,N_49974);
and UO_2430 (O_2430,N_49480,N_49779);
nand UO_2431 (O_2431,N_49083,N_49021);
nand UO_2432 (O_2432,N_49517,N_49676);
xor UO_2433 (O_2433,N_49693,N_49508);
xnor UO_2434 (O_2434,N_49914,N_49021);
nand UO_2435 (O_2435,N_49169,N_49120);
nand UO_2436 (O_2436,N_49073,N_49946);
xor UO_2437 (O_2437,N_49911,N_49482);
xnor UO_2438 (O_2438,N_49563,N_49875);
and UO_2439 (O_2439,N_49248,N_49768);
and UO_2440 (O_2440,N_49486,N_49572);
or UO_2441 (O_2441,N_49396,N_49593);
and UO_2442 (O_2442,N_49070,N_49915);
and UO_2443 (O_2443,N_49272,N_49524);
and UO_2444 (O_2444,N_49227,N_49474);
or UO_2445 (O_2445,N_49955,N_49879);
and UO_2446 (O_2446,N_49826,N_49335);
xnor UO_2447 (O_2447,N_49831,N_49658);
nor UO_2448 (O_2448,N_49401,N_49784);
nand UO_2449 (O_2449,N_49513,N_49360);
nand UO_2450 (O_2450,N_49891,N_49277);
and UO_2451 (O_2451,N_49408,N_49783);
or UO_2452 (O_2452,N_49757,N_49700);
xor UO_2453 (O_2453,N_49363,N_49411);
nor UO_2454 (O_2454,N_49652,N_49899);
xor UO_2455 (O_2455,N_49900,N_49918);
nor UO_2456 (O_2456,N_49926,N_49334);
nor UO_2457 (O_2457,N_49330,N_49586);
nand UO_2458 (O_2458,N_49521,N_49443);
nor UO_2459 (O_2459,N_49034,N_49697);
nand UO_2460 (O_2460,N_49943,N_49319);
xnor UO_2461 (O_2461,N_49777,N_49210);
or UO_2462 (O_2462,N_49952,N_49889);
xor UO_2463 (O_2463,N_49488,N_49387);
and UO_2464 (O_2464,N_49945,N_49579);
nor UO_2465 (O_2465,N_49056,N_49348);
nand UO_2466 (O_2466,N_49752,N_49259);
and UO_2467 (O_2467,N_49162,N_49425);
and UO_2468 (O_2468,N_49725,N_49393);
nor UO_2469 (O_2469,N_49311,N_49941);
nand UO_2470 (O_2470,N_49741,N_49554);
or UO_2471 (O_2471,N_49889,N_49426);
nor UO_2472 (O_2472,N_49529,N_49403);
xor UO_2473 (O_2473,N_49412,N_49884);
nor UO_2474 (O_2474,N_49300,N_49615);
nand UO_2475 (O_2475,N_49849,N_49695);
and UO_2476 (O_2476,N_49273,N_49004);
or UO_2477 (O_2477,N_49128,N_49181);
or UO_2478 (O_2478,N_49950,N_49788);
and UO_2479 (O_2479,N_49167,N_49863);
xor UO_2480 (O_2480,N_49089,N_49975);
nor UO_2481 (O_2481,N_49742,N_49125);
nand UO_2482 (O_2482,N_49624,N_49884);
xnor UO_2483 (O_2483,N_49803,N_49474);
and UO_2484 (O_2484,N_49617,N_49878);
or UO_2485 (O_2485,N_49465,N_49730);
nand UO_2486 (O_2486,N_49918,N_49468);
nand UO_2487 (O_2487,N_49947,N_49688);
nor UO_2488 (O_2488,N_49166,N_49325);
xnor UO_2489 (O_2489,N_49373,N_49320);
or UO_2490 (O_2490,N_49525,N_49375);
nor UO_2491 (O_2491,N_49652,N_49308);
nand UO_2492 (O_2492,N_49682,N_49407);
or UO_2493 (O_2493,N_49645,N_49367);
nor UO_2494 (O_2494,N_49229,N_49316);
nand UO_2495 (O_2495,N_49165,N_49558);
xnor UO_2496 (O_2496,N_49749,N_49493);
nor UO_2497 (O_2497,N_49233,N_49218);
or UO_2498 (O_2498,N_49185,N_49116);
and UO_2499 (O_2499,N_49412,N_49153);
xor UO_2500 (O_2500,N_49862,N_49261);
nand UO_2501 (O_2501,N_49474,N_49030);
xnor UO_2502 (O_2502,N_49965,N_49060);
and UO_2503 (O_2503,N_49002,N_49199);
xor UO_2504 (O_2504,N_49191,N_49420);
or UO_2505 (O_2505,N_49479,N_49980);
nand UO_2506 (O_2506,N_49339,N_49863);
nand UO_2507 (O_2507,N_49344,N_49979);
or UO_2508 (O_2508,N_49471,N_49172);
and UO_2509 (O_2509,N_49586,N_49441);
or UO_2510 (O_2510,N_49491,N_49886);
nand UO_2511 (O_2511,N_49008,N_49439);
xor UO_2512 (O_2512,N_49772,N_49043);
nand UO_2513 (O_2513,N_49622,N_49936);
nor UO_2514 (O_2514,N_49953,N_49303);
and UO_2515 (O_2515,N_49812,N_49584);
xnor UO_2516 (O_2516,N_49763,N_49232);
and UO_2517 (O_2517,N_49417,N_49573);
and UO_2518 (O_2518,N_49900,N_49740);
nor UO_2519 (O_2519,N_49561,N_49647);
nor UO_2520 (O_2520,N_49395,N_49946);
nor UO_2521 (O_2521,N_49584,N_49944);
and UO_2522 (O_2522,N_49301,N_49018);
and UO_2523 (O_2523,N_49085,N_49417);
nand UO_2524 (O_2524,N_49351,N_49331);
or UO_2525 (O_2525,N_49714,N_49220);
or UO_2526 (O_2526,N_49462,N_49475);
nand UO_2527 (O_2527,N_49240,N_49388);
or UO_2528 (O_2528,N_49841,N_49653);
or UO_2529 (O_2529,N_49786,N_49752);
nor UO_2530 (O_2530,N_49997,N_49503);
or UO_2531 (O_2531,N_49253,N_49388);
xor UO_2532 (O_2532,N_49737,N_49067);
or UO_2533 (O_2533,N_49871,N_49975);
or UO_2534 (O_2534,N_49176,N_49393);
nor UO_2535 (O_2535,N_49907,N_49388);
and UO_2536 (O_2536,N_49220,N_49438);
xor UO_2537 (O_2537,N_49322,N_49701);
xnor UO_2538 (O_2538,N_49907,N_49722);
or UO_2539 (O_2539,N_49805,N_49367);
or UO_2540 (O_2540,N_49472,N_49905);
nor UO_2541 (O_2541,N_49375,N_49580);
nand UO_2542 (O_2542,N_49180,N_49225);
nand UO_2543 (O_2543,N_49144,N_49229);
or UO_2544 (O_2544,N_49473,N_49707);
or UO_2545 (O_2545,N_49787,N_49131);
xnor UO_2546 (O_2546,N_49265,N_49237);
nor UO_2547 (O_2547,N_49804,N_49946);
xnor UO_2548 (O_2548,N_49688,N_49455);
xnor UO_2549 (O_2549,N_49119,N_49921);
or UO_2550 (O_2550,N_49903,N_49510);
xor UO_2551 (O_2551,N_49727,N_49399);
and UO_2552 (O_2552,N_49387,N_49530);
xor UO_2553 (O_2553,N_49272,N_49988);
nor UO_2554 (O_2554,N_49016,N_49182);
or UO_2555 (O_2555,N_49508,N_49841);
nand UO_2556 (O_2556,N_49123,N_49842);
nor UO_2557 (O_2557,N_49380,N_49364);
and UO_2558 (O_2558,N_49648,N_49944);
or UO_2559 (O_2559,N_49041,N_49004);
and UO_2560 (O_2560,N_49518,N_49847);
nand UO_2561 (O_2561,N_49908,N_49286);
and UO_2562 (O_2562,N_49101,N_49713);
xor UO_2563 (O_2563,N_49059,N_49931);
nor UO_2564 (O_2564,N_49271,N_49715);
or UO_2565 (O_2565,N_49541,N_49049);
nor UO_2566 (O_2566,N_49228,N_49825);
and UO_2567 (O_2567,N_49005,N_49234);
xor UO_2568 (O_2568,N_49975,N_49753);
xnor UO_2569 (O_2569,N_49801,N_49471);
or UO_2570 (O_2570,N_49398,N_49732);
and UO_2571 (O_2571,N_49581,N_49592);
nand UO_2572 (O_2572,N_49042,N_49746);
and UO_2573 (O_2573,N_49824,N_49561);
xor UO_2574 (O_2574,N_49503,N_49760);
and UO_2575 (O_2575,N_49349,N_49168);
nand UO_2576 (O_2576,N_49202,N_49019);
nand UO_2577 (O_2577,N_49798,N_49654);
nor UO_2578 (O_2578,N_49185,N_49507);
nor UO_2579 (O_2579,N_49304,N_49706);
or UO_2580 (O_2580,N_49058,N_49758);
xnor UO_2581 (O_2581,N_49645,N_49126);
and UO_2582 (O_2582,N_49273,N_49881);
or UO_2583 (O_2583,N_49926,N_49287);
nor UO_2584 (O_2584,N_49202,N_49721);
or UO_2585 (O_2585,N_49430,N_49557);
xor UO_2586 (O_2586,N_49674,N_49318);
and UO_2587 (O_2587,N_49643,N_49568);
nor UO_2588 (O_2588,N_49870,N_49766);
xor UO_2589 (O_2589,N_49194,N_49006);
nor UO_2590 (O_2590,N_49854,N_49452);
and UO_2591 (O_2591,N_49506,N_49405);
and UO_2592 (O_2592,N_49073,N_49650);
nor UO_2593 (O_2593,N_49437,N_49424);
and UO_2594 (O_2594,N_49682,N_49017);
or UO_2595 (O_2595,N_49452,N_49319);
or UO_2596 (O_2596,N_49620,N_49702);
nand UO_2597 (O_2597,N_49333,N_49176);
or UO_2598 (O_2598,N_49428,N_49130);
and UO_2599 (O_2599,N_49665,N_49092);
nand UO_2600 (O_2600,N_49336,N_49525);
or UO_2601 (O_2601,N_49250,N_49469);
and UO_2602 (O_2602,N_49901,N_49074);
or UO_2603 (O_2603,N_49842,N_49941);
nand UO_2604 (O_2604,N_49272,N_49819);
and UO_2605 (O_2605,N_49891,N_49998);
and UO_2606 (O_2606,N_49153,N_49704);
nor UO_2607 (O_2607,N_49507,N_49304);
or UO_2608 (O_2608,N_49608,N_49110);
or UO_2609 (O_2609,N_49583,N_49441);
nand UO_2610 (O_2610,N_49733,N_49996);
xor UO_2611 (O_2611,N_49594,N_49249);
xnor UO_2612 (O_2612,N_49755,N_49461);
xor UO_2613 (O_2613,N_49077,N_49866);
and UO_2614 (O_2614,N_49066,N_49655);
nand UO_2615 (O_2615,N_49506,N_49284);
xor UO_2616 (O_2616,N_49857,N_49230);
nand UO_2617 (O_2617,N_49545,N_49886);
xnor UO_2618 (O_2618,N_49025,N_49122);
nand UO_2619 (O_2619,N_49949,N_49385);
nor UO_2620 (O_2620,N_49303,N_49124);
or UO_2621 (O_2621,N_49959,N_49684);
nor UO_2622 (O_2622,N_49112,N_49750);
and UO_2623 (O_2623,N_49643,N_49839);
xnor UO_2624 (O_2624,N_49435,N_49481);
or UO_2625 (O_2625,N_49882,N_49755);
and UO_2626 (O_2626,N_49372,N_49106);
nand UO_2627 (O_2627,N_49229,N_49002);
xor UO_2628 (O_2628,N_49928,N_49926);
xor UO_2629 (O_2629,N_49205,N_49750);
nand UO_2630 (O_2630,N_49005,N_49489);
and UO_2631 (O_2631,N_49250,N_49311);
or UO_2632 (O_2632,N_49966,N_49253);
nor UO_2633 (O_2633,N_49096,N_49571);
and UO_2634 (O_2634,N_49195,N_49404);
or UO_2635 (O_2635,N_49329,N_49935);
and UO_2636 (O_2636,N_49817,N_49169);
nand UO_2637 (O_2637,N_49483,N_49319);
xor UO_2638 (O_2638,N_49590,N_49500);
nand UO_2639 (O_2639,N_49897,N_49318);
nor UO_2640 (O_2640,N_49562,N_49336);
nor UO_2641 (O_2641,N_49218,N_49315);
and UO_2642 (O_2642,N_49469,N_49899);
xor UO_2643 (O_2643,N_49341,N_49947);
and UO_2644 (O_2644,N_49925,N_49778);
or UO_2645 (O_2645,N_49468,N_49718);
xor UO_2646 (O_2646,N_49127,N_49573);
or UO_2647 (O_2647,N_49627,N_49545);
or UO_2648 (O_2648,N_49199,N_49506);
xor UO_2649 (O_2649,N_49907,N_49865);
and UO_2650 (O_2650,N_49601,N_49153);
nor UO_2651 (O_2651,N_49987,N_49719);
nand UO_2652 (O_2652,N_49867,N_49193);
xor UO_2653 (O_2653,N_49589,N_49579);
and UO_2654 (O_2654,N_49345,N_49563);
or UO_2655 (O_2655,N_49740,N_49375);
and UO_2656 (O_2656,N_49233,N_49736);
xor UO_2657 (O_2657,N_49427,N_49941);
and UO_2658 (O_2658,N_49869,N_49734);
and UO_2659 (O_2659,N_49114,N_49940);
xor UO_2660 (O_2660,N_49313,N_49492);
nand UO_2661 (O_2661,N_49324,N_49072);
and UO_2662 (O_2662,N_49165,N_49483);
or UO_2663 (O_2663,N_49112,N_49240);
nor UO_2664 (O_2664,N_49180,N_49741);
or UO_2665 (O_2665,N_49454,N_49843);
and UO_2666 (O_2666,N_49723,N_49781);
and UO_2667 (O_2667,N_49144,N_49335);
xor UO_2668 (O_2668,N_49694,N_49516);
nor UO_2669 (O_2669,N_49411,N_49804);
or UO_2670 (O_2670,N_49433,N_49946);
or UO_2671 (O_2671,N_49993,N_49542);
nand UO_2672 (O_2672,N_49895,N_49447);
nor UO_2673 (O_2673,N_49346,N_49379);
and UO_2674 (O_2674,N_49091,N_49183);
xor UO_2675 (O_2675,N_49300,N_49745);
nand UO_2676 (O_2676,N_49785,N_49687);
nand UO_2677 (O_2677,N_49677,N_49460);
and UO_2678 (O_2678,N_49790,N_49705);
nor UO_2679 (O_2679,N_49666,N_49623);
nand UO_2680 (O_2680,N_49508,N_49235);
and UO_2681 (O_2681,N_49247,N_49848);
nand UO_2682 (O_2682,N_49647,N_49376);
nand UO_2683 (O_2683,N_49175,N_49153);
nand UO_2684 (O_2684,N_49806,N_49931);
xnor UO_2685 (O_2685,N_49393,N_49485);
xnor UO_2686 (O_2686,N_49670,N_49089);
or UO_2687 (O_2687,N_49087,N_49229);
or UO_2688 (O_2688,N_49123,N_49630);
or UO_2689 (O_2689,N_49158,N_49508);
xnor UO_2690 (O_2690,N_49132,N_49090);
nand UO_2691 (O_2691,N_49359,N_49856);
or UO_2692 (O_2692,N_49965,N_49508);
or UO_2693 (O_2693,N_49832,N_49606);
xor UO_2694 (O_2694,N_49133,N_49499);
or UO_2695 (O_2695,N_49462,N_49850);
and UO_2696 (O_2696,N_49984,N_49134);
or UO_2697 (O_2697,N_49735,N_49947);
xnor UO_2698 (O_2698,N_49345,N_49198);
nor UO_2699 (O_2699,N_49018,N_49263);
nand UO_2700 (O_2700,N_49470,N_49761);
nor UO_2701 (O_2701,N_49140,N_49271);
or UO_2702 (O_2702,N_49324,N_49038);
nor UO_2703 (O_2703,N_49944,N_49935);
and UO_2704 (O_2704,N_49439,N_49754);
or UO_2705 (O_2705,N_49337,N_49985);
and UO_2706 (O_2706,N_49122,N_49197);
or UO_2707 (O_2707,N_49400,N_49211);
nor UO_2708 (O_2708,N_49042,N_49485);
xnor UO_2709 (O_2709,N_49100,N_49281);
xnor UO_2710 (O_2710,N_49398,N_49479);
and UO_2711 (O_2711,N_49766,N_49980);
and UO_2712 (O_2712,N_49942,N_49975);
or UO_2713 (O_2713,N_49334,N_49707);
or UO_2714 (O_2714,N_49704,N_49711);
and UO_2715 (O_2715,N_49737,N_49158);
nor UO_2716 (O_2716,N_49597,N_49412);
or UO_2717 (O_2717,N_49527,N_49500);
xnor UO_2718 (O_2718,N_49019,N_49853);
nor UO_2719 (O_2719,N_49117,N_49532);
xor UO_2720 (O_2720,N_49586,N_49536);
xnor UO_2721 (O_2721,N_49497,N_49263);
nor UO_2722 (O_2722,N_49294,N_49798);
xor UO_2723 (O_2723,N_49176,N_49500);
nor UO_2724 (O_2724,N_49329,N_49772);
and UO_2725 (O_2725,N_49738,N_49923);
or UO_2726 (O_2726,N_49757,N_49891);
or UO_2727 (O_2727,N_49036,N_49201);
xor UO_2728 (O_2728,N_49064,N_49672);
or UO_2729 (O_2729,N_49759,N_49568);
xor UO_2730 (O_2730,N_49574,N_49624);
xnor UO_2731 (O_2731,N_49112,N_49069);
nand UO_2732 (O_2732,N_49912,N_49704);
nand UO_2733 (O_2733,N_49932,N_49776);
or UO_2734 (O_2734,N_49636,N_49204);
nand UO_2735 (O_2735,N_49136,N_49057);
and UO_2736 (O_2736,N_49623,N_49843);
and UO_2737 (O_2737,N_49818,N_49164);
or UO_2738 (O_2738,N_49770,N_49350);
nand UO_2739 (O_2739,N_49292,N_49449);
nand UO_2740 (O_2740,N_49466,N_49602);
or UO_2741 (O_2741,N_49123,N_49026);
or UO_2742 (O_2742,N_49639,N_49537);
and UO_2743 (O_2743,N_49364,N_49383);
and UO_2744 (O_2744,N_49489,N_49566);
or UO_2745 (O_2745,N_49321,N_49989);
nor UO_2746 (O_2746,N_49263,N_49244);
and UO_2747 (O_2747,N_49447,N_49779);
and UO_2748 (O_2748,N_49058,N_49794);
and UO_2749 (O_2749,N_49437,N_49535);
or UO_2750 (O_2750,N_49666,N_49959);
nand UO_2751 (O_2751,N_49249,N_49248);
nand UO_2752 (O_2752,N_49135,N_49053);
or UO_2753 (O_2753,N_49088,N_49871);
xnor UO_2754 (O_2754,N_49953,N_49735);
or UO_2755 (O_2755,N_49829,N_49150);
and UO_2756 (O_2756,N_49375,N_49321);
nor UO_2757 (O_2757,N_49928,N_49224);
nand UO_2758 (O_2758,N_49675,N_49331);
and UO_2759 (O_2759,N_49581,N_49202);
nor UO_2760 (O_2760,N_49280,N_49095);
nand UO_2761 (O_2761,N_49461,N_49652);
and UO_2762 (O_2762,N_49243,N_49855);
nand UO_2763 (O_2763,N_49775,N_49361);
and UO_2764 (O_2764,N_49574,N_49649);
nand UO_2765 (O_2765,N_49975,N_49703);
or UO_2766 (O_2766,N_49398,N_49080);
nor UO_2767 (O_2767,N_49573,N_49273);
xnor UO_2768 (O_2768,N_49203,N_49495);
nand UO_2769 (O_2769,N_49137,N_49624);
xnor UO_2770 (O_2770,N_49327,N_49044);
xnor UO_2771 (O_2771,N_49554,N_49060);
and UO_2772 (O_2772,N_49729,N_49029);
and UO_2773 (O_2773,N_49355,N_49062);
and UO_2774 (O_2774,N_49708,N_49198);
and UO_2775 (O_2775,N_49915,N_49910);
xnor UO_2776 (O_2776,N_49376,N_49821);
nand UO_2777 (O_2777,N_49239,N_49109);
nand UO_2778 (O_2778,N_49929,N_49961);
nor UO_2779 (O_2779,N_49742,N_49980);
xor UO_2780 (O_2780,N_49522,N_49280);
nor UO_2781 (O_2781,N_49685,N_49565);
nand UO_2782 (O_2782,N_49827,N_49265);
and UO_2783 (O_2783,N_49591,N_49935);
or UO_2784 (O_2784,N_49988,N_49727);
or UO_2785 (O_2785,N_49307,N_49405);
nor UO_2786 (O_2786,N_49067,N_49243);
nor UO_2787 (O_2787,N_49578,N_49724);
xnor UO_2788 (O_2788,N_49042,N_49785);
nand UO_2789 (O_2789,N_49370,N_49034);
nor UO_2790 (O_2790,N_49980,N_49089);
or UO_2791 (O_2791,N_49744,N_49658);
xnor UO_2792 (O_2792,N_49666,N_49957);
or UO_2793 (O_2793,N_49453,N_49897);
and UO_2794 (O_2794,N_49182,N_49827);
and UO_2795 (O_2795,N_49705,N_49183);
nand UO_2796 (O_2796,N_49605,N_49644);
xor UO_2797 (O_2797,N_49318,N_49132);
and UO_2798 (O_2798,N_49602,N_49499);
or UO_2799 (O_2799,N_49933,N_49881);
nand UO_2800 (O_2800,N_49995,N_49787);
or UO_2801 (O_2801,N_49721,N_49502);
xor UO_2802 (O_2802,N_49130,N_49033);
and UO_2803 (O_2803,N_49758,N_49856);
or UO_2804 (O_2804,N_49443,N_49397);
or UO_2805 (O_2805,N_49780,N_49211);
nor UO_2806 (O_2806,N_49212,N_49837);
and UO_2807 (O_2807,N_49076,N_49682);
or UO_2808 (O_2808,N_49473,N_49316);
nor UO_2809 (O_2809,N_49716,N_49026);
nor UO_2810 (O_2810,N_49191,N_49224);
nand UO_2811 (O_2811,N_49754,N_49772);
or UO_2812 (O_2812,N_49917,N_49744);
nor UO_2813 (O_2813,N_49353,N_49463);
or UO_2814 (O_2814,N_49120,N_49761);
nand UO_2815 (O_2815,N_49363,N_49746);
nand UO_2816 (O_2816,N_49869,N_49022);
nand UO_2817 (O_2817,N_49731,N_49294);
nand UO_2818 (O_2818,N_49895,N_49977);
nor UO_2819 (O_2819,N_49244,N_49769);
or UO_2820 (O_2820,N_49754,N_49357);
xor UO_2821 (O_2821,N_49076,N_49045);
nor UO_2822 (O_2822,N_49540,N_49260);
nand UO_2823 (O_2823,N_49836,N_49870);
nand UO_2824 (O_2824,N_49234,N_49461);
nor UO_2825 (O_2825,N_49424,N_49559);
or UO_2826 (O_2826,N_49653,N_49978);
and UO_2827 (O_2827,N_49514,N_49083);
nand UO_2828 (O_2828,N_49895,N_49327);
and UO_2829 (O_2829,N_49245,N_49698);
nor UO_2830 (O_2830,N_49196,N_49372);
nor UO_2831 (O_2831,N_49076,N_49603);
nand UO_2832 (O_2832,N_49617,N_49296);
xor UO_2833 (O_2833,N_49504,N_49017);
nand UO_2834 (O_2834,N_49551,N_49721);
or UO_2835 (O_2835,N_49255,N_49496);
xor UO_2836 (O_2836,N_49752,N_49022);
nor UO_2837 (O_2837,N_49837,N_49132);
nor UO_2838 (O_2838,N_49426,N_49786);
or UO_2839 (O_2839,N_49006,N_49131);
or UO_2840 (O_2840,N_49621,N_49672);
xor UO_2841 (O_2841,N_49255,N_49017);
or UO_2842 (O_2842,N_49533,N_49538);
xnor UO_2843 (O_2843,N_49782,N_49529);
and UO_2844 (O_2844,N_49388,N_49604);
xnor UO_2845 (O_2845,N_49679,N_49920);
xor UO_2846 (O_2846,N_49585,N_49405);
nor UO_2847 (O_2847,N_49351,N_49200);
nand UO_2848 (O_2848,N_49889,N_49694);
and UO_2849 (O_2849,N_49951,N_49095);
nand UO_2850 (O_2850,N_49691,N_49023);
or UO_2851 (O_2851,N_49007,N_49129);
or UO_2852 (O_2852,N_49082,N_49646);
xnor UO_2853 (O_2853,N_49473,N_49727);
or UO_2854 (O_2854,N_49482,N_49196);
or UO_2855 (O_2855,N_49043,N_49619);
nand UO_2856 (O_2856,N_49208,N_49645);
nand UO_2857 (O_2857,N_49393,N_49225);
xnor UO_2858 (O_2858,N_49465,N_49043);
nand UO_2859 (O_2859,N_49057,N_49522);
nor UO_2860 (O_2860,N_49909,N_49972);
nand UO_2861 (O_2861,N_49953,N_49060);
nand UO_2862 (O_2862,N_49202,N_49993);
nand UO_2863 (O_2863,N_49228,N_49835);
or UO_2864 (O_2864,N_49624,N_49170);
or UO_2865 (O_2865,N_49985,N_49130);
or UO_2866 (O_2866,N_49250,N_49424);
xnor UO_2867 (O_2867,N_49107,N_49584);
nor UO_2868 (O_2868,N_49924,N_49300);
or UO_2869 (O_2869,N_49423,N_49267);
and UO_2870 (O_2870,N_49674,N_49692);
or UO_2871 (O_2871,N_49507,N_49087);
and UO_2872 (O_2872,N_49569,N_49389);
nand UO_2873 (O_2873,N_49012,N_49202);
nand UO_2874 (O_2874,N_49572,N_49138);
nand UO_2875 (O_2875,N_49044,N_49952);
nand UO_2876 (O_2876,N_49301,N_49172);
nand UO_2877 (O_2877,N_49312,N_49642);
nand UO_2878 (O_2878,N_49968,N_49904);
xor UO_2879 (O_2879,N_49756,N_49323);
xnor UO_2880 (O_2880,N_49435,N_49674);
or UO_2881 (O_2881,N_49471,N_49209);
or UO_2882 (O_2882,N_49217,N_49182);
nand UO_2883 (O_2883,N_49178,N_49030);
nor UO_2884 (O_2884,N_49070,N_49374);
nand UO_2885 (O_2885,N_49561,N_49707);
or UO_2886 (O_2886,N_49018,N_49162);
and UO_2887 (O_2887,N_49642,N_49821);
nor UO_2888 (O_2888,N_49288,N_49197);
nand UO_2889 (O_2889,N_49097,N_49729);
or UO_2890 (O_2890,N_49890,N_49741);
xnor UO_2891 (O_2891,N_49955,N_49376);
or UO_2892 (O_2892,N_49640,N_49633);
and UO_2893 (O_2893,N_49052,N_49744);
nor UO_2894 (O_2894,N_49991,N_49701);
nor UO_2895 (O_2895,N_49266,N_49369);
xnor UO_2896 (O_2896,N_49901,N_49588);
nor UO_2897 (O_2897,N_49927,N_49358);
nand UO_2898 (O_2898,N_49723,N_49579);
or UO_2899 (O_2899,N_49729,N_49356);
and UO_2900 (O_2900,N_49250,N_49965);
xor UO_2901 (O_2901,N_49464,N_49665);
nor UO_2902 (O_2902,N_49281,N_49546);
nor UO_2903 (O_2903,N_49175,N_49695);
xnor UO_2904 (O_2904,N_49202,N_49253);
and UO_2905 (O_2905,N_49178,N_49131);
and UO_2906 (O_2906,N_49883,N_49784);
nor UO_2907 (O_2907,N_49240,N_49293);
nor UO_2908 (O_2908,N_49830,N_49520);
or UO_2909 (O_2909,N_49887,N_49589);
xnor UO_2910 (O_2910,N_49897,N_49160);
or UO_2911 (O_2911,N_49427,N_49195);
and UO_2912 (O_2912,N_49178,N_49215);
nand UO_2913 (O_2913,N_49307,N_49984);
xnor UO_2914 (O_2914,N_49489,N_49053);
xnor UO_2915 (O_2915,N_49513,N_49115);
or UO_2916 (O_2916,N_49399,N_49573);
xor UO_2917 (O_2917,N_49365,N_49705);
and UO_2918 (O_2918,N_49088,N_49297);
nand UO_2919 (O_2919,N_49146,N_49382);
nor UO_2920 (O_2920,N_49851,N_49032);
nand UO_2921 (O_2921,N_49792,N_49282);
xnor UO_2922 (O_2922,N_49941,N_49948);
nand UO_2923 (O_2923,N_49535,N_49271);
or UO_2924 (O_2924,N_49184,N_49618);
xnor UO_2925 (O_2925,N_49887,N_49460);
or UO_2926 (O_2926,N_49878,N_49536);
nand UO_2927 (O_2927,N_49495,N_49111);
and UO_2928 (O_2928,N_49927,N_49831);
and UO_2929 (O_2929,N_49610,N_49312);
xor UO_2930 (O_2930,N_49652,N_49660);
nor UO_2931 (O_2931,N_49726,N_49297);
xor UO_2932 (O_2932,N_49808,N_49277);
xor UO_2933 (O_2933,N_49759,N_49484);
nand UO_2934 (O_2934,N_49233,N_49603);
and UO_2935 (O_2935,N_49468,N_49700);
nor UO_2936 (O_2936,N_49720,N_49571);
xor UO_2937 (O_2937,N_49339,N_49312);
or UO_2938 (O_2938,N_49560,N_49434);
xor UO_2939 (O_2939,N_49882,N_49049);
or UO_2940 (O_2940,N_49427,N_49082);
and UO_2941 (O_2941,N_49568,N_49048);
and UO_2942 (O_2942,N_49176,N_49651);
nor UO_2943 (O_2943,N_49216,N_49244);
and UO_2944 (O_2944,N_49242,N_49331);
xnor UO_2945 (O_2945,N_49516,N_49835);
or UO_2946 (O_2946,N_49799,N_49157);
nand UO_2947 (O_2947,N_49549,N_49665);
xor UO_2948 (O_2948,N_49575,N_49696);
or UO_2949 (O_2949,N_49766,N_49826);
xor UO_2950 (O_2950,N_49095,N_49486);
nor UO_2951 (O_2951,N_49455,N_49593);
nor UO_2952 (O_2952,N_49749,N_49093);
and UO_2953 (O_2953,N_49635,N_49530);
xor UO_2954 (O_2954,N_49599,N_49612);
or UO_2955 (O_2955,N_49224,N_49556);
and UO_2956 (O_2956,N_49374,N_49435);
or UO_2957 (O_2957,N_49544,N_49336);
and UO_2958 (O_2958,N_49534,N_49027);
and UO_2959 (O_2959,N_49805,N_49389);
or UO_2960 (O_2960,N_49669,N_49526);
nand UO_2961 (O_2961,N_49813,N_49225);
nand UO_2962 (O_2962,N_49969,N_49819);
nor UO_2963 (O_2963,N_49291,N_49457);
xnor UO_2964 (O_2964,N_49400,N_49734);
or UO_2965 (O_2965,N_49309,N_49622);
or UO_2966 (O_2966,N_49494,N_49905);
nand UO_2967 (O_2967,N_49792,N_49885);
xnor UO_2968 (O_2968,N_49093,N_49860);
nor UO_2969 (O_2969,N_49424,N_49815);
nand UO_2970 (O_2970,N_49991,N_49491);
nand UO_2971 (O_2971,N_49201,N_49307);
and UO_2972 (O_2972,N_49570,N_49576);
nor UO_2973 (O_2973,N_49208,N_49840);
or UO_2974 (O_2974,N_49588,N_49548);
xor UO_2975 (O_2975,N_49425,N_49621);
or UO_2976 (O_2976,N_49145,N_49848);
nor UO_2977 (O_2977,N_49935,N_49387);
xor UO_2978 (O_2978,N_49088,N_49903);
nand UO_2979 (O_2979,N_49341,N_49666);
and UO_2980 (O_2980,N_49990,N_49840);
xor UO_2981 (O_2981,N_49322,N_49477);
nor UO_2982 (O_2982,N_49478,N_49874);
and UO_2983 (O_2983,N_49905,N_49531);
and UO_2984 (O_2984,N_49688,N_49709);
nor UO_2985 (O_2985,N_49050,N_49876);
nor UO_2986 (O_2986,N_49832,N_49120);
nor UO_2987 (O_2987,N_49682,N_49316);
nor UO_2988 (O_2988,N_49625,N_49420);
and UO_2989 (O_2989,N_49641,N_49130);
xnor UO_2990 (O_2990,N_49925,N_49095);
nor UO_2991 (O_2991,N_49532,N_49910);
nand UO_2992 (O_2992,N_49019,N_49720);
xnor UO_2993 (O_2993,N_49000,N_49900);
nor UO_2994 (O_2994,N_49466,N_49307);
nor UO_2995 (O_2995,N_49082,N_49671);
or UO_2996 (O_2996,N_49642,N_49501);
or UO_2997 (O_2997,N_49251,N_49637);
or UO_2998 (O_2998,N_49727,N_49236);
and UO_2999 (O_2999,N_49496,N_49241);
nor UO_3000 (O_3000,N_49232,N_49135);
xor UO_3001 (O_3001,N_49521,N_49163);
nand UO_3002 (O_3002,N_49105,N_49996);
nand UO_3003 (O_3003,N_49766,N_49533);
nand UO_3004 (O_3004,N_49683,N_49995);
nand UO_3005 (O_3005,N_49168,N_49259);
nor UO_3006 (O_3006,N_49691,N_49616);
and UO_3007 (O_3007,N_49962,N_49327);
xor UO_3008 (O_3008,N_49414,N_49925);
nor UO_3009 (O_3009,N_49578,N_49100);
and UO_3010 (O_3010,N_49380,N_49212);
xor UO_3011 (O_3011,N_49804,N_49282);
nor UO_3012 (O_3012,N_49238,N_49761);
nor UO_3013 (O_3013,N_49165,N_49891);
nand UO_3014 (O_3014,N_49074,N_49772);
and UO_3015 (O_3015,N_49988,N_49699);
nor UO_3016 (O_3016,N_49960,N_49487);
or UO_3017 (O_3017,N_49698,N_49395);
and UO_3018 (O_3018,N_49732,N_49091);
xnor UO_3019 (O_3019,N_49509,N_49560);
or UO_3020 (O_3020,N_49390,N_49672);
nand UO_3021 (O_3021,N_49092,N_49088);
and UO_3022 (O_3022,N_49856,N_49553);
nand UO_3023 (O_3023,N_49505,N_49733);
or UO_3024 (O_3024,N_49526,N_49698);
and UO_3025 (O_3025,N_49502,N_49776);
xnor UO_3026 (O_3026,N_49846,N_49307);
nand UO_3027 (O_3027,N_49932,N_49854);
or UO_3028 (O_3028,N_49078,N_49471);
xor UO_3029 (O_3029,N_49955,N_49550);
nand UO_3030 (O_3030,N_49246,N_49702);
or UO_3031 (O_3031,N_49272,N_49952);
nand UO_3032 (O_3032,N_49985,N_49156);
nor UO_3033 (O_3033,N_49649,N_49906);
nand UO_3034 (O_3034,N_49923,N_49630);
nand UO_3035 (O_3035,N_49475,N_49908);
and UO_3036 (O_3036,N_49723,N_49459);
xor UO_3037 (O_3037,N_49750,N_49682);
nor UO_3038 (O_3038,N_49289,N_49177);
nor UO_3039 (O_3039,N_49200,N_49515);
nand UO_3040 (O_3040,N_49540,N_49309);
xor UO_3041 (O_3041,N_49457,N_49606);
nand UO_3042 (O_3042,N_49272,N_49482);
xnor UO_3043 (O_3043,N_49489,N_49313);
nor UO_3044 (O_3044,N_49336,N_49950);
or UO_3045 (O_3045,N_49329,N_49236);
nand UO_3046 (O_3046,N_49651,N_49554);
nand UO_3047 (O_3047,N_49913,N_49706);
nor UO_3048 (O_3048,N_49842,N_49930);
or UO_3049 (O_3049,N_49226,N_49695);
and UO_3050 (O_3050,N_49730,N_49156);
or UO_3051 (O_3051,N_49157,N_49469);
or UO_3052 (O_3052,N_49472,N_49953);
xor UO_3053 (O_3053,N_49375,N_49983);
nor UO_3054 (O_3054,N_49759,N_49963);
nand UO_3055 (O_3055,N_49395,N_49745);
nor UO_3056 (O_3056,N_49821,N_49985);
or UO_3057 (O_3057,N_49110,N_49172);
nand UO_3058 (O_3058,N_49585,N_49773);
and UO_3059 (O_3059,N_49541,N_49699);
or UO_3060 (O_3060,N_49124,N_49053);
and UO_3061 (O_3061,N_49827,N_49807);
nor UO_3062 (O_3062,N_49381,N_49918);
or UO_3063 (O_3063,N_49312,N_49014);
nor UO_3064 (O_3064,N_49626,N_49587);
xor UO_3065 (O_3065,N_49013,N_49576);
nor UO_3066 (O_3066,N_49695,N_49078);
nor UO_3067 (O_3067,N_49172,N_49159);
nor UO_3068 (O_3068,N_49402,N_49399);
xor UO_3069 (O_3069,N_49179,N_49685);
and UO_3070 (O_3070,N_49044,N_49735);
nor UO_3071 (O_3071,N_49426,N_49423);
nand UO_3072 (O_3072,N_49454,N_49641);
nand UO_3073 (O_3073,N_49585,N_49059);
and UO_3074 (O_3074,N_49984,N_49723);
or UO_3075 (O_3075,N_49545,N_49562);
nor UO_3076 (O_3076,N_49700,N_49546);
and UO_3077 (O_3077,N_49214,N_49278);
nand UO_3078 (O_3078,N_49843,N_49899);
or UO_3079 (O_3079,N_49419,N_49674);
xor UO_3080 (O_3080,N_49708,N_49018);
and UO_3081 (O_3081,N_49887,N_49851);
or UO_3082 (O_3082,N_49344,N_49072);
nand UO_3083 (O_3083,N_49047,N_49610);
xnor UO_3084 (O_3084,N_49919,N_49733);
nor UO_3085 (O_3085,N_49319,N_49921);
nor UO_3086 (O_3086,N_49306,N_49481);
xnor UO_3087 (O_3087,N_49772,N_49051);
xor UO_3088 (O_3088,N_49214,N_49592);
nand UO_3089 (O_3089,N_49876,N_49945);
nor UO_3090 (O_3090,N_49504,N_49687);
xor UO_3091 (O_3091,N_49074,N_49479);
and UO_3092 (O_3092,N_49559,N_49016);
nor UO_3093 (O_3093,N_49565,N_49100);
xor UO_3094 (O_3094,N_49244,N_49159);
or UO_3095 (O_3095,N_49159,N_49491);
xor UO_3096 (O_3096,N_49637,N_49222);
nor UO_3097 (O_3097,N_49125,N_49963);
or UO_3098 (O_3098,N_49212,N_49298);
nor UO_3099 (O_3099,N_49203,N_49228);
nand UO_3100 (O_3100,N_49961,N_49423);
nand UO_3101 (O_3101,N_49878,N_49244);
xor UO_3102 (O_3102,N_49720,N_49159);
and UO_3103 (O_3103,N_49246,N_49034);
nand UO_3104 (O_3104,N_49571,N_49247);
or UO_3105 (O_3105,N_49890,N_49176);
nand UO_3106 (O_3106,N_49877,N_49204);
or UO_3107 (O_3107,N_49879,N_49006);
and UO_3108 (O_3108,N_49011,N_49351);
nor UO_3109 (O_3109,N_49768,N_49206);
nand UO_3110 (O_3110,N_49553,N_49018);
xnor UO_3111 (O_3111,N_49130,N_49037);
or UO_3112 (O_3112,N_49600,N_49835);
and UO_3113 (O_3113,N_49712,N_49684);
nor UO_3114 (O_3114,N_49379,N_49870);
nor UO_3115 (O_3115,N_49869,N_49943);
or UO_3116 (O_3116,N_49683,N_49651);
and UO_3117 (O_3117,N_49830,N_49537);
nor UO_3118 (O_3118,N_49819,N_49030);
xor UO_3119 (O_3119,N_49011,N_49991);
and UO_3120 (O_3120,N_49333,N_49749);
nor UO_3121 (O_3121,N_49274,N_49801);
and UO_3122 (O_3122,N_49531,N_49463);
and UO_3123 (O_3123,N_49904,N_49683);
xnor UO_3124 (O_3124,N_49733,N_49391);
and UO_3125 (O_3125,N_49963,N_49229);
nand UO_3126 (O_3126,N_49414,N_49988);
and UO_3127 (O_3127,N_49378,N_49592);
and UO_3128 (O_3128,N_49404,N_49047);
or UO_3129 (O_3129,N_49494,N_49620);
or UO_3130 (O_3130,N_49366,N_49890);
nor UO_3131 (O_3131,N_49638,N_49452);
nand UO_3132 (O_3132,N_49181,N_49286);
nor UO_3133 (O_3133,N_49167,N_49815);
nor UO_3134 (O_3134,N_49420,N_49320);
xnor UO_3135 (O_3135,N_49178,N_49833);
nor UO_3136 (O_3136,N_49640,N_49070);
or UO_3137 (O_3137,N_49236,N_49180);
and UO_3138 (O_3138,N_49946,N_49441);
and UO_3139 (O_3139,N_49490,N_49072);
nor UO_3140 (O_3140,N_49079,N_49237);
or UO_3141 (O_3141,N_49748,N_49783);
and UO_3142 (O_3142,N_49660,N_49666);
nor UO_3143 (O_3143,N_49115,N_49070);
nand UO_3144 (O_3144,N_49305,N_49310);
nor UO_3145 (O_3145,N_49450,N_49774);
nor UO_3146 (O_3146,N_49392,N_49695);
and UO_3147 (O_3147,N_49235,N_49921);
and UO_3148 (O_3148,N_49990,N_49024);
xnor UO_3149 (O_3149,N_49414,N_49834);
or UO_3150 (O_3150,N_49177,N_49285);
and UO_3151 (O_3151,N_49976,N_49772);
xnor UO_3152 (O_3152,N_49942,N_49752);
or UO_3153 (O_3153,N_49430,N_49818);
nand UO_3154 (O_3154,N_49882,N_49944);
and UO_3155 (O_3155,N_49578,N_49748);
and UO_3156 (O_3156,N_49875,N_49928);
or UO_3157 (O_3157,N_49898,N_49382);
or UO_3158 (O_3158,N_49761,N_49378);
or UO_3159 (O_3159,N_49980,N_49877);
nor UO_3160 (O_3160,N_49127,N_49682);
nor UO_3161 (O_3161,N_49160,N_49791);
xor UO_3162 (O_3162,N_49370,N_49461);
xor UO_3163 (O_3163,N_49197,N_49821);
and UO_3164 (O_3164,N_49988,N_49079);
xor UO_3165 (O_3165,N_49855,N_49269);
nand UO_3166 (O_3166,N_49903,N_49584);
nand UO_3167 (O_3167,N_49105,N_49730);
xnor UO_3168 (O_3168,N_49003,N_49542);
and UO_3169 (O_3169,N_49338,N_49685);
nand UO_3170 (O_3170,N_49530,N_49624);
and UO_3171 (O_3171,N_49569,N_49517);
and UO_3172 (O_3172,N_49847,N_49555);
nor UO_3173 (O_3173,N_49507,N_49717);
xnor UO_3174 (O_3174,N_49711,N_49279);
and UO_3175 (O_3175,N_49444,N_49134);
and UO_3176 (O_3176,N_49452,N_49727);
nor UO_3177 (O_3177,N_49991,N_49817);
xor UO_3178 (O_3178,N_49560,N_49723);
nand UO_3179 (O_3179,N_49016,N_49219);
nor UO_3180 (O_3180,N_49292,N_49461);
xnor UO_3181 (O_3181,N_49272,N_49881);
xnor UO_3182 (O_3182,N_49818,N_49442);
nor UO_3183 (O_3183,N_49437,N_49268);
and UO_3184 (O_3184,N_49675,N_49189);
nor UO_3185 (O_3185,N_49208,N_49770);
and UO_3186 (O_3186,N_49137,N_49234);
or UO_3187 (O_3187,N_49870,N_49954);
xnor UO_3188 (O_3188,N_49645,N_49920);
or UO_3189 (O_3189,N_49903,N_49253);
nor UO_3190 (O_3190,N_49700,N_49350);
nor UO_3191 (O_3191,N_49636,N_49513);
nand UO_3192 (O_3192,N_49336,N_49486);
nand UO_3193 (O_3193,N_49503,N_49007);
or UO_3194 (O_3194,N_49740,N_49396);
nand UO_3195 (O_3195,N_49218,N_49791);
nor UO_3196 (O_3196,N_49062,N_49708);
nor UO_3197 (O_3197,N_49040,N_49468);
and UO_3198 (O_3198,N_49064,N_49288);
and UO_3199 (O_3199,N_49274,N_49348);
xor UO_3200 (O_3200,N_49836,N_49666);
and UO_3201 (O_3201,N_49277,N_49909);
xor UO_3202 (O_3202,N_49710,N_49303);
or UO_3203 (O_3203,N_49500,N_49122);
or UO_3204 (O_3204,N_49707,N_49842);
xor UO_3205 (O_3205,N_49841,N_49431);
xor UO_3206 (O_3206,N_49232,N_49381);
and UO_3207 (O_3207,N_49743,N_49671);
or UO_3208 (O_3208,N_49932,N_49173);
and UO_3209 (O_3209,N_49446,N_49822);
nor UO_3210 (O_3210,N_49013,N_49475);
or UO_3211 (O_3211,N_49336,N_49986);
and UO_3212 (O_3212,N_49717,N_49040);
xor UO_3213 (O_3213,N_49569,N_49604);
or UO_3214 (O_3214,N_49064,N_49436);
nand UO_3215 (O_3215,N_49653,N_49862);
nor UO_3216 (O_3216,N_49510,N_49753);
and UO_3217 (O_3217,N_49590,N_49696);
or UO_3218 (O_3218,N_49880,N_49292);
xnor UO_3219 (O_3219,N_49923,N_49486);
and UO_3220 (O_3220,N_49212,N_49233);
and UO_3221 (O_3221,N_49491,N_49692);
xnor UO_3222 (O_3222,N_49849,N_49929);
xor UO_3223 (O_3223,N_49300,N_49602);
nand UO_3224 (O_3224,N_49173,N_49319);
nor UO_3225 (O_3225,N_49834,N_49887);
nor UO_3226 (O_3226,N_49202,N_49674);
nand UO_3227 (O_3227,N_49104,N_49373);
or UO_3228 (O_3228,N_49706,N_49069);
nand UO_3229 (O_3229,N_49668,N_49777);
and UO_3230 (O_3230,N_49751,N_49319);
xor UO_3231 (O_3231,N_49153,N_49715);
nand UO_3232 (O_3232,N_49468,N_49097);
and UO_3233 (O_3233,N_49726,N_49428);
and UO_3234 (O_3234,N_49336,N_49907);
nor UO_3235 (O_3235,N_49871,N_49221);
or UO_3236 (O_3236,N_49686,N_49642);
and UO_3237 (O_3237,N_49971,N_49136);
and UO_3238 (O_3238,N_49338,N_49319);
nand UO_3239 (O_3239,N_49423,N_49767);
nor UO_3240 (O_3240,N_49335,N_49794);
nor UO_3241 (O_3241,N_49181,N_49098);
and UO_3242 (O_3242,N_49170,N_49919);
and UO_3243 (O_3243,N_49507,N_49073);
xor UO_3244 (O_3244,N_49714,N_49774);
and UO_3245 (O_3245,N_49749,N_49009);
nor UO_3246 (O_3246,N_49325,N_49652);
nor UO_3247 (O_3247,N_49872,N_49306);
nand UO_3248 (O_3248,N_49807,N_49248);
nor UO_3249 (O_3249,N_49096,N_49312);
nand UO_3250 (O_3250,N_49971,N_49960);
nor UO_3251 (O_3251,N_49462,N_49776);
nand UO_3252 (O_3252,N_49518,N_49816);
and UO_3253 (O_3253,N_49564,N_49718);
and UO_3254 (O_3254,N_49073,N_49586);
xnor UO_3255 (O_3255,N_49613,N_49009);
nor UO_3256 (O_3256,N_49140,N_49851);
and UO_3257 (O_3257,N_49187,N_49716);
xor UO_3258 (O_3258,N_49878,N_49956);
or UO_3259 (O_3259,N_49774,N_49885);
xnor UO_3260 (O_3260,N_49088,N_49212);
nand UO_3261 (O_3261,N_49230,N_49103);
and UO_3262 (O_3262,N_49423,N_49219);
and UO_3263 (O_3263,N_49098,N_49752);
or UO_3264 (O_3264,N_49344,N_49448);
xor UO_3265 (O_3265,N_49400,N_49294);
nand UO_3266 (O_3266,N_49469,N_49006);
nand UO_3267 (O_3267,N_49759,N_49691);
nor UO_3268 (O_3268,N_49455,N_49120);
and UO_3269 (O_3269,N_49435,N_49665);
nor UO_3270 (O_3270,N_49928,N_49779);
nand UO_3271 (O_3271,N_49444,N_49951);
nand UO_3272 (O_3272,N_49490,N_49706);
xnor UO_3273 (O_3273,N_49568,N_49810);
or UO_3274 (O_3274,N_49540,N_49484);
xor UO_3275 (O_3275,N_49964,N_49556);
xnor UO_3276 (O_3276,N_49379,N_49619);
and UO_3277 (O_3277,N_49525,N_49397);
nor UO_3278 (O_3278,N_49435,N_49327);
xnor UO_3279 (O_3279,N_49161,N_49936);
or UO_3280 (O_3280,N_49792,N_49442);
or UO_3281 (O_3281,N_49771,N_49477);
xnor UO_3282 (O_3282,N_49144,N_49113);
and UO_3283 (O_3283,N_49308,N_49026);
or UO_3284 (O_3284,N_49855,N_49279);
or UO_3285 (O_3285,N_49473,N_49340);
nor UO_3286 (O_3286,N_49630,N_49032);
nor UO_3287 (O_3287,N_49900,N_49356);
and UO_3288 (O_3288,N_49127,N_49876);
xor UO_3289 (O_3289,N_49806,N_49656);
nor UO_3290 (O_3290,N_49562,N_49507);
xnor UO_3291 (O_3291,N_49123,N_49198);
xor UO_3292 (O_3292,N_49293,N_49066);
or UO_3293 (O_3293,N_49029,N_49846);
nand UO_3294 (O_3294,N_49948,N_49602);
or UO_3295 (O_3295,N_49217,N_49631);
nand UO_3296 (O_3296,N_49451,N_49757);
and UO_3297 (O_3297,N_49590,N_49671);
xnor UO_3298 (O_3298,N_49308,N_49430);
or UO_3299 (O_3299,N_49060,N_49048);
or UO_3300 (O_3300,N_49924,N_49952);
or UO_3301 (O_3301,N_49958,N_49414);
xnor UO_3302 (O_3302,N_49787,N_49841);
or UO_3303 (O_3303,N_49918,N_49437);
nor UO_3304 (O_3304,N_49762,N_49213);
and UO_3305 (O_3305,N_49218,N_49167);
nor UO_3306 (O_3306,N_49870,N_49334);
xor UO_3307 (O_3307,N_49619,N_49570);
xor UO_3308 (O_3308,N_49262,N_49900);
nor UO_3309 (O_3309,N_49893,N_49478);
or UO_3310 (O_3310,N_49830,N_49389);
nor UO_3311 (O_3311,N_49115,N_49619);
nor UO_3312 (O_3312,N_49984,N_49168);
and UO_3313 (O_3313,N_49636,N_49723);
or UO_3314 (O_3314,N_49176,N_49737);
or UO_3315 (O_3315,N_49510,N_49923);
or UO_3316 (O_3316,N_49551,N_49288);
xnor UO_3317 (O_3317,N_49944,N_49175);
and UO_3318 (O_3318,N_49361,N_49954);
and UO_3319 (O_3319,N_49296,N_49634);
nand UO_3320 (O_3320,N_49034,N_49020);
nor UO_3321 (O_3321,N_49882,N_49002);
and UO_3322 (O_3322,N_49966,N_49405);
nand UO_3323 (O_3323,N_49688,N_49176);
or UO_3324 (O_3324,N_49414,N_49893);
or UO_3325 (O_3325,N_49338,N_49909);
nand UO_3326 (O_3326,N_49502,N_49743);
xnor UO_3327 (O_3327,N_49402,N_49686);
xnor UO_3328 (O_3328,N_49213,N_49156);
or UO_3329 (O_3329,N_49377,N_49380);
nor UO_3330 (O_3330,N_49968,N_49356);
or UO_3331 (O_3331,N_49959,N_49095);
nand UO_3332 (O_3332,N_49819,N_49319);
xnor UO_3333 (O_3333,N_49415,N_49841);
xnor UO_3334 (O_3334,N_49038,N_49348);
or UO_3335 (O_3335,N_49054,N_49874);
nor UO_3336 (O_3336,N_49729,N_49766);
and UO_3337 (O_3337,N_49903,N_49783);
or UO_3338 (O_3338,N_49408,N_49297);
and UO_3339 (O_3339,N_49297,N_49355);
and UO_3340 (O_3340,N_49535,N_49790);
or UO_3341 (O_3341,N_49006,N_49308);
or UO_3342 (O_3342,N_49261,N_49199);
nor UO_3343 (O_3343,N_49957,N_49133);
nor UO_3344 (O_3344,N_49488,N_49105);
and UO_3345 (O_3345,N_49598,N_49612);
or UO_3346 (O_3346,N_49016,N_49213);
nand UO_3347 (O_3347,N_49790,N_49217);
xnor UO_3348 (O_3348,N_49176,N_49980);
and UO_3349 (O_3349,N_49744,N_49891);
and UO_3350 (O_3350,N_49481,N_49441);
nor UO_3351 (O_3351,N_49435,N_49434);
or UO_3352 (O_3352,N_49793,N_49215);
nor UO_3353 (O_3353,N_49548,N_49651);
or UO_3354 (O_3354,N_49562,N_49759);
and UO_3355 (O_3355,N_49114,N_49364);
nand UO_3356 (O_3356,N_49440,N_49911);
or UO_3357 (O_3357,N_49707,N_49060);
nand UO_3358 (O_3358,N_49279,N_49439);
nand UO_3359 (O_3359,N_49849,N_49453);
nand UO_3360 (O_3360,N_49619,N_49816);
or UO_3361 (O_3361,N_49967,N_49961);
and UO_3362 (O_3362,N_49586,N_49298);
nor UO_3363 (O_3363,N_49522,N_49085);
nand UO_3364 (O_3364,N_49252,N_49773);
nand UO_3365 (O_3365,N_49474,N_49661);
nor UO_3366 (O_3366,N_49906,N_49786);
or UO_3367 (O_3367,N_49281,N_49415);
nor UO_3368 (O_3368,N_49955,N_49174);
nor UO_3369 (O_3369,N_49500,N_49072);
and UO_3370 (O_3370,N_49291,N_49376);
nand UO_3371 (O_3371,N_49836,N_49036);
nor UO_3372 (O_3372,N_49102,N_49556);
and UO_3373 (O_3373,N_49251,N_49149);
nor UO_3374 (O_3374,N_49510,N_49422);
xor UO_3375 (O_3375,N_49035,N_49206);
or UO_3376 (O_3376,N_49117,N_49826);
and UO_3377 (O_3377,N_49730,N_49418);
and UO_3378 (O_3378,N_49033,N_49861);
or UO_3379 (O_3379,N_49219,N_49920);
or UO_3380 (O_3380,N_49764,N_49561);
xor UO_3381 (O_3381,N_49703,N_49316);
xor UO_3382 (O_3382,N_49295,N_49276);
and UO_3383 (O_3383,N_49413,N_49671);
nand UO_3384 (O_3384,N_49583,N_49003);
xor UO_3385 (O_3385,N_49868,N_49612);
xnor UO_3386 (O_3386,N_49498,N_49405);
xnor UO_3387 (O_3387,N_49338,N_49479);
and UO_3388 (O_3388,N_49667,N_49890);
and UO_3389 (O_3389,N_49482,N_49562);
xnor UO_3390 (O_3390,N_49609,N_49500);
nand UO_3391 (O_3391,N_49341,N_49004);
nor UO_3392 (O_3392,N_49161,N_49201);
or UO_3393 (O_3393,N_49864,N_49953);
nor UO_3394 (O_3394,N_49170,N_49970);
nand UO_3395 (O_3395,N_49903,N_49844);
xor UO_3396 (O_3396,N_49213,N_49337);
xnor UO_3397 (O_3397,N_49756,N_49537);
and UO_3398 (O_3398,N_49512,N_49730);
nand UO_3399 (O_3399,N_49530,N_49037);
nor UO_3400 (O_3400,N_49431,N_49995);
nand UO_3401 (O_3401,N_49744,N_49342);
nand UO_3402 (O_3402,N_49673,N_49917);
or UO_3403 (O_3403,N_49636,N_49870);
and UO_3404 (O_3404,N_49567,N_49271);
nor UO_3405 (O_3405,N_49359,N_49602);
or UO_3406 (O_3406,N_49730,N_49978);
nand UO_3407 (O_3407,N_49775,N_49686);
or UO_3408 (O_3408,N_49622,N_49421);
nor UO_3409 (O_3409,N_49948,N_49518);
nand UO_3410 (O_3410,N_49187,N_49890);
nor UO_3411 (O_3411,N_49967,N_49726);
and UO_3412 (O_3412,N_49194,N_49952);
nand UO_3413 (O_3413,N_49300,N_49945);
and UO_3414 (O_3414,N_49858,N_49626);
or UO_3415 (O_3415,N_49882,N_49964);
nor UO_3416 (O_3416,N_49118,N_49885);
nor UO_3417 (O_3417,N_49739,N_49980);
or UO_3418 (O_3418,N_49459,N_49250);
xor UO_3419 (O_3419,N_49326,N_49148);
or UO_3420 (O_3420,N_49713,N_49081);
or UO_3421 (O_3421,N_49346,N_49196);
xor UO_3422 (O_3422,N_49662,N_49609);
nor UO_3423 (O_3423,N_49505,N_49536);
xnor UO_3424 (O_3424,N_49060,N_49813);
nor UO_3425 (O_3425,N_49339,N_49872);
and UO_3426 (O_3426,N_49629,N_49706);
or UO_3427 (O_3427,N_49989,N_49383);
or UO_3428 (O_3428,N_49711,N_49843);
and UO_3429 (O_3429,N_49532,N_49591);
and UO_3430 (O_3430,N_49963,N_49475);
or UO_3431 (O_3431,N_49235,N_49890);
or UO_3432 (O_3432,N_49241,N_49044);
nor UO_3433 (O_3433,N_49765,N_49304);
nor UO_3434 (O_3434,N_49041,N_49997);
or UO_3435 (O_3435,N_49389,N_49542);
nor UO_3436 (O_3436,N_49908,N_49379);
nor UO_3437 (O_3437,N_49371,N_49835);
or UO_3438 (O_3438,N_49075,N_49301);
and UO_3439 (O_3439,N_49652,N_49010);
xnor UO_3440 (O_3440,N_49615,N_49884);
xor UO_3441 (O_3441,N_49694,N_49124);
or UO_3442 (O_3442,N_49126,N_49636);
nor UO_3443 (O_3443,N_49969,N_49553);
or UO_3444 (O_3444,N_49480,N_49043);
or UO_3445 (O_3445,N_49064,N_49266);
and UO_3446 (O_3446,N_49063,N_49974);
xor UO_3447 (O_3447,N_49820,N_49047);
or UO_3448 (O_3448,N_49845,N_49692);
xor UO_3449 (O_3449,N_49312,N_49408);
xnor UO_3450 (O_3450,N_49893,N_49790);
and UO_3451 (O_3451,N_49456,N_49465);
nor UO_3452 (O_3452,N_49974,N_49491);
nand UO_3453 (O_3453,N_49168,N_49543);
or UO_3454 (O_3454,N_49250,N_49517);
and UO_3455 (O_3455,N_49218,N_49379);
nand UO_3456 (O_3456,N_49538,N_49915);
or UO_3457 (O_3457,N_49279,N_49908);
nor UO_3458 (O_3458,N_49387,N_49216);
nor UO_3459 (O_3459,N_49576,N_49707);
xnor UO_3460 (O_3460,N_49859,N_49719);
xnor UO_3461 (O_3461,N_49208,N_49234);
nand UO_3462 (O_3462,N_49665,N_49200);
xnor UO_3463 (O_3463,N_49063,N_49465);
xor UO_3464 (O_3464,N_49242,N_49892);
nand UO_3465 (O_3465,N_49350,N_49957);
nor UO_3466 (O_3466,N_49507,N_49854);
xor UO_3467 (O_3467,N_49025,N_49514);
nor UO_3468 (O_3468,N_49051,N_49104);
nor UO_3469 (O_3469,N_49385,N_49730);
xnor UO_3470 (O_3470,N_49009,N_49311);
and UO_3471 (O_3471,N_49933,N_49597);
or UO_3472 (O_3472,N_49167,N_49691);
or UO_3473 (O_3473,N_49948,N_49828);
and UO_3474 (O_3474,N_49175,N_49208);
nand UO_3475 (O_3475,N_49507,N_49023);
or UO_3476 (O_3476,N_49680,N_49199);
nand UO_3477 (O_3477,N_49899,N_49052);
nand UO_3478 (O_3478,N_49219,N_49217);
and UO_3479 (O_3479,N_49425,N_49847);
or UO_3480 (O_3480,N_49130,N_49285);
xnor UO_3481 (O_3481,N_49426,N_49492);
nand UO_3482 (O_3482,N_49673,N_49128);
or UO_3483 (O_3483,N_49492,N_49826);
nand UO_3484 (O_3484,N_49779,N_49418);
xnor UO_3485 (O_3485,N_49455,N_49825);
nor UO_3486 (O_3486,N_49421,N_49508);
or UO_3487 (O_3487,N_49406,N_49714);
nand UO_3488 (O_3488,N_49174,N_49641);
and UO_3489 (O_3489,N_49418,N_49825);
nor UO_3490 (O_3490,N_49868,N_49498);
nor UO_3491 (O_3491,N_49011,N_49318);
and UO_3492 (O_3492,N_49340,N_49639);
xnor UO_3493 (O_3493,N_49898,N_49652);
and UO_3494 (O_3494,N_49061,N_49288);
and UO_3495 (O_3495,N_49160,N_49411);
nand UO_3496 (O_3496,N_49149,N_49842);
or UO_3497 (O_3497,N_49319,N_49606);
and UO_3498 (O_3498,N_49202,N_49270);
nor UO_3499 (O_3499,N_49682,N_49564);
nand UO_3500 (O_3500,N_49737,N_49412);
or UO_3501 (O_3501,N_49301,N_49397);
or UO_3502 (O_3502,N_49540,N_49949);
nand UO_3503 (O_3503,N_49974,N_49954);
xor UO_3504 (O_3504,N_49532,N_49168);
nor UO_3505 (O_3505,N_49160,N_49660);
or UO_3506 (O_3506,N_49748,N_49665);
nand UO_3507 (O_3507,N_49903,N_49878);
nand UO_3508 (O_3508,N_49835,N_49756);
xor UO_3509 (O_3509,N_49784,N_49093);
nand UO_3510 (O_3510,N_49854,N_49310);
nor UO_3511 (O_3511,N_49469,N_49375);
or UO_3512 (O_3512,N_49021,N_49585);
or UO_3513 (O_3513,N_49313,N_49282);
nor UO_3514 (O_3514,N_49048,N_49808);
nand UO_3515 (O_3515,N_49692,N_49395);
xnor UO_3516 (O_3516,N_49345,N_49967);
or UO_3517 (O_3517,N_49562,N_49409);
or UO_3518 (O_3518,N_49062,N_49724);
xor UO_3519 (O_3519,N_49899,N_49211);
xor UO_3520 (O_3520,N_49647,N_49887);
and UO_3521 (O_3521,N_49078,N_49140);
nor UO_3522 (O_3522,N_49716,N_49632);
nor UO_3523 (O_3523,N_49449,N_49814);
or UO_3524 (O_3524,N_49421,N_49592);
xnor UO_3525 (O_3525,N_49026,N_49318);
xnor UO_3526 (O_3526,N_49874,N_49407);
xor UO_3527 (O_3527,N_49589,N_49509);
nor UO_3528 (O_3528,N_49462,N_49452);
nand UO_3529 (O_3529,N_49785,N_49165);
xor UO_3530 (O_3530,N_49321,N_49916);
or UO_3531 (O_3531,N_49368,N_49656);
and UO_3532 (O_3532,N_49218,N_49404);
xor UO_3533 (O_3533,N_49520,N_49674);
xnor UO_3534 (O_3534,N_49215,N_49396);
nor UO_3535 (O_3535,N_49436,N_49889);
nor UO_3536 (O_3536,N_49592,N_49508);
and UO_3537 (O_3537,N_49271,N_49241);
nor UO_3538 (O_3538,N_49157,N_49354);
xor UO_3539 (O_3539,N_49167,N_49964);
nand UO_3540 (O_3540,N_49332,N_49242);
and UO_3541 (O_3541,N_49431,N_49557);
or UO_3542 (O_3542,N_49113,N_49015);
and UO_3543 (O_3543,N_49991,N_49007);
xor UO_3544 (O_3544,N_49034,N_49116);
nor UO_3545 (O_3545,N_49921,N_49582);
or UO_3546 (O_3546,N_49626,N_49935);
nor UO_3547 (O_3547,N_49520,N_49880);
xor UO_3548 (O_3548,N_49603,N_49438);
nor UO_3549 (O_3549,N_49723,N_49061);
or UO_3550 (O_3550,N_49421,N_49209);
nand UO_3551 (O_3551,N_49981,N_49528);
and UO_3552 (O_3552,N_49490,N_49231);
and UO_3553 (O_3553,N_49030,N_49884);
nand UO_3554 (O_3554,N_49564,N_49284);
or UO_3555 (O_3555,N_49010,N_49226);
nand UO_3556 (O_3556,N_49585,N_49729);
xnor UO_3557 (O_3557,N_49538,N_49304);
nor UO_3558 (O_3558,N_49789,N_49440);
xor UO_3559 (O_3559,N_49616,N_49537);
and UO_3560 (O_3560,N_49411,N_49507);
nor UO_3561 (O_3561,N_49854,N_49139);
or UO_3562 (O_3562,N_49212,N_49338);
or UO_3563 (O_3563,N_49572,N_49220);
nand UO_3564 (O_3564,N_49376,N_49827);
xnor UO_3565 (O_3565,N_49979,N_49853);
and UO_3566 (O_3566,N_49947,N_49704);
nor UO_3567 (O_3567,N_49527,N_49206);
xnor UO_3568 (O_3568,N_49870,N_49942);
or UO_3569 (O_3569,N_49965,N_49993);
xor UO_3570 (O_3570,N_49404,N_49574);
nand UO_3571 (O_3571,N_49599,N_49774);
xor UO_3572 (O_3572,N_49664,N_49046);
nand UO_3573 (O_3573,N_49221,N_49952);
xor UO_3574 (O_3574,N_49124,N_49010);
xor UO_3575 (O_3575,N_49831,N_49562);
and UO_3576 (O_3576,N_49111,N_49815);
xnor UO_3577 (O_3577,N_49653,N_49169);
nand UO_3578 (O_3578,N_49859,N_49706);
and UO_3579 (O_3579,N_49339,N_49944);
or UO_3580 (O_3580,N_49654,N_49176);
nand UO_3581 (O_3581,N_49853,N_49544);
xnor UO_3582 (O_3582,N_49997,N_49071);
or UO_3583 (O_3583,N_49897,N_49748);
or UO_3584 (O_3584,N_49191,N_49201);
or UO_3585 (O_3585,N_49494,N_49593);
nor UO_3586 (O_3586,N_49200,N_49000);
nand UO_3587 (O_3587,N_49920,N_49483);
or UO_3588 (O_3588,N_49407,N_49513);
nand UO_3589 (O_3589,N_49412,N_49036);
and UO_3590 (O_3590,N_49497,N_49103);
and UO_3591 (O_3591,N_49625,N_49478);
xnor UO_3592 (O_3592,N_49236,N_49523);
xor UO_3593 (O_3593,N_49860,N_49551);
nand UO_3594 (O_3594,N_49395,N_49511);
nor UO_3595 (O_3595,N_49032,N_49561);
nor UO_3596 (O_3596,N_49542,N_49999);
or UO_3597 (O_3597,N_49603,N_49389);
nor UO_3598 (O_3598,N_49148,N_49032);
xor UO_3599 (O_3599,N_49785,N_49741);
and UO_3600 (O_3600,N_49945,N_49598);
xor UO_3601 (O_3601,N_49122,N_49261);
nand UO_3602 (O_3602,N_49889,N_49447);
xor UO_3603 (O_3603,N_49479,N_49550);
and UO_3604 (O_3604,N_49107,N_49922);
and UO_3605 (O_3605,N_49539,N_49331);
or UO_3606 (O_3606,N_49386,N_49061);
xor UO_3607 (O_3607,N_49443,N_49969);
xor UO_3608 (O_3608,N_49213,N_49202);
nand UO_3609 (O_3609,N_49605,N_49866);
xnor UO_3610 (O_3610,N_49171,N_49888);
or UO_3611 (O_3611,N_49938,N_49964);
xor UO_3612 (O_3612,N_49496,N_49523);
xnor UO_3613 (O_3613,N_49546,N_49508);
or UO_3614 (O_3614,N_49816,N_49311);
xor UO_3615 (O_3615,N_49460,N_49985);
xnor UO_3616 (O_3616,N_49702,N_49896);
or UO_3617 (O_3617,N_49967,N_49114);
nand UO_3618 (O_3618,N_49896,N_49824);
xnor UO_3619 (O_3619,N_49141,N_49189);
and UO_3620 (O_3620,N_49116,N_49700);
nor UO_3621 (O_3621,N_49580,N_49232);
nand UO_3622 (O_3622,N_49118,N_49942);
or UO_3623 (O_3623,N_49608,N_49758);
nor UO_3624 (O_3624,N_49463,N_49340);
or UO_3625 (O_3625,N_49056,N_49101);
xor UO_3626 (O_3626,N_49017,N_49580);
nor UO_3627 (O_3627,N_49580,N_49120);
xnor UO_3628 (O_3628,N_49656,N_49548);
nand UO_3629 (O_3629,N_49444,N_49424);
and UO_3630 (O_3630,N_49402,N_49595);
nand UO_3631 (O_3631,N_49139,N_49460);
and UO_3632 (O_3632,N_49088,N_49983);
and UO_3633 (O_3633,N_49093,N_49130);
nor UO_3634 (O_3634,N_49028,N_49519);
xnor UO_3635 (O_3635,N_49967,N_49377);
or UO_3636 (O_3636,N_49746,N_49913);
and UO_3637 (O_3637,N_49341,N_49675);
xor UO_3638 (O_3638,N_49433,N_49556);
nand UO_3639 (O_3639,N_49999,N_49170);
nand UO_3640 (O_3640,N_49512,N_49857);
nand UO_3641 (O_3641,N_49175,N_49615);
and UO_3642 (O_3642,N_49196,N_49940);
xnor UO_3643 (O_3643,N_49432,N_49986);
xnor UO_3644 (O_3644,N_49469,N_49763);
nand UO_3645 (O_3645,N_49106,N_49494);
and UO_3646 (O_3646,N_49274,N_49718);
nand UO_3647 (O_3647,N_49226,N_49173);
and UO_3648 (O_3648,N_49512,N_49345);
nand UO_3649 (O_3649,N_49352,N_49585);
nand UO_3650 (O_3650,N_49471,N_49225);
or UO_3651 (O_3651,N_49463,N_49163);
and UO_3652 (O_3652,N_49058,N_49417);
nor UO_3653 (O_3653,N_49724,N_49120);
nand UO_3654 (O_3654,N_49339,N_49682);
and UO_3655 (O_3655,N_49152,N_49073);
nand UO_3656 (O_3656,N_49779,N_49457);
nor UO_3657 (O_3657,N_49892,N_49714);
and UO_3658 (O_3658,N_49807,N_49474);
nor UO_3659 (O_3659,N_49089,N_49357);
or UO_3660 (O_3660,N_49090,N_49458);
xor UO_3661 (O_3661,N_49492,N_49312);
or UO_3662 (O_3662,N_49355,N_49928);
nor UO_3663 (O_3663,N_49774,N_49017);
and UO_3664 (O_3664,N_49980,N_49388);
and UO_3665 (O_3665,N_49192,N_49209);
nand UO_3666 (O_3666,N_49808,N_49846);
and UO_3667 (O_3667,N_49612,N_49936);
nor UO_3668 (O_3668,N_49195,N_49173);
nand UO_3669 (O_3669,N_49018,N_49647);
nand UO_3670 (O_3670,N_49650,N_49160);
or UO_3671 (O_3671,N_49060,N_49854);
nor UO_3672 (O_3672,N_49443,N_49739);
nand UO_3673 (O_3673,N_49936,N_49900);
and UO_3674 (O_3674,N_49121,N_49226);
nand UO_3675 (O_3675,N_49983,N_49131);
and UO_3676 (O_3676,N_49090,N_49691);
or UO_3677 (O_3677,N_49842,N_49748);
and UO_3678 (O_3678,N_49800,N_49841);
nand UO_3679 (O_3679,N_49756,N_49216);
xor UO_3680 (O_3680,N_49600,N_49330);
xnor UO_3681 (O_3681,N_49261,N_49500);
xor UO_3682 (O_3682,N_49575,N_49127);
nand UO_3683 (O_3683,N_49263,N_49060);
and UO_3684 (O_3684,N_49038,N_49014);
or UO_3685 (O_3685,N_49642,N_49635);
or UO_3686 (O_3686,N_49405,N_49865);
nand UO_3687 (O_3687,N_49423,N_49013);
nor UO_3688 (O_3688,N_49362,N_49283);
xor UO_3689 (O_3689,N_49077,N_49796);
and UO_3690 (O_3690,N_49731,N_49992);
xor UO_3691 (O_3691,N_49900,N_49275);
or UO_3692 (O_3692,N_49512,N_49368);
or UO_3693 (O_3693,N_49185,N_49343);
nor UO_3694 (O_3694,N_49235,N_49190);
or UO_3695 (O_3695,N_49318,N_49204);
nand UO_3696 (O_3696,N_49100,N_49977);
or UO_3697 (O_3697,N_49933,N_49010);
xnor UO_3698 (O_3698,N_49536,N_49624);
nand UO_3699 (O_3699,N_49402,N_49238);
xor UO_3700 (O_3700,N_49487,N_49721);
or UO_3701 (O_3701,N_49429,N_49618);
or UO_3702 (O_3702,N_49886,N_49002);
xor UO_3703 (O_3703,N_49244,N_49577);
or UO_3704 (O_3704,N_49750,N_49654);
xnor UO_3705 (O_3705,N_49921,N_49769);
or UO_3706 (O_3706,N_49082,N_49831);
xor UO_3707 (O_3707,N_49971,N_49705);
or UO_3708 (O_3708,N_49336,N_49307);
and UO_3709 (O_3709,N_49433,N_49374);
nand UO_3710 (O_3710,N_49062,N_49202);
and UO_3711 (O_3711,N_49172,N_49398);
and UO_3712 (O_3712,N_49708,N_49607);
xnor UO_3713 (O_3713,N_49221,N_49722);
nor UO_3714 (O_3714,N_49011,N_49749);
or UO_3715 (O_3715,N_49002,N_49945);
nand UO_3716 (O_3716,N_49599,N_49519);
and UO_3717 (O_3717,N_49626,N_49062);
or UO_3718 (O_3718,N_49105,N_49172);
nand UO_3719 (O_3719,N_49588,N_49559);
nand UO_3720 (O_3720,N_49824,N_49048);
nand UO_3721 (O_3721,N_49942,N_49182);
nor UO_3722 (O_3722,N_49497,N_49221);
or UO_3723 (O_3723,N_49359,N_49932);
nand UO_3724 (O_3724,N_49750,N_49580);
and UO_3725 (O_3725,N_49152,N_49370);
or UO_3726 (O_3726,N_49442,N_49811);
and UO_3727 (O_3727,N_49528,N_49309);
xor UO_3728 (O_3728,N_49910,N_49672);
nor UO_3729 (O_3729,N_49038,N_49804);
nand UO_3730 (O_3730,N_49018,N_49931);
and UO_3731 (O_3731,N_49744,N_49882);
nor UO_3732 (O_3732,N_49362,N_49331);
nand UO_3733 (O_3733,N_49169,N_49024);
nand UO_3734 (O_3734,N_49593,N_49865);
nor UO_3735 (O_3735,N_49138,N_49112);
nand UO_3736 (O_3736,N_49576,N_49327);
and UO_3737 (O_3737,N_49273,N_49535);
or UO_3738 (O_3738,N_49081,N_49522);
nor UO_3739 (O_3739,N_49570,N_49477);
or UO_3740 (O_3740,N_49099,N_49732);
nor UO_3741 (O_3741,N_49826,N_49322);
nand UO_3742 (O_3742,N_49655,N_49868);
xor UO_3743 (O_3743,N_49258,N_49435);
or UO_3744 (O_3744,N_49254,N_49031);
or UO_3745 (O_3745,N_49578,N_49677);
or UO_3746 (O_3746,N_49498,N_49308);
or UO_3747 (O_3747,N_49953,N_49494);
nor UO_3748 (O_3748,N_49739,N_49779);
nor UO_3749 (O_3749,N_49054,N_49318);
and UO_3750 (O_3750,N_49755,N_49484);
nor UO_3751 (O_3751,N_49730,N_49364);
and UO_3752 (O_3752,N_49256,N_49303);
nand UO_3753 (O_3753,N_49458,N_49585);
xnor UO_3754 (O_3754,N_49766,N_49458);
xnor UO_3755 (O_3755,N_49217,N_49483);
and UO_3756 (O_3756,N_49882,N_49095);
and UO_3757 (O_3757,N_49800,N_49915);
and UO_3758 (O_3758,N_49456,N_49176);
and UO_3759 (O_3759,N_49464,N_49822);
nor UO_3760 (O_3760,N_49752,N_49426);
nor UO_3761 (O_3761,N_49671,N_49731);
xnor UO_3762 (O_3762,N_49507,N_49817);
xor UO_3763 (O_3763,N_49109,N_49390);
nand UO_3764 (O_3764,N_49055,N_49922);
nand UO_3765 (O_3765,N_49702,N_49657);
or UO_3766 (O_3766,N_49159,N_49194);
or UO_3767 (O_3767,N_49685,N_49415);
and UO_3768 (O_3768,N_49748,N_49477);
and UO_3769 (O_3769,N_49243,N_49444);
nand UO_3770 (O_3770,N_49178,N_49474);
or UO_3771 (O_3771,N_49466,N_49473);
or UO_3772 (O_3772,N_49412,N_49660);
and UO_3773 (O_3773,N_49101,N_49592);
nor UO_3774 (O_3774,N_49011,N_49395);
nand UO_3775 (O_3775,N_49462,N_49715);
or UO_3776 (O_3776,N_49899,N_49190);
or UO_3777 (O_3777,N_49143,N_49533);
or UO_3778 (O_3778,N_49856,N_49738);
or UO_3779 (O_3779,N_49435,N_49528);
nand UO_3780 (O_3780,N_49554,N_49675);
or UO_3781 (O_3781,N_49325,N_49745);
xnor UO_3782 (O_3782,N_49404,N_49342);
nand UO_3783 (O_3783,N_49644,N_49641);
nand UO_3784 (O_3784,N_49417,N_49764);
nand UO_3785 (O_3785,N_49949,N_49787);
and UO_3786 (O_3786,N_49514,N_49623);
nor UO_3787 (O_3787,N_49334,N_49244);
xnor UO_3788 (O_3788,N_49201,N_49583);
and UO_3789 (O_3789,N_49440,N_49968);
nand UO_3790 (O_3790,N_49725,N_49758);
xor UO_3791 (O_3791,N_49607,N_49934);
nand UO_3792 (O_3792,N_49441,N_49292);
nor UO_3793 (O_3793,N_49396,N_49497);
xor UO_3794 (O_3794,N_49277,N_49783);
and UO_3795 (O_3795,N_49164,N_49527);
xnor UO_3796 (O_3796,N_49248,N_49245);
or UO_3797 (O_3797,N_49185,N_49554);
or UO_3798 (O_3798,N_49545,N_49833);
or UO_3799 (O_3799,N_49129,N_49419);
xnor UO_3800 (O_3800,N_49351,N_49868);
and UO_3801 (O_3801,N_49363,N_49753);
nand UO_3802 (O_3802,N_49807,N_49210);
xnor UO_3803 (O_3803,N_49090,N_49875);
or UO_3804 (O_3804,N_49978,N_49050);
nor UO_3805 (O_3805,N_49889,N_49479);
or UO_3806 (O_3806,N_49432,N_49041);
xor UO_3807 (O_3807,N_49490,N_49368);
xor UO_3808 (O_3808,N_49784,N_49363);
or UO_3809 (O_3809,N_49692,N_49413);
and UO_3810 (O_3810,N_49814,N_49665);
or UO_3811 (O_3811,N_49981,N_49435);
nand UO_3812 (O_3812,N_49325,N_49666);
and UO_3813 (O_3813,N_49780,N_49207);
and UO_3814 (O_3814,N_49369,N_49750);
and UO_3815 (O_3815,N_49657,N_49139);
xor UO_3816 (O_3816,N_49796,N_49755);
xnor UO_3817 (O_3817,N_49809,N_49636);
xor UO_3818 (O_3818,N_49979,N_49859);
and UO_3819 (O_3819,N_49630,N_49940);
or UO_3820 (O_3820,N_49171,N_49523);
or UO_3821 (O_3821,N_49974,N_49264);
nand UO_3822 (O_3822,N_49856,N_49160);
nor UO_3823 (O_3823,N_49949,N_49254);
xor UO_3824 (O_3824,N_49421,N_49980);
xnor UO_3825 (O_3825,N_49412,N_49560);
xnor UO_3826 (O_3826,N_49401,N_49903);
nor UO_3827 (O_3827,N_49710,N_49581);
nor UO_3828 (O_3828,N_49717,N_49984);
or UO_3829 (O_3829,N_49623,N_49419);
nor UO_3830 (O_3830,N_49161,N_49840);
or UO_3831 (O_3831,N_49957,N_49997);
xnor UO_3832 (O_3832,N_49806,N_49594);
or UO_3833 (O_3833,N_49100,N_49487);
and UO_3834 (O_3834,N_49628,N_49795);
nor UO_3835 (O_3835,N_49456,N_49450);
xnor UO_3836 (O_3836,N_49709,N_49027);
nor UO_3837 (O_3837,N_49809,N_49582);
and UO_3838 (O_3838,N_49466,N_49634);
xnor UO_3839 (O_3839,N_49590,N_49890);
nand UO_3840 (O_3840,N_49517,N_49832);
and UO_3841 (O_3841,N_49251,N_49380);
nand UO_3842 (O_3842,N_49986,N_49399);
nor UO_3843 (O_3843,N_49016,N_49215);
nand UO_3844 (O_3844,N_49137,N_49784);
and UO_3845 (O_3845,N_49364,N_49768);
or UO_3846 (O_3846,N_49522,N_49682);
nor UO_3847 (O_3847,N_49860,N_49046);
xor UO_3848 (O_3848,N_49260,N_49516);
or UO_3849 (O_3849,N_49500,N_49048);
or UO_3850 (O_3850,N_49686,N_49103);
nor UO_3851 (O_3851,N_49088,N_49661);
xor UO_3852 (O_3852,N_49520,N_49249);
nor UO_3853 (O_3853,N_49439,N_49972);
xor UO_3854 (O_3854,N_49708,N_49035);
and UO_3855 (O_3855,N_49227,N_49535);
or UO_3856 (O_3856,N_49322,N_49183);
or UO_3857 (O_3857,N_49040,N_49953);
xor UO_3858 (O_3858,N_49860,N_49180);
and UO_3859 (O_3859,N_49268,N_49791);
nor UO_3860 (O_3860,N_49634,N_49373);
or UO_3861 (O_3861,N_49553,N_49820);
nor UO_3862 (O_3862,N_49598,N_49030);
nand UO_3863 (O_3863,N_49607,N_49391);
and UO_3864 (O_3864,N_49322,N_49543);
xnor UO_3865 (O_3865,N_49697,N_49244);
and UO_3866 (O_3866,N_49160,N_49378);
nand UO_3867 (O_3867,N_49254,N_49835);
nand UO_3868 (O_3868,N_49913,N_49040);
and UO_3869 (O_3869,N_49071,N_49575);
or UO_3870 (O_3870,N_49935,N_49811);
nand UO_3871 (O_3871,N_49291,N_49428);
or UO_3872 (O_3872,N_49624,N_49870);
xnor UO_3873 (O_3873,N_49755,N_49694);
and UO_3874 (O_3874,N_49179,N_49709);
nand UO_3875 (O_3875,N_49835,N_49545);
xnor UO_3876 (O_3876,N_49553,N_49548);
and UO_3877 (O_3877,N_49525,N_49871);
or UO_3878 (O_3878,N_49949,N_49147);
and UO_3879 (O_3879,N_49868,N_49031);
nor UO_3880 (O_3880,N_49509,N_49427);
and UO_3881 (O_3881,N_49416,N_49336);
xnor UO_3882 (O_3882,N_49841,N_49798);
and UO_3883 (O_3883,N_49432,N_49246);
or UO_3884 (O_3884,N_49045,N_49495);
and UO_3885 (O_3885,N_49381,N_49548);
xor UO_3886 (O_3886,N_49786,N_49260);
nand UO_3887 (O_3887,N_49111,N_49007);
or UO_3888 (O_3888,N_49160,N_49559);
nor UO_3889 (O_3889,N_49708,N_49477);
nand UO_3890 (O_3890,N_49864,N_49436);
or UO_3891 (O_3891,N_49485,N_49255);
or UO_3892 (O_3892,N_49987,N_49630);
or UO_3893 (O_3893,N_49987,N_49299);
nand UO_3894 (O_3894,N_49039,N_49258);
or UO_3895 (O_3895,N_49406,N_49361);
xor UO_3896 (O_3896,N_49560,N_49142);
or UO_3897 (O_3897,N_49253,N_49908);
or UO_3898 (O_3898,N_49547,N_49246);
xor UO_3899 (O_3899,N_49036,N_49549);
nand UO_3900 (O_3900,N_49036,N_49117);
nor UO_3901 (O_3901,N_49836,N_49376);
xnor UO_3902 (O_3902,N_49048,N_49665);
xor UO_3903 (O_3903,N_49424,N_49996);
nor UO_3904 (O_3904,N_49708,N_49114);
and UO_3905 (O_3905,N_49256,N_49090);
or UO_3906 (O_3906,N_49867,N_49920);
and UO_3907 (O_3907,N_49796,N_49350);
nor UO_3908 (O_3908,N_49571,N_49362);
xnor UO_3909 (O_3909,N_49177,N_49241);
nor UO_3910 (O_3910,N_49655,N_49714);
xor UO_3911 (O_3911,N_49893,N_49773);
xor UO_3912 (O_3912,N_49492,N_49795);
and UO_3913 (O_3913,N_49497,N_49496);
nor UO_3914 (O_3914,N_49327,N_49877);
nor UO_3915 (O_3915,N_49811,N_49425);
and UO_3916 (O_3916,N_49815,N_49098);
or UO_3917 (O_3917,N_49748,N_49074);
and UO_3918 (O_3918,N_49738,N_49276);
nand UO_3919 (O_3919,N_49230,N_49202);
or UO_3920 (O_3920,N_49753,N_49658);
nor UO_3921 (O_3921,N_49625,N_49804);
nand UO_3922 (O_3922,N_49254,N_49506);
nor UO_3923 (O_3923,N_49504,N_49966);
nor UO_3924 (O_3924,N_49590,N_49491);
nor UO_3925 (O_3925,N_49118,N_49461);
and UO_3926 (O_3926,N_49564,N_49889);
and UO_3927 (O_3927,N_49792,N_49728);
or UO_3928 (O_3928,N_49467,N_49811);
nor UO_3929 (O_3929,N_49773,N_49445);
nor UO_3930 (O_3930,N_49296,N_49056);
or UO_3931 (O_3931,N_49622,N_49762);
nor UO_3932 (O_3932,N_49253,N_49483);
nor UO_3933 (O_3933,N_49821,N_49156);
xnor UO_3934 (O_3934,N_49549,N_49227);
or UO_3935 (O_3935,N_49368,N_49406);
and UO_3936 (O_3936,N_49537,N_49111);
nand UO_3937 (O_3937,N_49127,N_49040);
nor UO_3938 (O_3938,N_49568,N_49846);
xor UO_3939 (O_3939,N_49747,N_49768);
nor UO_3940 (O_3940,N_49712,N_49477);
xor UO_3941 (O_3941,N_49148,N_49103);
xor UO_3942 (O_3942,N_49594,N_49508);
xor UO_3943 (O_3943,N_49079,N_49186);
or UO_3944 (O_3944,N_49952,N_49457);
and UO_3945 (O_3945,N_49628,N_49052);
nand UO_3946 (O_3946,N_49544,N_49751);
nand UO_3947 (O_3947,N_49237,N_49054);
or UO_3948 (O_3948,N_49124,N_49343);
xor UO_3949 (O_3949,N_49337,N_49192);
or UO_3950 (O_3950,N_49195,N_49747);
xnor UO_3951 (O_3951,N_49094,N_49183);
and UO_3952 (O_3952,N_49049,N_49512);
or UO_3953 (O_3953,N_49060,N_49042);
nand UO_3954 (O_3954,N_49195,N_49226);
nor UO_3955 (O_3955,N_49179,N_49281);
or UO_3956 (O_3956,N_49540,N_49596);
xor UO_3957 (O_3957,N_49451,N_49426);
or UO_3958 (O_3958,N_49375,N_49567);
xor UO_3959 (O_3959,N_49919,N_49983);
xnor UO_3960 (O_3960,N_49135,N_49120);
and UO_3961 (O_3961,N_49830,N_49522);
xor UO_3962 (O_3962,N_49074,N_49916);
and UO_3963 (O_3963,N_49211,N_49479);
xor UO_3964 (O_3964,N_49869,N_49326);
xnor UO_3965 (O_3965,N_49072,N_49295);
nand UO_3966 (O_3966,N_49348,N_49385);
xnor UO_3967 (O_3967,N_49791,N_49845);
nand UO_3968 (O_3968,N_49187,N_49286);
and UO_3969 (O_3969,N_49219,N_49213);
or UO_3970 (O_3970,N_49988,N_49758);
xor UO_3971 (O_3971,N_49411,N_49640);
nand UO_3972 (O_3972,N_49499,N_49374);
nor UO_3973 (O_3973,N_49574,N_49843);
and UO_3974 (O_3974,N_49079,N_49693);
and UO_3975 (O_3975,N_49998,N_49125);
nand UO_3976 (O_3976,N_49503,N_49034);
and UO_3977 (O_3977,N_49097,N_49526);
and UO_3978 (O_3978,N_49864,N_49662);
xnor UO_3979 (O_3979,N_49669,N_49116);
and UO_3980 (O_3980,N_49619,N_49995);
xor UO_3981 (O_3981,N_49691,N_49972);
xor UO_3982 (O_3982,N_49855,N_49313);
and UO_3983 (O_3983,N_49591,N_49091);
nor UO_3984 (O_3984,N_49092,N_49049);
and UO_3985 (O_3985,N_49371,N_49370);
nand UO_3986 (O_3986,N_49014,N_49265);
and UO_3987 (O_3987,N_49873,N_49674);
xnor UO_3988 (O_3988,N_49411,N_49309);
or UO_3989 (O_3989,N_49699,N_49214);
or UO_3990 (O_3990,N_49793,N_49533);
and UO_3991 (O_3991,N_49695,N_49303);
or UO_3992 (O_3992,N_49831,N_49992);
nor UO_3993 (O_3993,N_49283,N_49656);
xnor UO_3994 (O_3994,N_49450,N_49346);
nor UO_3995 (O_3995,N_49760,N_49718);
nand UO_3996 (O_3996,N_49656,N_49895);
nand UO_3997 (O_3997,N_49401,N_49971);
xnor UO_3998 (O_3998,N_49975,N_49931);
nor UO_3999 (O_3999,N_49022,N_49861);
xor UO_4000 (O_4000,N_49740,N_49318);
and UO_4001 (O_4001,N_49739,N_49312);
xor UO_4002 (O_4002,N_49593,N_49539);
and UO_4003 (O_4003,N_49373,N_49450);
xnor UO_4004 (O_4004,N_49578,N_49987);
nor UO_4005 (O_4005,N_49645,N_49698);
and UO_4006 (O_4006,N_49257,N_49611);
xnor UO_4007 (O_4007,N_49748,N_49661);
or UO_4008 (O_4008,N_49156,N_49096);
or UO_4009 (O_4009,N_49151,N_49876);
xnor UO_4010 (O_4010,N_49476,N_49286);
nor UO_4011 (O_4011,N_49108,N_49131);
nor UO_4012 (O_4012,N_49670,N_49493);
or UO_4013 (O_4013,N_49520,N_49471);
or UO_4014 (O_4014,N_49646,N_49265);
and UO_4015 (O_4015,N_49394,N_49612);
xnor UO_4016 (O_4016,N_49696,N_49419);
or UO_4017 (O_4017,N_49771,N_49809);
nor UO_4018 (O_4018,N_49572,N_49722);
xnor UO_4019 (O_4019,N_49898,N_49735);
nand UO_4020 (O_4020,N_49720,N_49507);
and UO_4021 (O_4021,N_49261,N_49049);
and UO_4022 (O_4022,N_49233,N_49694);
or UO_4023 (O_4023,N_49421,N_49336);
xor UO_4024 (O_4024,N_49389,N_49928);
xnor UO_4025 (O_4025,N_49147,N_49132);
xnor UO_4026 (O_4026,N_49151,N_49180);
nor UO_4027 (O_4027,N_49312,N_49941);
and UO_4028 (O_4028,N_49971,N_49223);
xor UO_4029 (O_4029,N_49462,N_49837);
nor UO_4030 (O_4030,N_49654,N_49417);
or UO_4031 (O_4031,N_49170,N_49327);
nand UO_4032 (O_4032,N_49550,N_49460);
xor UO_4033 (O_4033,N_49483,N_49704);
and UO_4034 (O_4034,N_49101,N_49027);
nor UO_4035 (O_4035,N_49601,N_49661);
xor UO_4036 (O_4036,N_49194,N_49904);
and UO_4037 (O_4037,N_49826,N_49435);
nor UO_4038 (O_4038,N_49216,N_49656);
or UO_4039 (O_4039,N_49112,N_49752);
nand UO_4040 (O_4040,N_49097,N_49126);
nand UO_4041 (O_4041,N_49940,N_49059);
or UO_4042 (O_4042,N_49276,N_49367);
nand UO_4043 (O_4043,N_49096,N_49381);
nor UO_4044 (O_4044,N_49354,N_49780);
and UO_4045 (O_4045,N_49714,N_49616);
or UO_4046 (O_4046,N_49538,N_49739);
or UO_4047 (O_4047,N_49498,N_49018);
xor UO_4048 (O_4048,N_49567,N_49870);
nor UO_4049 (O_4049,N_49558,N_49380);
nand UO_4050 (O_4050,N_49245,N_49303);
or UO_4051 (O_4051,N_49992,N_49866);
nor UO_4052 (O_4052,N_49440,N_49771);
or UO_4053 (O_4053,N_49686,N_49282);
xor UO_4054 (O_4054,N_49119,N_49050);
xnor UO_4055 (O_4055,N_49506,N_49038);
and UO_4056 (O_4056,N_49039,N_49975);
xor UO_4057 (O_4057,N_49127,N_49491);
xor UO_4058 (O_4058,N_49261,N_49129);
and UO_4059 (O_4059,N_49591,N_49216);
and UO_4060 (O_4060,N_49560,N_49708);
xor UO_4061 (O_4061,N_49930,N_49368);
or UO_4062 (O_4062,N_49040,N_49046);
xor UO_4063 (O_4063,N_49964,N_49726);
nand UO_4064 (O_4064,N_49791,N_49121);
nor UO_4065 (O_4065,N_49010,N_49082);
nor UO_4066 (O_4066,N_49333,N_49458);
and UO_4067 (O_4067,N_49444,N_49837);
nor UO_4068 (O_4068,N_49723,N_49323);
xor UO_4069 (O_4069,N_49628,N_49959);
and UO_4070 (O_4070,N_49824,N_49579);
and UO_4071 (O_4071,N_49212,N_49418);
nor UO_4072 (O_4072,N_49704,N_49930);
and UO_4073 (O_4073,N_49584,N_49099);
and UO_4074 (O_4074,N_49654,N_49244);
nand UO_4075 (O_4075,N_49209,N_49733);
and UO_4076 (O_4076,N_49208,N_49683);
xor UO_4077 (O_4077,N_49018,N_49425);
and UO_4078 (O_4078,N_49739,N_49589);
or UO_4079 (O_4079,N_49602,N_49916);
or UO_4080 (O_4080,N_49947,N_49013);
nand UO_4081 (O_4081,N_49295,N_49173);
or UO_4082 (O_4082,N_49435,N_49065);
nor UO_4083 (O_4083,N_49963,N_49252);
xor UO_4084 (O_4084,N_49983,N_49062);
nor UO_4085 (O_4085,N_49291,N_49711);
and UO_4086 (O_4086,N_49248,N_49254);
or UO_4087 (O_4087,N_49502,N_49024);
and UO_4088 (O_4088,N_49701,N_49525);
and UO_4089 (O_4089,N_49087,N_49147);
xnor UO_4090 (O_4090,N_49725,N_49826);
and UO_4091 (O_4091,N_49544,N_49949);
xnor UO_4092 (O_4092,N_49045,N_49838);
and UO_4093 (O_4093,N_49318,N_49882);
or UO_4094 (O_4094,N_49871,N_49431);
nand UO_4095 (O_4095,N_49795,N_49602);
xnor UO_4096 (O_4096,N_49734,N_49510);
and UO_4097 (O_4097,N_49096,N_49833);
nor UO_4098 (O_4098,N_49685,N_49002);
and UO_4099 (O_4099,N_49602,N_49997);
or UO_4100 (O_4100,N_49103,N_49358);
nand UO_4101 (O_4101,N_49455,N_49290);
and UO_4102 (O_4102,N_49410,N_49771);
or UO_4103 (O_4103,N_49478,N_49185);
and UO_4104 (O_4104,N_49975,N_49948);
and UO_4105 (O_4105,N_49894,N_49312);
nand UO_4106 (O_4106,N_49065,N_49221);
xnor UO_4107 (O_4107,N_49585,N_49704);
or UO_4108 (O_4108,N_49042,N_49767);
nand UO_4109 (O_4109,N_49861,N_49153);
or UO_4110 (O_4110,N_49234,N_49190);
nor UO_4111 (O_4111,N_49637,N_49586);
or UO_4112 (O_4112,N_49897,N_49081);
xnor UO_4113 (O_4113,N_49539,N_49040);
and UO_4114 (O_4114,N_49318,N_49031);
xor UO_4115 (O_4115,N_49406,N_49539);
or UO_4116 (O_4116,N_49904,N_49324);
nor UO_4117 (O_4117,N_49679,N_49939);
or UO_4118 (O_4118,N_49378,N_49794);
nor UO_4119 (O_4119,N_49225,N_49614);
and UO_4120 (O_4120,N_49528,N_49070);
nand UO_4121 (O_4121,N_49562,N_49368);
xnor UO_4122 (O_4122,N_49571,N_49458);
xnor UO_4123 (O_4123,N_49959,N_49597);
xor UO_4124 (O_4124,N_49783,N_49592);
or UO_4125 (O_4125,N_49454,N_49455);
or UO_4126 (O_4126,N_49723,N_49137);
xor UO_4127 (O_4127,N_49735,N_49970);
and UO_4128 (O_4128,N_49877,N_49982);
nor UO_4129 (O_4129,N_49178,N_49620);
or UO_4130 (O_4130,N_49487,N_49158);
nand UO_4131 (O_4131,N_49939,N_49754);
nand UO_4132 (O_4132,N_49456,N_49897);
xnor UO_4133 (O_4133,N_49028,N_49320);
xor UO_4134 (O_4134,N_49516,N_49496);
nand UO_4135 (O_4135,N_49120,N_49181);
xor UO_4136 (O_4136,N_49854,N_49718);
xor UO_4137 (O_4137,N_49895,N_49860);
nand UO_4138 (O_4138,N_49663,N_49722);
nor UO_4139 (O_4139,N_49089,N_49747);
nor UO_4140 (O_4140,N_49803,N_49575);
xor UO_4141 (O_4141,N_49190,N_49575);
nor UO_4142 (O_4142,N_49845,N_49686);
nand UO_4143 (O_4143,N_49633,N_49897);
nand UO_4144 (O_4144,N_49033,N_49841);
nand UO_4145 (O_4145,N_49131,N_49815);
and UO_4146 (O_4146,N_49951,N_49346);
and UO_4147 (O_4147,N_49483,N_49964);
nor UO_4148 (O_4148,N_49716,N_49676);
nor UO_4149 (O_4149,N_49249,N_49958);
xnor UO_4150 (O_4150,N_49477,N_49377);
nor UO_4151 (O_4151,N_49552,N_49004);
nand UO_4152 (O_4152,N_49625,N_49882);
xor UO_4153 (O_4153,N_49515,N_49812);
nand UO_4154 (O_4154,N_49282,N_49608);
xnor UO_4155 (O_4155,N_49008,N_49301);
xor UO_4156 (O_4156,N_49277,N_49129);
or UO_4157 (O_4157,N_49552,N_49162);
and UO_4158 (O_4158,N_49452,N_49444);
nand UO_4159 (O_4159,N_49349,N_49283);
nand UO_4160 (O_4160,N_49305,N_49643);
nor UO_4161 (O_4161,N_49859,N_49515);
or UO_4162 (O_4162,N_49665,N_49701);
and UO_4163 (O_4163,N_49310,N_49872);
nor UO_4164 (O_4164,N_49511,N_49894);
or UO_4165 (O_4165,N_49666,N_49642);
nor UO_4166 (O_4166,N_49152,N_49440);
or UO_4167 (O_4167,N_49795,N_49791);
xnor UO_4168 (O_4168,N_49575,N_49858);
nor UO_4169 (O_4169,N_49537,N_49944);
and UO_4170 (O_4170,N_49148,N_49310);
nand UO_4171 (O_4171,N_49219,N_49535);
and UO_4172 (O_4172,N_49071,N_49852);
nand UO_4173 (O_4173,N_49950,N_49680);
nor UO_4174 (O_4174,N_49349,N_49927);
and UO_4175 (O_4175,N_49080,N_49648);
and UO_4176 (O_4176,N_49606,N_49048);
nand UO_4177 (O_4177,N_49868,N_49751);
nand UO_4178 (O_4178,N_49479,N_49456);
xor UO_4179 (O_4179,N_49438,N_49363);
nor UO_4180 (O_4180,N_49232,N_49241);
or UO_4181 (O_4181,N_49237,N_49408);
and UO_4182 (O_4182,N_49985,N_49782);
and UO_4183 (O_4183,N_49175,N_49301);
and UO_4184 (O_4184,N_49808,N_49598);
nor UO_4185 (O_4185,N_49056,N_49313);
nor UO_4186 (O_4186,N_49346,N_49371);
nand UO_4187 (O_4187,N_49036,N_49587);
and UO_4188 (O_4188,N_49119,N_49156);
or UO_4189 (O_4189,N_49410,N_49357);
and UO_4190 (O_4190,N_49199,N_49918);
or UO_4191 (O_4191,N_49727,N_49194);
xor UO_4192 (O_4192,N_49475,N_49892);
or UO_4193 (O_4193,N_49236,N_49602);
nand UO_4194 (O_4194,N_49029,N_49927);
or UO_4195 (O_4195,N_49073,N_49198);
nand UO_4196 (O_4196,N_49525,N_49169);
and UO_4197 (O_4197,N_49348,N_49332);
xor UO_4198 (O_4198,N_49661,N_49722);
or UO_4199 (O_4199,N_49699,N_49918);
xor UO_4200 (O_4200,N_49540,N_49879);
and UO_4201 (O_4201,N_49021,N_49874);
or UO_4202 (O_4202,N_49236,N_49548);
nand UO_4203 (O_4203,N_49764,N_49013);
nor UO_4204 (O_4204,N_49646,N_49698);
nor UO_4205 (O_4205,N_49763,N_49713);
nand UO_4206 (O_4206,N_49058,N_49750);
nor UO_4207 (O_4207,N_49883,N_49376);
and UO_4208 (O_4208,N_49919,N_49482);
xnor UO_4209 (O_4209,N_49858,N_49480);
or UO_4210 (O_4210,N_49079,N_49459);
or UO_4211 (O_4211,N_49172,N_49653);
nand UO_4212 (O_4212,N_49392,N_49671);
nand UO_4213 (O_4213,N_49783,N_49055);
nand UO_4214 (O_4214,N_49819,N_49552);
xnor UO_4215 (O_4215,N_49993,N_49918);
nor UO_4216 (O_4216,N_49976,N_49342);
or UO_4217 (O_4217,N_49803,N_49163);
xor UO_4218 (O_4218,N_49778,N_49077);
xnor UO_4219 (O_4219,N_49950,N_49145);
nand UO_4220 (O_4220,N_49081,N_49498);
and UO_4221 (O_4221,N_49205,N_49644);
nand UO_4222 (O_4222,N_49427,N_49857);
nor UO_4223 (O_4223,N_49037,N_49572);
or UO_4224 (O_4224,N_49509,N_49905);
xnor UO_4225 (O_4225,N_49055,N_49959);
xor UO_4226 (O_4226,N_49570,N_49709);
nor UO_4227 (O_4227,N_49587,N_49130);
nand UO_4228 (O_4228,N_49001,N_49698);
nor UO_4229 (O_4229,N_49593,N_49779);
nor UO_4230 (O_4230,N_49891,N_49280);
or UO_4231 (O_4231,N_49785,N_49608);
nor UO_4232 (O_4232,N_49976,N_49993);
xnor UO_4233 (O_4233,N_49997,N_49276);
nor UO_4234 (O_4234,N_49857,N_49850);
or UO_4235 (O_4235,N_49433,N_49948);
xnor UO_4236 (O_4236,N_49197,N_49193);
nor UO_4237 (O_4237,N_49906,N_49202);
xnor UO_4238 (O_4238,N_49892,N_49788);
xor UO_4239 (O_4239,N_49939,N_49384);
nand UO_4240 (O_4240,N_49849,N_49303);
or UO_4241 (O_4241,N_49805,N_49352);
or UO_4242 (O_4242,N_49686,N_49562);
nor UO_4243 (O_4243,N_49918,N_49877);
xnor UO_4244 (O_4244,N_49708,N_49338);
or UO_4245 (O_4245,N_49362,N_49550);
nand UO_4246 (O_4246,N_49825,N_49721);
xnor UO_4247 (O_4247,N_49178,N_49354);
xor UO_4248 (O_4248,N_49369,N_49647);
and UO_4249 (O_4249,N_49213,N_49734);
and UO_4250 (O_4250,N_49388,N_49206);
or UO_4251 (O_4251,N_49233,N_49087);
or UO_4252 (O_4252,N_49607,N_49414);
and UO_4253 (O_4253,N_49077,N_49926);
xnor UO_4254 (O_4254,N_49699,N_49272);
nor UO_4255 (O_4255,N_49323,N_49532);
nand UO_4256 (O_4256,N_49613,N_49866);
nor UO_4257 (O_4257,N_49634,N_49880);
or UO_4258 (O_4258,N_49562,N_49921);
nor UO_4259 (O_4259,N_49093,N_49405);
xor UO_4260 (O_4260,N_49923,N_49282);
and UO_4261 (O_4261,N_49921,N_49285);
nand UO_4262 (O_4262,N_49423,N_49728);
xnor UO_4263 (O_4263,N_49315,N_49700);
nor UO_4264 (O_4264,N_49121,N_49037);
or UO_4265 (O_4265,N_49203,N_49693);
nor UO_4266 (O_4266,N_49227,N_49777);
and UO_4267 (O_4267,N_49243,N_49316);
and UO_4268 (O_4268,N_49311,N_49831);
xnor UO_4269 (O_4269,N_49789,N_49797);
nor UO_4270 (O_4270,N_49086,N_49092);
nand UO_4271 (O_4271,N_49656,N_49735);
and UO_4272 (O_4272,N_49700,N_49688);
nor UO_4273 (O_4273,N_49304,N_49824);
or UO_4274 (O_4274,N_49534,N_49485);
nand UO_4275 (O_4275,N_49730,N_49671);
or UO_4276 (O_4276,N_49367,N_49139);
nand UO_4277 (O_4277,N_49028,N_49920);
nor UO_4278 (O_4278,N_49048,N_49477);
xor UO_4279 (O_4279,N_49244,N_49028);
or UO_4280 (O_4280,N_49230,N_49055);
nand UO_4281 (O_4281,N_49197,N_49113);
nor UO_4282 (O_4282,N_49512,N_49369);
nand UO_4283 (O_4283,N_49279,N_49627);
and UO_4284 (O_4284,N_49254,N_49548);
nand UO_4285 (O_4285,N_49411,N_49339);
or UO_4286 (O_4286,N_49386,N_49439);
and UO_4287 (O_4287,N_49984,N_49812);
or UO_4288 (O_4288,N_49413,N_49945);
and UO_4289 (O_4289,N_49710,N_49499);
nor UO_4290 (O_4290,N_49056,N_49428);
xnor UO_4291 (O_4291,N_49769,N_49393);
nor UO_4292 (O_4292,N_49893,N_49374);
and UO_4293 (O_4293,N_49381,N_49726);
or UO_4294 (O_4294,N_49607,N_49342);
nor UO_4295 (O_4295,N_49734,N_49190);
and UO_4296 (O_4296,N_49393,N_49074);
nand UO_4297 (O_4297,N_49224,N_49247);
or UO_4298 (O_4298,N_49494,N_49036);
or UO_4299 (O_4299,N_49921,N_49178);
xor UO_4300 (O_4300,N_49196,N_49905);
or UO_4301 (O_4301,N_49776,N_49123);
nand UO_4302 (O_4302,N_49389,N_49232);
and UO_4303 (O_4303,N_49710,N_49146);
nand UO_4304 (O_4304,N_49953,N_49073);
nor UO_4305 (O_4305,N_49822,N_49694);
nor UO_4306 (O_4306,N_49927,N_49682);
or UO_4307 (O_4307,N_49799,N_49289);
xnor UO_4308 (O_4308,N_49317,N_49023);
nand UO_4309 (O_4309,N_49187,N_49457);
nand UO_4310 (O_4310,N_49882,N_49741);
nand UO_4311 (O_4311,N_49029,N_49985);
nor UO_4312 (O_4312,N_49058,N_49006);
nand UO_4313 (O_4313,N_49070,N_49347);
xnor UO_4314 (O_4314,N_49567,N_49486);
xnor UO_4315 (O_4315,N_49019,N_49517);
or UO_4316 (O_4316,N_49100,N_49666);
or UO_4317 (O_4317,N_49663,N_49411);
nor UO_4318 (O_4318,N_49195,N_49661);
nor UO_4319 (O_4319,N_49596,N_49421);
xor UO_4320 (O_4320,N_49986,N_49773);
or UO_4321 (O_4321,N_49327,N_49373);
nand UO_4322 (O_4322,N_49579,N_49713);
nor UO_4323 (O_4323,N_49801,N_49943);
nand UO_4324 (O_4324,N_49893,N_49497);
xor UO_4325 (O_4325,N_49717,N_49710);
nand UO_4326 (O_4326,N_49822,N_49664);
nor UO_4327 (O_4327,N_49906,N_49656);
and UO_4328 (O_4328,N_49153,N_49676);
xnor UO_4329 (O_4329,N_49996,N_49067);
nor UO_4330 (O_4330,N_49138,N_49752);
or UO_4331 (O_4331,N_49224,N_49537);
nand UO_4332 (O_4332,N_49966,N_49556);
nand UO_4333 (O_4333,N_49237,N_49045);
nor UO_4334 (O_4334,N_49559,N_49298);
nor UO_4335 (O_4335,N_49710,N_49833);
nor UO_4336 (O_4336,N_49584,N_49618);
and UO_4337 (O_4337,N_49263,N_49966);
or UO_4338 (O_4338,N_49205,N_49266);
xnor UO_4339 (O_4339,N_49383,N_49779);
or UO_4340 (O_4340,N_49239,N_49170);
and UO_4341 (O_4341,N_49865,N_49602);
nor UO_4342 (O_4342,N_49435,N_49007);
nand UO_4343 (O_4343,N_49640,N_49965);
xnor UO_4344 (O_4344,N_49770,N_49631);
nor UO_4345 (O_4345,N_49699,N_49268);
and UO_4346 (O_4346,N_49926,N_49076);
or UO_4347 (O_4347,N_49791,N_49861);
nand UO_4348 (O_4348,N_49307,N_49210);
or UO_4349 (O_4349,N_49067,N_49888);
nand UO_4350 (O_4350,N_49274,N_49164);
nor UO_4351 (O_4351,N_49913,N_49382);
or UO_4352 (O_4352,N_49179,N_49294);
and UO_4353 (O_4353,N_49995,N_49192);
or UO_4354 (O_4354,N_49149,N_49286);
and UO_4355 (O_4355,N_49731,N_49061);
nor UO_4356 (O_4356,N_49006,N_49665);
nor UO_4357 (O_4357,N_49695,N_49916);
or UO_4358 (O_4358,N_49122,N_49286);
xnor UO_4359 (O_4359,N_49551,N_49089);
or UO_4360 (O_4360,N_49990,N_49320);
nor UO_4361 (O_4361,N_49158,N_49226);
xor UO_4362 (O_4362,N_49890,N_49150);
and UO_4363 (O_4363,N_49867,N_49705);
and UO_4364 (O_4364,N_49965,N_49881);
nor UO_4365 (O_4365,N_49858,N_49083);
xor UO_4366 (O_4366,N_49228,N_49623);
nand UO_4367 (O_4367,N_49377,N_49727);
nand UO_4368 (O_4368,N_49806,N_49429);
nor UO_4369 (O_4369,N_49450,N_49850);
or UO_4370 (O_4370,N_49279,N_49818);
or UO_4371 (O_4371,N_49144,N_49629);
nor UO_4372 (O_4372,N_49816,N_49109);
nor UO_4373 (O_4373,N_49974,N_49041);
and UO_4374 (O_4374,N_49721,N_49593);
and UO_4375 (O_4375,N_49922,N_49685);
nor UO_4376 (O_4376,N_49230,N_49342);
xor UO_4377 (O_4377,N_49810,N_49782);
or UO_4378 (O_4378,N_49286,N_49894);
xnor UO_4379 (O_4379,N_49244,N_49376);
nor UO_4380 (O_4380,N_49319,N_49450);
nor UO_4381 (O_4381,N_49286,N_49177);
or UO_4382 (O_4382,N_49972,N_49023);
and UO_4383 (O_4383,N_49272,N_49401);
and UO_4384 (O_4384,N_49997,N_49213);
and UO_4385 (O_4385,N_49959,N_49754);
and UO_4386 (O_4386,N_49567,N_49604);
and UO_4387 (O_4387,N_49897,N_49672);
nand UO_4388 (O_4388,N_49322,N_49934);
or UO_4389 (O_4389,N_49679,N_49680);
xnor UO_4390 (O_4390,N_49262,N_49742);
xnor UO_4391 (O_4391,N_49923,N_49917);
nand UO_4392 (O_4392,N_49136,N_49429);
nor UO_4393 (O_4393,N_49069,N_49218);
or UO_4394 (O_4394,N_49820,N_49026);
xnor UO_4395 (O_4395,N_49459,N_49389);
and UO_4396 (O_4396,N_49608,N_49650);
nand UO_4397 (O_4397,N_49354,N_49704);
xnor UO_4398 (O_4398,N_49876,N_49706);
and UO_4399 (O_4399,N_49506,N_49526);
or UO_4400 (O_4400,N_49038,N_49627);
and UO_4401 (O_4401,N_49696,N_49403);
nor UO_4402 (O_4402,N_49529,N_49275);
xnor UO_4403 (O_4403,N_49928,N_49477);
nand UO_4404 (O_4404,N_49081,N_49511);
or UO_4405 (O_4405,N_49858,N_49970);
nor UO_4406 (O_4406,N_49201,N_49633);
and UO_4407 (O_4407,N_49071,N_49609);
and UO_4408 (O_4408,N_49214,N_49720);
nand UO_4409 (O_4409,N_49629,N_49263);
or UO_4410 (O_4410,N_49626,N_49441);
nand UO_4411 (O_4411,N_49097,N_49596);
nor UO_4412 (O_4412,N_49615,N_49585);
or UO_4413 (O_4413,N_49586,N_49778);
and UO_4414 (O_4414,N_49936,N_49794);
nand UO_4415 (O_4415,N_49663,N_49761);
nand UO_4416 (O_4416,N_49614,N_49658);
nand UO_4417 (O_4417,N_49689,N_49592);
xor UO_4418 (O_4418,N_49514,N_49607);
nand UO_4419 (O_4419,N_49288,N_49786);
nand UO_4420 (O_4420,N_49064,N_49996);
nand UO_4421 (O_4421,N_49620,N_49133);
xnor UO_4422 (O_4422,N_49866,N_49916);
and UO_4423 (O_4423,N_49656,N_49409);
nor UO_4424 (O_4424,N_49951,N_49081);
nor UO_4425 (O_4425,N_49666,N_49273);
or UO_4426 (O_4426,N_49154,N_49394);
xor UO_4427 (O_4427,N_49163,N_49424);
and UO_4428 (O_4428,N_49536,N_49871);
and UO_4429 (O_4429,N_49194,N_49167);
or UO_4430 (O_4430,N_49941,N_49129);
and UO_4431 (O_4431,N_49370,N_49784);
xor UO_4432 (O_4432,N_49209,N_49130);
nand UO_4433 (O_4433,N_49753,N_49852);
nand UO_4434 (O_4434,N_49006,N_49616);
nor UO_4435 (O_4435,N_49258,N_49607);
xnor UO_4436 (O_4436,N_49458,N_49563);
or UO_4437 (O_4437,N_49210,N_49190);
nor UO_4438 (O_4438,N_49131,N_49410);
nand UO_4439 (O_4439,N_49933,N_49430);
nand UO_4440 (O_4440,N_49424,N_49150);
or UO_4441 (O_4441,N_49010,N_49638);
and UO_4442 (O_4442,N_49581,N_49745);
and UO_4443 (O_4443,N_49017,N_49694);
or UO_4444 (O_4444,N_49012,N_49568);
nand UO_4445 (O_4445,N_49198,N_49231);
nor UO_4446 (O_4446,N_49372,N_49505);
nor UO_4447 (O_4447,N_49632,N_49700);
nand UO_4448 (O_4448,N_49727,N_49413);
nand UO_4449 (O_4449,N_49753,N_49611);
xor UO_4450 (O_4450,N_49590,N_49008);
nor UO_4451 (O_4451,N_49255,N_49077);
nor UO_4452 (O_4452,N_49958,N_49708);
and UO_4453 (O_4453,N_49372,N_49181);
nand UO_4454 (O_4454,N_49464,N_49952);
or UO_4455 (O_4455,N_49719,N_49761);
or UO_4456 (O_4456,N_49113,N_49274);
xor UO_4457 (O_4457,N_49946,N_49253);
and UO_4458 (O_4458,N_49690,N_49348);
or UO_4459 (O_4459,N_49218,N_49350);
nor UO_4460 (O_4460,N_49170,N_49262);
and UO_4461 (O_4461,N_49487,N_49404);
and UO_4462 (O_4462,N_49467,N_49315);
or UO_4463 (O_4463,N_49835,N_49830);
and UO_4464 (O_4464,N_49873,N_49028);
nand UO_4465 (O_4465,N_49932,N_49260);
xor UO_4466 (O_4466,N_49506,N_49476);
nor UO_4467 (O_4467,N_49075,N_49573);
nor UO_4468 (O_4468,N_49932,N_49921);
or UO_4469 (O_4469,N_49868,N_49836);
or UO_4470 (O_4470,N_49909,N_49953);
and UO_4471 (O_4471,N_49105,N_49869);
or UO_4472 (O_4472,N_49790,N_49763);
nand UO_4473 (O_4473,N_49065,N_49621);
xor UO_4474 (O_4474,N_49357,N_49538);
xor UO_4475 (O_4475,N_49874,N_49752);
xnor UO_4476 (O_4476,N_49229,N_49747);
nor UO_4477 (O_4477,N_49043,N_49401);
nand UO_4478 (O_4478,N_49834,N_49795);
nor UO_4479 (O_4479,N_49706,N_49050);
and UO_4480 (O_4480,N_49590,N_49200);
xor UO_4481 (O_4481,N_49852,N_49666);
nand UO_4482 (O_4482,N_49582,N_49537);
or UO_4483 (O_4483,N_49764,N_49656);
and UO_4484 (O_4484,N_49071,N_49418);
or UO_4485 (O_4485,N_49102,N_49522);
or UO_4486 (O_4486,N_49005,N_49480);
xnor UO_4487 (O_4487,N_49539,N_49234);
and UO_4488 (O_4488,N_49582,N_49672);
and UO_4489 (O_4489,N_49357,N_49175);
or UO_4490 (O_4490,N_49788,N_49455);
nand UO_4491 (O_4491,N_49624,N_49614);
or UO_4492 (O_4492,N_49510,N_49114);
xor UO_4493 (O_4493,N_49095,N_49392);
xnor UO_4494 (O_4494,N_49496,N_49530);
nor UO_4495 (O_4495,N_49119,N_49600);
and UO_4496 (O_4496,N_49233,N_49111);
or UO_4497 (O_4497,N_49555,N_49027);
or UO_4498 (O_4498,N_49786,N_49684);
nand UO_4499 (O_4499,N_49761,N_49934);
xnor UO_4500 (O_4500,N_49313,N_49286);
nand UO_4501 (O_4501,N_49387,N_49574);
xor UO_4502 (O_4502,N_49693,N_49441);
nor UO_4503 (O_4503,N_49093,N_49850);
xnor UO_4504 (O_4504,N_49256,N_49634);
or UO_4505 (O_4505,N_49068,N_49019);
nor UO_4506 (O_4506,N_49561,N_49086);
nand UO_4507 (O_4507,N_49382,N_49550);
nor UO_4508 (O_4508,N_49891,N_49651);
or UO_4509 (O_4509,N_49790,N_49588);
nor UO_4510 (O_4510,N_49460,N_49027);
xnor UO_4511 (O_4511,N_49649,N_49179);
xor UO_4512 (O_4512,N_49376,N_49046);
nor UO_4513 (O_4513,N_49319,N_49119);
nand UO_4514 (O_4514,N_49887,N_49769);
and UO_4515 (O_4515,N_49092,N_49720);
and UO_4516 (O_4516,N_49154,N_49561);
xor UO_4517 (O_4517,N_49701,N_49865);
and UO_4518 (O_4518,N_49417,N_49519);
nor UO_4519 (O_4519,N_49421,N_49510);
and UO_4520 (O_4520,N_49143,N_49959);
xnor UO_4521 (O_4521,N_49572,N_49028);
and UO_4522 (O_4522,N_49752,N_49726);
and UO_4523 (O_4523,N_49398,N_49606);
nand UO_4524 (O_4524,N_49258,N_49675);
nor UO_4525 (O_4525,N_49069,N_49571);
nand UO_4526 (O_4526,N_49292,N_49969);
xnor UO_4527 (O_4527,N_49325,N_49278);
or UO_4528 (O_4528,N_49124,N_49710);
xor UO_4529 (O_4529,N_49302,N_49948);
and UO_4530 (O_4530,N_49355,N_49272);
and UO_4531 (O_4531,N_49614,N_49069);
or UO_4532 (O_4532,N_49280,N_49440);
and UO_4533 (O_4533,N_49401,N_49815);
and UO_4534 (O_4534,N_49176,N_49264);
nor UO_4535 (O_4535,N_49615,N_49405);
or UO_4536 (O_4536,N_49283,N_49737);
xnor UO_4537 (O_4537,N_49581,N_49086);
nand UO_4538 (O_4538,N_49759,N_49716);
or UO_4539 (O_4539,N_49995,N_49290);
nand UO_4540 (O_4540,N_49012,N_49036);
nor UO_4541 (O_4541,N_49028,N_49062);
nor UO_4542 (O_4542,N_49239,N_49731);
nand UO_4543 (O_4543,N_49328,N_49697);
and UO_4544 (O_4544,N_49576,N_49656);
nand UO_4545 (O_4545,N_49051,N_49417);
xor UO_4546 (O_4546,N_49975,N_49384);
and UO_4547 (O_4547,N_49017,N_49916);
xor UO_4548 (O_4548,N_49480,N_49864);
nand UO_4549 (O_4549,N_49649,N_49392);
xnor UO_4550 (O_4550,N_49644,N_49023);
nor UO_4551 (O_4551,N_49611,N_49211);
xor UO_4552 (O_4552,N_49013,N_49298);
xnor UO_4553 (O_4553,N_49378,N_49393);
and UO_4554 (O_4554,N_49201,N_49623);
nor UO_4555 (O_4555,N_49298,N_49818);
nand UO_4556 (O_4556,N_49867,N_49511);
nand UO_4557 (O_4557,N_49450,N_49714);
nor UO_4558 (O_4558,N_49684,N_49969);
or UO_4559 (O_4559,N_49204,N_49966);
and UO_4560 (O_4560,N_49934,N_49526);
and UO_4561 (O_4561,N_49965,N_49165);
xnor UO_4562 (O_4562,N_49599,N_49116);
nand UO_4563 (O_4563,N_49422,N_49115);
or UO_4564 (O_4564,N_49753,N_49430);
and UO_4565 (O_4565,N_49277,N_49569);
and UO_4566 (O_4566,N_49403,N_49747);
nand UO_4567 (O_4567,N_49402,N_49442);
nand UO_4568 (O_4568,N_49063,N_49203);
nor UO_4569 (O_4569,N_49711,N_49841);
and UO_4570 (O_4570,N_49904,N_49023);
xor UO_4571 (O_4571,N_49319,N_49098);
nor UO_4572 (O_4572,N_49020,N_49178);
and UO_4573 (O_4573,N_49493,N_49365);
and UO_4574 (O_4574,N_49301,N_49914);
nand UO_4575 (O_4575,N_49054,N_49144);
or UO_4576 (O_4576,N_49626,N_49883);
xor UO_4577 (O_4577,N_49844,N_49980);
and UO_4578 (O_4578,N_49563,N_49241);
or UO_4579 (O_4579,N_49426,N_49996);
nor UO_4580 (O_4580,N_49159,N_49505);
nand UO_4581 (O_4581,N_49524,N_49643);
and UO_4582 (O_4582,N_49882,N_49275);
nand UO_4583 (O_4583,N_49345,N_49845);
nand UO_4584 (O_4584,N_49432,N_49125);
nor UO_4585 (O_4585,N_49267,N_49622);
and UO_4586 (O_4586,N_49468,N_49405);
or UO_4587 (O_4587,N_49209,N_49513);
and UO_4588 (O_4588,N_49966,N_49169);
xnor UO_4589 (O_4589,N_49826,N_49138);
nand UO_4590 (O_4590,N_49238,N_49021);
xor UO_4591 (O_4591,N_49118,N_49621);
nor UO_4592 (O_4592,N_49884,N_49330);
xor UO_4593 (O_4593,N_49351,N_49403);
nand UO_4594 (O_4594,N_49654,N_49903);
xor UO_4595 (O_4595,N_49786,N_49552);
or UO_4596 (O_4596,N_49097,N_49897);
or UO_4597 (O_4597,N_49419,N_49507);
xor UO_4598 (O_4598,N_49916,N_49676);
xor UO_4599 (O_4599,N_49505,N_49071);
or UO_4600 (O_4600,N_49245,N_49922);
and UO_4601 (O_4601,N_49603,N_49351);
and UO_4602 (O_4602,N_49299,N_49365);
and UO_4603 (O_4603,N_49342,N_49370);
or UO_4604 (O_4604,N_49797,N_49970);
nor UO_4605 (O_4605,N_49835,N_49035);
or UO_4606 (O_4606,N_49646,N_49701);
nand UO_4607 (O_4607,N_49024,N_49295);
nand UO_4608 (O_4608,N_49679,N_49090);
xor UO_4609 (O_4609,N_49571,N_49773);
nor UO_4610 (O_4610,N_49488,N_49554);
nor UO_4611 (O_4611,N_49628,N_49058);
nand UO_4612 (O_4612,N_49697,N_49555);
and UO_4613 (O_4613,N_49466,N_49948);
nor UO_4614 (O_4614,N_49687,N_49367);
nand UO_4615 (O_4615,N_49641,N_49065);
or UO_4616 (O_4616,N_49528,N_49445);
nor UO_4617 (O_4617,N_49723,N_49184);
and UO_4618 (O_4618,N_49643,N_49252);
and UO_4619 (O_4619,N_49181,N_49191);
xnor UO_4620 (O_4620,N_49519,N_49474);
or UO_4621 (O_4621,N_49285,N_49447);
or UO_4622 (O_4622,N_49689,N_49078);
or UO_4623 (O_4623,N_49503,N_49373);
or UO_4624 (O_4624,N_49961,N_49326);
and UO_4625 (O_4625,N_49508,N_49364);
nor UO_4626 (O_4626,N_49825,N_49444);
or UO_4627 (O_4627,N_49794,N_49088);
nor UO_4628 (O_4628,N_49090,N_49510);
and UO_4629 (O_4629,N_49086,N_49339);
xnor UO_4630 (O_4630,N_49904,N_49696);
and UO_4631 (O_4631,N_49745,N_49269);
xnor UO_4632 (O_4632,N_49964,N_49942);
and UO_4633 (O_4633,N_49996,N_49069);
nand UO_4634 (O_4634,N_49387,N_49558);
xnor UO_4635 (O_4635,N_49173,N_49312);
or UO_4636 (O_4636,N_49293,N_49195);
nand UO_4637 (O_4637,N_49073,N_49807);
xnor UO_4638 (O_4638,N_49761,N_49669);
nand UO_4639 (O_4639,N_49839,N_49622);
xor UO_4640 (O_4640,N_49487,N_49189);
xor UO_4641 (O_4641,N_49073,N_49042);
nand UO_4642 (O_4642,N_49534,N_49851);
nor UO_4643 (O_4643,N_49893,N_49717);
or UO_4644 (O_4644,N_49998,N_49021);
xnor UO_4645 (O_4645,N_49399,N_49247);
xnor UO_4646 (O_4646,N_49188,N_49988);
nand UO_4647 (O_4647,N_49281,N_49337);
xor UO_4648 (O_4648,N_49937,N_49084);
or UO_4649 (O_4649,N_49705,N_49064);
nor UO_4650 (O_4650,N_49414,N_49124);
nor UO_4651 (O_4651,N_49211,N_49901);
or UO_4652 (O_4652,N_49988,N_49287);
nor UO_4653 (O_4653,N_49217,N_49810);
xnor UO_4654 (O_4654,N_49497,N_49868);
xnor UO_4655 (O_4655,N_49542,N_49099);
and UO_4656 (O_4656,N_49256,N_49170);
nor UO_4657 (O_4657,N_49003,N_49501);
or UO_4658 (O_4658,N_49748,N_49412);
xnor UO_4659 (O_4659,N_49563,N_49384);
nand UO_4660 (O_4660,N_49247,N_49607);
or UO_4661 (O_4661,N_49874,N_49096);
nor UO_4662 (O_4662,N_49353,N_49271);
and UO_4663 (O_4663,N_49321,N_49422);
nand UO_4664 (O_4664,N_49873,N_49334);
nand UO_4665 (O_4665,N_49819,N_49591);
nand UO_4666 (O_4666,N_49668,N_49746);
and UO_4667 (O_4667,N_49591,N_49546);
xnor UO_4668 (O_4668,N_49717,N_49879);
nor UO_4669 (O_4669,N_49704,N_49174);
xnor UO_4670 (O_4670,N_49819,N_49783);
xor UO_4671 (O_4671,N_49701,N_49861);
and UO_4672 (O_4672,N_49163,N_49382);
nand UO_4673 (O_4673,N_49989,N_49760);
xor UO_4674 (O_4674,N_49589,N_49102);
nand UO_4675 (O_4675,N_49466,N_49779);
and UO_4676 (O_4676,N_49979,N_49128);
nand UO_4677 (O_4677,N_49026,N_49770);
and UO_4678 (O_4678,N_49238,N_49905);
or UO_4679 (O_4679,N_49434,N_49846);
or UO_4680 (O_4680,N_49200,N_49530);
and UO_4681 (O_4681,N_49691,N_49850);
or UO_4682 (O_4682,N_49885,N_49829);
or UO_4683 (O_4683,N_49135,N_49955);
and UO_4684 (O_4684,N_49349,N_49284);
nor UO_4685 (O_4685,N_49002,N_49023);
and UO_4686 (O_4686,N_49049,N_49225);
or UO_4687 (O_4687,N_49531,N_49334);
and UO_4688 (O_4688,N_49879,N_49720);
xor UO_4689 (O_4689,N_49929,N_49023);
nor UO_4690 (O_4690,N_49918,N_49251);
or UO_4691 (O_4691,N_49395,N_49937);
xor UO_4692 (O_4692,N_49870,N_49856);
nor UO_4693 (O_4693,N_49718,N_49120);
or UO_4694 (O_4694,N_49809,N_49464);
or UO_4695 (O_4695,N_49073,N_49817);
or UO_4696 (O_4696,N_49360,N_49956);
nor UO_4697 (O_4697,N_49961,N_49452);
nand UO_4698 (O_4698,N_49777,N_49757);
nand UO_4699 (O_4699,N_49863,N_49228);
xnor UO_4700 (O_4700,N_49586,N_49013);
and UO_4701 (O_4701,N_49367,N_49837);
nand UO_4702 (O_4702,N_49999,N_49039);
or UO_4703 (O_4703,N_49304,N_49246);
nor UO_4704 (O_4704,N_49688,N_49531);
and UO_4705 (O_4705,N_49684,N_49184);
xor UO_4706 (O_4706,N_49973,N_49371);
or UO_4707 (O_4707,N_49679,N_49079);
and UO_4708 (O_4708,N_49664,N_49553);
xor UO_4709 (O_4709,N_49327,N_49704);
nor UO_4710 (O_4710,N_49590,N_49495);
xnor UO_4711 (O_4711,N_49147,N_49628);
xnor UO_4712 (O_4712,N_49406,N_49555);
nor UO_4713 (O_4713,N_49060,N_49212);
and UO_4714 (O_4714,N_49960,N_49565);
and UO_4715 (O_4715,N_49136,N_49323);
and UO_4716 (O_4716,N_49211,N_49691);
nor UO_4717 (O_4717,N_49298,N_49073);
or UO_4718 (O_4718,N_49223,N_49170);
nand UO_4719 (O_4719,N_49964,N_49553);
xnor UO_4720 (O_4720,N_49641,N_49718);
nand UO_4721 (O_4721,N_49423,N_49801);
or UO_4722 (O_4722,N_49474,N_49408);
nor UO_4723 (O_4723,N_49681,N_49178);
xor UO_4724 (O_4724,N_49540,N_49908);
xnor UO_4725 (O_4725,N_49317,N_49637);
and UO_4726 (O_4726,N_49878,N_49891);
or UO_4727 (O_4727,N_49462,N_49638);
nor UO_4728 (O_4728,N_49876,N_49024);
xor UO_4729 (O_4729,N_49748,N_49939);
nand UO_4730 (O_4730,N_49044,N_49449);
nand UO_4731 (O_4731,N_49437,N_49191);
xnor UO_4732 (O_4732,N_49751,N_49706);
nor UO_4733 (O_4733,N_49476,N_49207);
xor UO_4734 (O_4734,N_49537,N_49319);
and UO_4735 (O_4735,N_49376,N_49601);
nor UO_4736 (O_4736,N_49484,N_49101);
xor UO_4737 (O_4737,N_49201,N_49663);
xor UO_4738 (O_4738,N_49993,N_49155);
xor UO_4739 (O_4739,N_49032,N_49722);
xor UO_4740 (O_4740,N_49720,N_49608);
nor UO_4741 (O_4741,N_49628,N_49993);
xnor UO_4742 (O_4742,N_49139,N_49527);
xor UO_4743 (O_4743,N_49867,N_49789);
nor UO_4744 (O_4744,N_49913,N_49316);
or UO_4745 (O_4745,N_49827,N_49000);
nand UO_4746 (O_4746,N_49129,N_49714);
nor UO_4747 (O_4747,N_49459,N_49676);
xor UO_4748 (O_4748,N_49977,N_49991);
and UO_4749 (O_4749,N_49439,N_49730);
nand UO_4750 (O_4750,N_49212,N_49976);
or UO_4751 (O_4751,N_49004,N_49108);
xor UO_4752 (O_4752,N_49175,N_49134);
and UO_4753 (O_4753,N_49938,N_49404);
or UO_4754 (O_4754,N_49247,N_49561);
xor UO_4755 (O_4755,N_49837,N_49361);
and UO_4756 (O_4756,N_49696,N_49740);
nand UO_4757 (O_4757,N_49136,N_49055);
xor UO_4758 (O_4758,N_49260,N_49252);
xnor UO_4759 (O_4759,N_49664,N_49801);
and UO_4760 (O_4760,N_49476,N_49261);
or UO_4761 (O_4761,N_49350,N_49214);
xnor UO_4762 (O_4762,N_49752,N_49742);
nor UO_4763 (O_4763,N_49446,N_49897);
xnor UO_4764 (O_4764,N_49007,N_49323);
and UO_4765 (O_4765,N_49208,N_49527);
xor UO_4766 (O_4766,N_49859,N_49914);
xnor UO_4767 (O_4767,N_49346,N_49222);
or UO_4768 (O_4768,N_49972,N_49782);
or UO_4769 (O_4769,N_49059,N_49079);
and UO_4770 (O_4770,N_49122,N_49707);
nand UO_4771 (O_4771,N_49846,N_49177);
and UO_4772 (O_4772,N_49186,N_49570);
and UO_4773 (O_4773,N_49688,N_49454);
nor UO_4774 (O_4774,N_49308,N_49506);
nor UO_4775 (O_4775,N_49941,N_49316);
xor UO_4776 (O_4776,N_49850,N_49087);
or UO_4777 (O_4777,N_49035,N_49240);
or UO_4778 (O_4778,N_49522,N_49163);
xor UO_4779 (O_4779,N_49463,N_49971);
nor UO_4780 (O_4780,N_49449,N_49645);
and UO_4781 (O_4781,N_49752,N_49680);
nand UO_4782 (O_4782,N_49889,N_49467);
nand UO_4783 (O_4783,N_49241,N_49660);
and UO_4784 (O_4784,N_49682,N_49201);
and UO_4785 (O_4785,N_49837,N_49017);
nor UO_4786 (O_4786,N_49452,N_49711);
xor UO_4787 (O_4787,N_49960,N_49089);
nor UO_4788 (O_4788,N_49216,N_49312);
or UO_4789 (O_4789,N_49427,N_49892);
nor UO_4790 (O_4790,N_49627,N_49563);
nor UO_4791 (O_4791,N_49397,N_49011);
xnor UO_4792 (O_4792,N_49508,N_49452);
and UO_4793 (O_4793,N_49160,N_49209);
xor UO_4794 (O_4794,N_49081,N_49384);
nand UO_4795 (O_4795,N_49110,N_49390);
or UO_4796 (O_4796,N_49509,N_49644);
nand UO_4797 (O_4797,N_49824,N_49149);
nor UO_4798 (O_4798,N_49093,N_49057);
or UO_4799 (O_4799,N_49805,N_49761);
nor UO_4800 (O_4800,N_49495,N_49736);
and UO_4801 (O_4801,N_49589,N_49288);
and UO_4802 (O_4802,N_49267,N_49777);
nand UO_4803 (O_4803,N_49750,N_49933);
and UO_4804 (O_4804,N_49624,N_49340);
or UO_4805 (O_4805,N_49827,N_49519);
or UO_4806 (O_4806,N_49671,N_49479);
and UO_4807 (O_4807,N_49309,N_49498);
and UO_4808 (O_4808,N_49000,N_49266);
xor UO_4809 (O_4809,N_49219,N_49880);
xnor UO_4810 (O_4810,N_49485,N_49802);
or UO_4811 (O_4811,N_49766,N_49955);
or UO_4812 (O_4812,N_49791,N_49288);
nand UO_4813 (O_4813,N_49350,N_49139);
and UO_4814 (O_4814,N_49406,N_49769);
and UO_4815 (O_4815,N_49267,N_49723);
nor UO_4816 (O_4816,N_49539,N_49163);
nand UO_4817 (O_4817,N_49135,N_49975);
or UO_4818 (O_4818,N_49963,N_49437);
nor UO_4819 (O_4819,N_49251,N_49829);
and UO_4820 (O_4820,N_49243,N_49455);
nand UO_4821 (O_4821,N_49384,N_49125);
and UO_4822 (O_4822,N_49661,N_49537);
xor UO_4823 (O_4823,N_49029,N_49161);
and UO_4824 (O_4824,N_49049,N_49764);
nand UO_4825 (O_4825,N_49118,N_49251);
nor UO_4826 (O_4826,N_49729,N_49485);
nand UO_4827 (O_4827,N_49008,N_49818);
nand UO_4828 (O_4828,N_49356,N_49753);
and UO_4829 (O_4829,N_49872,N_49096);
nor UO_4830 (O_4830,N_49328,N_49720);
nand UO_4831 (O_4831,N_49030,N_49066);
xnor UO_4832 (O_4832,N_49092,N_49679);
nor UO_4833 (O_4833,N_49370,N_49019);
and UO_4834 (O_4834,N_49526,N_49339);
and UO_4835 (O_4835,N_49634,N_49589);
nand UO_4836 (O_4836,N_49113,N_49873);
or UO_4837 (O_4837,N_49785,N_49247);
or UO_4838 (O_4838,N_49531,N_49145);
or UO_4839 (O_4839,N_49667,N_49884);
and UO_4840 (O_4840,N_49450,N_49690);
nand UO_4841 (O_4841,N_49797,N_49658);
nand UO_4842 (O_4842,N_49652,N_49741);
nor UO_4843 (O_4843,N_49968,N_49196);
and UO_4844 (O_4844,N_49187,N_49176);
and UO_4845 (O_4845,N_49110,N_49491);
nand UO_4846 (O_4846,N_49671,N_49845);
or UO_4847 (O_4847,N_49052,N_49579);
xor UO_4848 (O_4848,N_49871,N_49619);
or UO_4849 (O_4849,N_49135,N_49917);
and UO_4850 (O_4850,N_49755,N_49252);
nor UO_4851 (O_4851,N_49839,N_49037);
or UO_4852 (O_4852,N_49086,N_49711);
xor UO_4853 (O_4853,N_49270,N_49298);
nand UO_4854 (O_4854,N_49041,N_49825);
nor UO_4855 (O_4855,N_49893,N_49549);
xor UO_4856 (O_4856,N_49581,N_49653);
nand UO_4857 (O_4857,N_49567,N_49358);
or UO_4858 (O_4858,N_49058,N_49286);
xnor UO_4859 (O_4859,N_49429,N_49985);
or UO_4860 (O_4860,N_49723,N_49249);
or UO_4861 (O_4861,N_49867,N_49074);
or UO_4862 (O_4862,N_49045,N_49465);
and UO_4863 (O_4863,N_49595,N_49077);
xor UO_4864 (O_4864,N_49679,N_49516);
xnor UO_4865 (O_4865,N_49767,N_49285);
nor UO_4866 (O_4866,N_49750,N_49493);
xor UO_4867 (O_4867,N_49130,N_49498);
nor UO_4868 (O_4868,N_49745,N_49504);
and UO_4869 (O_4869,N_49045,N_49157);
and UO_4870 (O_4870,N_49845,N_49234);
nand UO_4871 (O_4871,N_49130,N_49795);
and UO_4872 (O_4872,N_49782,N_49274);
and UO_4873 (O_4873,N_49325,N_49611);
or UO_4874 (O_4874,N_49341,N_49061);
nand UO_4875 (O_4875,N_49208,N_49540);
or UO_4876 (O_4876,N_49486,N_49348);
xor UO_4877 (O_4877,N_49658,N_49534);
xnor UO_4878 (O_4878,N_49908,N_49269);
xnor UO_4879 (O_4879,N_49622,N_49122);
nor UO_4880 (O_4880,N_49338,N_49993);
and UO_4881 (O_4881,N_49542,N_49256);
or UO_4882 (O_4882,N_49063,N_49758);
nand UO_4883 (O_4883,N_49146,N_49905);
nand UO_4884 (O_4884,N_49478,N_49019);
nor UO_4885 (O_4885,N_49537,N_49891);
xnor UO_4886 (O_4886,N_49883,N_49711);
nor UO_4887 (O_4887,N_49327,N_49937);
nor UO_4888 (O_4888,N_49618,N_49180);
and UO_4889 (O_4889,N_49807,N_49339);
and UO_4890 (O_4890,N_49034,N_49216);
nand UO_4891 (O_4891,N_49622,N_49847);
xnor UO_4892 (O_4892,N_49737,N_49533);
nand UO_4893 (O_4893,N_49946,N_49645);
xor UO_4894 (O_4894,N_49908,N_49640);
and UO_4895 (O_4895,N_49287,N_49829);
xnor UO_4896 (O_4896,N_49450,N_49846);
xor UO_4897 (O_4897,N_49122,N_49362);
and UO_4898 (O_4898,N_49437,N_49471);
or UO_4899 (O_4899,N_49868,N_49085);
or UO_4900 (O_4900,N_49398,N_49863);
nor UO_4901 (O_4901,N_49452,N_49499);
or UO_4902 (O_4902,N_49653,N_49507);
or UO_4903 (O_4903,N_49964,N_49116);
nor UO_4904 (O_4904,N_49772,N_49625);
nand UO_4905 (O_4905,N_49619,N_49567);
and UO_4906 (O_4906,N_49556,N_49971);
nor UO_4907 (O_4907,N_49789,N_49224);
nand UO_4908 (O_4908,N_49627,N_49353);
and UO_4909 (O_4909,N_49482,N_49385);
nand UO_4910 (O_4910,N_49024,N_49678);
xnor UO_4911 (O_4911,N_49460,N_49397);
and UO_4912 (O_4912,N_49238,N_49438);
nand UO_4913 (O_4913,N_49668,N_49672);
xor UO_4914 (O_4914,N_49776,N_49318);
or UO_4915 (O_4915,N_49815,N_49934);
nor UO_4916 (O_4916,N_49396,N_49417);
and UO_4917 (O_4917,N_49188,N_49982);
and UO_4918 (O_4918,N_49531,N_49876);
and UO_4919 (O_4919,N_49077,N_49151);
nand UO_4920 (O_4920,N_49159,N_49758);
nand UO_4921 (O_4921,N_49019,N_49857);
nor UO_4922 (O_4922,N_49015,N_49802);
or UO_4923 (O_4923,N_49066,N_49076);
nor UO_4924 (O_4924,N_49117,N_49460);
xor UO_4925 (O_4925,N_49281,N_49216);
and UO_4926 (O_4926,N_49849,N_49347);
or UO_4927 (O_4927,N_49955,N_49170);
xnor UO_4928 (O_4928,N_49605,N_49776);
and UO_4929 (O_4929,N_49454,N_49538);
nand UO_4930 (O_4930,N_49000,N_49181);
nor UO_4931 (O_4931,N_49130,N_49573);
nor UO_4932 (O_4932,N_49482,N_49020);
nor UO_4933 (O_4933,N_49136,N_49369);
or UO_4934 (O_4934,N_49460,N_49587);
nor UO_4935 (O_4935,N_49232,N_49875);
nand UO_4936 (O_4936,N_49399,N_49942);
and UO_4937 (O_4937,N_49262,N_49691);
nand UO_4938 (O_4938,N_49334,N_49750);
and UO_4939 (O_4939,N_49607,N_49974);
and UO_4940 (O_4940,N_49087,N_49135);
xnor UO_4941 (O_4941,N_49033,N_49173);
xor UO_4942 (O_4942,N_49234,N_49726);
nand UO_4943 (O_4943,N_49127,N_49677);
or UO_4944 (O_4944,N_49037,N_49521);
xnor UO_4945 (O_4945,N_49416,N_49021);
xor UO_4946 (O_4946,N_49334,N_49854);
nor UO_4947 (O_4947,N_49656,N_49781);
or UO_4948 (O_4948,N_49821,N_49058);
xor UO_4949 (O_4949,N_49546,N_49479);
xor UO_4950 (O_4950,N_49760,N_49985);
or UO_4951 (O_4951,N_49075,N_49213);
and UO_4952 (O_4952,N_49368,N_49969);
xnor UO_4953 (O_4953,N_49940,N_49868);
nand UO_4954 (O_4954,N_49414,N_49692);
nor UO_4955 (O_4955,N_49495,N_49296);
nand UO_4956 (O_4956,N_49062,N_49857);
xor UO_4957 (O_4957,N_49317,N_49613);
xor UO_4958 (O_4958,N_49191,N_49660);
nand UO_4959 (O_4959,N_49596,N_49994);
nand UO_4960 (O_4960,N_49317,N_49497);
xor UO_4961 (O_4961,N_49379,N_49840);
or UO_4962 (O_4962,N_49966,N_49095);
nand UO_4963 (O_4963,N_49390,N_49302);
or UO_4964 (O_4964,N_49666,N_49774);
nor UO_4965 (O_4965,N_49719,N_49462);
or UO_4966 (O_4966,N_49776,N_49802);
nor UO_4967 (O_4967,N_49061,N_49967);
and UO_4968 (O_4968,N_49436,N_49434);
nor UO_4969 (O_4969,N_49683,N_49934);
nand UO_4970 (O_4970,N_49589,N_49924);
xor UO_4971 (O_4971,N_49830,N_49704);
nor UO_4972 (O_4972,N_49742,N_49452);
or UO_4973 (O_4973,N_49955,N_49217);
nor UO_4974 (O_4974,N_49340,N_49929);
nand UO_4975 (O_4975,N_49600,N_49117);
and UO_4976 (O_4976,N_49047,N_49622);
and UO_4977 (O_4977,N_49338,N_49780);
and UO_4978 (O_4978,N_49690,N_49518);
nor UO_4979 (O_4979,N_49732,N_49314);
nand UO_4980 (O_4980,N_49064,N_49025);
nand UO_4981 (O_4981,N_49067,N_49929);
nand UO_4982 (O_4982,N_49323,N_49049);
nand UO_4983 (O_4983,N_49420,N_49244);
xnor UO_4984 (O_4984,N_49891,N_49341);
nand UO_4985 (O_4985,N_49844,N_49322);
nand UO_4986 (O_4986,N_49599,N_49704);
xnor UO_4987 (O_4987,N_49361,N_49514);
nand UO_4988 (O_4988,N_49469,N_49059);
and UO_4989 (O_4989,N_49143,N_49326);
xor UO_4990 (O_4990,N_49322,N_49648);
or UO_4991 (O_4991,N_49072,N_49863);
and UO_4992 (O_4992,N_49304,N_49656);
and UO_4993 (O_4993,N_49977,N_49202);
or UO_4994 (O_4994,N_49470,N_49391);
nand UO_4995 (O_4995,N_49220,N_49428);
nand UO_4996 (O_4996,N_49974,N_49255);
nand UO_4997 (O_4997,N_49153,N_49332);
and UO_4998 (O_4998,N_49712,N_49515);
nand UO_4999 (O_4999,N_49150,N_49255);
endmodule